
module fpSqrt(rst, clk, ce, ld, \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] , \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] , \o[24] , \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] , \o[32] , \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] , \o[40] , \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] , \o[48] , \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] , \o[56] , \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63] , \o[64] , \o[65] , \o[66] , \o[67] , \o[68] , \o[69] , \o[70] , \o[71] , \o[72] , \o[73] , \o[74] , \o[75] , \o[76] , \o[77] , \o[78] , \o[79] , \o[80] , \o[81] , \o[82] , \o[83] , \o[84] , \o[85] , \o[86] , \o[87] , \o[88] , \o[89] , \o[90] , \o[91] , \o[92] , \o[93] , \o[94] , \o[95] , \o[96] , \o[97] , \o[98] , \o[99] , \o[100] , \o[101] , \o[102] , \o[103] , \o[104] , \o[105] , \o[106] , \o[107] , \o[108] , \o[109] , \o[110] , \o[111] , \o[112] , \o[113] , \o[114] , \o[115] , \o[116] , \o[117] , \o[118] , \o[119] , \o[120] , \o[121] , \o[122] , \o[123] , \o[124] , \o[125] , \o[126] , \o[127] , \o[128] , \o[129] , \o[130] , \o[131] , \o[132] , \o[133] , \o[134] , \o[135] , \o[136] , \o[137] , \o[138] , \o[139] , \o[140] , \o[141] , \o[142] , \o[143] , \o[144] , \o[145] , \o[146] , \o[147] , \o[148] , \o[149] , \o[150] , \o[151] , \o[152] , \o[153] , \o[154] , \o[155] , \o[156] , \o[157] , \o[158] , \o[159] , \o[160] , \o[161] , \o[162] , \o[163] , \o[164] , \o[165] , \o[166] , \o[167] , \o[168] , \o[169] , \o[170] , \o[171] , \o[172] , \o[173] , \o[174] , \o[175] , \o[176] , \o[177] , \o[178] , \o[179] , \o[180] , \o[181] , \o[182] , \o[183] , \o[184] , \o[185] , \o[186] , \o[187] , \o[188] , \o[189] , \o[190] , \o[191] , \o[192] , \o[193] , \o[194] , \o[195] , \o[196] , \o[197] , \o[198] , \o[199] , \o[200] , \o[201] , \o[202] , \o[203] , \o[204] , \o[205] , \o[206] , \o[207] , \o[208] , \o[209] , \o[210] , \o[211] , \o[212] , \o[213] , \o[214] , \o[215] , \o[216] , \o[217] , \o[218] , \o[219] , \o[220] , \o[221] , \o[222] , \o[223] , \o[224] , \o[225] , \o[226] , \o[227] , \o[228] , \o[229] , \o[230] , \o[231] , \o[232] , \o[233] , \o[234] , \o[235] , \o[236] , \o[237] , \o[238] , \o[239] , \o[240] , \o[241] , done);
  wire _abc_64468_n1001;
  wire _abc_64468_n1002;
  wire _abc_64468_n1004;
  wire _abc_64468_n1005;
  wire _abc_64468_n1007;
  wire _abc_64468_n1008;
  wire _abc_64468_n1010;
  wire _abc_64468_n1011;
  wire _abc_64468_n1013;
  wire _abc_64468_n1014;
  wire _abc_64468_n1016;
  wire _abc_64468_n1017;
  wire _abc_64468_n1019;
  wire _abc_64468_n1020;
  wire _abc_64468_n1022;
  wire _abc_64468_n1023;
  wire _abc_64468_n1025;
  wire _abc_64468_n1026;
  wire _abc_64468_n1028;
  wire _abc_64468_n1029;
  wire _abc_64468_n1031;
  wire _abc_64468_n1032;
  wire _abc_64468_n1034;
  wire _abc_64468_n1035;
  wire _abc_64468_n1037;
  wire _abc_64468_n1038;
  wire _abc_64468_n1040;
  wire _abc_64468_n1041;
  wire _abc_64468_n1043;
  wire _abc_64468_n1044;
  wire _abc_64468_n1046;
  wire _abc_64468_n1047;
  wire _abc_64468_n1049;
  wire _abc_64468_n1050;
  wire _abc_64468_n1052;
  wire _abc_64468_n1053;
  wire _abc_64468_n1055;
  wire _abc_64468_n1056;
  wire _abc_64468_n1058;
  wire _abc_64468_n1059;
  wire _abc_64468_n1061;
  wire _abc_64468_n1062;
  wire _abc_64468_n1064;
  wire _abc_64468_n1065;
  wire _abc_64468_n1067;
  wire _abc_64468_n1068;
  wire _abc_64468_n1070;
  wire _abc_64468_n1071;
  wire _abc_64468_n1073;
  wire _abc_64468_n1074;
  wire _abc_64468_n1076;
  wire _abc_64468_n1077;
  wire _abc_64468_n1079;
  wire _abc_64468_n1080;
  wire _abc_64468_n1082;
  wire _abc_64468_n1083;
  wire _abc_64468_n1085;
  wire _abc_64468_n1086;
  wire _abc_64468_n1088;
  wire _abc_64468_n1089;
  wire _abc_64468_n1091;
  wire _abc_64468_n1092;
  wire _abc_64468_n1094;
  wire _abc_64468_n1095;
  wire _abc_64468_n1097;
  wire _abc_64468_n1098;
  wire _abc_64468_n1100;
  wire _abc_64468_n1101;
  wire _abc_64468_n1103;
  wire _abc_64468_n1104;
  wire _abc_64468_n1106;
  wire _abc_64468_n1107;
  wire _abc_64468_n1109;
  wire _abc_64468_n1110;
  wire _abc_64468_n1112;
  wire _abc_64468_n1113;
  wire _abc_64468_n1115;
  wire _abc_64468_n1116;
  wire _abc_64468_n1118;
  wire _abc_64468_n1119;
  wire _abc_64468_n1121;
  wire _abc_64468_n1122;
  wire _abc_64468_n1124;
  wire _abc_64468_n1125;
  wire _abc_64468_n1127;
  wire _abc_64468_n1128;
  wire _abc_64468_n1130;
  wire _abc_64468_n1131;
  wire _abc_64468_n1133;
  wire _abc_64468_n1134;
  wire _abc_64468_n1136;
  wire _abc_64468_n1137;
  wire _abc_64468_n1139;
  wire _abc_64468_n1140;
  wire _abc_64468_n1142;
  wire _abc_64468_n1143;
  wire _abc_64468_n1145;
  wire _abc_64468_n1146;
  wire _abc_64468_n1148;
  wire _abc_64468_n1149;
  wire _abc_64468_n1151;
  wire _abc_64468_n1152;
  wire _abc_64468_n1154;
  wire _abc_64468_n1155;
  wire _abc_64468_n1157;
  wire _abc_64468_n1158;
  wire _abc_64468_n1160;
  wire _abc_64468_n1161;
  wire _abc_64468_n1163;
  wire _abc_64468_n1164;
  wire _abc_64468_n1169;
  wire _abc_64468_n1170;
  wire _abc_64468_n1170_bF_buf0;
  wire _abc_64468_n1170_bF_buf1;
  wire _abc_64468_n1170_bF_buf2;
  wire _abc_64468_n1170_bF_buf3;
  wire _abc_64468_n1170_bF_buf4;
  wire _abc_64468_n1170_bF_buf5;
  wire _abc_64468_n1170_bF_buf6;
  wire _abc_64468_n1170_bF_buf7;
  wire _abc_64468_n1170_bF_buf8;
  wire _abc_64468_n1170_bF_buf9;
  wire _abc_64468_n1171;
  wire _abc_64468_n1173;
  wire _abc_64468_n1174;
  wire _abc_64468_n1176;
  wire _abc_64468_n1177;
  wire _abc_64468_n1179;
  wire _abc_64468_n1180;
  wire _abc_64468_n1182;
  wire _abc_64468_n1183;
  wire _abc_64468_n1185;
  wire _abc_64468_n1186;
  wire _abc_64468_n1188;
  wire _abc_64468_n1189;
  wire _abc_64468_n1191;
  wire _abc_64468_n1192;
  wire _abc_64468_n1194;
  wire _abc_64468_n1195;
  wire _abc_64468_n1197;
  wire _abc_64468_n1198;
  wire _abc_64468_n1200;
  wire _abc_64468_n1201;
  wire _abc_64468_n1203;
  wire _abc_64468_n1204;
  wire _abc_64468_n1206;
  wire _abc_64468_n1207;
  wire _abc_64468_n1209;
  wire _abc_64468_n1210;
  wire _abc_64468_n1212;
  wire _abc_64468_n1213;
  wire _abc_64468_n1215;
  wire _abc_64468_n1216;
  wire _abc_64468_n1218;
  wire _abc_64468_n1219;
  wire _abc_64468_n1221;
  wire _abc_64468_n1222;
  wire _abc_64468_n1224;
  wire _abc_64468_n1225;
  wire _abc_64468_n1227;
  wire _abc_64468_n1228;
  wire _abc_64468_n1230;
  wire _abc_64468_n1231;
  wire _abc_64468_n1233;
  wire _abc_64468_n1234;
  wire _abc_64468_n1236;
  wire _abc_64468_n1237;
  wire _abc_64468_n1239;
  wire _abc_64468_n1240;
  wire _abc_64468_n1242;
  wire _abc_64468_n1243;
  wire _abc_64468_n1245;
  wire _abc_64468_n1246;
  wire _abc_64468_n1248;
  wire _abc_64468_n1249;
  wire _abc_64468_n1251;
  wire _abc_64468_n1252;
  wire _abc_64468_n1254;
  wire _abc_64468_n1255;
  wire _abc_64468_n1257;
  wire _abc_64468_n1258;
  wire _abc_64468_n1260;
  wire _abc_64468_n1261;
  wire _abc_64468_n1263;
  wire _abc_64468_n1264;
  wire _abc_64468_n1266;
  wire _abc_64468_n1267;
  wire _abc_64468_n1269;
  wire _abc_64468_n1270;
  wire _abc_64468_n1272;
  wire _abc_64468_n1273;
  wire _abc_64468_n1275;
  wire _abc_64468_n1276;
  wire _abc_64468_n1278;
  wire _abc_64468_n1279;
  wire _abc_64468_n1281;
  wire _abc_64468_n1282;
  wire _abc_64468_n1284;
  wire _abc_64468_n1285;
  wire _abc_64468_n1287;
  wire _abc_64468_n1288;
  wire _abc_64468_n1290;
  wire _abc_64468_n1291;
  wire _abc_64468_n1293;
  wire _abc_64468_n1294;
  wire _abc_64468_n1296;
  wire _abc_64468_n1297;
  wire _abc_64468_n1299;
  wire _abc_64468_n1300;
  wire _abc_64468_n1302;
  wire _abc_64468_n1303;
  wire _abc_64468_n1305;
  wire _abc_64468_n1306;
  wire _abc_64468_n1308;
  wire _abc_64468_n1309;
  wire _abc_64468_n1311;
  wire _abc_64468_n1312;
  wire _abc_64468_n1314;
  wire _abc_64468_n1315;
  wire _abc_64468_n1317;
  wire _abc_64468_n1318;
  wire _abc_64468_n1320;
  wire _abc_64468_n1321;
  wire _abc_64468_n1323;
  wire _abc_64468_n1324;
  wire _abc_64468_n1326;
  wire _abc_64468_n1327;
  wire _abc_64468_n1329;
  wire _abc_64468_n1330;
  wire _abc_64468_n1332;
  wire _abc_64468_n1333;
  wire _abc_64468_n1335;
  wire _abc_64468_n1336;
  wire _abc_64468_n1338;
  wire _abc_64468_n1339;
  wire _abc_64468_n1341;
  wire _abc_64468_n1342;
  wire _abc_64468_n1344;
  wire _abc_64468_n1345;
  wire _abc_64468_n1347;
  wire _abc_64468_n1348;
  wire _abc_64468_n1350;
  wire _abc_64468_n1351;
  wire _abc_64468_n1353;
  wire _abc_64468_n1354;
  wire _abc_64468_n1356;
  wire _abc_64468_n1357;
  wire _abc_64468_n1359;
  wire _abc_64468_n1360;
  wire _abc_64468_n1362;
  wire _abc_64468_n1363;
  wire _abc_64468_n1365;
  wire _abc_64468_n1366;
  wire _abc_64468_n1368;
  wire _abc_64468_n1369;
  wire _abc_64468_n1371;
  wire _abc_64468_n1372;
  wire _abc_64468_n1374;
  wire _abc_64468_n1375;
  wire _abc_64468_n1377;
  wire _abc_64468_n1378;
  wire _abc_64468_n1380;
  wire _abc_64468_n1381;
  wire _abc_64468_n1383;
  wire _abc_64468_n1384;
  wire _abc_64468_n1386;
  wire _abc_64468_n1387;
  wire _abc_64468_n1389;
  wire _abc_64468_n1390;
  wire _abc_64468_n1392;
  wire _abc_64468_n1393;
  wire _abc_64468_n1395;
  wire _abc_64468_n1396;
  wire _abc_64468_n1398;
  wire _abc_64468_n1399;
  wire _abc_64468_n1401;
  wire _abc_64468_n1402;
  wire _abc_64468_n1404;
  wire _abc_64468_n1405;
  wire _abc_64468_n1407;
  wire _abc_64468_n1408;
  wire _abc_64468_n1410;
  wire _abc_64468_n1411;
  wire _abc_64468_n1413;
  wire _abc_64468_n1414;
  wire _abc_64468_n1416;
  wire _abc_64468_n1417;
  wire _abc_64468_n1419;
  wire _abc_64468_n1420;
  wire _abc_64468_n1422;
  wire _abc_64468_n1423;
  wire _abc_64468_n1425;
  wire _abc_64468_n1426;
  wire _abc_64468_n1428;
  wire _abc_64468_n1429;
  wire _abc_64468_n1431;
  wire _abc_64468_n1432;
  wire _abc_64468_n1434;
  wire _abc_64468_n1435;
  wire _abc_64468_n1437;
  wire _abc_64468_n1438;
  wire _abc_64468_n1440;
  wire _abc_64468_n1441;
  wire _abc_64468_n1443;
  wire _abc_64468_n1444;
  wire _abc_64468_n1446;
  wire _abc_64468_n1447;
  wire _abc_64468_n1449;
  wire _abc_64468_n1450;
  wire _abc_64468_n1452;
  wire _abc_64468_n1453;
  wire _abc_64468_n1455;
  wire _abc_64468_n1456;
  wire _abc_64468_n1458;
  wire _abc_64468_n1459;
  wire _abc_64468_n1461;
  wire _abc_64468_n1462;
  wire _abc_64468_n1464;
  wire _abc_64468_n1465;
  wire _abc_64468_n1467;
  wire _abc_64468_n1468;
  wire _abc_64468_n1470;
  wire _abc_64468_n1471;
  wire _abc_64468_n1473;
  wire _abc_64468_n1474;
  wire _abc_64468_n1476;
  wire _abc_64468_n1477;
  wire _abc_64468_n1479;
  wire _abc_64468_n1480;
  wire _abc_64468_n1482;
  wire _abc_64468_n1483;
  wire _abc_64468_n1485;
  wire _abc_64468_n1486;
  wire _abc_64468_n1488;
  wire _abc_64468_n1489;
  wire _abc_64468_n1491;
  wire _abc_64468_n1492;
  wire _abc_64468_n1494;
  wire _abc_64468_n1495;
  wire _abc_64468_n1497;
  wire _abc_64468_n1498;
  wire _abc_64468_n1500;
  wire _abc_64468_n1501;
  wire _abc_64468_n1503;
  wire _abc_64468_n1504;
  wire _abc_64468_n1507;
  wire _abc_64468_n1508;
  wire _abc_64468_n1509;
  wire _abc_64468_n1510;
  wire _abc_64468_n1511;
  wire _abc_64468_n1512;
  wire _abc_64468_n1514;
  wire _abc_64468_n1515;
  wire _abc_64468_n1516;
  wire _abc_64468_n1517;
  wire _abc_64468_n1518;
  wire _abc_64468_n1519;
  wire _abc_64468_n1520;
  wire _abc_64468_n1521;
  wire _abc_64468_n1523;
  wire _abc_64468_n1524;
  wire _abc_64468_n1525;
  wire _abc_64468_n1526;
  wire _abc_64468_n1527;
  wire _abc_64468_n1528;
  wire _abc_64468_n1529;
  wire _abc_64468_n1530;
  wire _abc_64468_n1531;
  wire _abc_64468_n1532;
  wire _abc_64468_n1533;
  wire _abc_64468_n1534;
  wire _abc_64468_n1535;
  wire _abc_64468_n1536;
  wire _abc_64468_n1538;
  wire _abc_64468_n1539;
  wire _abc_64468_n1540;
  wire _abc_64468_n1541;
  wire _abc_64468_n1542;
  wire _abc_64468_n1543;
  wire _abc_64468_n1544;
  wire _abc_64468_n1545;
  wire _abc_64468_n1546;
  wire _abc_64468_n1547;
  wire _abc_64468_n1548;
  wire _abc_64468_n1549;
  wire _abc_64468_n1550;
  wire _abc_64468_n1552;
  wire _abc_64468_n1553;
  wire _abc_64468_n1554;
  wire _abc_64468_n1555;
  wire _abc_64468_n1556;
  wire _abc_64468_n1557;
  wire _abc_64468_n1558;
  wire _abc_64468_n1559;
  wire _abc_64468_n1560;
  wire _abc_64468_n1561;
  wire _abc_64468_n1562;
  wire _abc_64468_n1563;
  wire _abc_64468_n1564;
  wire _abc_64468_n1566;
  wire _abc_64468_n1567;
  wire _abc_64468_n1568;
  wire _abc_64468_n1569;
  wire _abc_64468_n1570;
  wire _abc_64468_n1571;
  wire _abc_64468_n1572;
  wire _abc_64468_n1573;
  wire _abc_64468_n1574;
  wire _abc_64468_n1575;
  wire _abc_64468_n1576;
  wire _abc_64468_n1577;
  wire _abc_64468_n1579;
  wire _abc_64468_n1580;
  wire _abc_64468_n1581;
  wire _abc_64468_n1582;
  wire _abc_64468_n1583;
  wire _abc_64468_n1584;
  wire _abc_64468_n1585;
  wire _abc_64468_n1586;
  wire _abc_64468_n1587;
  wire _abc_64468_n1588;
  wire _abc_64468_n1589;
  wire _abc_64468_n1590;
  wire _abc_64468_n1591;
  wire _abc_64468_n1593;
  wire _abc_64468_n1594;
  wire _abc_64468_n1595;
  wire _abc_64468_n1596;
  wire _abc_64468_n1597;
  wire _abc_64468_n1598;
  wire _abc_64468_n1599;
  wire _abc_64468_n1600;
  wire _abc_64468_n1601;
  wire _abc_64468_n1602;
  wire _abc_64468_n1603;
  wire _abc_64468_n1604;
  wire _abc_64468_n1605;
  wire _abc_64468_n1607;
  wire _abc_64468_n1608;
  wire _abc_64468_n1609;
  wire _abc_64468_n1610;
  wire _abc_64468_n1611;
  wire _abc_64468_n1612;
  wire _abc_64468_n1613;
  wire _abc_64468_n1614;
  wire _abc_64468_n1615;
  wire _abc_64468_n1616;
  wire _abc_64468_n1617;
  wire _abc_64468_n1618;
  wire _abc_64468_n1619;
  wire _abc_64468_n1621;
  wire _abc_64468_n1622;
  wire _abc_64468_n1623;
  wire _abc_64468_n1624;
  wire _abc_64468_n1625;
  wire _abc_64468_n1626;
  wire _abc_64468_n1627;
  wire _abc_64468_n1628;
  wire _abc_64468_n1629;
  wire _abc_64468_n1630;
  wire _abc_64468_n1631;
  wire _abc_64468_n1632;
  wire _abc_64468_n1633;
  wire _abc_64468_n1635;
  wire _abc_64468_n1636;
  wire _abc_64468_n1637;
  wire _abc_64468_n1638;
  wire _abc_64468_n1639;
  wire _abc_64468_n1640;
  wire _abc_64468_n1641;
  wire _abc_64468_n1642;
  wire _abc_64468_n1643;
  wire _abc_64468_n1644;
  wire _abc_64468_n1645;
  wire _abc_64468_n1646;
  wire _abc_64468_n1647;
  wire _abc_64468_n1649;
  wire _abc_64468_n1650;
  wire _abc_64468_n1651;
  wire _abc_64468_n1652;
  wire _abc_64468_n1653;
  wire _abc_64468_n1654;
  wire _abc_64468_n1655;
  wire _abc_64468_n1656;
  wire _abc_64468_n1657;
  wire _abc_64468_n1658;
  wire _abc_64468_n1659;
  wire _abc_64468_n1660;
  wire _abc_64468_n1661;
  wire _abc_64468_n1663;
  wire _abc_64468_n1664;
  wire _abc_64468_n1665;
  wire _abc_64468_n1666;
  wire _abc_64468_n1667;
  wire _abc_64468_n1668;
  wire _abc_64468_n1669;
  wire _abc_64468_n1670;
  wire _abc_64468_n1671;
  wire _abc_64468_n1672;
  wire _abc_64468_n1673;
  wire _abc_64468_n1674;
  wire _abc_64468_n1675;
  wire _abc_64468_n1677;
  wire _abc_64468_n1678;
  wire _abc_64468_n1679;
  wire _abc_64468_n1680;
  wire _abc_64468_n1681;
  wire _abc_64468_n1682;
  wire _abc_64468_n1683;
  wire _abc_64468_n1684;
  wire _abc_64468_n1685;
  wire _abc_64468_n1686;
  wire _abc_64468_n1687;
  wire _abc_64468_n1688;
  wire _abc_64468_n1690;
  wire _abc_64468_n1691;
  wire _abc_64468_n1692;
  wire _abc_64468_n1693;
  wire _abc_64468_n753;
  wire _abc_64468_n753_bF_buf0;
  wire _abc_64468_n753_bF_buf1;
  wire _abc_64468_n753_bF_buf10;
  wire _abc_64468_n753_bF_buf11;
  wire _abc_64468_n753_bF_buf12;
  wire _abc_64468_n753_bF_buf13;
  wire _abc_64468_n753_bF_buf2;
  wire _abc_64468_n753_bF_buf3;
  wire _abc_64468_n753_bF_buf4;
  wire _abc_64468_n753_bF_buf5;
  wire _abc_64468_n753_bF_buf6;
  wire _abc_64468_n753_bF_buf7;
  wire _abc_64468_n753_bF_buf8;
  wire _abc_64468_n753_bF_buf9;
  wire _abc_64468_n830;
  wire _abc_64468_n831_1;
  wire _abc_64468_n833;
  wire _abc_64468_n834;
  wire _abc_64468_n836;
  wire _abc_64468_n837;
  wire _abc_64468_n839_1;
  wire _abc_64468_n840_1;
  wire _abc_64468_n842;
  wire _abc_64468_n843;
  wire _abc_64468_n845;
  wire _abc_64468_n846;
  wire _abc_64468_n848;
  wire _abc_64468_n849;
  wire _abc_64468_n851;
  wire _abc_64468_n852;
  wire _abc_64468_n854;
  wire _abc_64468_n855;
  wire _abc_64468_n857;
  wire _abc_64468_n858;
  wire _abc_64468_n860;
  wire _abc_64468_n861;
  wire _abc_64468_n863;
  wire _abc_64468_n864;
  wire _abc_64468_n866;
  wire _abc_64468_n867;
  wire _abc_64468_n869;
  wire _abc_64468_n870;
  wire _abc_64468_n872;
  wire _abc_64468_n873;
  wire _abc_64468_n875;
  wire _abc_64468_n876;
  wire _abc_64468_n878;
  wire _abc_64468_n879;
  wire _abc_64468_n881;
  wire _abc_64468_n882;
  wire _abc_64468_n884;
  wire _abc_64468_n885;
  wire _abc_64468_n887;
  wire _abc_64468_n888;
  wire _abc_64468_n890;
  wire _abc_64468_n891;
  wire _abc_64468_n893;
  wire _abc_64468_n894;
  wire _abc_64468_n896;
  wire _abc_64468_n897;
  wire _abc_64468_n899;
  wire _abc_64468_n900;
  wire _abc_64468_n902;
  wire _abc_64468_n903;
  wire _abc_64468_n905;
  wire _abc_64468_n906;
  wire _abc_64468_n908;
  wire _abc_64468_n909;
  wire _abc_64468_n911;
  wire _abc_64468_n912;
  wire _abc_64468_n914;
  wire _abc_64468_n915;
  wire _abc_64468_n917;
  wire _abc_64468_n918;
  wire _abc_64468_n920;
  wire _abc_64468_n921;
  wire _abc_64468_n923;
  wire _abc_64468_n924;
  wire _abc_64468_n926;
  wire _abc_64468_n927;
  wire _abc_64468_n929;
  wire _abc_64468_n930;
  wire _abc_64468_n932;
  wire _abc_64468_n933;
  wire _abc_64468_n935;
  wire _abc_64468_n936;
  wire _abc_64468_n938;
  wire _abc_64468_n939;
  wire _abc_64468_n941;
  wire _abc_64468_n942;
  wire _abc_64468_n944;
  wire _abc_64468_n945;
  wire _abc_64468_n947;
  wire _abc_64468_n948;
  wire _abc_64468_n950;
  wire _abc_64468_n951;
  wire _abc_64468_n953;
  wire _abc_64468_n954;
  wire _abc_64468_n956;
  wire _abc_64468_n957;
  wire _abc_64468_n959;
  wire _abc_64468_n960;
  wire _abc_64468_n962;
  wire _abc_64468_n963;
  wire _abc_64468_n965;
  wire _abc_64468_n966;
  wire _abc_64468_n968;
  wire _abc_64468_n969;
  wire _abc_64468_n971;
  wire _abc_64468_n972;
  wire _abc_64468_n974;
  wire _abc_64468_n975;
  wire _abc_64468_n977;
  wire _abc_64468_n978;
  wire _abc_64468_n980;
  wire _abc_64468_n981;
  wire _abc_64468_n983;
  wire _abc_64468_n984;
  wire _abc_64468_n986;
  wire _abc_64468_n987;
  wire _abc_64468_n989;
  wire _abc_64468_n990;
  wire _abc_64468_n992;
  wire _abc_64468_n993;
  wire _abc_64468_n995;
  wire _abc_64468_n996;
  wire _abc_64468_n998;
  wire _abc_64468_n999;
  wire _auto_iopadmap_cc_313_execute_65412;
  wire _auto_iopadmap_cc_313_execute_65414_100_;
  wire _auto_iopadmap_cc_313_execute_65414_101_;
  wire _auto_iopadmap_cc_313_execute_65414_102_;
  wire _auto_iopadmap_cc_313_execute_65414_103_;
  wire _auto_iopadmap_cc_313_execute_65414_104_;
  wire _auto_iopadmap_cc_313_execute_65414_105_;
  wire _auto_iopadmap_cc_313_execute_65414_106_;
  wire _auto_iopadmap_cc_313_execute_65414_107_;
  wire _auto_iopadmap_cc_313_execute_65414_108_;
  wire _auto_iopadmap_cc_313_execute_65414_109_;
  wire _auto_iopadmap_cc_313_execute_65414_110_;
  wire _auto_iopadmap_cc_313_execute_65414_111_;
  wire _auto_iopadmap_cc_313_execute_65414_112_;
  wire _auto_iopadmap_cc_313_execute_65414_113_;
  wire _auto_iopadmap_cc_313_execute_65414_114_;
  wire _auto_iopadmap_cc_313_execute_65414_115_;
  wire _auto_iopadmap_cc_313_execute_65414_116_;
  wire _auto_iopadmap_cc_313_execute_65414_117_;
  wire _auto_iopadmap_cc_313_execute_65414_118_;
  wire _auto_iopadmap_cc_313_execute_65414_119_;
  wire _auto_iopadmap_cc_313_execute_65414_120_;
  wire _auto_iopadmap_cc_313_execute_65414_121_;
  wire _auto_iopadmap_cc_313_execute_65414_122_;
  wire _auto_iopadmap_cc_313_execute_65414_123_;
  wire _auto_iopadmap_cc_313_execute_65414_124_;
  wire _auto_iopadmap_cc_313_execute_65414_125_;
  wire _auto_iopadmap_cc_313_execute_65414_126_;
  wire _auto_iopadmap_cc_313_execute_65414_127_;
  wire _auto_iopadmap_cc_313_execute_65414_128_;
  wire _auto_iopadmap_cc_313_execute_65414_129_;
  wire _auto_iopadmap_cc_313_execute_65414_130_;
  wire _auto_iopadmap_cc_313_execute_65414_131_;
  wire _auto_iopadmap_cc_313_execute_65414_132_;
  wire _auto_iopadmap_cc_313_execute_65414_133_;
  wire _auto_iopadmap_cc_313_execute_65414_134_;
  wire _auto_iopadmap_cc_313_execute_65414_135_;
  wire _auto_iopadmap_cc_313_execute_65414_136_;
  wire _auto_iopadmap_cc_313_execute_65414_137_;
  wire _auto_iopadmap_cc_313_execute_65414_138_;
  wire _auto_iopadmap_cc_313_execute_65414_139_;
  wire _auto_iopadmap_cc_313_execute_65414_140_;
  wire _auto_iopadmap_cc_313_execute_65414_141_;
  wire _auto_iopadmap_cc_313_execute_65414_142_;
  wire _auto_iopadmap_cc_313_execute_65414_143_;
  wire _auto_iopadmap_cc_313_execute_65414_144_;
  wire _auto_iopadmap_cc_313_execute_65414_145_;
  wire _auto_iopadmap_cc_313_execute_65414_146_;
  wire _auto_iopadmap_cc_313_execute_65414_147_;
  wire _auto_iopadmap_cc_313_execute_65414_148_;
  wire _auto_iopadmap_cc_313_execute_65414_149_;
  wire _auto_iopadmap_cc_313_execute_65414_150_;
  wire _auto_iopadmap_cc_313_execute_65414_151_;
  wire _auto_iopadmap_cc_313_execute_65414_152_;
  wire _auto_iopadmap_cc_313_execute_65414_153_;
  wire _auto_iopadmap_cc_313_execute_65414_154_;
  wire _auto_iopadmap_cc_313_execute_65414_155_;
  wire _auto_iopadmap_cc_313_execute_65414_156_;
  wire _auto_iopadmap_cc_313_execute_65414_157_;
  wire _auto_iopadmap_cc_313_execute_65414_158_;
  wire _auto_iopadmap_cc_313_execute_65414_159_;
  wire _auto_iopadmap_cc_313_execute_65414_160_;
  wire _auto_iopadmap_cc_313_execute_65414_161_;
  wire _auto_iopadmap_cc_313_execute_65414_162_;
  wire _auto_iopadmap_cc_313_execute_65414_163_;
  wire _auto_iopadmap_cc_313_execute_65414_164_;
  wire _auto_iopadmap_cc_313_execute_65414_165_;
  wire _auto_iopadmap_cc_313_execute_65414_166_;
  wire _auto_iopadmap_cc_313_execute_65414_167_;
  wire _auto_iopadmap_cc_313_execute_65414_168_;
  wire _auto_iopadmap_cc_313_execute_65414_169_;
  wire _auto_iopadmap_cc_313_execute_65414_170_;
  wire _auto_iopadmap_cc_313_execute_65414_171_;
  wire _auto_iopadmap_cc_313_execute_65414_172_;
  wire _auto_iopadmap_cc_313_execute_65414_173_;
  wire _auto_iopadmap_cc_313_execute_65414_174_;
  wire _auto_iopadmap_cc_313_execute_65414_175_;
  wire _auto_iopadmap_cc_313_execute_65414_176_;
  wire _auto_iopadmap_cc_313_execute_65414_177_;
  wire _auto_iopadmap_cc_313_execute_65414_178_;
  wire _auto_iopadmap_cc_313_execute_65414_179_;
  wire _auto_iopadmap_cc_313_execute_65414_180_;
  wire _auto_iopadmap_cc_313_execute_65414_181_;
  wire _auto_iopadmap_cc_313_execute_65414_182_;
  wire _auto_iopadmap_cc_313_execute_65414_183_;
  wire _auto_iopadmap_cc_313_execute_65414_184_;
  wire _auto_iopadmap_cc_313_execute_65414_185_;
  wire _auto_iopadmap_cc_313_execute_65414_186_;
  wire _auto_iopadmap_cc_313_execute_65414_187_;
  wire _auto_iopadmap_cc_313_execute_65414_188_;
  wire _auto_iopadmap_cc_313_execute_65414_189_;
  wire _auto_iopadmap_cc_313_execute_65414_190_;
  wire _auto_iopadmap_cc_313_execute_65414_191_;
  wire _auto_iopadmap_cc_313_execute_65414_192_;
  wire _auto_iopadmap_cc_313_execute_65414_193_;
  wire _auto_iopadmap_cc_313_execute_65414_194_;
  wire _auto_iopadmap_cc_313_execute_65414_195_;
  wire _auto_iopadmap_cc_313_execute_65414_196_;
  wire _auto_iopadmap_cc_313_execute_65414_197_;
  wire _auto_iopadmap_cc_313_execute_65414_198_;
  wire _auto_iopadmap_cc_313_execute_65414_199_;
  wire _auto_iopadmap_cc_313_execute_65414_200_;
  wire _auto_iopadmap_cc_313_execute_65414_201_;
  wire _auto_iopadmap_cc_313_execute_65414_202_;
  wire _auto_iopadmap_cc_313_execute_65414_203_;
  wire _auto_iopadmap_cc_313_execute_65414_204_;
  wire _auto_iopadmap_cc_313_execute_65414_205_;
  wire _auto_iopadmap_cc_313_execute_65414_206_;
  wire _auto_iopadmap_cc_313_execute_65414_207_;
  wire _auto_iopadmap_cc_313_execute_65414_208_;
  wire _auto_iopadmap_cc_313_execute_65414_209_;
  wire _auto_iopadmap_cc_313_execute_65414_210_;
  wire _auto_iopadmap_cc_313_execute_65414_211_;
  wire _auto_iopadmap_cc_313_execute_65414_212_;
  wire _auto_iopadmap_cc_313_execute_65414_213_;
  wire _auto_iopadmap_cc_313_execute_65414_214_;
  wire _auto_iopadmap_cc_313_execute_65414_215_;
  wire _auto_iopadmap_cc_313_execute_65414_216_;
  wire _auto_iopadmap_cc_313_execute_65414_217_;
  wire _auto_iopadmap_cc_313_execute_65414_218_;
  wire _auto_iopadmap_cc_313_execute_65414_219_;
  wire _auto_iopadmap_cc_313_execute_65414_220_;
  wire _auto_iopadmap_cc_313_execute_65414_221_;
  wire _auto_iopadmap_cc_313_execute_65414_222_;
  wire _auto_iopadmap_cc_313_execute_65414_223_;
  wire _auto_iopadmap_cc_313_execute_65414_224_;
  wire _auto_iopadmap_cc_313_execute_65414_225_;
  wire _auto_iopadmap_cc_313_execute_65414_226_;
  wire _auto_iopadmap_cc_313_execute_65414_227_;
  wire _auto_iopadmap_cc_313_execute_65414_228_;
  wire _auto_iopadmap_cc_313_execute_65414_229_;
  wire _auto_iopadmap_cc_313_execute_65414_230_;
  wire _auto_iopadmap_cc_313_execute_65414_231_;
  wire _auto_iopadmap_cc_313_execute_65414_232_;
  wire _auto_iopadmap_cc_313_execute_65414_233_;
  wire _auto_iopadmap_cc_313_execute_65414_234_;
  wire _auto_iopadmap_cc_313_execute_65414_235_;
  wire _auto_iopadmap_cc_313_execute_65414_236_;
  wire _auto_iopadmap_cc_313_execute_65414_237_;
  wire _auto_iopadmap_cc_313_execute_65414_238_;
  wire _auto_iopadmap_cc_313_execute_65414_239_;
  wire _auto_iopadmap_cc_313_execute_65414_240_;
  wire _auto_iopadmap_cc_313_execute_65414_241_;
  wire _auto_iopadmap_cc_313_execute_65414_36_;
  wire _auto_iopadmap_cc_313_execute_65414_37_;
  wire _auto_iopadmap_cc_313_execute_65414_38_;
  wire _auto_iopadmap_cc_313_execute_65414_39_;
  wire _auto_iopadmap_cc_313_execute_65414_40_;
  wire _auto_iopadmap_cc_313_execute_65414_41_;
  wire _auto_iopadmap_cc_313_execute_65414_42_;
  wire _auto_iopadmap_cc_313_execute_65414_43_;
  wire _auto_iopadmap_cc_313_execute_65414_44_;
  wire _auto_iopadmap_cc_313_execute_65414_45_;
  wire _auto_iopadmap_cc_313_execute_65414_46_;
  wire _auto_iopadmap_cc_313_execute_65414_47_;
  wire _auto_iopadmap_cc_313_execute_65414_48_;
  wire _auto_iopadmap_cc_313_execute_65414_49_;
  wire _auto_iopadmap_cc_313_execute_65414_50_;
  wire _auto_iopadmap_cc_313_execute_65414_51_;
  wire _auto_iopadmap_cc_313_execute_65414_52_;
  wire _auto_iopadmap_cc_313_execute_65414_53_;
  wire _auto_iopadmap_cc_313_execute_65414_54_;
  wire _auto_iopadmap_cc_313_execute_65414_55_;
  wire _auto_iopadmap_cc_313_execute_65414_56_;
  wire _auto_iopadmap_cc_313_execute_65414_57_;
  wire _auto_iopadmap_cc_313_execute_65414_58_;
  wire _auto_iopadmap_cc_313_execute_65414_59_;
  wire _auto_iopadmap_cc_313_execute_65414_60_;
  wire _auto_iopadmap_cc_313_execute_65414_61_;
  wire _auto_iopadmap_cc_313_execute_65414_62_;
  wire _auto_iopadmap_cc_313_execute_65414_63_;
  wire _auto_iopadmap_cc_313_execute_65414_64_;
  wire _auto_iopadmap_cc_313_execute_65414_65_;
  wire _auto_iopadmap_cc_313_execute_65414_66_;
  wire _auto_iopadmap_cc_313_execute_65414_67_;
  wire _auto_iopadmap_cc_313_execute_65414_68_;
  wire _auto_iopadmap_cc_313_execute_65414_69_;
  wire _auto_iopadmap_cc_313_execute_65414_70_;
  wire _auto_iopadmap_cc_313_execute_65414_71_;
  wire _auto_iopadmap_cc_313_execute_65414_72_;
  wire _auto_iopadmap_cc_313_execute_65414_73_;
  wire _auto_iopadmap_cc_313_execute_65414_74_;
  wire _auto_iopadmap_cc_313_execute_65414_75_;
  wire _auto_iopadmap_cc_313_execute_65414_76_;
  wire _auto_iopadmap_cc_313_execute_65414_77_;
  wire _auto_iopadmap_cc_313_execute_65414_78_;
  wire _auto_iopadmap_cc_313_execute_65414_79_;
  wire _auto_iopadmap_cc_313_execute_65414_80_;
  wire _auto_iopadmap_cc_313_execute_65414_81_;
  wire _auto_iopadmap_cc_313_execute_65414_82_;
  wire _auto_iopadmap_cc_313_execute_65414_83_;
  wire _auto_iopadmap_cc_313_execute_65414_84_;
  wire _auto_iopadmap_cc_313_execute_65414_85_;
  wire _auto_iopadmap_cc_313_execute_65414_86_;
  wire _auto_iopadmap_cc_313_execute_65414_87_;
  wire _auto_iopadmap_cc_313_execute_65414_88_;
  wire _auto_iopadmap_cc_313_execute_65414_89_;
  wire _auto_iopadmap_cc_313_execute_65414_90_;
  wire _auto_iopadmap_cc_313_execute_65414_91_;
  wire _auto_iopadmap_cc_313_execute_65414_92_;
  wire _auto_iopadmap_cc_313_execute_65414_93_;
  wire _auto_iopadmap_cc_313_execute_65414_94_;
  wire _auto_iopadmap_cc_313_execute_65414_95_;
  wire _auto_iopadmap_cc_313_execute_65414_96_;
  wire _auto_iopadmap_cc_313_execute_65414_97_;
  wire _auto_iopadmap_cc_313_execute_65414_98_;
  wire _auto_iopadmap_cc_313_execute_65414_99_;
  wire aNan;
  wire aNan_bF_buf0;
  wire aNan_bF_buf1;
  wire aNan_bF_buf10;
  wire aNan_bF_buf2;
  wire aNan_bF_buf3;
  wire aNan_bF_buf4;
  wire aNan_bF_buf5;
  wire aNan_bF_buf6;
  wire aNan_bF_buf7;
  wire aNan_bF_buf8;
  wire aNan_bF_buf9;
  input \a[0] ;
  input \a[100] ;
  input \a[101] ;
  input \a[102] ;
  input \a[103] ;
  input \a[104] ;
  input \a[105] ;
  input \a[106] ;
  input \a[107] ;
  input \a[108] ;
  input \a[109] ;
  input \a[10] ;
  input \a[110] ;
  input \a[111] ;
  input \a[112] ;
  input \a[113] ;
  input \a[114] ;
  input \a[115] ;
  input \a[116] ;
  input \a[117] ;
  input \a[118] ;
  input \a[119] ;
  input \a[11] ;
  input \a[120] ;
  input \a[121] ;
  input \a[122] ;
  input \a[123] ;
  input \a[124] ;
  input \a[125] ;
  input \a[126] ;
  input \a[127] ;
  input \a[12] ;
  input \a[13] ;
  input \a[14] ;
  input \a[15] ;
  input \a[16] ;
  input \a[17] ;
  input \a[18] ;
  input \a[19] ;
  input \a[1] ;
  input \a[20] ;
  input \a[21] ;
  input \a[22] ;
  input \a[23] ;
  input \a[24] ;
  input \a[25] ;
  input \a[26] ;
  input \a[27] ;
  input \a[28] ;
  input \a[29] ;
  input \a[2] ;
  input \a[30] ;
  input \a[31] ;
  input \a[32] ;
  input \a[33] ;
  input \a[34] ;
  input \a[35] ;
  input \a[36] ;
  input \a[37] ;
  input \a[38] ;
  input \a[39] ;
  input \a[3] ;
  input \a[40] ;
  input \a[41] ;
  input \a[42] ;
  input \a[43] ;
  input \a[44] ;
  input \a[45] ;
  input \a[46] ;
  input \a[47] ;
  input \a[48] ;
  input \a[49] ;
  input \a[4] ;
  input \a[50] ;
  input \a[51] ;
  input \a[52] ;
  input \a[53] ;
  input \a[54] ;
  input \a[55] ;
  input \a[56] ;
  input \a[57] ;
  input \a[58] ;
  input \a[59] ;
  input \a[5] ;
  input \a[60] ;
  input \a[61] ;
  input \a[62] ;
  input \a[63] ;
  input \a[64] ;
  input \a[65] ;
  input \a[66] ;
  input \a[67] ;
  input \a[68] ;
  input \a[69] ;
  input \a[6] ;
  input \a[70] ;
  input \a[71] ;
  input \a[72] ;
  input \a[73] ;
  input \a[74] ;
  input \a[75] ;
  input \a[76] ;
  input \a[77] ;
  input \a[78] ;
  input \a[79] ;
  input \a[7] ;
  input \a[80] ;
  input \a[81] ;
  input \a[82] ;
  input \a[83] ;
  input \a[84] ;
  input \a[85] ;
  input \a[86] ;
  input \a[87] ;
  input \a[88] ;
  input \a[89] ;
  input \a[8] ;
  input \a[90] ;
  input \a[91] ;
  input \a[92] ;
  input \a[93] ;
  input \a[94] ;
  input \a[95] ;
  input \a[96] ;
  input \a[97] ;
  input \a[98] ;
  input \a[99] ;
  input \a[9] ;
  wire a_112_bF_buf0;
  wire a_112_bF_buf1;
  wire a_112_bF_buf2;
  wire a_112_bF_buf3;
  wire a_112_bF_buf4;
  wire a_112_bF_buf5;
  wire a_112_bF_buf6;
  wire a_112_bF_buf7;
  wire a_112_bF_buf8;
  wire a_112_bF_buf9;
  input ce;
  input clk;
  wire clk_bF_buf0;
  wire clk_bF_buf1;
  wire clk_bF_buf10;
  wire clk_bF_buf100;
  wire clk_bF_buf101;
  wire clk_bF_buf102;
  wire clk_bF_buf103;
  wire clk_bF_buf104;
  wire clk_bF_buf105;
  wire clk_bF_buf106;
  wire clk_bF_buf107;
  wire clk_bF_buf108;
  wire clk_bF_buf109;
  wire clk_bF_buf11;
  wire clk_bF_buf110;
  wire clk_bF_buf111;
  wire clk_bF_buf112;
  wire clk_bF_buf113;
  wire clk_bF_buf114;
  wire clk_bF_buf115;
  wire clk_bF_buf116;
  wire clk_bF_buf117;
  wire clk_bF_buf118;
  wire clk_bF_buf119;
  wire clk_bF_buf12;
  wire clk_bF_buf120;
  wire clk_bF_buf121;
  wire clk_bF_buf13;
  wire clk_bF_buf14;
  wire clk_bF_buf15;
  wire clk_bF_buf16;
  wire clk_bF_buf17;
  wire clk_bF_buf18;
  wire clk_bF_buf19;
  wire clk_bF_buf2;
  wire clk_bF_buf20;
  wire clk_bF_buf21;
  wire clk_bF_buf22;
  wire clk_bF_buf23;
  wire clk_bF_buf24;
  wire clk_bF_buf25;
  wire clk_bF_buf26;
  wire clk_bF_buf27;
  wire clk_bF_buf28;
  wire clk_bF_buf29;
  wire clk_bF_buf3;
  wire clk_bF_buf30;
  wire clk_bF_buf31;
  wire clk_bF_buf32;
  wire clk_bF_buf33;
  wire clk_bF_buf34;
  wire clk_bF_buf35;
  wire clk_bF_buf36;
  wire clk_bF_buf37;
  wire clk_bF_buf38;
  wire clk_bF_buf39;
  wire clk_bF_buf4;
  wire clk_bF_buf40;
  wire clk_bF_buf41;
  wire clk_bF_buf42;
  wire clk_bF_buf43;
  wire clk_bF_buf44;
  wire clk_bF_buf45;
  wire clk_bF_buf46;
  wire clk_bF_buf47;
  wire clk_bF_buf48;
  wire clk_bF_buf49;
  wire clk_bF_buf5;
  wire clk_bF_buf50;
  wire clk_bF_buf51;
  wire clk_bF_buf52;
  wire clk_bF_buf53;
  wire clk_bF_buf54;
  wire clk_bF_buf55;
  wire clk_bF_buf56;
  wire clk_bF_buf57;
  wire clk_bF_buf58;
  wire clk_bF_buf59;
  wire clk_bF_buf6;
  wire clk_bF_buf60;
  wire clk_bF_buf61;
  wire clk_bF_buf62;
  wire clk_bF_buf63;
  wire clk_bF_buf64;
  wire clk_bF_buf65;
  wire clk_bF_buf66;
  wire clk_bF_buf67;
  wire clk_bF_buf68;
  wire clk_bF_buf69;
  wire clk_bF_buf7;
  wire clk_bF_buf70;
  wire clk_bF_buf71;
  wire clk_bF_buf72;
  wire clk_bF_buf73;
  wire clk_bF_buf74;
  wire clk_bF_buf75;
  wire clk_bF_buf76;
  wire clk_bF_buf77;
  wire clk_bF_buf78;
  wire clk_bF_buf79;
  wire clk_bF_buf8;
  wire clk_bF_buf80;
  wire clk_bF_buf81;
  wire clk_bF_buf82;
  wire clk_bF_buf83;
  wire clk_bF_buf84;
  wire clk_bF_buf85;
  wire clk_bF_buf86;
  wire clk_bF_buf87;
  wire clk_bF_buf88;
  wire clk_bF_buf89;
  wire clk_bF_buf9;
  wire clk_bF_buf90;
  wire clk_bF_buf91;
  wire clk_bF_buf92;
  wire clk_bF_buf93;
  wire clk_bF_buf94;
  wire clk_bF_buf95;
  wire clk_bF_buf96;
  wire clk_bF_buf97;
  wire clk_bF_buf98;
  wire clk_bF_buf99;
  wire clk_hier0_bF_buf0;
  wire clk_hier0_bF_buf1;
  wire clk_hier0_bF_buf10;
  wire clk_hier0_bF_buf2;
  wire clk_hier0_bF_buf3;
  wire clk_hier0_bF_buf4;
  wire clk_hier0_bF_buf5;
  wire clk_hier0_bF_buf6;
  wire clk_hier0_bF_buf7;
  wire clk_hier0_bF_buf8;
  wire clk_hier0_bF_buf9;
  output done;
  wire fracta1_0_;
  wire fracta1_100_;
  wire fracta1_101_;
  wire fracta1_102_;
  wire fracta1_103_;
  wire fracta1_104_;
  wire fracta1_105_;
  wire fracta1_106_;
  wire fracta1_107_;
  wire fracta1_108_;
  wire fracta1_109_;
  wire fracta1_10_;
  wire fracta1_110_;
  wire fracta1_111_;
  wire fracta1_112_;
  wire fracta1_113_;
  wire fracta1_11_;
  wire fracta1_12_;
  wire fracta1_13_;
  wire fracta1_14_;
  wire fracta1_15_;
  wire fracta1_16_;
  wire fracta1_17_;
  wire fracta1_18_;
  wire fracta1_19_;
  wire fracta1_1_;
  wire fracta1_20_;
  wire fracta1_21_;
  wire fracta1_22_;
  wire fracta1_23_;
  wire fracta1_24_;
  wire fracta1_25_;
  wire fracta1_26_;
  wire fracta1_27_;
  wire fracta1_28_;
  wire fracta1_29_;
  wire fracta1_2_;
  wire fracta1_30_;
  wire fracta1_31_;
  wire fracta1_32_;
  wire fracta1_33_;
  wire fracta1_34_;
  wire fracta1_35_;
  wire fracta1_36_;
  wire fracta1_37_;
  wire fracta1_38_;
  wire fracta1_39_;
  wire fracta1_3_;
  wire fracta1_40_;
  wire fracta1_41_;
  wire fracta1_42_;
  wire fracta1_43_;
  wire fracta1_44_;
  wire fracta1_45_;
  wire fracta1_46_;
  wire fracta1_47_;
  wire fracta1_48_;
  wire fracta1_49_;
  wire fracta1_4_;
  wire fracta1_50_;
  wire fracta1_51_;
  wire fracta1_52_;
  wire fracta1_53_;
  wire fracta1_54_;
  wire fracta1_55_;
  wire fracta1_56_;
  wire fracta1_57_;
  wire fracta1_58_;
  wire fracta1_59_;
  wire fracta1_5_;
  wire fracta1_60_;
  wire fracta1_61_;
  wire fracta1_62_;
  wire fracta1_63_;
  wire fracta1_64_;
  wire fracta1_65_;
  wire fracta1_66_;
  wire fracta1_67_;
  wire fracta1_68_;
  wire fracta1_69_;
  wire fracta1_6_;
  wire fracta1_70_;
  wire fracta1_71_;
  wire fracta1_72_;
  wire fracta1_73_;
  wire fracta1_74_;
  wire fracta1_75_;
  wire fracta1_76_;
  wire fracta1_77_;
  wire fracta1_78_;
  wire fracta1_79_;
  wire fracta1_7_;
  wire fracta1_80_;
  wire fracta1_81_;
  wire fracta1_82_;
  wire fracta1_83_;
  wire fracta1_84_;
  wire fracta1_85_;
  wire fracta1_86_;
  wire fracta1_87_;
  wire fracta1_88_;
  wire fracta1_89_;
  wire fracta1_8_;
  wire fracta1_90_;
  wire fracta1_91_;
  wire fracta1_92_;
  wire fracta1_93_;
  wire fracta1_94_;
  wire fracta1_95_;
  wire fracta1_96_;
  wire fracta1_97_;
  wire fracta1_98_;
  wire fracta1_99_;
  wire fracta1_9_;
  wire fracta_112_;
  input ld;
  output \o[0] ;
  output \o[100] ;
  output \o[101] ;
  output \o[102] ;
  output \o[103] ;
  output \o[104] ;
  output \o[105] ;
  output \o[106] ;
  output \o[107] ;
  output \o[108] ;
  output \o[109] ;
  output \o[10] ;
  output \o[110] ;
  output \o[111] ;
  output \o[112] ;
  output \o[113] ;
  output \o[114] ;
  output \o[115] ;
  output \o[116] ;
  output \o[117] ;
  output \o[118] ;
  output \o[119] ;
  output \o[11] ;
  output \o[120] ;
  output \o[121] ;
  output \o[122] ;
  output \o[123] ;
  output \o[124] ;
  output \o[125] ;
  output \o[126] ;
  output \o[127] ;
  output \o[128] ;
  output \o[129] ;
  output \o[12] ;
  output \o[130] ;
  output \o[131] ;
  output \o[132] ;
  output \o[133] ;
  output \o[134] ;
  output \o[135] ;
  output \o[136] ;
  output \o[137] ;
  output \o[138] ;
  output \o[139] ;
  output \o[13] ;
  output \o[140] ;
  output \o[141] ;
  output \o[142] ;
  output \o[143] ;
  output \o[144] ;
  output \o[145] ;
  output \o[146] ;
  output \o[147] ;
  output \o[148] ;
  output \o[149] ;
  output \o[14] ;
  output \o[150] ;
  output \o[151] ;
  output \o[152] ;
  output \o[153] ;
  output \o[154] ;
  output \o[155] ;
  output \o[156] ;
  output \o[157] ;
  output \o[158] ;
  output \o[159] ;
  output \o[15] ;
  output \o[160] ;
  output \o[161] ;
  output \o[162] ;
  output \o[163] ;
  output \o[164] ;
  output \o[165] ;
  output \o[166] ;
  output \o[167] ;
  output \o[168] ;
  output \o[169] ;
  output \o[16] ;
  output \o[170] ;
  output \o[171] ;
  output \o[172] ;
  output \o[173] ;
  output \o[174] ;
  output \o[175] ;
  output \o[176] ;
  output \o[177] ;
  output \o[178] ;
  output \o[179] ;
  output \o[17] ;
  output \o[180] ;
  output \o[181] ;
  output \o[182] ;
  output \o[183] ;
  output \o[184] ;
  output \o[185] ;
  output \o[186] ;
  output \o[187] ;
  output \o[188] ;
  output \o[189] ;
  output \o[18] ;
  output \o[190] ;
  output \o[191] ;
  output \o[192] ;
  output \o[193] ;
  output \o[194] ;
  output \o[195] ;
  output \o[196] ;
  output \o[197] ;
  output \o[198] ;
  output \o[199] ;
  output \o[19] ;
  output \o[1] ;
  output \o[200] ;
  output \o[201] ;
  output \o[202] ;
  output \o[203] ;
  output \o[204] ;
  output \o[205] ;
  output \o[206] ;
  output \o[207] ;
  output \o[208] ;
  output \o[209] ;
  output \o[20] ;
  output \o[210] ;
  output \o[211] ;
  output \o[212] ;
  output \o[213] ;
  output \o[214] ;
  output \o[215] ;
  output \o[216] ;
  output \o[217] ;
  output \o[218] ;
  output \o[219] ;
  output \o[21] ;
  output \o[220] ;
  output \o[221] ;
  output \o[222] ;
  output \o[223] ;
  output \o[224] ;
  output \o[225] ;
  output \o[226] ;
  output \o[227] ;
  output \o[228] ;
  output \o[229] ;
  output \o[22] ;
  output \o[230] ;
  output \o[231] ;
  output \o[232] ;
  output \o[233] ;
  output \o[234] ;
  output \o[235] ;
  output \o[236] ;
  output \o[237] ;
  output \o[238] ;
  output \o[239] ;
  output \o[23] ;
  output \o[240] ;
  output \o[241] ;
  output \o[24] ;
  output \o[25] ;
  output \o[26] ;
  output \o[27] ;
  output \o[28] ;
  output \o[29] ;
  output \o[2] ;
  output \o[30] ;
  output \o[31] ;
  output \o[32] ;
  output \o[33] ;
  output \o[34] ;
  output \o[35] ;
  output \o[36] ;
  output \o[37] ;
  output \o[38] ;
  output \o[39] ;
  output \o[3] ;
  output \o[40] ;
  output \o[41] ;
  output \o[42] ;
  output \o[43] ;
  output \o[44] ;
  output \o[45] ;
  output \o[46] ;
  output \o[47] ;
  output \o[48] ;
  output \o[49] ;
  output \o[4] ;
  output \o[50] ;
  output \o[51] ;
  output \o[52] ;
  output \o[53] ;
  output \o[54] ;
  output \o[55] ;
  output \o[56] ;
  output \o[57] ;
  output \o[58] ;
  output \o[59] ;
  output \o[5] ;
  output \o[60] ;
  output \o[61] ;
  output \o[62] ;
  output \o[63] ;
  output \o[64] ;
  output \o[65] ;
  output \o[66] ;
  output \o[67] ;
  output \o[68] ;
  output \o[69] ;
  output \o[6] ;
  output \o[70] ;
  output \o[71] ;
  output \o[72] ;
  output \o[73] ;
  output \o[74] ;
  output \o[75] ;
  output \o[76] ;
  output \o[77] ;
  output \o[78] ;
  output \o[79] ;
  output \o[7] ;
  output \o[80] ;
  output \o[81] ;
  output \o[82] ;
  output \o[83] ;
  output \o[84] ;
  output \o[85] ;
  output \o[86] ;
  output \o[87] ;
  output \o[88] ;
  output \o[89] ;
  output \o[8] ;
  output \o[90] ;
  output \o[91] ;
  output \o[92] ;
  output \o[93] ;
  output \o[94] ;
  output \o[95] ;
  output \o[96] ;
  output \o[97] ;
  output \o[98] ;
  output \o[99] ;
  output \o[9] ;
  input rst;
  wire sqrto_0_;
  wire sqrto_100_;
  wire sqrto_101_;
  wire sqrto_102_;
  wire sqrto_103_;
  wire sqrto_104_;
  wire sqrto_105_;
  wire sqrto_106_;
  wire sqrto_107_;
  wire sqrto_108_;
  wire sqrto_109_;
  wire sqrto_10_;
  wire sqrto_110_;
  wire sqrto_111_;
  wire sqrto_112_;
  wire sqrto_113_;
  wire sqrto_114_;
  wire sqrto_115_;
  wire sqrto_116_;
  wire sqrto_117_;
  wire sqrto_118_;
  wire sqrto_119_;
  wire sqrto_11_;
  wire sqrto_120_;
  wire sqrto_121_;
  wire sqrto_122_;
  wire sqrto_123_;
  wire sqrto_124_;
  wire sqrto_125_;
  wire sqrto_126_;
  wire sqrto_127_;
  wire sqrto_128_;
  wire sqrto_129_;
  wire sqrto_12_;
  wire sqrto_130_;
  wire sqrto_131_;
  wire sqrto_132_;
  wire sqrto_133_;
  wire sqrto_134_;
  wire sqrto_135_;
  wire sqrto_136_;
  wire sqrto_137_;
  wire sqrto_138_;
  wire sqrto_139_;
  wire sqrto_13_;
  wire sqrto_140_;
  wire sqrto_141_;
  wire sqrto_142_;
  wire sqrto_143_;
  wire sqrto_144_;
  wire sqrto_145_;
  wire sqrto_146_;
  wire sqrto_147_;
  wire sqrto_148_;
  wire sqrto_149_;
  wire sqrto_14_;
  wire sqrto_150_;
  wire sqrto_151_;
  wire sqrto_152_;
  wire sqrto_153_;
  wire sqrto_154_;
  wire sqrto_155_;
  wire sqrto_156_;
  wire sqrto_157_;
  wire sqrto_158_;
  wire sqrto_159_;
  wire sqrto_15_;
  wire sqrto_160_;
  wire sqrto_161_;
  wire sqrto_162_;
  wire sqrto_163_;
  wire sqrto_164_;
  wire sqrto_165_;
  wire sqrto_166_;
  wire sqrto_167_;
  wire sqrto_168_;
  wire sqrto_169_;
  wire sqrto_16_;
  wire sqrto_170_;
  wire sqrto_171_;
  wire sqrto_172_;
  wire sqrto_173_;
  wire sqrto_174_;
  wire sqrto_175_;
  wire sqrto_176_;
  wire sqrto_177_;
  wire sqrto_178_;
  wire sqrto_179_;
  wire sqrto_17_;
  wire sqrto_180_;
  wire sqrto_181_;
  wire sqrto_182_;
  wire sqrto_183_;
  wire sqrto_184_;
  wire sqrto_185_;
  wire sqrto_186_;
  wire sqrto_187_;
  wire sqrto_188_;
  wire sqrto_189_;
  wire sqrto_18_;
  wire sqrto_190_;
  wire sqrto_191_;
  wire sqrto_192_;
  wire sqrto_193_;
  wire sqrto_194_;
  wire sqrto_195_;
  wire sqrto_196_;
  wire sqrto_197_;
  wire sqrto_198_;
  wire sqrto_199_;
  wire sqrto_19_;
  wire sqrto_1_;
  wire sqrto_200_;
  wire sqrto_201_;
  wire sqrto_202_;
  wire sqrto_203_;
  wire sqrto_204_;
  wire sqrto_205_;
  wire sqrto_206_;
  wire sqrto_207_;
  wire sqrto_208_;
  wire sqrto_209_;
  wire sqrto_20_;
  wire sqrto_210_;
  wire sqrto_211_;
  wire sqrto_212_;
  wire sqrto_213_;
  wire sqrto_214_;
  wire sqrto_215_;
  wire sqrto_216_;
  wire sqrto_217_;
  wire sqrto_218_;
  wire sqrto_219_;
  wire sqrto_21_;
  wire sqrto_220_;
  wire sqrto_221_;
  wire sqrto_222_;
  wire sqrto_223_;
  wire sqrto_224_;
  wire sqrto_225_;
  wire sqrto_22_;
  wire sqrto_23_;
  wire sqrto_24_;
  wire sqrto_25_;
  wire sqrto_26_;
  wire sqrto_27_;
  wire sqrto_28_;
  wire sqrto_29_;
  wire sqrto_2_;
  wire sqrto_30_;
  wire sqrto_31_;
  wire sqrto_32_;
  wire sqrto_33_;
  wire sqrto_34_;
  wire sqrto_35_;
  wire sqrto_36_;
  wire sqrto_37_;
  wire sqrto_38_;
  wire sqrto_39_;
  wire sqrto_3_;
  wire sqrto_40_;
  wire sqrto_41_;
  wire sqrto_42_;
  wire sqrto_43_;
  wire sqrto_44_;
  wire sqrto_45_;
  wire sqrto_46_;
  wire sqrto_47_;
  wire sqrto_48_;
  wire sqrto_49_;
  wire sqrto_4_;
  wire sqrto_50_;
  wire sqrto_51_;
  wire sqrto_52_;
  wire sqrto_53_;
  wire sqrto_54_;
  wire sqrto_55_;
  wire sqrto_56_;
  wire sqrto_57_;
  wire sqrto_58_;
  wire sqrto_59_;
  wire sqrto_5_;
  wire sqrto_60_;
  wire sqrto_61_;
  wire sqrto_62_;
  wire sqrto_63_;
  wire sqrto_64_;
  wire sqrto_65_;
  wire sqrto_66_;
  wire sqrto_67_;
  wire sqrto_68_;
  wire sqrto_69_;
  wire sqrto_6_;
  wire sqrto_70_;
  wire sqrto_71_;
  wire sqrto_72_;
  wire sqrto_73_;
  wire sqrto_74_;
  wire sqrto_75_;
  wire sqrto_76_;
  wire sqrto_77_;
  wire sqrto_78_;
  wire sqrto_79_;
  wire sqrto_7_;
  wire sqrto_80_;
  wire sqrto_81_;
  wire sqrto_82_;
  wire sqrto_83_;
  wire sqrto_84_;
  wire sqrto_85_;
  wire sqrto_86_;
  wire sqrto_87_;
  wire sqrto_88_;
  wire sqrto_89_;
  wire sqrto_8_;
  wire sqrto_90_;
  wire sqrto_91_;
  wire sqrto_92_;
  wire sqrto_93_;
  wire sqrto_94_;
  wire sqrto_95_;
  wire sqrto_96_;
  wire sqrto_97_;
  wire sqrto_98_;
  wire sqrto_99_;
  wire sqrto_9_;
  wire u1__abc_43968_n137;
  wire u1__abc_43968_n138;
  wire u1__abc_43968_n139_1;
  wire u1__abc_43968_n140_1;
  wire u1__abc_43968_n141;
  wire u1__abc_43968_n142_1;
  wire u1__abc_43968_n143_1;
  wire u1__abc_43968_n144;
  wire u1__abc_43968_n145;
  wire u1__abc_43968_n146_1;
  wire u1__abc_43968_n147_1;
  wire u1__abc_43968_n148;
  wire u1__abc_43968_n149_1;
  wire u1__abc_43968_n152;
  wire u1__abc_43968_n153;
  wire u1__abc_43968_n154_1;
  wire u1__abc_43968_n155_1;
  wire u1__abc_43968_n156;
  wire u1__abc_43968_n157_1;
  wire u1__abc_43968_n158_1;
  wire u1__abc_43968_n159;
  wire u1__abc_43968_n160;
  wire u1__abc_43968_n161_1;
  wire u1__abc_43968_n162_1;
  wire u1__abc_43968_n163;
  wire u1__abc_43968_n164_1;
  wire u1__abc_43968_n166;
  wire u1__abc_43968_n167;
  wire u1__abc_43968_n168;
  wire u1__abc_43968_n169;
  wire u1__abc_43968_n170_1;
  wire u1__abc_43968_n171_1;
  wire u1__abc_43968_n172;
  wire u1__abc_43968_n173_1;
  wire u1__abc_43968_n174_1;
  wire u1__abc_43968_n175;
  wire u1__abc_43968_n176;
  wire u1__abc_43968_n177_1;
  wire u1__abc_43968_n178_1;
  wire u1__abc_43968_n179;
  wire u1__abc_43968_n180_1;
  wire u1__abc_43968_n181_1;
  wire u1__abc_43968_n182;
  wire u1__abc_43968_n183;
  wire u1__abc_43968_n184;
  wire u1__abc_43968_n185_1;
  wire u1__abc_43968_n186_1;
  wire u1__abc_43968_n187;
  wire u1__abc_43968_n188_1;
  wire u1__abc_43968_n189_1;
  wire u1__abc_43968_n190;
  wire u1__abc_43968_n191;
  wire u1__abc_43968_n192_1;
  wire u1__abc_43968_n193_1;
  wire u1__abc_43968_n194;
  wire u1__abc_43968_n195_1;
  wire u1__abc_43968_n196_1;
  wire u1__abc_43968_n197;
  wire u1__abc_43968_n198;
  wire u1__abc_43968_n199;
  wire u1__abc_43968_n200;
  wire u1__abc_43968_n201;
  wire u1__abc_43968_n202_1;
  wire u1__abc_43968_n203_1;
  wire u1__abc_43968_n204;
  wire u1__abc_43968_n205_1;
  wire u1__abc_43968_n206_1;
  wire u1__abc_43968_n207;
  wire u1__abc_43968_n208;
  wire u1__abc_43968_n209_1;
  wire u1__abc_43968_n210_1;
  wire u1__abc_43968_n211;
  wire u1__abc_43968_n212_1;
  wire u1__abc_43968_n213_1;
  wire u1__abc_43968_n214;
  wire u1__abc_43968_n215;
  wire u1__abc_43968_n216;
  wire u1__abc_43968_n217_1;
  wire u1__abc_43968_n218_1;
  wire u1__abc_43968_n219;
  wire u1__abc_43968_n220_1;
  wire u1__abc_43968_n221_1;
  wire u1__abc_43968_n222;
  wire u1__abc_43968_n223;
  wire u1__abc_43968_n224_1;
  wire u1__abc_43968_n225_1;
  wire u1__abc_43968_n226;
  wire u1__abc_43968_n227_1;
  wire u1__abc_43968_n228_1;
  wire u1__abc_43968_n229;
  wire u1__abc_43968_n230;
  wire u1__abc_43968_n231;
  wire u1__abc_43968_n232;
  wire u1__abc_43968_n233_1;
  wire u1__abc_43968_n234_1;
  wire u1__abc_43968_n235;
  wire u1__abc_43968_n236_1;
  wire u1__abc_43968_n237_1;
  wire u1__abc_43968_n238;
  wire u1__abc_43968_n239;
  wire u1__abc_43968_n240_1;
  wire u1__abc_43968_n241_1;
  wire u1__abc_43968_n242;
  wire u1__abc_43968_n243_1;
  wire u1__abc_43968_n244_1;
  wire u1__abc_43968_n245;
  wire u1__abc_43968_n246;
  wire u1__abc_43968_n247;
  wire u1__abc_43968_n248_1;
  wire u1__abc_43968_n249_1;
  wire u1__abc_43968_n250;
  wire u1__abc_43968_n251_1;
  wire u1__abc_43968_n252_1;
  wire u1__abc_43968_n253;
  wire u1__abc_43968_n254;
  wire u1__abc_43968_n255_1;
  wire u1__abc_43968_n256_1;
  wire u1__abc_43968_n257;
  wire u1__abc_43968_n258_1;
  wire u1__abc_43968_n259_1;
  wire u1__abc_43968_n260;
  wire u1__abc_43968_n261;
  wire u1__abc_43968_n262;
  wire u1__abc_43968_n263;
  wire u1__abc_43968_n264;
  wire u1__abc_43968_n265;
  wire u1__abc_43968_n266_1;
  wire u1__abc_43968_n267_1;
  wire u1__abc_43968_n268_1;
  wire u1__abc_43968_n269_1;
  wire u1__abc_43968_n270;
  wire u1__abc_43968_n271;
  wire u1__abc_43968_n272_1;
  wire u1__abc_43968_n273_1;
  wire u1__abc_43968_n274;
  wire u1__abc_43968_n275;
  wire u1__abc_43968_n276;
  wire u1__abc_43968_n277;
  wire u1__abc_43968_n278;
  wire u1__abc_43968_n279;
  wire u1__abc_43968_n280;
  wire u1__abc_43968_n281;
  wire u1__abc_43968_n282;
  wire u1__abc_43968_n283;
  wire u1__abc_43968_n284;
  wire u1__abc_43968_n285;
  wire u1__abc_43968_n286;
  wire u1__abc_43968_n287;
  wire u1__abc_43968_n288;
  wire u1__abc_43968_n289;
  wire u1__abc_43968_n290;
  wire u1__abc_43968_n291;
  wire u1__abc_43968_n292;
  wire u1__abc_43968_n293;
  wire u1__abc_43968_n294;
  wire u1__abc_43968_n295;
  wire u1__abc_43968_n296;
  wire u1__abc_43968_n297;
  wire u1__abc_43968_n298;
  wire u1__abc_43968_n299;
  wire u1__abc_43968_n300;
  wire u1__abc_43968_n301;
  wire u1__abc_43968_n302;
  wire u1__abc_43968_n303;
  wire u1__abc_43968_n304;
  wire u1__abc_43968_n305;
  wire u1__abc_43968_n306;
  wire u1__abc_43968_n307;
  wire u1__abc_43968_n308;
  wire u1__abc_43968_n309;
  wire u1__abc_43968_n310;
  wire u1__abc_43968_n311;
  wire u1__abc_43968_n312;
  wire u1__abc_43968_n313;
  wire u1__abc_43968_n314;
  wire u1__abc_43968_n315;
  wire u1__abc_43968_n316;
  wire u1__abc_43968_n317;
  wire u1__abc_43968_n318;
  wire u1__abc_43968_n319;
  wire u1__abc_43968_n320;
  wire u1__abc_43968_n321;
  wire u1__abc_43968_n322;
  wire u1__abc_43968_n323;
  wire u1__abc_43968_n324;
  wire u1__abc_43968_n325;
  wire u1__abc_43968_n326;
  wire u1__abc_43968_n327;
  wire u1__abc_43968_n328;
  wire u1__abc_43968_n329;
  wire u1__abc_43968_n330;
  wire u1__abc_43968_n331;
  wire u1__abc_43968_n332;
  wire u1__abc_43968_n333;
  wire u1__abc_43968_n334;
  wire u1__abc_43968_n335;
  wire u1__abc_43968_n336;
  wire u1__abc_43968_n337;
  wire u1__abc_43968_n338;
  wire u1__abc_43968_n339;
  wire u1__abc_43968_n340;
  wire u1__abc_43968_n341;
  wire u1__abc_43968_n342;
  wire u1__abc_43968_n343;
  wire u1__abc_43968_n344;
  wire u1__abc_43968_n345;
  wire u1__abc_43968_n346;
  wire u1__abc_43968_n347;
  wire u1__abc_43968_n348;
  wire u1__abc_43968_n349;
  wire u1__abc_43968_n350;
  wire u1__abc_43968_n351;
  wire u1__abc_43968_n352;
  wire u1__abc_43968_n353;
  wire u1__abc_43968_n354;
  wire u1__abc_43968_n355;
  wire u1__abc_43968_n356;
  wire u1__abc_43968_n357;
  wire u1__abc_43968_n358;
  wire u1__abc_43968_n359;
  wire u1__abc_43968_n360;
  wire u1__abc_43968_n361;
  wire u1__abc_43968_n362;
  wire u1__abc_43968_n363;
  wire u1__abc_43968_n364;
  wire u1__abc_43968_n365;
  wire u1__abc_43968_n366;
  wire u1__abc_43968_n367;
  wire u1__abc_43968_n368;
  wire u1__abc_43968_n369;
  wire u1__abc_43968_n370;
  wire u1__abc_43968_n371;
  wire u1__abc_43968_n372;
  wire u1__abc_43968_n373;
  wire u1__abc_43968_n374;
  wire u1__abc_43968_n375;
  wire u1__abc_43968_n376;
  wire u1__abc_43968_n377;
  wire u1__abc_43968_n378;
  wire u1__abc_43968_n379;
  wire u1__abc_43968_n380;
  wire u1__abc_43968_n381;
  wire u1__abc_43968_n382;
  wire u1__abc_43968_n383;
  wire u1__abc_43968_n384;
  wire u1__abc_43968_n385;
  wire u1__abc_43968_n386;
  wire u1__abc_43968_n387;
  wire u1__abc_43968_n392;
  wire u1_mz;
  wire u1_xinf;
  wire u2__abc_29664_n1191;
  wire u2__abc_29664_n3922;
  wire u2__abc_29664_n3927;
  wire u2__abc_44228_n10000;
  wire u2__abc_44228_n10001_1;
  wire u2__abc_44228_n10002;
  wire u2__abc_44228_n10003;
  wire u2__abc_44228_n10004;
  wire u2__abc_44228_n10005;
  wire u2__abc_44228_n10006_1;
  wire u2__abc_44228_n10007_1;
  wire u2__abc_44228_n10008;
  wire u2__abc_44228_n10009;
  wire u2__abc_44228_n10010;
  wire u2__abc_44228_n10011;
  wire u2__abc_44228_n10012_1;
  wire u2__abc_44228_n10013;
  wire u2__abc_44228_n10014;
  wire u2__abc_44228_n10015;
  wire u2__abc_44228_n10017_1;
  wire u2__abc_44228_n10018_1;
  wire u2__abc_44228_n10019;
  wire u2__abc_44228_n10020;
  wire u2__abc_44228_n10021;
  wire u2__abc_44228_n10022;
  wire u2__abc_44228_n10023_1;
  wire u2__abc_44228_n10024;
  wire u2__abc_44228_n10025;
  wire u2__abc_44228_n10026;
  wire u2__abc_44228_n10027;
  wire u2__abc_44228_n10028_1;
  wire u2__abc_44228_n10029_1;
  wire u2__abc_44228_n10030;
  wire u2__abc_44228_n10031;
  wire u2__abc_44228_n10032;
  wire u2__abc_44228_n10034_1;
  wire u2__abc_44228_n10035;
  wire u2__abc_44228_n10036;
  wire u2__abc_44228_n10037;
  wire u2__abc_44228_n10038;
  wire u2__abc_44228_n10039_1;
  wire u2__abc_44228_n10040_1;
  wire u2__abc_44228_n10041;
  wire u2__abc_44228_n10042;
  wire u2__abc_44228_n10043;
  wire u2__abc_44228_n10044;
  wire u2__abc_44228_n10045_1;
  wire u2__abc_44228_n10046;
  wire u2__abc_44228_n10047;
  wire u2__abc_44228_n10048;
  wire u2__abc_44228_n10049;
  wire u2__abc_44228_n10051_1;
  wire u2__abc_44228_n10052;
  wire u2__abc_44228_n10053;
  wire u2__abc_44228_n10054;
  wire u2__abc_44228_n10055;
  wire u2__abc_44228_n10056_1;
  wire u2__abc_44228_n10057;
  wire u2__abc_44228_n10058;
  wire u2__abc_44228_n10059;
  wire u2__abc_44228_n10060;
  wire u2__abc_44228_n10061_1;
  wire u2__abc_44228_n10062_1;
  wire u2__abc_44228_n10063;
  wire u2__abc_44228_n10064;
  wire u2__abc_44228_n10065;
  wire u2__abc_44228_n10066;
  wire u2__abc_44228_n10068;
  wire u2__abc_44228_n10069;
  wire u2__abc_44228_n10070;
  wire u2__abc_44228_n10071;
  wire u2__abc_44228_n10072_1;
  wire u2__abc_44228_n10073_1;
  wire u2__abc_44228_n10074;
  wire u2__abc_44228_n10075;
  wire u2__abc_44228_n10076;
  wire u2__abc_44228_n10077;
  wire u2__abc_44228_n10078_1;
  wire u2__abc_44228_n10079;
  wire u2__abc_44228_n10080;
  wire u2__abc_44228_n10081;
  wire u2__abc_44228_n10082;
  wire u2__abc_44228_n10083_1;
  wire u2__abc_44228_n10084_1;
  wire u2__abc_44228_n10086;
  wire u2__abc_44228_n10087;
  wire u2__abc_44228_n10088;
  wire u2__abc_44228_n10089_1;
  wire u2__abc_44228_n10090;
  wire u2__abc_44228_n10091;
  wire u2__abc_44228_n10092;
  wire u2__abc_44228_n10093;
  wire u2__abc_44228_n10094_1;
  wire u2__abc_44228_n10095_1;
  wire u2__abc_44228_n10096;
  wire u2__abc_44228_n10097;
  wire u2__abc_44228_n10098;
  wire u2__abc_44228_n10099;
  wire u2__abc_44228_n10100_1;
  wire u2__abc_44228_n10101;
  wire u2__abc_44228_n10103;
  wire u2__abc_44228_n10104;
  wire u2__abc_44228_n10105_1;
  wire u2__abc_44228_n10106_1;
  wire u2__abc_44228_n10107;
  wire u2__abc_44228_n10108;
  wire u2__abc_44228_n10109;
  wire u2__abc_44228_n10110;
  wire u2__abc_44228_n10111_1;
  wire u2__abc_44228_n10112;
  wire u2__abc_44228_n10113;
  wire u2__abc_44228_n10114;
  wire u2__abc_44228_n10115;
  wire u2__abc_44228_n10116_1;
  wire u2__abc_44228_n10117_1;
  wire u2__abc_44228_n10118;
  wire u2__abc_44228_n10119;
  wire u2__abc_44228_n10121;
  wire u2__abc_44228_n10122_1;
  wire u2__abc_44228_n10123;
  wire u2__abc_44228_n10124;
  wire u2__abc_44228_n10125;
  wire u2__abc_44228_n10126;
  wire u2__abc_44228_n10127_1;
  wire u2__abc_44228_n10128_1;
  wire u2__abc_44228_n10129;
  wire u2__abc_44228_n10130;
  wire u2__abc_44228_n10131;
  wire u2__abc_44228_n10132;
  wire u2__abc_44228_n10133_1;
  wire u2__abc_44228_n10134;
  wire u2__abc_44228_n10135;
  wire u2__abc_44228_n10136;
  wire u2__abc_44228_n10138_1;
  wire u2__abc_44228_n10139_1;
  wire u2__abc_44228_n10140;
  wire u2__abc_44228_n10141;
  wire u2__abc_44228_n10142;
  wire u2__abc_44228_n10143;
  wire u2__abc_44228_n10144_1;
  wire u2__abc_44228_n10145;
  wire u2__abc_44228_n10146;
  wire u2__abc_44228_n10147;
  wire u2__abc_44228_n10148;
  wire u2__abc_44228_n10149_1;
  wire u2__abc_44228_n10150_1;
  wire u2__abc_44228_n10151;
  wire u2__abc_44228_n10152;
  wire u2__abc_44228_n10153;
  wire u2__abc_44228_n10155_1;
  wire u2__abc_44228_n10156;
  wire u2__abc_44228_n10157;
  wire u2__abc_44228_n10158;
  wire u2__abc_44228_n10159;
  wire u2__abc_44228_n10160_1;
  wire u2__abc_44228_n10161_1;
  wire u2__abc_44228_n10162;
  wire u2__abc_44228_n10163;
  wire u2__abc_44228_n10164;
  wire u2__abc_44228_n10165;
  wire u2__abc_44228_n10166_1;
  wire u2__abc_44228_n10167;
  wire u2__abc_44228_n10168;
  wire u2__abc_44228_n10169;
  wire u2__abc_44228_n10170;
  wire u2__abc_44228_n10172_1;
  wire u2__abc_44228_n10173;
  wire u2__abc_44228_n10174;
  wire u2__abc_44228_n10175;
  wire u2__abc_44228_n10176;
  wire u2__abc_44228_n10177_1;
  wire u2__abc_44228_n10178;
  wire u2__abc_44228_n10179;
  wire u2__abc_44228_n10180;
  wire u2__abc_44228_n10181;
  wire u2__abc_44228_n10182_1;
  wire u2__abc_44228_n10183_1;
  wire u2__abc_44228_n10184;
  wire u2__abc_44228_n10185;
  wire u2__abc_44228_n10186;
  wire u2__abc_44228_n10187;
  wire u2__abc_44228_n10188_1;
  wire u2__abc_44228_n10190;
  wire u2__abc_44228_n10191;
  wire u2__abc_44228_n10192;
  wire u2__abc_44228_n10193_1;
  wire u2__abc_44228_n10194_1;
  wire u2__abc_44228_n10195;
  wire u2__abc_44228_n10196;
  wire u2__abc_44228_n10197;
  wire u2__abc_44228_n10198;
  wire u2__abc_44228_n10199_1;
  wire u2__abc_44228_n10200;
  wire u2__abc_44228_n10201;
  wire u2__abc_44228_n10202;
  wire u2__abc_44228_n10203;
  wire u2__abc_44228_n10204_1;
  wire u2__abc_44228_n10205_1;
  wire u2__abc_44228_n10207;
  wire u2__abc_44228_n10208;
  wire u2__abc_44228_n10209;
  wire u2__abc_44228_n10210_1;
  wire u2__abc_44228_n10211;
  wire u2__abc_44228_n10212;
  wire u2__abc_44228_n10213;
  wire u2__abc_44228_n10214;
  wire u2__abc_44228_n10215_1;
  wire u2__abc_44228_n10216_1;
  wire u2__abc_44228_n10217;
  wire u2__abc_44228_n10218;
  wire u2__abc_44228_n10219;
  wire u2__abc_44228_n10220;
  wire u2__abc_44228_n10221_1;
  wire u2__abc_44228_n10222;
  wire u2__abc_44228_n10224;
  wire u2__abc_44228_n10225;
  wire u2__abc_44228_n10226_1;
  wire u2__abc_44228_n10227_1;
  wire u2__abc_44228_n10228;
  wire u2__abc_44228_n10229;
  wire u2__abc_44228_n10230;
  wire u2__abc_44228_n10231;
  wire u2__abc_44228_n10232_1;
  wire u2__abc_44228_n10233;
  wire u2__abc_44228_n10234;
  wire u2__abc_44228_n10235;
  wire u2__abc_44228_n10236;
  wire u2__abc_44228_n10237_1;
  wire u2__abc_44228_n10238_1;
  wire u2__abc_44228_n10239;
  wire u2__abc_44228_n10241;
  wire u2__abc_44228_n10242;
  wire u2__abc_44228_n10243_1;
  wire u2__abc_44228_n10244;
  wire u2__abc_44228_n10245;
  wire u2__abc_44228_n10246;
  wire u2__abc_44228_n10247;
  wire u2__abc_44228_n10248_1;
  wire u2__abc_44228_n10249_1;
  wire u2__abc_44228_n10250;
  wire u2__abc_44228_n10251;
  wire u2__abc_44228_n10252;
  wire u2__abc_44228_n10253;
  wire u2__abc_44228_n10254_1;
  wire u2__abc_44228_n10255;
  wire u2__abc_44228_n10256;
  wire u2__abc_44228_n10258;
  wire u2__abc_44228_n10259_1;
  wire u2__abc_44228_n10260_1;
  wire u2__abc_44228_n10261;
  wire u2__abc_44228_n10262;
  wire u2__abc_44228_n10263;
  wire u2__abc_44228_n10264;
  wire u2__abc_44228_n10265_1;
  wire u2__abc_44228_n10266;
  wire u2__abc_44228_n10267;
  wire u2__abc_44228_n10268;
  wire u2__abc_44228_n10269;
  wire u2__abc_44228_n10270_1;
  wire u2__abc_44228_n10271_1;
  wire u2__abc_44228_n10272;
  wire u2__abc_44228_n10273;
  wire u2__abc_44228_n10275;
  wire u2__abc_44228_n10276_1;
  wire u2__abc_44228_n10277;
  wire u2__abc_44228_n10278;
  wire u2__abc_44228_n10279;
  wire u2__abc_44228_n10280;
  wire u2__abc_44228_n10281_1;
  wire u2__abc_44228_n10282_1;
  wire u2__abc_44228_n10283;
  wire u2__abc_44228_n10284;
  wire u2__abc_44228_n10285;
  wire u2__abc_44228_n10286;
  wire u2__abc_44228_n10287_1;
  wire u2__abc_44228_n10288;
  wire u2__abc_44228_n10289;
  wire u2__abc_44228_n10290;
  wire u2__abc_44228_n10292_1;
  wire u2__abc_44228_n10293_1;
  wire u2__abc_44228_n10294;
  wire u2__abc_44228_n10295;
  wire u2__abc_44228_n10296;
  wire u2__abc_44228_n10297;
  wire u2__abc_44228_n10298_1;
  wire u2__abc_44228_n10299;
  wire u2__abc_44228_n10300;
  wire u2__abc_44228_n10301;
  wire u2__abc_44228_n10302;
  wire u2__abc_44228_n10303_1;
  wire u2__abc_44228_n10304_1;
  wire u2__abc_44228_n10305;
  wire u2__abc_44228_n10306;
  wire u2__abc_44228_n10307;
  wire u2__abc_44228_n10309_1;
  wire u2__abc_44228_n10310;
  wire u2__abc_44228_n10311;
  wire u2__abc_44228_n10312;
  wire u2__abc_44228_n10313;
  wire u2__abc_44228_n10314_1;
  wire u2__abc_44228_n10315_1;
  wire u2__abc_44228_n10316;
  wire u2__abc_44228_n10317;
  wire u2__abc_44228_n10318;
  wire u2__abc_44228_n10319;
  wire u2__abc_44228_n10320_1;
  wire u2__abc_44228_n10321;
  wire u2__abc_44228_n10322;
  wire u2__abc_44228_n10323;
  wire u2__abc_44228_n10324;
  wire u2__abc_44228_n10326_1;
  wire u2__abc_44228_n10327;
  wire u2__abc_44228_n10328;
  wire u2__abc_44228_n10329;
  wire u2__abc_44228_n10330;
  wire u2__abc_44228_n10331;
  wire u2__abc_44228_n10332_1;
  wire u2__abc_44228_n10333_1;
  wire u2__abc_44228_n10334;
  wire u2__abc_44228_n10335;
  wire u2__abc_44228_n10336;
  wire u2__abc_44228_n10337;
  wire u2__abc_44228_n10338;
  wire u2__abc_44228_n10339_1;
  wire u2__abc_44228_n10340_1;
  wire u2__abc_44228_n10341;
  wire u2__abc_44228_n10343;
  wire u2__abc_44228_n10344;
  wire u2__abc_44228_n10345;
  wire u2__abc_44228_n10346_1;
  wire u2__abc_44228_n10347_1;
  wire u2__abc_44228_n10348;
  wire u2__abc_44228_n10349;
  wire u2__abc_44228_n10350;
  wire u2__abc_44228_n10351;
  wire u2__abc_44228_n10352;
  wire u2__abc_44228_n10353_1;
  wire u2__abc_44228_n10354_1;
  wire u2__abc_44228_n10355;
  wire u2__abc_44228_n10356;
  wire u2__abc_44228_n10357;
  wire u2__abc_44228_n10358;
  wire u2__abc_44228_n10360_1;
  wire u2__abc_44228_n10361_1;
  wire u2__abc_44228_n10362;
  wire u2__abc_44228_n10363;
  wire u2__abc_44228_n10364;
  wire u2__abc_44228_n10365;
  wire u2__abc_44228_n10366;
  wire u2__abc_44228_n10367_1;
  wire u2__abc_44228_n10368_1;
  wire u2__abc_44228_n10369;
  wire u2__abc_44228_n10370;
  wire u2__abc_44228_n10371;
  wire u2__abc_44228_n10372;
  wire u2__abc_44228_n10373;
  wire u2__abc_44228_n10374_1;
  wire u2__abc_44228_n10375_1;
  wire u2__abc_44228_n10377;
  wire u2__abc_44228_n10378;
  wire u2__abc_44228_n10379;
  wire u2__abc_44228_n10380;
  wire u2__abc_44228_n10381_1;
  wire u2__abc_44228_n10382_1;
  wire u2__abc_44228_n10383;
  wire u2__abc_44228_n10384;
  wire u2__abc_44228_n10385;
  wire u2__abc_44228_n10386;
  wire u2__abc_44228_n10387;
  wire u2__abc_44228_n10388_1;
  wire u2__abc_44228_n10389_1;
  wire u2__abc_44228_n10390;
  wire u2__abc_44228_n10391;
  wire u2__abc_44228_n10392;
  wire u2__abc_44228_n10393;
  wire u2__abc_44228_n10395_1;
  wire u2__abc_44228_n10396_1;
  wire u2__abc_44228_n10397;
  wire u2__abc_44228_n10398;
  wire u2__abc_44228_n10399;
  wire u2__abc_44228_n10400;
  wire u2__abc_44228_n10401;
  wire u2__abc_44228_n10402_1;
  wire u2__abc_44228_n10403_1;
  wire u2__abc_44228_n10404;
  wire u2__abc_44228_n10405;
  wire u2__abc_44228_n10406;
  wire u2__abc_44228_n10407;
  wire u2__abc_44228_n10408;
  wire u2__abc_44228_n10409_1;
  wire u2__abc_44228_n10410_1;
  wire u2__abc_44228_n10412;
  wire u2__abc_44228_n10413;
  wire u2__abc_44228_n10414;
  wire u2__abc_44228_n10415;
  wire u2__abc_44228_n10416_1;
  wire u2__abc_44228_n10417_1;
  wire u2__abc_44228_n10418;
  wire u2__abc_44228_n10419;
  wire u2__abc_44228_n10420;
  wire u2__abc_44228_n10421;
  wire u2__abc_44228_n10422;
  wire u2__abc_44228_n10423_1;
  wire u2__abc_44228_n10424_1;
  wire u2__abc_44228_n10425;
  wire u2__abc_44228_n10426;
  wire u2__abc_44228_n10427;
  wire u2__abc_44228_n10429;
  wire u2__abc_44228_n10430_1;
  wire u2__abc_44228_n10431_1;
  wire u2__abc_44228_n10432;
  wire u2__abc_44228_n10433;
  wire u2__abc_44228_n10434;
  wire u2__abc_44228_n10435;
  wire u2__abc_44228_n10436;
  wire u2__abc_44228_n10437_1;
  wire u2__abc_44228_n10438_1;
  wire u2__abc_44228_n10439;
  wire u2__abc_44228_n10440;
  wire u2__abc_44228_n10441;
  wire u2__abc_44228_n10442;
  wire u2__abc_44228_n10443;
  wire u2__abc_44228_n10444_1;
  wire u2__abc_44228_n10446;
  wire u2__abc_44228_n10447;
  wire u2__abc_44228_n10448;
  wire u2__abc_44228_n10449;
  wire u2__abc_44228_n10450;
  wire u2__abc_44228_n10451_1;
  wire u2__abc_44228_n10452_1;
  wire u2__abc_44228_n10453;
  wire u2__abc_44228_n10454;
  wire u2__abc_44228_n10455;
  wire u2__abc_44228_n10456;
  wire u2__abc_44228_n10457;
  wire u2__abc_44228_n10458_1;
  wire u2__abc_44228_n10459_1;
  wire u2__abc_44228_n10460;
  wire u2__abc_44228_n10461;
  wire u2__abc_44228_n10462;
  wire u2__abc_44228_n10464;
  wire u2__abc_44228_n10465_1;
  wire u2__abc_44228_n10466_1;
  wire u2__abc_44228_n10467;
  wire u2__abc_44228_n10468;
  wire u2__abc_44228_n10469;
  wire u2__abc_44228_n10470;
  wire u2__abc_44228_n10471;
  wire u2__abc_44228_n10472_1;
  wire u2__abc_44228_n10473_1;
  wire u2__abc_44228_n10474;
  wire u2__abc_44228_n10475;
  wire u2__abc_44228_n10476;
  wire u2__abc_44228_n10477;
  wire u2__abc_44228_n10478;
  wire u2__abc_44228_n10479_1;
  wire u2__abc_44228_n10481;
  wire u2__abc_44228_n10482;
  wire u2__abc_44228_n10483;
  wire u2__abc_44228_n10484;
  wire u2__abc_44228_n10485;
  wire u2__abc_44228_n10486_1;
  wire u2__abc_44228_n10487_1;
  wire u2__abc_44228_n10488;
  wire u2__abc_44228_n10489;
  wire u2__abc_44228_n10490;
  wire u2__abc_44228_n10491;
  wire u2__abc_44228_n10492;
  wire u2__abc_44228_n10493_1;
  wire u2__abc_44228_n10494_1;
  wire u2__abc_44228_n10495;
  wire u2__abc_44228_n10496;
  wire u2__abc_44228_n10498;
  wire u2__abc_44228_n10499;
  wire u2__abc_44228_n10500_1;
  wire u2__abc_44228_n10501_1;
  wire u2__abc_44228_n10502;
  wire u2__abc_44228_n10503;
  wire u2__abc_44228_n10504;
  wire u2__abc_44228_n10505;
  wire u2__abc_44228_n10506;
  wire u2__abc_44228_n10507_1;
  wire u2__abc_44228_n10508_1;
  wire u2__abc_44228_n10509;
  wire u2__abc_44228_n10510;
  wire u2__abc_44228_n10511;
  wire u2__abc_44228_n10512;
  wire u2__abc_44228_n10513;
  wire u2__abc_44228_n10515_1;
  wire u2__abc_44228_n10516;
  wire u2__abc_44228_n10517;
  wire u2__abc_44228_n10518;
  wire u2__abc_44228_n10519;
  wire u2__abc_44228_n10520;
  wire u2__abc_44228_n10521_1;
  wire u2__abc_44228_n10522_1;
  wire u2__abc_44228_n10523;
  wire u2__abc_44228_n10524;
  wire u2__abc_44228_n10525;
  wire u2__abc_44228_n10526;
  wire u2__abc_44228_n10527;
  wire u2__abc_44228_n10528_1;
  wire u2__abc_44228_n10529_1;
  wire u2__abc_44228_n10530;
  wire u2__abc_44228_n10531;
  wire u2__abc_44228_n10533;
  wire u2__abc_44228_n10534;
  wire u2__abc_44228_n10535_1;
  wire u2__abc_44228_n10536_1;
  wire u2__abc_44228_n10537;
  wire u2__abc_44228_n10538;
  wire u2__abc_44228_n10539;
  wire u2__abc_44228_n10540;
  wire u2__abc_44228_n10541;
  wire u2__abc_44228_n10542_1;
  wire u2__abc_44228_n10543_1;
  wire u2__abc_44228_n10544;
  wire u2__abc_44228_n10545;
  wire u2__abc_44228_n10546;
  wire u2__abc_44228_n10547;
  wire u2__abc_44228_n10548;
  wire u2__abc_44228_n10550_1;
  wire u2__abc_44228_n10551;
  wire u2__abc_44228_n10552;
  wire u2__abc_44228_n10553;
  wire u2__abc_44228_n10554;
  wire u2__abc_44228_n10555;
  wire u2__abc_44228_n10556_1;
  wire u2__abc_44228_n10557_1;
  wire u2__abc_44228_n10558;
  wire u2__abc_44228_n10559;
  wire u2__abc_44228_n10560;
  wire u2__abc_44228_n10561;
  wire u2__abc_44228_n10562;
  wire u2__abc_44228_n10563_1;
  wire u2__abc_44228_n10564_1;
  wire u2__abc_44228_n10565;
  wire u2__abc_44228_n10567;
  wire u2__abc_44228_n10568;
  wire u2__abc_44228_n10569;
  wire u2__abc_44228_n10570_1;
  wire u2__abc_44228_n10571_1;
  wire u2__abc_44228_n10572;
  wire u2__abc_44228_n10573;
  wire u2__abc_44228_n10574;
  wire u2__abc_44228_n10575;
  wire u2__abc_44228_n10576;
  wire u2__abc_44228_n10577_1;
  wire u2__abc_44228_n10578_1;
  wire u2__abc_44228_n10579;
  wire u2__abc_44228_n10580;
  wire u2__abc_44228_n10581;
  wire u2__abc_44228_n10582;
  wire u2__abc_44228_n10584_1;
  wire u2__abc_44228_n10585_1;
  wire u2__abc_44228_n10586;
  wire u2__abc_44228_n10587;
  wire u2__abc_44228_n10588;
  wire u2__abc_44228_n10589;
  wire u2__abc_44228_n10590;
  wire u2__abc_44228_n10591_1;
  wire u2__abc_44228_n10592_1;
  wire u2__abc_44228_n10593;
  wire u2__abc_44228_n10594;
  wire u2__abc_44228_n10595;
  wire u2__abc_44228_n10596;
  wire u2__abc_44228_n10597;
  wire u2__abc_44228_n10598_1;
  wire u2__abc_44228_n10599_1;
  wire u2__abc_44228_n10601;
  wire u2__abc_44228_n10602;
  wire u2__abc_44228_n10603;
  wire u2__abc_44228_n10604;
  wire u2__abc_44228_n10605_1;
  wire u2__abc_44228_n10606_1;
  wire u2__abc_44228_n10607;
  wire u2__abc_44228_n10608;
  wire u2__abc_44228_n10609;
  wire u2__abc_44228_n10610;
  wire u2__abc_44228_n10611;
  wire u2__abc_44228_n10612_1;
  wire u2__abc_44228_n10613_1;
  wire u2__abc_44228_n10614;
  wire u2__abc_44228_n10615;
  wire u2__abc_44228_n10616;
  wire u2__abc_44228_n10618;
  wire u2__abc_44228_n10619_1;
  wire u2__abc_44228_n10620_1;
  wire u2__abc_44228_n10621;
  wire u2__abc_44228_n10622;
  wire u2__abc_44228_n10623;
  wire u2__abc_44228_n10624;
  wire u2__abc_44228_n10625;
  wire u2__abc_44228_n10626_1;
  wire u2__abc_44228_n10627_1;
  wire u2__abc_44228_n10628;
  wire u2__abc_44228_n10629;
  wire u2__abc_44228_n10630;
  wire u2__abc_44228_n10631;
  wire u2__abc_44228_n10632;
  wire u2__abc_44228_n10633_1;
  wire u2__abc_44228_n10635;
  wire u2__abc_44228_n10636;
  wire u2__abc_44228_n10637;
  wire u2__abc_44228_n10638;
  wire u2__abc_44228_n10639;
  wire u2__abc_44228_n10640_1;
  wire u2__abc_44228_n10641_1;
  wire u2__abc_44228_n10642;
  wire u2__abc_44228_n10643;
  wire u2__abc_44228_n10644;
  wire u2__abc_44228_n10645;
  wire u2__abc_44228_n10646;
  wire u2__abc_44228_n10647_1;
  wire u2__abc_44228_n10648_1;
  wire u2__abc_44228_n10649;
  wire u2__abc_44228_n10650;
  wire u2__abc_44228_n10652;
  wire u2__abc_44228_n10653;
  wire u2__abc_44228_n10654_1;
  wire u2__abc_44228_n10655_1;
  wire u2__abc_44228_n10656;
  wire u2__abc_44228_n10657;
  wire u2__abc_44228_n10658;
  wire u2__abc_44228_n10659;
  wire u2__abc_44228_n10660;
  wire u2__abc_44228_n10661_1;
  wire u2__abc_44228_n10662_1;
  wire u2__abc_44228_n10663;
  wire u2__abc_44228_n10664;
  wire u2__abc_44228_n10665;
  wire u2__abc_44228_n10666;
  wire u2__abc_44228_n10667;
  wire u2__abc_44228_n10669_1;
  wire u2__abc_44228_n10670;
  wire u2__abc_44228_n10671;
  wire u2__abc_44228_n10672;
  wire u2__abc_44228_n10673;
  wire u2__abc_44228_n10674;
  wire u2__abc_44228_n10675_1;
  wire u2__abc_44228_n10676_1;
  wire u2__abc_44228_n10677;
  wire u2__abc_44228_n10678;
  wire u2__abc_44228_n10679;
  wire u2__abc_44228_n10680;
  wire u2__abc_44228_n10681;
  wire u2__abc_44228_n10682_1;
  wire u2__abc_44228_n10683_1;
  wire u2__abc_44228_n10684;
  wire u2__abc_44228_n10686;
  wire u2__abc_44228_n10687;
  wire u2__abc_44228_n10688;
  wire u2__abc_44228_n10689_1;
  wire u2__abc_44228_n10690_1;
  wire u2__abc_44228_n10691;
  wire u2__abc_44228_n10692;
  wire u2__abc_44228_n10693;
  wire u2__abc_44228_n10694;
  wire u2__abc_44228_n10695;
  wire u2__abc_44228_n10696_1;
  wire u2__abc_44228_n10697_1;
  wire u2__abc_44228_n10698;
  wire u2__abc_44228_n10699;
  wire u2__abc_44228_n10700;
  wire u2__abc_44228_n10701;
  wire u2__abc_44228_n10703_1;
  wire u2__abc_44228_n10704_1;
  wire u2__abc_44228_n10705;
  wire u2__abc_44228_n10706;
  wire u2__abc_44228_n10707;
  wire u2__abc_44228_n10708;
  wire u2__abc_44228_n10709;
  wire u2__abc_44228_n10710_1;
  wire u2__abc_44228_n10711_1;
  wire u2__abc_44228_n10712;
  wire u2__abc_44228_n10713;
  wire u2__abc_44228_n10714;
  wire u2__abc_44228_n10715;
  wire u2__abc_44228_n10716;
  wire u2__abc_44228_n10717_1;
  wire u2__abc_44228_n10718_1;
  wire u2__abc_44228_n10720;
  wire u2__abc_44228_n10721;
  wire u2__abc_44228_n10722;
  wire u2__abc_44228_n10723;
  wire u2__abc_44228_n10724_1;
  wire u2__abc_44228_n10725_1;
  wire u2__abc_44228_n10726;
  wire u2__abc_44228_n10727;
  wire u2__abc_44228_n10728;
  wire u2__abc_44228_n10729;
  wire u2__abc_44228_n10730;
  wire u2__abc_44228_n10731_1;
  wire u2__abc_44228_n10732_1;
  wire u2__abc_44228_n10733;
  wire u2__abc_44228_n10734;
  wire u2__abc_44228_n10735;
  wire u2__abc_44228_n10737;
  wire u2__abc_44228_n10738_1;
  wire u2__abc_44228_n10739_1;
  wire u2__abc_44228_n10740;
  wire u2__abc_44228_n10741;
  wire u2__abc_44228_n10742;
  wire u2__abc_44228_n10743;
  wire u2__abc_44228_n10744;
  wire u2__abc_44228_n10745_1;
  wire u2__abc_44228_n10746_1;
  wire u2__abc_44228_n10747;
  wire u2__abc_44228_n10748;
  wire u2__abc_44228_n10749;
  wire u2__abc_44228_n10750;
  wire u2__abc_44228_n10751;
  wire u2__abc_44228_n10752_1;
  wire u2__abc_44228_n10754;
  wire u2__abc_44228_n10755;
  wire u2__abc_44228_n10756;
  wire u2__abc_44228_n10757;
  wire u2__abc_44228_n10758;
  wire u2__abc_44228_n10759_1;
  wire u2__abc_44228_n10760_1;
  wire u2__abc_44228_n10761;
  wire u2__abc_44228_n10762;
  wire u2__abc_44228_n10763;
  wire u2__abc_44228_n10764;
  wire u2__abc_44228_n10765;
  wire u2__abc_44228_n10766_1;
  wire u2__abc_44228_n10767_1;
  wire u2__abc_44228_n10768;
  wire u2__abc_44228_n10769;
  wire u2__abc_44228_n10770;
  wire u2__abc_44228_n10772;
  wire u2__abc_44228_n10773_1;
  wire u2__abc_44228_n10774_1;
  wire u2__abc_44228_n10775;
  wire u2__abc_44228_n10776;
  wire u2__abc_44228_n10777;
  wire u2__abc_44228_n10778;
  wire u2__abc_44228_n10779;
  wire u2__abc_44228_n10780_1;
  wire u2__abc_44228_n10781_1;
  wire u2__abc_44228_n10782;
  wire u2__abc_44228_n10783;
  wire u2__abc_44228_n10784;
  wire u2__abc_44228_n10785;
  wire u2__abc_44228_n10786;
  wire u2__abc_44228_n10787_1;
  wire u2__abc_44228_n10789;
  wire u2__abc_44228_n10790;
  wire u2__abc_44228_n10791;
  wire u2__abc_44228_n10792;
  wire u2__abc_44228_n10793;
  wire u2__abc_44228_n10794_1;
  wire u2__abc_44228_n10795_1;
  wire u2__abc_44228_n10796;
  wire u2__abc_44228_n10797;
  wire u2__abc_44228_n10798;
  wire u2__abc_44228_n10799;
  wire u2__abc_44228_n10800;
  wire u2__abc_44228_n10801_1;
  wire u2__abc_44228_n10802_1;
  wire u2__abc_44228_n10803;
  wire u2__abc_44228_n10804;
  wire u2__abc_44228_n10806;
  wire u2__abc_44228_n10807;
  wire u2__abc_44228_n10808_1;
  wire u2__abc_44228_n10809_1;
  wire u2__abc_44228_n10810;
  wire u2__abc_44228_n10811;
  wire u2__abc_44228_n10812;
  wire u2__abc_44228_n10813;
  wire u2__abc_44228_n10814;
  wire u2__abc_44228_n10815_1;
  wire u2__abc_44228_n10816_1;
  wire u2__abc_44228_n10817;
  wire u2__abc_44228_n10818;
  wire u2__abc_44228_n10819;
  wire u2__abc_44228_n10820;
  wire u2__abc_44228_n10821;
  wire u2__abc_44228_n10823_1;
  wire u2__abc_44228_n10824;
  wire u2__abc_44228_n10825;
  wire u2__abc_44228_n10826;
  wire u2__abc_44228_n10827;
  wire u2__abc_44228_n10828;
  wire u2__abc_44228_n10829_1;
  wire u2__abc_44228_n10830_1;
  wire u2__abc_44228_n10831;
  wire u2__abc_44228_n10832;
  wire u2__abc_44228_n10833;
  wire u2__abc_44228_n10834;
  wire u2__abc_44228_n10835;
  wire u2__abc_44228_n10836_1;
  wire u2__abc_44228_n10837_1;
  wire u2__abc_44228_n10838;
  wire u2__abc_44228_n10840;
  wire u2__abc_44228_n10841;
  wire u2__abc_44228_n10842;
  wire u2__abc_44228_n10843_1;
  wire u2__abc_44228_n10844_1;
  wire u2__abc_44228_n10845;
  wire u2__abc_44228_n10846;
  wire u2__abc_44228_n10847;
  wire u2__abc_44228_n10848;
  wire u2__abc_44228_n10849;
  wire u2__abc_44228_n10850_1;
  wire u2__abc_44228_n10851_1;
  wire u2__abc_44228_n10852;
  wire u2__abc_44228_n10853;
  wire u2__abc_44228_n10854;
  wire u2__abc_44228_n10855;
  wire u2__abc_44228_n10857_1;
  wire u2__abc_44228_n10858_1;
  wire u2__abc_44228_n10859;
  wire u2__abc_44228_n10860;
  wire u2__abc_44228_n10861;
  wire u2__abc_44228_n10862;
  wire u2__abc_44228_n10863;
  wire u2__abc_44228_n10864_1;
  wire u2__abc_44228_n10865_1;
  wire u2__abc_44228_n10866;
  wire u2__abc_44228_n10867;
  wire u2__abc_44228_n10868;
  wire u2__abc_44228_n10869;
  wire u2__abc_44228_n10870;
  wire u2__abc_44228_n10871_1;
  wire u2__abc_44228_n10872_1;
  wire u2__abc_44228_n10874;
  wire u2__abc_44228_n10875;
  wire u2__abc_44228_n10876;
  wire u2__abc_44228_n10877;
  wire u2__abc_44228_n10878_1;
  wire u2__abc_44228_n10879_1;
  wire u2__abc_44228_n10880;
  wire u2__abc_44228_n10881;
  wire u2__abc_44228_n10882;
  wire u2__abc_44228_n10883;
  wire u2__abc_44228_n10884;
  wire u2__abc_44228_n10885_1;
  wire u2__abc_44228_n10886_1;
  wire u2__abc_44228_n10887;
  wire u2__abc_44228_n10888;
  wire u2__abc_44228_n10889;
  wire u2__abc_44228_n10891;
  wire u2__abc_44228_n10892_1;
  wire u2__abc_44228_n10893_1;
  wire u2__abc_44228_n10894;
  wire u2__abc_44228_n10895;
  wire u2__abc_44228_n10896;
  wire u2__abc_44228_n10897;
  wire u2__abc_44228_n10898;
  wire u2__abc_44228_n10899_1;
  wire u2__abc_44228_n10900_1;
  wire u2__abc_44228_n10901;
  wire u2__abc_44228_n10902;
  wire u2__abc_44228_n10903;
  wire u2__abc_44228_n10904;
  wire u2__abc_44228_n10905;
  wire u2__abc_44228_n10906_1;
  wire u2__abc_44228_n10908;
  wire u2__abc_44228_n10909;
  wire u2__abc_44228_n10910;
  wire u2__abc_44228_n10911;
  wire u2__abc_44228_n10912;
  wire u2__abc_44228_n10913_1;
  wire u2__abc_44228_n10914_1;
  wire u2__abc_44228_n10915;
  wire u2__abc_44228_n10916;
  wire u2__abc_44228_n10917;
  wire u2__abc_44228_n10918;
  wire u2__abc_44228_n10919;
  wire u2__abc_44228_n10920_1;
  wire u2__abc_44228_n10921_1;
  wire u2__abc_44228_n10922;
  wire u2__abc_44228_n10923;
  wire u2__abc_44228_n10925;
  wire u2__abc_44228_n10926;
  wire u2__abc_44228_n10927_1;
  wire u2__abc_44228_n10928_1;
  wire u2__abc_44228_n10929;
  wire u2__abc_44228_n10930;
  wire u2__abc_44228_n10931;
  wire u2__abc_44228_n10932;
  wire u2__abc_44228_n10933;
  wire u2__abc_44228_n10934_1;
  wire u2__abc_44228_n10935_1;
  wire u2__abc_44228_n10936;
  wire u2__abc_44228_n10937;
  wire u2__abc_44228_n10938;
  wire u2__abc_44228_n10939;
  wire u2__abc_44228_n10940;
  wire u2__abc_44228_n10942_1;
  wire u2__abc_44228_n10943;
  wire u2__abc_44228_n10944;
  wire u2__abc_44228_n10945;
  wire u2__abc_44228_n10946;
  wire u2__abc_44228_n10947;
  wire u2__abc_44228_n10948_1;
  wire u2__abc_44228_n10949_1;
  wire u2__abc_44228_n10950;
  wire u2__abc_44228_n10951;
  wire u2__abc_44228_n10952;
  wire u2__abc_44228_n10953;
  wire u2__abc_44228_n10954;
  wire u2__abc_44228_n10955_1;
  wire u2__abc_44228_n10956_1;
  wire u2__abc_44228_n10957;
  wire u2__abc_44228_n10959;
  wire u2__abc_44228_n10960;
  wire u2__abc_44228_n10961;
  wire u2__abc_44228_n10962_1;
  wire u2__abc_44228_n10963_1;
  wire u2__abc_44228_n10964;
  wire u2__abc_44228_n10965;
  wire u2__abc_44228_n10966;
  wire u2__abc_44228_n10967;
  wire u2__abc_44228_n10968;
  wire u2__abc_44228_n10969_1;
  wire u2__abc_44228_n10970_1;
  wire u2__abc_44228_n10971;
  wire u2__abc_44228_n10972;
  wire u2__abc_44228_n10973;
  wire u2__abc_44228_n10974;
  wire u2__abc_44228_n10976_1;
  wire u2__abc_44228_n10977_1;
  wire u2__abc_44228_n10978;
  wire u2__abc_44228_n10979;
  wire u2__abc_44228_n10980;
  wire u2__abc_44228_n10981;
  wire u2__abc_44228_n10982;
  wire u2__abc_44228_n10983_1;
  wire u2__abc_44228_n10984_1;
  wire u2__abc_44228_n10985;
  wire u2__abc_44228_n10986;
  wire u2__abc_44228_n10987;
  wire u2__abc_44228_n10988;
  wire u2__abc_44228_n10989;
  wire u2__abc_44228_n10990_1;
  wire u2__abc_44228_n10991_1;
  wire u2__abc_44228_n10993;
  wire u2__abc_44228_n10994;
  wire u2__abc_44228_n10995;
  wire u2__abc_44228_n10996;
  wire u2__abc_44228_n10997_1;
  wire u2__abc_44228_n10998_1;
  wire u2__abc_44228_n10999;
  wire u2__abc_44228_n11000;
  wire u2__abc_44228_n11001;
  wire u2__abc_44228_n11002;
  wire u2__abc_44228_n11003;
  wire u2__abc_44228_n11004_1;
  wire u2__abc_44228_n11005_1;
  wire u2__abc_44228_n11006;
  wire u2__abc_44228_n11007;
  wire u2__abc_44228_n11008;
  wire u2__abc_44228_n11009;
  wire u2__abc_44228_n11011_1;
  wire u2__abc_44228_n11012_1;
  wire u2__abc_44228_n11013;
  wire u2__abc_44228_n11014;
  wire u2__abc_44228_n11015;
  wire u2__abc_44228_n11016;
  wire u2__abc_44228_n11017;
  wire u2__abc_44228_n11018_1;
  wire u2__abc_44228_n11019_1;
  wire u2__abc_44228_n11020;
  wire u2__abc_44228_n11021;
  wire u2__abc_44228_n11022;
  wire u2__abc_44228_n11023;
  wire u2__abc_44228_n11024;
  wire u2__abc_44228_n11025_1;
  wire u2__abc_44228_n11026_1;
  wire u2__abc_44228_n11028;
  wire u2__abc_44228_n11029;
  wire u2__abc_44228_n11030;
  wire u2__abc_44228_n11031;
  wire u2__abc_44228_n11032_1;
  wire u2__abc_44228_n11033_1;
  wire u2__abc_44228_n11034;
  wire u2__abc_44228_n11035;
  wire u2__abc_44228_n11036;
  wire u2__abc_44228_n11037;
  wire u2__abc_44228_n11038;
  wire u2__abc_44228_n11039_1;
  wire u2__abc_44228_n11040_1;
  wire u2__abc_44228_n11041;
  wire u2__abc_44228_n11042;
  wire u2__abc_44228_n11043;
  wire u2__abc_44228_n11045;
  wire u2__abc_44228_n11046_1;
  wire u2__abc_44228_n11047_1;
  wire u2__abc_44228_n11048;
  wire u2__abc_44228_n11049;
  wire u2__abc_44228_n11050;
  wire u2__abc_44228_n11051;
  wire u2__abc_44228_n11052;
  wire u2__abc_44228_n11053_1;
  wire u2__abc_44228_n11054_1;
  wire u2__abc_44228_n11055;
  wire u2__abc_44228_n11056;
  wire u2__abc_44228_n11057;
  wire u2__abc_44228_n11058;
  wire u2__abc_44228_n11059;
  wire u2__abc_44228_n11060_1;
  wire u2__abc_44228_n11062;
  wire u2__abc_44228_n11063;
  wire u2__abc_44228_n11064;
  wire u2__abc_44228_n11065;
  wire u2__abc_44228_n11066;
  wire u2__abc_44228_n11067_1;
  wire u2__abc_44228_n11068_1;
  wire u2__abc_44228_n11069;
  wire u2__abc_44228_n11070;
  wire u2__abc_44228_n11071;
  wire u2__abc_44228_n11072;
  wire u2__abc_44228_n11073;
  wire u2__abc_44228_n11074_1;
  wire u2__abc_44228_n11075_1;
  wire u2__abc_44228_n11076;
  wire u2__abc_44228_n11077;
  wire u2__abc_44228_n11079;
  wire u2__abc_44228_n11080;
  wire u2__abc_44228_n11081_1;
  wire u2__abc_44228_n11082_1;
  wire u2__abc_44228_n11083;
  wire u2__abc_44228_n11084;
  wire u2__abc_44228_n11085;
  wire u2__abc_44228_n11086;
  wire u2__abc_44228_n11087;
  wire u2__abc_44228_n11088_1;
  wire u2__abc_44228_n11089_1;
  wire u2__abc_44228_n11090;
  wire u2__abc_44228_n11091;
  wire u2__abc_44228_n11092;
  wire u2__abc_44228_n11093;
  wire u2__abc_44228_n11094;
  wire u2__abc_44228_n11096_1;
  wire u2__abc_44228_n11097;
  wire u2__abc_44228_n11098;
  wire u2__abc_44228_n11099;
  wire u2__abc_44228_n11100;
  wire u2__abc_44228_n11101;
  wire u2__abc_44228_n11102_1;
  wire u2__abc_44228_n11103_1;
  wire u2__abc_44228_n11104;
  wire u2__abc_44228_n11105;
  wire u2__abc_44228_n11106;
  wire u2__abc_44228_n11107;
  wire u2__abc_44228_n11108;
  wire u2__abc_44228_n11109_1;
  wire u2__abc_44228_n11110_1;
  wire u2__abc_44228_n11111;
  wire u2__abc_44228_n11113;
  wire u2__abc_44228_n11114;
  wire u2__abc_44228_n11115;
  wire u2__abc_44228_n11116_1;
  wire u2__abc_44228_n11117_1;
  wire u2__abc_44228_n11118;
  wire u2__abc_44228_n11119;
  wire u2__abc_44228_n11120;
  wire u2__abc_44228_n11121;
  wire u2__abc_44228_n11122;
  wire u2__abc_44228_n11123_1;
  wire u2__abc_44228_n11124_1;
  wire u2__abc_44228_n11125;
  wire u2__abc_44228_n11126;
  wire u2__abc_44228_n11127;
  wire u2__abc_44228_n11128;
  wire u2__abc_44228_n11130_1;
  wire u2__abc_44228_n11131_1;
  wire u2__abc_44228_n11132;
  wire u2__abc_44228_n11133;
  wire u2__abc_44228_n11134;
  wire u2__abc_44228_n11135;
  wire u2__abc_44228_n11136;
  wire u2__abc_44228_n11137_1;
  wire u2__abc_44228_n11138_1;
  wire u2__abc_44228_n11139;
  wire u2__abc_44228_n11140;
  wire u2__abc_44228_n11141;
  wire u2__abc_44228_n11142;
  wire u2__abc_44228_n11143;
  wire u2__abc_44228_n11144_1;
  wire u2__abc_44228_n11145_1;
  wire u2__abc_44228_n11147;
  wire u2__abc_44228_n11148;
  wire u2__abc_44228_n11149;
  wire u2__abc_44228_n11150;
  wire u2__abc_44228_n11151_1;
  wire u2__abc_44228_n11152_1;
  wire u2__abc_44228_n11153;
  wire u2__abc_44228_n11154;
  wire u2__abc_44228_n11155;
  wire u2__abc_44228_n11156;
  wire u2__abc_44228_n11157;
  wire u2__abc_44228_n11158_1;
  wire u2__abc_44228_n11159_1;
  wire u2__abc_44228_n11160;
  wire u2__abc_44228_n11161;
  wire u2__abc_44228_n11162;
  wire u2__abc_44228_n11164;
  wire u2__abc_44228_n11165_1;
  wire u2__abc_44228_n11166_1;
  wire u2__abc_44228_n11167;
  wire u2__abc_44228_n11168;
  wire u2__abc_44228_n11169;
  wire u2__abc_44228_n11170;
  wire u2__abc_44228_n11171;
  wire u2__abc_44228_n11172_1;
  wire u2__abc_44228_n11173_1;
  wire u2__abc_44228_n11174;
  wire u2__abc_44228_n11175;
  wire u2__abc_44228_n11176;
  wire u2__abc_44228_n11177;
  wire u2__abc_44228_n11178;
  wire u2__abc_44228_n11179_1;
  wire u2__abc_44228_n11181;
  wire u2__abc_44228_n11182;
  wire u2__abc_44228_n11183;
  wire u2__abc_44228_n11184;
  wire u2__abc_44228_n11185;
  wire u2__abc_44228_n11186_1;
  wire u2__abc_44228_n11187_1;
  wire u2__abc_44228_n11188;
  wire u2__abc_44228_n11189;
  wire u2__abc_44228_n11190;
  wire u2__abc_44228_n11191;
  wire u2__abc_44228_n11192;
  wire u2__abc_44228_n11193_1;
  wire u2__abc_44228_n11194_1;
  wire u2__abc_44228_n11195;
  wire u2__abc_44228_n11196;
  wire u2__abc_44228_n11198;
  wire u2__abc_44228_n11199;
  wire u2__abc_44228_n11200_1;
  wire u2__abc_44228_n11201_1;
  wire u2__abc_44228_n11202;
  wire u2__abc_44228_n11203;
  wire u2__abc_44228_n11204;
  wire u2__abc_44228_n11205;
  wire u2__abc_44228_n11206;
  wire u2__abc_44228_n11207_1;
  wire u2__abc_44228_n11208_1;
  wire u2__abc_44228_n11209;
  wire u2__abc_44228_n11210;
  wire u2__abc_44228_n11211;
  wire u2__abc_44228_n11212;
  wire u2__abc_44228_n11213;
  wire u2__abc_44228_n11214_1;
  wire u2__abc_44228_n11216;
  wire u2__abc_44228_n11217;
  wire u2__abc_44228_n11218;
  wire u2__abc_44228_n11219;
  wire u2__abc_44228_n11220;
  wire u2__abc_44228_n11221_1;
  wire u2__abc_44228_n11222_1;
  wire u2__abc_44228_n11223;
  wire u2__abc_44228_n11224;
  wire u2__abc_44228_n11225;
  wire u2__abc_44228_n11226;
  wire u2__abc_44228_n11227;
  wire u2__abc_44228_n11228_1;
  wire u2__abc_44228_n11229_1;
  wire u2__abc_44228_n11230;
  wire u2__abc_44228_n11231;
  wire u2__abc_44228_n11233;
  wire u2__abc_44228_n11234;
  wire u2__abc_44228_n11235_1;
  wire u2__abc_44228_n11236_1;
  wire u2__abc_44228_n11237;
  wire u2__abc_44228_n11238;
  wire u2__abc_44228_n11239;
  wire u2__abc_44228_n11240;
  wire u2__abc_44228_n11241;
  wire u2__abc_44228_n11242_1;
  wire u2__abc_44228_n11243_1;
  wire u2__abc_44228_n11244;
  wire u2__abc_44228_n11245;
  wire u2__abc_44228_n11246;
  wire u2__abc_44228_n11247;
  wire u2__abc_44228_n11248;
  wire u2__abc_44228_n11250_1;
  wire u2__abc_44228_n11251;
  wire u2__abc_44228_n11252;
  wire u2__abc_44228_n11253;
  wire u2__abc_44228_n11254;
  wire u2__abc_44228_n11255;
  wire u2__abc_44228_n11256_1;
  wire u2__abc_44228_n11257_1;
  wire u2__abc_44228_n11258;
  wire u2__abc_44228_n11259;
  wire u2__abc_44228_n11260;
  wire u2__abc_44228_n11261;
  wire u2__abc_44228_n11262;
  wire u2__abc_44228_n11263_1;
  wire u2__abc_44228_n11264_1;
  wire u2__abc_44228_n11265;
  wire u2__abc_44228_n11267;
  wire u2__abc_44228_n11268;
  wire u2__abc_44228_n11269;
  wire u2__abc_44228_n11270_1;
  wire u2__abc_44228_n11271_1;
  wire u2__abc_44228_n11272;
  wire u2__abc_44228_n11273;
  wire u2__abc_44228_n11274;
  wire u2__abc_44228_n11275;
  wire u2__abc_44228_n11276;
  wire u2__abc_44228_n11277_1;
  wire u2__abc_44228_n11278_1;
  wire u2__abc_44228_n11279;
  wire u2__abc_44228_n11280;
  wire u2__abc_44228_n11281;
  wire u2__abc_44228_n11282;
  wire u2__abc_44228_n11283;
  wire u2__abc_44228_n11285_1;
  wire u2__abc_44228_n11286;
  wire u2__abc_44228_n11287;
  wire u2__abc_44228_n11288;
  wire u2__abc_44228_n11289;
  wire u2__abc_44228_n11290;
  wire u2__abc_44228_n11291_1;
  wire u2__abc_44228_n11292_1;
  wire u2__abc_44228_n11293;
  wire u2__abc_44228_n11294;
  wire u2__abc_44228_n11295;
  wire u2__abc_44228_n11296;
  wire u2__abc_44228_n11297;
  wire u2__abc_44228_n11298_1;
  wire u2__abc_44228_n11299_1;
  wire u2__abc_44228_n11300;
  wire u2__abc_44228_n11302;
  wire u2__abc_44228_n11303;
  wire u2__abc_44228_n11304;
  wire u2__abc_44228_n11305_1;
  wire u2__abc_44228_n11306_1;
  wire u2__abc_44228_n11307;
  wire u2__abc_44228_n11308;
  wire u2__abc_44228_n11309;
  wire u2__abc_44228_n11310;
  wire u2__abc_44228_n11311;
  wire u2__abc_44228_n11312_1;
  wire u2__abc_44228_n11313_1;
  wire u2__abc_44228_n11314;
  wire u2__abc_44228_n11315;
  wire u2__abc_44228_n11316;
  wire u2__abc_44228_n11317;
  wire u2__abc_44228_n11319_1;
  wire u2__abc_44228_n11320_1;
  wire u2__abc_44228_n11321;
  wire u2__abc_44228_n11322;
  wire u2__abc_44228_n11323;
  wire u2__abc_44228_n11324;
  wire u2__abc_44228_n11325;
  wire u2__abc_44228_n11326_1;
  wire u2__abc_44228_n11327_1;
  wire u2__abc_44228_n11328;
  wire u2__abc_44228_n11329;
  wire u2__abc_44228_n11330;
  wire u2__abc_44228_n11331;
  wire u2__abc_44228_n11332;
  wire u2__abc_44228_n11333_1;
  wire u2__abc_44228_n11334_1;
  wire u2__abc_44228_n11336;
  wire u2__abc_44228_n11337;
  wire u2__abc_44228_n11338;
  wire u2__abc_44228_n11339;
  wire u2__abc_44228_n11340_1;
  wire u2__abc_44228_n11341_1;
  wire u2__abc_44228_n11342;
  wire u2__abc_44228_n11343;
  wire u2__abc_44228_n11344;
  wire u2__abc_44228_n11345;
  wire u2__abc_44228_n11346;
  wire u2__abc_44228_n11347_1;
  wire u2__abc_44228_n11348_1;
  wire u2__abc_44228_n11349;
  wire u2__abc_44228_n11350;
  wire u2__abc_44228_n11351;
  wire u2__abc_44228_n11352;
  wire u2__abc_44228_n11354_1;
  wire u2__abc_44228_n11355_1;
  wire u2__abc_44228_n11356;
  wire u2__abc_44228_n11357;
  wire u2__abc_44228_n11358;
  wire u2__abc_44228_n11359;
  wire u2__abc_44228_n11360;
  wire u2__abc_44228_n11361_1;
  wire u2__abc_44228_n11362_1;
  wire u2__abc_44228_n11363;
  wire u2__abc_44228_n11364;
  wire u2__abc_44228_n11365;
  wire u2__abc_44228_n11366;
  wire u2__abc_44228_n11367;
  wire u2__abc_44228_n11368_1;
  wire u2__abc_44228_n11369_1;
  wire u2__abc_44228_n11371;
  wire u2__abc_44228_n11372;
  wire u2__abc_44228_n11373;
  wire u2__abc_44228_n11374;
  wire u2__abc_44228_n11375_1;
  wire u2__abc_44228_n11376_1;
  wire u2__abc_44228_n11377;
  wire u2__abc_44228_n11378;
  wire u2__abc_44228_n11379;
  wire u2__abc_44228_n11380;
  wire u2__abc_44228_n11381;
  wire u2__abc_44228_n11382_1;
  wire u2__abc_44228_n11383_1;
  wire u2__abc_44228_n11384;
  wire u2__abc_44228_n11385;
  wire u2__abc_44228_n11386;
  wire u2__abc_44228_n11388;
  wire u2__abc_44228_n11389_1;
  wire u2__abc_44228_n11390_1;
  wire u2__abc_44228_n11391;
  wire u2__abc_44228_n11392;
  wire u2__abc_44228_n11393;
  wire u2__abc_44228_n11394;
  wire u2__abc_44228_n11395;
  wire u2__abc_44228_n11396_1;
  wire u2__abc_44228_n11397_1;
  wire u2__abc_44228_n11398;
  wire u2__abc_44228_n11399;
  wire u2__abc_44228_n11400;
  wire u2__abc_44228_n11401;
  wire u2__abc_44228_n11402;
  wire u2__abc_44228_n11403_1;
  wire u2__abc_44228_n11405;
  wire u2__abc_44228_n11406;
  wire u2__abc_44228_n11407;
  wire u2__abc_44228_n11408;
  wire u2__abc_44228_n11409;
  wire u2__abc_44228_n11410_1;
  wire u2__abc_44228_n11411_1;
  wire u2__abc_44228_n11412;
  wire u2__abc_44228_n11413;
  wire u2__abc_44228_n11414;
  wire u2__abc_44228_n11415;
  wire u2__abc_44228_n11416;
  wire u2__abc_44228_n11417_1;
  wire u2__abc_44228_n11418_1;
  wire u2__abc_44228_n11419;
  wire u2__abc_44228_n11420;
  wire u2__abc_44228_n11422;
  wire u2__abc_44228_n11423;
  wire u2__abc_44228_n11424_1;
  wire u2__abc_44228_n11425_1;
  wire u2__abc_44228_n11426;
  wire u2__abc_44228_n11427;
  wire u2__abc_44228_n11428;
  wire u2__abc_44228_n11429;
  wire u2__abc_44228_n11430;
  wire u2__abc_44228_n11431_1;
  wire u2__abc_44228_n11432_1;
  wire u2__abc_44228_n11433;
  wire u2__abc_44228_n11434;
  wire u2__abc_44228_n11435;
  wire u2__abc_44228_n11436;
  wire u2__abc_44228_n11437;
  wire u2__abc_44228_n11439_1;
  wire u2__abc_44228_n11440;
  wire u2__abc_44228_n11441;
  wire u2__abc_44228_n11442;
  wire u2__abc_44228_n11443;
  wire u2__abc_44228_n11444;
  wire u2__abc_44228_n11445_1;
  wire u2__abc_44228_n11446_1;
  wire u2__abc_44228_n11447;
  wire u2__abc_44228_n11448;
  wire u2__abc_44228_n11449;
  wire u2__abc_44228_n11450;
  wire u2__abc_44228_n11451;
  wire u2__abc_44228_n11452_1;
  wire u2__abc_44228_n11453_1;
  wire u2__abc_44228_n11454;
  wire u2__abc_44228_n11456;
  wire u2__abc_44228_n11457;
  wire u2__abc_44228_n11458;
  wire u2__abc_44228_n11459_1;
  wire u2__abc_44228_n11460_1;
  wire u2__abc_44228_n11461;
  wire u2__abc_44228_n11462;
  wire u2__abc_44228_n11463;
  wire u2__abc_44228_n11464;
  wire u2__abc_44228_n11465;
  wire u2__abc_44228_n11466_1;
  wire u2__abc_44228_n11467_1;
  wire u2__abc_44228_n11468;
  wire u2__abc_44228_n11469;
  wire u2__abc_44228_n11470;
  wire u2__abc_44228_n11471;
  wire u2__abc_44228_n11473_1;
  wire u2__abc_44228_n11474_1;
  wire u2__abc_44228_n11475;
  wire u2__abc_44228_n11476;
  wire u2__abc_44228_n11477;
  wire u2__abc_44228_n11478;
  wire u2__abc_44228_n11479;
  wire u2__abc_44228_n11480_1;
  wire u2__abc_44228_n11481_1;
  wire u2__abc_44228_n11482;
  wire u2__abc_44228_n11483;
  wire u2__abc_44228_n11484;
  wire u2__abc_44228_n11485;
  wire u2__abc_44228_n11486;
  wire u2__abc_44228_n11487_1;
  wire u2__abc_44228_n11488_1;
  wire u2__abc_44228_n11489;
  wire u2__abc_44228_n11491;
  wire u2__abc_44228_n11492;
  wire u2__abc_44228_n11493;
  wire u2__abc_44228_n11494_1;
  wire u2__abc_44228_n11495_1;
  wire u2__abc_44228_n11496;
  wire u2__abc_44228_n11497;
  wire u2__abc_44228_n11498;
  wire u2__abc_44228_n11499;
  wire u2__abc_44228_n11500;
  wire u2__abc_44228_n11501_1;
  wire u2__abc_44228_n11502_1;
  wire u2__abc_44228_n11503;
  wire u2__abc_44228_n11504;
  wire u2__abc_44228_n11505;
  wire u2__abc_44228_n11506;
  wire u2__abc_44228_n11508_1;
  wire u2__abc_44228_n11509_1;
  wire u2__abc_44228_n11510;
  wire u2__abc_44228_n11511;
  wire u2__abc_44228_n11512;
  wire u2__abc_44228_n11513;
  wire u2__abc_44228_n11514;
  wire u2__abc_44228_n11515_1;
  wire u2__abc_44228_n11516_1;
  wire u2__abc_44228_n11517;
  wire u2__abc_44228_n11518;
  wire u2__abc_44228_n11519;
  wire u2__abc_44228_n11520;
  wire u2__abc_44228_n11521;
  wire u2__abc_44228_n11522_1;
  wire u2__abc_44228_n11523_1;
  wire u2__abc_44228_n11525;
  wire u2__abc_44228_n11526;
  wire u2__abc_44228_n11527;
  wire u2__abc_44228_n11528;
  wire u2__abc_44228_n11529_1;
  wire u2__abc_44228_n11530_1;
  wire u2__abc_44228_n11531;
  wire u2__abc_44228_n11532;
  wire u2__abc_44228_n11533;
  wire u2__abc_44228_n11534;
  wire u2__abc_44228_n11535;
  wire u2__abc_44228_n11536_1;
  wire u2__abc_44228_n11537_1;
  wire u2__abc_44228_n11538;
  wire u2__abc_44228_n11539;
  wire u2__abc_44228_n11540;
  wire u2__abc_44228_n11542;
  wire u2__abc_44228_n11543_1;
  wire u2__abc_44228_n11544_1;
  wire u2__abc_44228_n11545;
  wire u2__abc_44228_n11546;
  wire u2__abc_44228_n11547;
  wire u2__abc_44228_n11548;
  wire u2__abc_44228_n11549;
  wire u2__abc_44228_n11550_1;
  wire u2__abc_44228_n11551_1;
  wire u2__abc_44228_n11552;
  wire u2__abc_44228_n11553;
  wire u2__abc_44228_n11554;
  wire u2__abc_44228_n11555;
  wire u2__abc_44228_n11556;
  wire u2__abc_44228_n11557_1;
  wire u2__abc_44228_n11559;
  wire u2__abc_44228_n11560;
  wire u2__abc_44228_n11561;
  wire u2__abc_44228_n11562;
  wire u2__abc_44228_n11563;
  wire u2__abc_44228_n11564_1;
  wire u2__abc_44228_n11565_1;
  wire u2__abc_44228_n11566;
  wire u2__abc_44228_n11567;
  wire u2__abc_44228_n11568;
  wire u2__abc_44228_n11569;
  wire u2__abc_44228_n11570;
  wire u2__abc_44228_n11571_1;
  wire u2__abc_44228_n11572_1;
  wire u2__abc_44228_n11573;
  wire u2__abc_44228_n11574;
  wire u2__abc_44228_n11576;
  wire u2__abc_44228_n11577;
  wire u2__abc_44228_n11578_1;
  wire u2__abc_44228_n11579_1;
  wire u2__abc_44228_n11580;
  wire u2__abc_44228_n11581;
  wire u2__abc_44228_n11582;
  wire u2__abc_44228_n11583;
  wire u2__abc_44228_n11584;
  wire u2__abc_44228_n11585_1;
  wire u2__abc_44228_n11586_1;
  wire u2__abc_44228_n11587;
  wire u2__abc_44228_n11588;
  wire u2__abc_44228_n11589;
  wire u2__abc_44228_n11590;
  wire u2__abc_44228_n11591;
  wire u2__abc_44228_n11592_1;
  wire u2__abc_44228_n11594;
  wire u2__abc_44228_n11595;
  wire u2__abc_44228_n11596;
  wire u2__abc_44228_n11597;
  wire u2__abc_44228_n11598;
  wire u2__abc_44228_n11599_1;
  wire u2__abc_44228_n11600_1;
  wire u2__abc_44228_n11601;
  wire u2__abc_44228_n11602;
  wire u2__abc_44228_n11603;
  wire u2__abc_44228_n11604;
  wire u2__abc_44228_n11605;
  wire u2__abc_44228_n11606_1;
  wire u2__abc_44228_n11607_1;
  wire u2__abc_44228_n11608;
  wire u2__abc_44228_n11609;
  wire u2__abc_44228_n11611;
  wire u2__abc_44228_n11612;
  wire u2__abc_44228_n11613_1;
  wire u2__abc_44228_n11614_1;
  wire u2__abc_44228_n11615;
  wire u2__abc_44228_n11616;
  wire u2__abc_44228_n11617;
  wire u2__abc_44228_n11618;
  wire u2__abc_44228_n11619;
  wire u2__abc_44228_n11620_1;
  wire u2__abc_44228_n11621_1;
  wire u2__abc_44228_n11622;
  wire u2__abc_44228_n11623;
  wire u2__abc_44228_n11624;
  wire u2__abc_44228_n11625;
  wire u2__abc_44228_n11626;
  wire u2__abc_44228_n11627_1;
  wire u2__abc_44228_n11629;
  wire u2__abc_44228_n11630;
  wire u2__abc_44228_n11631;
  wire u2__abc_44228_n11632;
  wire u2__abc_44228_n11633;
  wire u2__abc_44228_n11634_1;
  wire u2__abc_44228_n11635_1;
  wire u2__abc_44228_n11636;
  wire u2__abc_44228_n11637;
  wire u2__abc_44228_n11638;
  wire u2__abc_44228_n11639;
  wire u2__abc_44228_n11640;
  wire u2__abc_44228_n11641_1;
  wire u2__abc_44228_n11642_1;
  wire u2__abc_44228_n11643;
  wire u2__abc_44228_n11644;
  wire u2__abc_44228_n11646;
  wire u2__abc_44228_n11647;
  wire u2__abc_44228_n11648_1;
  wire u2__abc_44228_n11649_1;
  wire u2__abc_44228_n11650;
  wire u2__abc_44228_n11651;
  wire u2__abc_44228_n11652;
  wire u2__abc_44228_n11653;
  wire u2__abc_44228_n11654;
  wire u2__abc_44228_n11655_1;
  wire u2__abc_44228_n11656_1;
  wire u2__abc_44228_n11657;
  wire u2__abc_44228_n11658;
  wire u2__abc_44228_n11659;
  wire u2__abc_44228_n11660;
  wire u2__abc_44228_n11661;
  wire u2__abc_44228_n11663_1;
  wire u2__abc_44228_n11664;
  wire u2__abc_44228_n11665;
  wire u2__abc_44228_n11666;
  wire u2__abc_44228_n11667;
  wire u2__abc_44228_n11668;
  wire u2__abc_44228_n11669_1;
  wire u2__abc_44228_n11670;
  wire u2__abc_44228_n11671;
  wire u2__abc_44228_n11672;
  wire u2__abc_44228_n11673;
  wire u2__abc_44228_n11674_1;
  wire u2__abc_44228_n11675;
  wire u2__abc_44228_n11676;
  wire u2__abc_44228_n11677;
  wire u2__abc_44228_n11678;
  wire u2__abc_44228_n11680;
  wire u2__abc_44228_n11681;
  wire u2__abc_44228_n11682;
  wire u2__abc_44228_n11683;
  wire u2__abc_44228_n11684_1;
  wire u2__abc_44228_n11685;
  wire u2__abc_44228_n11686;
  wire u2__abc_44228_n11687;
  wire u2__abc_44228_n11688;
  wire u2__abc_44228_n11689;
  wire u2__abc_44228_n11690_1;
  wire u2__abc_44228_n11691;
  wire u2__abc_44228_n11692;
  wire u2__abc_44228_n11693;
  wire u2__abc_44228_n11694;
  wire u2__abc_44228_n11695;
  wire u2__abc_44228_n11696;
  wire u2__abc_44228_n11698;
  wire u2__abc_44228_n11699;
  wire u2__abc_44228_n11700;
  wire u2__abc_44228_n11701;
  wire u2__abc_44228_n11702;
  wire u2__abc_44228_n11703;
  wire u2__abc_44228_n11704_1;
  wire u2__abc_44228_n11705;
  wire u2__abc_44228_n11706;
  wire u2__abc_44228_n11707;
  wire u2__abc_44228_n11708;
  wire u2__abc_44228_n11709;
  wire u2__abc_44228_n11710;
  wire u2__abc_44228_n11711_1;
  wire u2__abc_44228_n11712;
  wire u2__abc_44228_n11713;
  wire u2__abc_44228_n11715;
  wire u2__abc_44228_n11716;
  wire u2__abc_44228_n11717;
  wire u2__abc_44228_n11718;
  wire u2__abc_44228_n11719_1;
  wire u2__abc_44228_n11720;
  wire u2__abc_44228_n11721;
  wire u2__abc_44228_n11722;
  wire u2__abc_44228_n11723;
  wire u2__abc_44228_n11724;
  wire u2__abc_44228_n11725;
  wire u2__abc_44228_n11726_1;
  wire u2__abc_44228_n11727;
  wire u2__abc_44228_n11728;
  wire u2__abc_44228_n11729;
  wire u2__abc_44228_n11730;
  wire u2__abc_44228_n11732;
  wire u2__abc_44228_n11733;
  wire u2__abc_44228_n11734_1;
  wire u2__abc_44228_n11735;
  wire u2__abc_44228_n11736;
  wire u2__abc_44228_n11737;
  wire u2__abc_44228_n11738;
  wire u2__abc_44228_n11739;
  wire u2__abc_44228_n11740;
  wire u2__abc_44228_n11741_1;
  wire u2__abc_44228_n11742;
  wire u2__abc_44228_n11743;
  wire u2__abc_44228_n11744;
  wire u2__abc_44228_n11745;
  wire u2__abc_44228_n11746;
  wire u2__abc_44228_n11747;
  wire u2__abc_44228_n11749;
  wire u2__abc_44228_n11750_1;
  wire u2__abc_44228_n11751;
  wire u2__abc_44228_n11752;
  wire u2__abc_44228_n11753;
  wire u2__abc_44228_n11754;
  wire u2__abc_44228_n11755;
  wire u2__abc_44228_n11756;
  wire u2__abc_44228_n11757_1;
  wire u2__abc_44228_n11758;
  wire u2__abc_44228_n11759;
  wire u2__abc_44228_n11760;
  wire u2__abc_44228_n11761;
  wire u2__abc_44228_n11762;
  wire u2__abc_44228_n11763;
  wire u2__abc_44228_n11764;
  wire u2__abc_44228_n11765_1;
  wire u2__abc_44228_n11767;
  wire u2__abc_44228_n11768;
  wire u2__abc_44228_n11769;
  wire u2__abc_44228_n11770;
  wire u2__abc_44228_n11771;
  wire u2__abc_44228_n11772_1;
  wire u2__abc_44228_n11773;
  wire u2__abc_44228_n11774;
  wire u2__abc_44228_n11775;
  wire u2__abc_44228_n11776;
  wire u2__abc_44228_n11777;
  wire u2__abc_44228_n11778;
  wire u2__abc_44228_n11779;
  wire u2__abc_44228_n11780;
  wire u2__abc_44228_n11781_1;
  wire u2__abc_44228_n11782;
  wire u2__abc_44228_n11784;
  wire u2__abc_44228_n11785;
  wire u2__abc_44228_n11786;
  wire u2__abc_44228_n11787;
  wire u2__abc_44228_n11788_1;
  wire u2__abc_44228_n11789;
  wire u2__abc_44228_n11790;
  wire u2__abc_44228_n11791;
  wire u2__abc_44228_n11792;
  wire u2__abc_44228_n11793;
  wire u2__abc_44228_n11794;
  wire u2__abc_44228_n11795;
  wire u2__abc_44228_n11796_1;
  wire u2__abc_44228_n11797;
  wire u2__abc_44228_n11798;
  wire u2__abc_44228_n11799;
  wire u2__abc_44228_n11801;
  wire u2__abc_44228_n11802;
  wire u2__abc_44228_n11803_1;
  wire u2__abc_44228_n11804;
  wire u2__abc_44228_n11805;
  wire u2__abc_44228_n11806;
  wire u2__abc_44228_n11807;
  wire u2__abc_44228_n11808;
  wire u2__abc_44228_n11809;
  wire u2__abc_44228_n11810;
  wire u2__abc_44228_n11811;
  wire u2__abc_44228_n11812;
  wire u2__abc_44228_n11813_1;
  wire u2__abc_44228_n11814;
  wire u2__abc_44228_n11815;
  wire u2__abc_44228_n11816;
  wire u2__abc_44228_n11818;
  wire u2__abc_44228_n11819;
  wire u2__abc_44228_n11820_1;
  wire u2__abc_44228_n11821;
  wire u2__abc_44228_n11822;
  wire u2__abc_44228_n11823;
  wire u2__abc_44228_n11824;
  wire u2__abc_44228_n11825;
  wire u2__abc_44228_n11826;
  wire u2__abc_44228_n11827;
  wire u2__abc_44228_n11828_1;
  wire u2__abc_44228_n11829;
  wire u2__abc_44228_n11830;
  wire u2__abc_44228_n11831;
  wire u2__abc_44228_n11832;
  wire u2__abc_44228_n11833;
  wire u2__abc_44228_n11834;
  wire u2__abc_44228_n11836;
  wire u2__abc_44228_n11837;
  wire u2__abc_44228_n11838;
  wire u2__abc_44228_n11839;
  wire u2__abc_44228_n11840;
  wire u2__abc_44228_n11841;
  wire u2__abc_44228_n11842;
  wire u2__abc_44228_n11843;
  wire u2__abc_44228_n11844_1;
  wire u2__abc_44228_n11845;
  wire u2__abc_44228_n11846;
  wire u2__abc_44228_n11847;
  wire u2__abc_44228_n11848;
  wire u2__abc_44228_n11849;
  wire u2__abc_44228_n11850;
  wire u2__abc_44228_n11851_1;
  wire u2__abc_44228_n11853;
  wire u2__abc_44228_n11854;
  wire u2__abc_44228_n11855;
  wire u2__abc_44228_n11856;
  wire u2__abc_44228_n11857;
  wire u2__abc_44228_n11858;
  wire u2__abc_44228_n11859_1;
  wire u2__abc_44228_n11860;
  wire u2__abc_44228_n11861;
  wire u2__abc_44228_n11862;
  wire u2__abc_44228_n11863;
  wire u2__abc_44228_n11864;
  wire u2__abc_44228_n11865;
  wire u2__abc_44228_n11866_1;
  wire u2__abc_44228_n11867;
  wire u2__abc_44228_n11868;
  wire u2__abc_44228_n11870;
  wire u2__abc_44228_n11871;
  wire u2__abc_44228_n11872;
  wire u2__abc_44228_n11873;
  wire u2__abc_44228_n11874;
  wire u2__abc_44228_n11875;
  wire u2__abc_44228_n11876_1;
  wire u2__abc_44228_n11877;
  wire u2__abc_44228_n11878;
  wire u2__abc_44228_n11879;
  wire u2__abc_44228_n11880;
  wire u2__abc_44228_n11881;
  wire u2__abc_44228_n11882;
  wire u2__abc_44228_n11883_1;
  wire u2__abc_44228_n11884;
  wire u2__abc_44228_n11885;
  wire u2__abc_44228_n11887;
  wire u2__abc_44228_n11888;
  wire u2__abc_44228_n11889;
  wire u2__abc_44228_n11890;
  wire u2__abc_44228_n11891_1;
  wire u2__abc_44228_n11892;
  wire u2__abc_44228_n11893;
  wire u2__abc_44228_n11894;
  wire u2__abc_44228_n11895;
  wire u2__abc_44228_n11896;
  wire u2__abc_44228_n11897;
  wire u2__abc_44228_n11898_1;
  wire u2__abc_44228_n11899;
  wire u2__abc_44228_n11900;
  wire u2__abc_44228_n11901;
  wire u2__abc_44228_n11902;
  wire u2__abc_44228_n11903;
  wire u2__abc_44228_n11905;
  wire u2__abc_44228_n11906;
  wire u2__abc_44228_n11907_1;
  wire u2__abc_44228_n11908;
  wire u2__abc_44228_n11909;
  wire u2__abc_44228_n11910;
  wire u2__abc_44228_n11911;
  wire u2__abc_44228_n11912;
  wire u2__abc_44228_n11913;
  wire u2__abc_44228_n11914_1;
  wire u2__abc_44228_n11915;
  wire u2__abc_44228_n11916;
  wire u2__abc_44228_n11917;
  wire u2__abc_44228_n11918;
  wire u2__abc_44228_n11919;
  wire u2__abc_44228_n11920;
  wire u2__abc_44228_n11922_1;
  wire u2__abc_44228_n11923;
  wire u2__abc_44228_n11924;
  wire u2__abc_44228_n11925;
  wire u2__abc_44228_n11926;
  wire u2__abc_44228_n11927;
  wire u2__abc_44228_n11928;
  wire u2__abc_44228_n11929_1;
  wire u2__abc_44228_n11930;
  wire u2__abc_44228_n11931;
  wire u2__abc_44228_n11932;
  wire u2__abc_44228_n11933;
  wire u2__abc_44228_n11934;
  wire u2__abc_44228_n11935;
  wire u2__abc_44228_n11937;
  wire u2__abc_44228_n11938;
  wire u2__abc_44228_n11939;
  wire u2__abc_44228_n11940_1;
  wire u2__abc_44228_n11941;
  wire u2__abc_44228_n11942;
  wire u2__abc_44228_n11943;
  wire u2__abc_44228_n11944;
  wire u2__abc_44228_n11945;
  wire u2__abc_44228_n11946;
  wire u2__abc_44228_n11947_1;
  wire u2__abc_44228_n11948;
  wire u2__abc_44228_n11949;
  wire u2__abc_44228_n11950;
  wire u2__abc_44228_n11951;
  wire u2__abc_44228_n11952;
  wire u2__abc_44228_n11954;
  wire u2__abc_44228_n11955_1;
  wire u2__abc_44228_n11956;
  wire u2__abc_44228_n11957;
  wire u2__abc_44228_n11958;
  wire u2__abc_44228_n11959;
  wire u2__abc_44228_n11960;
  wire u2__abc_44228_n11961;
  wire u2__abc_44228_n11962_1;
  wire u2__abc_44228_n11963;
  wire u2__abc_44228_n11964;
  wire u2__abc_44228_n11965;
  wire u2__abc_44228_n11966;
  wire u2__abc_44228_n11967;
  wire u2__abc_44228_n11968;
  wire u2__abc_44228_n11969;
  wire u2__abc_44228_n11971_1;
  wire u2__abc_44228_n11972;
  wire u2__abc_44228_n11973;
  wire u2__abc_44228_n11974;
  wire u2__abc_44228_n11975;
  wire u2__abc_44228_n11976;
  wire u2__abc_44228_n11977;
  wire u2__abc_44228_n11978_1;
  wire u2__abc_44228_n11979;
  wire u2__abc_44228_n11980;
  wire u2__abc_44228_n11981;
  wire u2__abc_44228_n11982;
  wire u2__abc_44228_n11983;
  wire u2__abc_44228_n11984;
  wire u2__abc_44228_n11985;
  wire u2__abc_44228_n11986_1;
  wire u2__abc_44228_n11988;
  wire u2__abc_44228_n11989;
  wire u2__abc_44228_n11990;
  wire u2__abc_44228_n11991;
  wire u2__abc_44228_n11992;
  wire u2__abc_44228_n11993_1;
  wire u2__abc_44228_n11994;
  wire u2__abc_44228_n11995;
  wire u2__abc_44228_n11996;
  wire u2__abc_44228_n11997;
  wire u2__abc_44228_n11998;
  wire u2__abc_44228_n11999;
  wire u2__abc_44228_n12000;
  wire u2__abc_44228_n12001;
  wire u2__abc_44228_n12002;
  wire u2__abc_44228_n12003_1;
  wire u2__abc_44228_n12005;
  wire u2__abc_44228_n12006;
  wire u2__abc_44228_n12007;
  wire u2__abc_44228_n12008;
  wire u2__abc_44228_n12009;
  wire u2__abc_44228_n12010_1;
  wire u2__abc_44228_n12011;
  wire u2__abc_44228_n12012;
  wire u2__abc_44228_n12013;
  wire u2__abc_44228_n12014;
  wire u2__abc_44228_n12015;
  wire u2__abc_44228_n12016;
  wire u2__abc_44228_n12017;
  wire u2__abc_44228_n12018_1;
  wire u2__abc_44228_n12019;
  wire u2__abc_44228_n12020;
  wire u2__abc_44228_n12022;
  wire u2__abc_44228_n12023;
  wire u2__abc_44228_n12024;
  wire u2__abc_44228_n12025_1;
  wire u2__abc_44228_n12026;
  wire u2__abc_44228_n12027;
  wire u2__abc_44228_n12028;
  wire u2__abc_44228_n12029;
  wire u2__abc_44228_n12030;
  wire u2__abc_44228_n12031;
  wire u2__abc_44228_n12032;
  wire u2__abc_44228_n12033;
  wire u2__abc_44228_n12034_1;
  wire u2__abc_44228_n12035;
  wire u2__abc_44228_n12036;
  wire u2__abc_44228_n12037;
  wire u2__abc_44228_n12039;
  wire u2__abc_44228_n12040;
  wire u2__abc_44228_n12041_1;
  wire u2__abc_44228_n12042;
  wire u2__abc_44228_n12043;
  wire u2__abc_44228_n12044;
  wire u2__abc_44228_n12045;
  wire u2__abc_44228_n12046;
  wire u2__abc_44228_n12047;
  wire u2__abc_44228_n12048;
  wire u2__abc_44228_n12049_1;
  wire u2__abc_44228_n12050;
  wire u2__abc_44228_n12051;
  wire u2__abc_44228_n12052;
  wire u2__abc_44228_n12053;
  wire u2__abc_44228_n12054;
  wire u2__abc_44228_n12056_1;
  wire u2__abc_44228_n12057;
  wire u2__abc_44228_n12058;
  wire u2__abc_44228_n12059;
  wire u2__abc_44228_n12060;
  wire u2__abc_44228_n12061;
  wire u2__abc_44228_n12062;
  wire u2__abc_44228_n12063;
  wire u2__abc_44228_n12064;
  wire u2__abc_44228_n12065;
  wire u2__abc_44228_n12066;
  wire u2__abc_44228_n12067_1;
  wire u2__abc_44228_n12068;
  wire u2__abc_44228_n12069;
  wire u2__abc_44228_n12070;
  wire u2__abc_44228_n12071;
  wire u2__abc_44228_n12073;
  wire u2__abc_44228_n12074_1;
  wire u2__abc_44228_n12075;
  wire u2__abc_44228_n12076;
  wire u2__abc_44228_n12077;
  wire u2__abc_44228_n12078;
  wire u2__abc_44228_n12079;
  wire u2__abc_44228_n12080;
  wire u2__abc_44228_n12081;
  wire u2__abc_44228_n12082_1;
  wire u2__abc_44228_n12083;
  wire u2__abc_44228_n12084;
  wire u2__abc_44228_n12085;
  wire u2__abc_44228_n12086;
  wire u2__abc_44228_n12087;
  wire u2__abc_44228_n12088;
  wire u2__abc_44228_n12090;
  wire u2__abc_44228_n12091;
  wire u2__abc_44228_n12092;
  wire u2__abc_44228_n12093;
  wire u2__abc_44228_n12094;
  wire u2__abc_44228_n12095;
  wire u2__abc_44228_n12096;
  wire u2__abc_44228_n12097;
  wire u2__abc_44228_n12098_1;
  wire u2__abc_44228_n12099;
  wire u2__abc_44228_n12100;
  wire u2__abc_44228_n12101;
  wire u2__abc_44228_n12102;
  wire u2__abc_44228_n12103;
  wire u2__abc_44228_n12104;
  wire u2__abc_44228_n12105_1;
  wire u2__abc_44228_n12106;
  wire u2__abc_44228_n12108;
  wire u2__abc_44228_n12109;
  wire u2__abc_44228_n12110;
  wire u2__abc_44228_n12111;
  wire u2__abc_44228_n12112;
  wire u2__abc_44228_n12113_1;
  wire u2__abc_44228_n12114;
  wire u2__abc_44228_n12115;
  wire u2__abc_44228_n12116;
  wire u2__abc_44228_n12117;
  wire u2__abc_44228_n12118;
  wire u2__abc_44228_n12119;
  wire u2__abc_44228_n12120_1;
  wire u2__abc_44228_n12121;
  wire u2__abc_44228_n12122;
  wire u2__abc_44228_n12123;
  wire u2__abc_44228_n12125;
  wire u2__abc_44228_n12126;
  wire u2__abc_44228_n12127;
  wire u2__abc_44228_n12128;
  wire u2__abc_44228_n12129;
  wire u2__abc_44228_n12130_1;
  wire u2__abc_44228_n12131;
  wire u2__abc_44228_n12132;
  wire u2__abc_44228_n12133;
  wire u2__abc_44228_n12134;
  wire u2__abc_44228_n12135;
  wire u2__abc_44228_n12136;
  wire u2__abc_44228_n12137_1;
  wire u2__abc_44228_n12138;
  wire u2__abc_44228_n12139;
  wire u2__abc_44228_n12140;
  wire u2__abc_44228_n12142;
  wire u2__abc_44228_n12143;
  wire u2__abc_44228_n12144;
  wire u2__abc_44228_n12145_1;
  wire u2__abc_44228_n12146;
  wire u2__abc_44228_n12147;
  wire u2__abc_44228_n12148;
  wire u2__abc_44228_n12149;
  wire u2__abc_44228_n12150;
  wire u2__abc_44228_n12151;
  wire u2__abc_44228_n12152_1;
  wire u2__abc_44228_n12153;
  wire u2__abc_44228_n12154;
  wire u2__abc_44228_n12155;
  wire u2__abc_44228_n12156;
  wire u2__abc_44228_n12157;
  wire u2__abc_44228_n12159;
  wire u2__abc_44228_n12160;
  wire u2__abc_44228_n12161_1;
  wire u2__abc_44228_n12162;
  wire u2__abc_44228_n12163;
  wire u2__abc_44228_n12164;
  wire u2__abc_44228_n12165;
  wire u2__abc_44228_n12166;
  wire u2__abc_44228_n12167;
  wire u2__abc_44228_n12168_1;
  wire u2__abc_44228_n12169;
  wire u2__abc_44228_n12170;
  wire u2__abc_44228_n12171;
  wire u2__abc_44228_n12172;
  wire u2__abc_44228_n12173;
  wire u2__abc_44228_n12174;
  wire u2__abc_44228_n12176_1;
  wire u2__abc_44228_n12177;
  wire u2__abc_44228_n12178;
  wire u2__abc_44228_n12179;
  wire u2__abc_44228_n12180;
  wire u2__abc_44228_n12181;
  wire u2__abc_44228_n12182;
  wire u2__abc_44228_n12183_1;
  wire u2__abc_44228_n12184;
  wire u2__abc_44228_n12185;
  wire u2__abc_44228_n12186;
  wire u2__abc_44228_n12187;
  wire u2__abc_44228_n12188;
  wire u2__abc_44228_n12189;
  wire u2__abc_44228_n12190;
  wire u2__abc_44228_n12191;
  wire u2__abc_44228_n12193;
  wire u2__abc_44228_n12194;
  wire u2__abc_44228_n12195_1;
  wire u2__abc_44228_n12196;
  wire u2__abc_44228_n12197;
  wire u2__abc_44228_n12198;
  wire u2__abc_44228_n12199;
  wire u2__abc_44228_n12200;
  wire u2__abc_44228_n12201;
  wire u2__abc_44228_n12202_1;
  wire u2__abc_44228_n12203;
  wire u2__abc_44228_n12204;
  wire u2__abc_44228_n12205;
  wire u2__abc_44228_n12206;
  wire u2__abc_44228_n12207;
  wire u2__abc_44228_n12208;
  wire u2__abc_44228_n12210_1;
  wire u2__abc_44228_n12211;
  wire u2__abc_44228_n12212;
  wire u2__abc_44228_n12213;
  wire u2__abc_44228_n12214;
  wire u2__abc_44228_n12215;
  wire u2__abc_44228_n12216;
  wire u2__abc_44228_n12217_1;
  wire u2__abc_44228_n12218;
  wire u2__abc_44228_n12219;
  wire u2__abc_44228_n12220;
  wire u2__abc_44228_n12221;
  wire u2__abc_44228_n12222;
  wire u2__abc_44228_n12223;
  wire u2__abc_44228_n12224;
  wire u2__abc_44228_n12225;
  wire u2__abc_44228_n12227;
  wire u2__abc_44228_n12228;
  wire u2__abc_44228_n12229;
  wire u2__abc_44228_n12230;
  wire u2__abc_44228_n12231;
  wire u2__abc_44228_n12232;
  wire u2__abc_44228_n12233_1;
  wire u2__abc_44228_n12234;
  wire u2__abc_44228_n12235;
  wire u2__abc_44228_n12236;
  wire u2__abc_44228_n12237;
  wire u2__abc_44228_n12238;
  wire u2__abc_44228_n12239;
  wire u2__abc_44228_n12240;
  wire u2__abc_44228_n12241_1;
  wire u2__abc_44228_n12242;
  wire u2__abc_44228_n12243;
  wire u2__abc_44228_n12245;
  wire u2__abc_44228_n12246;
  wire u2__abc_44228_n12247;
  wire u2__abc_44228_n12248_1;
  wire u2__abc_44228_n12249;
  wire u2__abc_44228_n12250;
  wire u2__abc_44228_n12251;
  wire u2__abc_44228_n12252;
  wire u2__abc_44228_n12253;
  wire u2__abc_44228_n12254;
  wire u2__abc_44228_n12255;
  wire u2__abc_44228_n12256;
  wire u2__abc_44228_n12257;
  wire u2__abc_44228_n12258_1;
  wire u2__abc_44228_n12259;
  wire u2__abc_44228_n12260;
  wire u2__abc_44228_n12262;
  wire u2__abc_44228_n12263;
  wire u2__abc_44228_n12264;
  wire u2__abc_44228_n12265_1;
  wire u2__abc_44228_n12266;
  wire u2__abc_44228_n12267;
  wire u2__abc_44228_n12268;
  wire u2__abc_44228_n12269;
  wire u2__abc_44228_n12270;
  wire u2__abc_44228_n12271;
  wire u2__abc_44228_n12272;
  wire u2__abc_44228_n12273_1;
  wire u2__abc_44228_n12274;
  wire u2__abc_44228_n12275;
  wire u2__abc_44228_n12276;
  wire u2__abc_44228_n12277;
  wire u2__abc_44228_n12279;
  wire u2__abc_44228_n12280_1;
  wire u2__abc_44228_n12281;
  wire u2__abc_44228_n12282;
  wire u2__abc_44228_n12283;
  wire u2__abc_44228_n12284;
  wire u2__abc_44228_n12285;
  wire u2__abc_44228_n12286;
  wire u2__abc_44228_n12287;
  wire u2__abc_44228_n12288;
  wire u2__abc_44228_n12289_1;
  wire u2__abc_44228_n12290;
  wire u2__abc_44228_n12291;
  wire u2__abc_44228_n12292;
  wire u2__abc_44228_n12293;
  wire u2__abc_44228_n12294;
  wire u2__abc_44228_n12296_1;
  wire u2__abc_44228_n12297;
  wire u2__abc_44228_n12298;
  wire u2__abc_44228_n12299;
  wire u2__abc_44228_n12300;
  wire u2__abc_44228_n12301;
  wire u2__abc_44228_n12302;
  wire u2__abc_44228_n12303;
  wire u2__abc_44228_n12304_1;
  wire u2__abc_44228_n12305;
  wire u2__abc_44228_n12306;
  wire u2__abc_44228_n12307;
  wire u2__abc_44228_n12308;
  wire u2__abc_44228_n12309;
  wire u2__abc_44228_n12310;
  wire u2__abc_44228_n12311_1;
  wire u2__abc_44228_n12313;
  wire u2__abc_44228_n12314;
  wire u2__abc_44228_n12315;
  wire u2__abc_44228_n12316;
  wire u2__abc_44228_n12317;
  wire u2__abc_44228_n12318;
  wire u2__abc_44228_n12319;
  wire u2__abc_44228_n12320;
  wire u2__abc_44228_n12321;
  wire u2__abc_44228_n12322_1;
  wire u2__abc_44228_n12323;
  wire u2__abc_44228_n12324;
  wire u2__abc_44228_n12325;
  wire u2__abc_44228_n12326;
  wire u2__abc_44228_n12327;
  wire u2__abc_44228_n12328;
  wire u2__abc_44228_n12330;
  wire u2__abc_44228_n12331;
  wire u2__abc_44228_n12332;
  wire u2__abc_44228_n12333;
  wire u2__abc_44228_n12334;
  wire u2__abc_44228_n12335;
  wire u2__abc_44228_n12336;
  wire u2__abc_44228_n12337_1;
  wire u2__abc_44228_n12338;
  wire u2__abc_44228_n12339;
  wire u2__abc_44228_n12340;
  wire u2__abc_44228_n12341;
  wire u2__abc_44228_n12342;
  wire u2__abc_44228_n12343;
  wire u2__abc_44228_n12344_1;
  wire u2__abc_44228_n12345;
  wire u2__abc_44228_n12347;
  wire u2__abc_44228_n12348;
  wire u2__abc_44228_n12349;
  wire u2__abc_44228_n12350;
  wire u2__abc_44228_n12351;
  wire u2__abc_44228_n12352;
  wire u2__abc_44228_n12353_1;
  wire u2__abc_44228_n12354;
  wire u2__abc_44228_n12355;
  wire u2__abc_44228_n12356;
  wire u2__abc_44228_n12357;
  wire u2__abc_44228_n12358;
  wire u2__abc_44228_n12359;
  wire u2__abc_44228_n12360_1;
  wire u2__abc_44228_n12361;
  wire u2__abc_44228_n12362;
  wire u2__abc_44228_n12364;
  wire u2__abc_44228_n12365;
  wire u2__abc_44228_n12366;
  wire u2__abc_44228_n12367;
  wire u2__abc_44228_n12368_1;
  wire u2__abc_44228_n12369;
  wire u2__abc_44228_n12370;
  wire u2__abc_44228_n12371;
  wire u2__abc_44228_n12372;
  wire u2__abc_44228_n12373;
  wire u2__abc_44228_n12374;
  wire u2__abc_44228_n12375_1;
  wire u2__abc_44228_n12376;
  wire u2__abc_44228_n12377;
  wire u2__abc_44228_n12378;
  wire u2__abc_44228_n12379;
  wire u2__abc_44228_n12381;
  wire u2__abc_44228_n12382;
  wire u2__abc_44228_n12383;
  wire u2__abc_44228_n12384;
  wire u2__abc_44228_n12385_1;
  wire u2__abc_44228_n12386;
  wire u2__abc_44228_n12387;
  wire u2__abc_44228_n12388;
  wire u2__abc_44228_n12389;
  wire u2__abc_44228_n12390;
  wire u2__abc_44228_n12391;
  wire u2__abc_44228_n12392_1;
  wire u2__abc_44228_n12393;
  wire u2__abc_44228_n12394;
  wire u2__abc_44228_n12395;
  wire u2__abc_44228_n12396;
  wire u2__abc_44228_n12398;
  wire u2__abc_44228_n12399;
  wire u2__abc_44228_n12400_1;
  wire u2__abc_44228_n12401;
  wire u2__abc_44228_n12402;
  wire u2__abc_44228_n12403;
  wire u2__abc_44228_n12404;
  wire u2__abc_44228_n12405;
  wire u2__abc_44228_n12406;
  wire u2__abc_44228_n12407_1;
  wire u2__abc_44228_n12408;
  wire u2__abc_44228_n12409;
  wire u2__abc_44228_n12410;
  wire u2__abc_44228_n12411;
  wire u2__abc_44228_n12412;
  wire u2__abc_44228_n12413;
  wire u2__abc_44228_n12414;
  wire u2__abc_44228_n12416_1;
  wire u2__abc_44228_n12417;
  wire u2__abc_44228_n12418;
  wire u2__abc_44228_n12419;
  wire u2__abc_44228_n12420;
  wire u2__abc_44228_n12421;
  wire u2__abc_44228_n12422;
  wire u2__abc_44228_n12423_1;
  wire u2__abc_44228_n12424;
  wire u2__abc_44228_n12425;
  wire u2__abc_44228_n12426;
  wire u2__abc_44228_n12427;
  wire u2__abc_44228_n12428;
  wire u2__abc_44228_n12429;
  wire u2__abc_44228_n12430;
  wire u2__abc_44228_n12431_1;
  wire u2__abc_44228_n12433;
  wire u2__abc_44228_n12434;
  wire u2__abc_44228_n12435;
  wire u2__abc_44228_n12436;
  wire u2__abc_44228_n12437;
  wire u2__abc_44228_n12438_1;
  wire u2__abc_44228_n12439;
  wire u2__abc_44228_n12440;
  wire u2__abc_44228_n12441;
  wire u2__abc_44228_n12442;
  wire u2__abc_44228_n12443;
  wire u2__abc_44228_n12444;
  wire u2__abc_44228_n12445;
  wire u2__abc_44228_n12446;
  wire u2__abc_44228_n12447;
  wire u2__abc_44228_n12448;
  wire u2__abc_44228_n12449;
  wire u2__abc_44228_n12451;
  wire u2__abc_44228_n12452;
  wire u2__abc_44228_n12453;
  wire u2__abc_44228_n12454;
  wire u2__abc_44228_n12455;
  wire u2__abc_44228_n12456;
  wire u2__abc_44228_n12457_1;
  wire u2__abc_44228_n12458;
  wire u2__abc_44228_n12459;
  wire u2__abc_44228_n12460;
  wire u2__abc_44228_n12461;
  wire u2__abc_44228_n12462;
  wire u2__abc_44228_n12463;
  wire u2__abc_44228_n12464;
  wire u2__abc_44228_n12465_1;
  wire u2__abc_44228_n12466;
  wire u2__abc_44228_n12468;
  wire u2__abc_44228_n12469;
  wire u2__abc_44228_n12470;
  wire u2__abc_44228_n12471;
  wire u2__abc_44228_n12472_1;
  wire u2__abc_44228_n12473;
  wire u2__abc_44228_n12474;
  wire u2__abc_44228_n12475;
  wire u2__abc_44228_n12476;
  wire u2__abc_44228_n12477;
  wire u2__abc_44228_n12478;
  wire u2__abc_44228_n12479;
  wire u2__abc_44228_n12480;
  wire u2__abc_44228_n12481_1;
  wire u2__abc_44228_n12482;
  wire u2__abc_44228_n12483;
  wire u2__abc_44228_n12485;
  wire u2__abc_44228_n12486;
  wire u2__abc_44228_n12487;
  wire u2__abc_44228_n12488_1;
  wire u2__abc_44228_n12489;
  wire u2__abc_44228_n12490;
  wire u2__abc_44228_n12491;
  wire u2__abc_44228_n12492;
  wire u2__abc_44228_n12493;
  wire u2__abc_44228_n12494;
  wire u2__abc_44228_n12495;
  wire u2__abc_44228_n12496_1;
  wire u2__abc_44228_n12497;
  wire u2__abc_44228_n12498;
  wire u2__abc_44228_n12499;
  wire u2__abc_44228_n12500;
  wire u2__abc_44228_n12502;
  wire u2__abc_44228_n12503_1;
  wire u2__abc_44228_n12504;
  wire u2__abc_44228_n12505;
  wire u2__abc_44228_n12506;
  wire u2__abc_44228_n12507;
  wire u2__abc_44228_n12508;
  wire u2__abc_44228_n12509;
  wire u2__abc_44228_n12510;
  wire u2__abc_44228_n12511;
  wire u2__abc_44228_n12512;
  wire u2__abc_44228_n12513_1;
  wire u2__abc_44228_n12514;
  wire u2__abc_44228_n12515;
  wire u2__abc_44228_n12516;
  wire u2__abc_44228_n12517;
  wire u2__abc_44228_n12519;
  wire u2__abc_44228_n12520_1;
  wire u2__abc_44228_n12521;
  wire u2__abc_44228_n12522;
  wire u2__abc_44228_n12523;
  wire u2__abc_44228_n12524;
  wire u2__abc_44228_n12525;
  wire u2__abc_44228_n12526;
  wire u2__abc_44228_n12527;
  wire u2__abc_44228_n12528_1;
  wire u2__abc_44228_n12529;
  wire u2__abc_44228_n12530;
  wire u2__abc_44228_n12531;
  wire u2__abc_44228_n12532;
  wire u2__abc_44228_n12533;
  wire u2__abc_44228_n12534;
  wire u2__abc_44228_n12536;
  wire u2__abc_44228_n12537;
  wire u2__abc_44228_n12538;
  wire u2__abc_44228_n12539;
  wire u2__abc_44228_n12540;
  wire u2__abc_44228_n12541;
  wire u2__abc_44228_n12542;
  wire u2__abc_44228_n12543;
  wire u2__abc_44228_n12544_1;
  wire u2__abc_44228_n12545;
  wire u2__abc_44228_n12546;
  wire u2__abc_44228_n12547;
  wire u2__abc_44228_n12548;
  wire u2__abc_44228_n12549;
  wire u2__abc_44228_n12550;
  wire u2__abc_44228_n12551_1;
  wire u2__abc_44228_n12553;
  wire u2__abc_44228_n12554;
  wire u2__abc_44228_n12555;
  wire u2__abc_44228_n12556;
  wire u2__abc_44228_n12557;
  wire u2__abc_44228_n12558;
  wire u2__abc_44228_n12559_1;
  wire u2__abc_44228_n12560;
  wire u2__abc_44228_n12561;
  wire u2__abc_44228_n12562;
  wire u2__abc_44228_n12563;
  wire u2__abc_44228_n12564;
  wire u2__abc_44228_n12565;
  wire u2__abc_44228_n12566_1;
  wire u2__abc_44228_n12567;
  wire u2__abc_44228_n12568;
  wire u2__abc_44228_n12570;
  wire u2__abc_44228_n12571;
  wire u2__abc_44228_n12572;
  wire u2__abc_44228_n12573;
  wire u2__abc_44228_n12574;
  wire u2__abc_44228_n12575;
  wire u2__abc_44228_n12576;
  wire u2__abc_44228_n12577_1;
  wire u2__abc_44228_n12578;
  wire u2__abc_44228_n12579;
  wire u2__abc_44228_n12580;
  wire u2__abc_44228_n12581;
  wire u2__abc_44228_n12582;
  wire u2__abc_44228_n12583;
  wire u2__abc_44228_n12584_1;
  wire u2__abc_44228_n12585;
  wire u2__abc_44228_n12587;
  wire u2__abc_44228_n12588;
  wire u2__abc_44228_n12589;
  wire u2__abc_44228_n12590;
  wire u2__abc_44228_n12591;
  wire u2__abc_44228_n12592_1;
  wire u2__abc_44228_n12593;
  wire u2__abc_44228_n12594;
  wire u2__abc_44228_n12595;
  wire u2__abc_44228_n12596;
  wire u2__abc_44228_n12597;
  wire u2__abc_44228_n12598;
  wire u2__abc_44228_n12599_1;
  wire u2__abc_44228_n12600;
  wire u2__abc_44228_n12601;
  wire u2__abc_44228_n12602;
  wire u2__abc_44228_n12604;
  wire u2__abc_44228_n12605;
  wire u2__abc_44228_n12606;
  wire u2__abc_44228_n12607;
  wire u2__abc_44228_n12608_1;
  wire u2__abc_44228_n12609;
  wire u2__abc_44228_n12610;
  wire u2__abc_44228_n12611;
  wire u2__abc_44228_n12612;
  wire u2__abc_44228_n12613;
  wire u2__abc_44228_n12614;
  wire u2__abc_44228_n12615_1;
  wire u2__abc_44228_n12616;
  wire u2__abc_44228_n12617;
  wire u2__abc_44228_n12618;
  wire u2__abc_44228_n12619;
  wire u2__abc_44228_n12621;
  wire u2__abc_44228_n12622;
  wire u2__abc_44228_n12623_1;
  wire u2__abc_44228_n12624;
  wire u2__abc_44228_n12625;
  wire u2__abc_44228_n12626;
  wire u2__abc_44228_n12627;
  wire u2__abc_44228_n12628;
  wire u2__abc_44228_n12629;
  wire u2__abc_44228_n12630_1;
  wire u2__abc_44228_n12631;
  wire u2__abc_44228_n12632;
  wire u2__abc_44228_n12633;
  wire u2__abc_44228_n12634;
  wire u2__abc_44228_n12635;
  wire u2__abc_44228_n12636;
  wire u2__abc_44228_n12638;
  wire u2__abc_44228_n12639;
  wire u2__abc_44228_n12640_1;
  wire u2__abc_44228_n12641;
  wire u2__abc_44228_n12642;
  wire u2__abc_44228_n12643;
  wire u2__abc_44228_n12644;
  wire u2__abc_44228_n12645;
  wire u2__abc_44228_n12646;
  wire u2__abc_44228_n12647_1;
  wire u2__abc_44228_n12648;
  wire u2__abc_44228_n12649;
  wire u2__abc_44228_n12650;
  wire u2__abc_44228_n12651;
  wire u2__abc_44228_n12652;
  wire u2__abc_44228_n12653;
  wire u2__abc_44228_n12655_1;
  wire u2__abc_44228_n12656;
  wire u2__abc_44228_n12657;
  wire u2__abc_44228_n12658;
  wire u2__abc_44228_n12659;
  wire u2__abc_44228_n12660;
  wire u2__abc_44228_n12661;
  wire u2__abc_44228_n12662_1;
  wire u2__abc_44228_n12663;
  wire u2__abc_44228_n12664;
  wire u2__abc_44228_n12665;
  wire u2__abc_44228_n12666;
  wire u2__abc_44228_n12667;
  wire u2__abc_44228_n12668;
  wire u2__abc_44228_n12669;
  wire u2__abc_44228_n12670;
  wire u2__abc_44228_n12672;
  wire u2__abc_44228_n12673;
  wire u2__abc_44228_n12674;
  wire u2__abc_44228_n12675;
  wire u2__abc_44228_n12676;
  wire u2__abc_44228_n12677;
  wire u2__abc_44228_n12678_1;
  wire u2__abc_44228_n12679;
  wire u2__abc_44228_n12680;
  wire u2__abc_44228_n12681;
  wire u2__abc_44228_n12682;
  wire u2__abc_44228_n12683;
  wire u2__abc_44228_n12684;
  wire u2__abc_44228_n12685;
  wire u2__abc_44228_n12686_1;
  wire u2__abc_44228_n12687;
  wire u2__abc_44228_n12688;
  wire u2__abc_44228_n12690;
  wire u2__abc_44228_n12691;
  wire u2__abc_44228_n12692;
  wire u2__abc_44228_n12693_1;
  wire u2__abc_44228_n12694;
  wire u2__abc_44228_n12695;
  wire u2__abc_44228_n12696;
  wire u2__abc_44228_n12697;
  wire u2__abc_44228_n12698;
  wire u2__abc_44228_n12699;
  wire u2__abc_44228_n12700;
  wire u2__abc_44228_n12701;
  wire u2__abc_44228_n12702;
  wire u2__abc_44228_n12703;
  wire u2__abc_44228_n12704;
  wire u2__abc_44228_n12705;
  wire u2__abc_44228_n12707;
  wire u2__abc_44228_n12708;
  wire u2__abc_44228_n12709;
  wire u2__abc_44228_n12710;
  wire u2__abc_44228_n12711;
  wire u2__abc_44228_n12712;
  wire u2__abc_44228_n12713_1;
  wire u2__abc_44228_n12714;
  wire u2__abc_44228_n12715;
  wire u2__abc_44228_n12716;
  wire u2__abc_44228_n12717;
  wire u2__abc_44228_n12718;
  wire u2__abc_44228_n12719;
  wire u2__abc_44228_n12720;
  wire u2__abc_44228_n12721_1;
  wire u2__abc_44228_n12722;
  wire u2__abc_44228_n12723;
  wire u2__abc_44228_n12725;
  wire u2__abc_44228_n12726;
  wire u2__abc_44228_n12727;
  wire u2__abc_44228_n12728_1;
  wire u2__abc_44228_n12729;
  wire u2__abc_44228_n12730;
  wire u2__abc_44228_n12731;
  wire u2__abc_44228_n12732;
  wire u2__abc_44228_n12733;
  wire u2__abc_44228_n12734;
  wire u2__abc_44228_n12735;
  wire u2__abc_44228_n12736;
  wire u2__abc_44228_n12737_1;
  wire u2__abc_44228_n12738;
  wire u2__abc_44228_n12739;
  wire u2__abc_44228_n12740;
  wire u2__abc_44228_n12742;
  wire u2__abc_44228_n12743;
  wire u2__abc_44228_n12744_1;
  wire u2__abc_44228_n12745;
  wire u2__abc_44228_n12746;
  wire u2__abc_44228_n12747;
  wire u2__abc_44228_n12748;
  wire u2__abc_44228_n12749;
  wire u2__abc_44228_n12750;
  wire u2__abc_44228_n12751;
  wire u2__abc_44228_n12752_1;
  wire u2__abc_44228_n12753;
  wire u2__abc_44228_n12754;
  wire u2__abc_44228_n12755;
  wire u2__abc_44228_n12756;
  wire u2__abc_44228_n12757;
  wire u2__abc_44228_n12759_1;
  wire u2__abc_44228_n12760;
  wire u2__abc_44228_n12761;
  wire u2__abc_44228_n12762;
  wire u2__abc_44228_n12763;
  wire u2__abc_44228_n12764;
  wire u2__abc_44228_n12765;
  wire u2__abc_44228_n12766;
  wire u2__abc_44228_n12767;
  wire u2__abc_44228_n12768;
  wire u2__abc_44228_n12769_1;
  wire u2__abc_44228_n12770;
  wire u2__abc_44228_n12771;
  wire u2__abc_44228_n12772;
  wire u2__abc_44228_n12773;
  wire u2__abc_44228_n12774;
  wire u2__abc_44228_n12776_1;
  wire u2__abc_44228_n12777;
  wire u2__abc_44228_n12778;
  wire u2__abc_44228_n12779;
  wire u2__abc_44228_n12780;
  wire u2__abc_44228_n12781;
  wire u2__abc_44228_n12782;
  wire u2__abc_44228_n12783;
  wire u2__abc_44228_n12784_1;
  wire u2__abc_44228_n12785;
  wire u2__abc_44228_n12786;
  wire u2__abc_44228_n12787;
  wire u2__abc_44228_n12788;
  wire u2__abc_44228_n12789;
  wire u2__abc_44228_n12790;
  wire u2__abc_44228_n12791_1;
  wire u2__abc_44228_n12793;
  wire u2__abc_44228_n12794;
  wire u2__abc_44228_n12795;
  wire u2__abc_44228_n12796;
  wire u2__abc_44228_n12797;
  wire u2__abc_44228_n12798;
  wire u2__abc_44228_n12799;
  wire u2__abc_44228_n12800_1;
  wire u2__abc_44228_n12801;
  wire u2__abc_44228_n12802;
  wire u2__abc_44228_n12803;
  wire u2__abc_44228_n12804;
  wire u2__abc_44228_n12805;
  wire u2__abc_44228_n12806;
  wire u2__abc_44228_n12807_1;
  wire u2__abc_44228_n12808;
  wire u2__abc_44228_n12810;
  wire u2__abc_44228_n12811;
  wire u2__abc_44228_n12812;
  wire u2__abc_44228_n12813;
  wire u2__abc_44228_n12814;
  wire u2__abc_44228_n12815_1;
  wire u2__abc_44228_n12816;
  wire u2__abc_44228_n12817;
  wire u2__abc_44228_n12818;
  wire u2__abc_44228_n12819;
  wire u2__abc_44228_n12820;
  wire u2__abc_44228_n12821;
  wire u2__abc_44228_n12822_1;
  wire u2__abc_44228_n12823;
  wire u2__abc_44228_n12824;
  wire u2__abc_44228_n12825;
  wire u2__abc_44228_n12827;
  wire u2__abc_44228_n12828;
  wire u2__abc_44228_n12829;
  wire u2__abc_44228_n12830;
  wire u2__abc_44228_n12831;
  wire u2__abc_44228_n12832;
  wire u2__abc_44228_n12833_1;
  wire u2__abc_44228_n12834;
  wire u2__abc_44228_n12835;
  wire u2__abc_44228_n12836;
  wire u2__abc_44228_n12837;
  wire u2__abc_44228_n12838;
  wire u2__abc_44228_n12839;
  wire u2__abc_44228_n12840_1;
  wire u2__abc_44228_n12841;
  wire u2__abc_44228_n12842;
  wire u2__abc_44228_n12844;
  wire u2__abc_44228_n12845;
  wire u2__abc_44228_n12846;
  wire u2__abc_44228_n12847;
  wire u2__abc_44228_n12848_1;
  wire u2__abc_44228_n12849;
  wire u2__abc_44228_n12850;
  wire u2__abc_44228_n12851;
  wire u2__abc_44228_n12852;
  wire u2__abc_44228_n12853;
  wire u2__abc_44228_n12854;
  wire u2__abc_44228_n12855_1;
  wire u2__abc_44228_n12856;
  wire u2__abc_44228_n12857;
  wire u2__abc_44228_n12858;
  wire u2__abc_44228_n12859;
  wire u2__abc_44228_n12861;
  wire u2__abc_44228_n12862;
  wire u2__abc_44228_n12863;
  wire u2__abc_44228_n12864_1;
  wire u2__abc_44228_n12865;
  wire u2__abc_44228_n12866;
  wire u2__abc_44228_n12867;
  wire u2__abc_44228_n12868;
  wire u2__abc_44228_n12869;
  wire u2__abc_44228_n12870;
  wire u2__abc_44228_n12871_1;
  wire u2__abc_44228_n12872;
  wire u2__abc_44228_n12873;
  wire u2__abc_44228_n12874;
  wire u2__abc_44228_n12875;
  wire u2__abc_44228_n12876;
  wire u2__abc_44228_n12878;
  wire u2__abc_44228_n12879_1;
  wire u2__abc_44228_n12880;
  wire u2__abc_44228_n12881;
  wire u2__abc_44228_n12882;
  wire u2__abc_44228_n12883;
  wire u2__abc_44228_n12884;
  wire u2__abc_44228_n12885;
  wire u2__abc_44228_n12886_1;
  wire u2__abc_44228_n12887;
  wire u2__abc_44228_n12888;
  wire u2__abc_44228_n12889;
  wire u2__abc_44228_n12890;
  wire u2__abc_44228_n12891;
  wire u2__abc_44228_n12892;
  wire u2__abc_44228_n12893;
  wire u2__abc_44228_n12895;
  wire u2__abc_44228_n12896_1;
  wire u2__abc_44228_n12897;
  wire u2__abc_44228_n12898;
  wire u2__abc_44228_n12899;
  wire u2__abc_44228_n12900;
  wire u2__abc_44228_n12901;
  wire u2__abc_44228_n12902;
  wire u2__abc_44228_n12903_1;
  wire u2__abc_44228_n12904;
  wire u2__abc_44228_n12905;
  wire u2__abc_44228_n12906;
  wire u2__abc_44228_n12907;
  wire u2__abc_44228_n12908;
  wire u2__abc_44228_n12909;
  wire u2__abc_44228_n12910;
  wire u2__abc_44228_n12912;
  wire u2__abc_44228_n12913;
  wire u2__abc_44228_n12914;
  wire u2__abc_44228_n12915;
  wire u2__abc_44228_n12916;
  wire u2__abc_44228_n12917;
  wire u2__abc_44228_n12918_1;
  wire u2__abc_44228_n12919;
  wire u2__abc_44228_n12920;
  wire u2__abc_44228_n12921;
  wire u2__abc_44228_n12922;
  wire u2__abc_44228_n12923;
  wire u2__abc_44228_n12924;
  wire u2__abc_44228_n12925;
  wire u2__abc_44228_n12926;
  wire u2__abc_44228_n12927_1;
  wire u2__abc_44228_n12929;
  wire u2__abc_44228_n12930;
  wire u2__abc_44228_n12931;
  wire u2__abc_44228_n12932;
  wire u2__abc_44228_n12933;
  wire u2__abc_44228_n12934_1;
  wire u2__abc_44228_n12935;
  wire u2__abc_44228_n12936;
  wire u2__abc_44228_n12937;
  wire u2__abc_44228_n12938;
  wire u2__abc_44228_n12939;
  wire u2__abc_44228_n12940;
  wire u2__abc_44228_n12941;
  wire u2__abc_44228_n12942_1;
  wire u2__abc_44228_n12943;
  wire u2__abc_44228_n12944;
  wire u2__abc_44228_n12946;
  wire u2__abc_44228_n12947;
  wire u2__abc_44228_n12948;
  wire u2__abc_44228_n12949_1;
  wire u2__abc_44228_n12950;
  wire u2__abc_44228_n12951;
  wire u2__abc_44228_n12952;
  wire u2__abc_44228_n12953;
  wire u2__abc_44228_n12954;
  wire u2__abc_44228_n12955;
  wire u2__abc_44228_n12956;
  wire u2__abc_44228_n12957;
  wire u2__abc_44228_n12958;
  wire u2__abc_44228_n12959;
  wire u2__abc_44228_n12960;
  wire u2__abc_44228_n12961_1;
  wire u2__abc_44228_n12962;
  wire u2__abc_44228_n12964;
  wire u2__abc_44228_n12965;
  wire u2__abc_44228_n12966;
  wire u2__abc_44228_n12967;
  wire u2__abc_44228_n12968_1;
  wire u2__abc_44228_n12969;
  wire u2__abc_44228_n12970;
  wire u2__abc_44228_n12971;
  wire u2__abc_44228_n12972;
  wire u2__abc_44228_n12973;
  wire u2__abc_44228_n12974;
  wire u2__abc_44228_n12975;
  wire u2__abc_44228_n12976_1;
  wire u2__abc_44228_n12977;
  wire u2__abc_44228_n12978;
  wire u2__abc_44228_n12979;
  wire u2__abc_44228_n12981;
  wire u2__abc_44228_n12982;
  wire u2__abc_44228_n12983_1;
  wire u2__abc_44228_n12984;
  wire u2__abc_44228_n12985;
  wire u2__abc_44228_n12986;
  wire u2__abc_44228_n12987;
  wire u2__abc_44228_n12988;
  wire u2__abc_44228_n12989;
  wire u2__abc_44228_n12990;
  wire u2__abc_44228_n12991;
  wire u2__abc_44228_n12992_1;
  wire u2__abc_44228_n12993;
  wire u2__abc_44228_n12994;
  wire u2__abc_44228_n12995;
  wire u2__abc_44228_n12996;
  wire u2__abc_44228_n12998;
  wire u2__abc_44228_n12999_1;
  wire u2__abc_44228_n13000;
  wire u2__abc_44228_n13001;
  wire u2__abc_44228_n13002;
  wire u2__abc_44228_n13003;
  wire u2__abc_44228_n13004;
  wire u2__abc_44228_n13005;
  wire u2__abc_44228_n13006;
  wire u2__abc_44228_n13007_1;
  wire u2__abc_44228_n13008;
  wire u2__abc_44228_n13009;
  wire u2__abc_44228_n13010;
  wire u2__abc_44228_n13011;
  wire u2__abc_44228_n13012;
  wire u2__abc_44228_n13013;
  wire u2__abc_44228_n13015;
  wire u2__abc_44228_n13016;
  wire u2__abc_44228_n13017;
  wire u2__abc_44228_n13018;
  wire u2__abc_44228_n13019;
  wire u2__abc_44228_n13020;
  wire u2__abc_44228_n13021;
  wire u2__abc_44228_n13022;
  wire u2__abc_44228_n13023;
  wire u2__abc_44228_n13024_1;
  wire u2__abc_44228_n13025;
  wire u2__abc_44228_n13026;
  wire u2__abc_44228_n13027;
  wire u2__abc_44228_n13028;
  wire u2__abc_44228_n13029;
  wire u2__abc_44228_n13030;
  wire u2__abc_44228_n13032;
  wire u2__abc_44228_n13033;
  wire u2__abc_44228_n13034;
  wire u2__abc_44228_n13035;
  wire u2__abc_44228_n13036;
  wire u2__abc_44228_n13037;
  wire u2__abc_44228_n13038;
  wire u2__abc_44228_n13039_1;
  wire u2__abc_44228_n13040;
  wire u2__abc_44228_n13041;
  wire u2__abc_44228_n13042;
  wire u2__abc_44228_n13043;
  wire u2__abc_44228_n13044;
  wire u2__abc_44228_n13045;
  wire u2__abc_44228_n13046_1;
  wire u2__abc_44228_n13047;
  wire u2__abc_44228_n13049;
  wire u2__abc_44228_n13050;
  wire u2__abc_44228_n13051;
  wire u2__abc_44228_n13052;
  wire u2__abc_44228_n13053;
  wire u2__abc_44228_n13054;
  wire u2__abc_44228_n13055_1;
  wire u2__abc_44228_n13056;
  wire u2__abc_44228_n13057;
  wire u2__abc_44228_n13058;
  wire u2__abc_44228_n13059;
  wire u2__abc_44228_n13060;
  wire u2__abc_44228_n13061;
  wire u2__abc_44228_n13062_1;
  wire u2__abc_44228_n13063;
  wire u2__abc_44228_n13064;
  wire u2__abc_44228_n13065;
  wire u2__abc_44228_n13067;
  wire u2__abc_44228_n13068;
  wire u2__abc_44228_n13069;
  wire u2__abc_44228_n13070_1;
  wire u2__abc_44228_n13071;
  wire u2__abc_44228_n13072;
  wire u2__abc_44228_n13073;
  wire u2__abc_44228_n13074;
  wire u2__abc_44228_n13075;
  wire u2__abc_44228_n13076;
  wire u2__abc_44228_n13077_1;
  wire u2__abc_44228_n13078;
  wire u2__abc_44228_n13079;
  wire u2__abc_44228_n13080;
  wire u2__abc_44228_n13081;
  wire u2__abc_44228_n13082;
  wire u2__abc_44228_n13084;
  wire u2__abc_44228_n13085;
  wire u2__abc_44228_n13086;
  wire u2__abc_44228_n13087;
  wire u2__abc_44228_n13088_1;
  wire u2__abc_44228_n13089;
  wire u2__abc_44228_n13090;
  wire u2__abc_44228_n13091;
  wire u2__abc_44228_n13092;
  wire u2__abc_44228_n13093;
  wire u2__abc_44228_n13094;
  wire u2__abc_44228_n13095_1;
  wire u2__abc_44228_n13096;
  wire u2__abc_44228_n13097;
  wire u2__abc_44228_n13098;
  wire u2__abc_44228_n13099;
  wire u2__abc_44228_n13101;
  wire u2__abc_44228_n13102;
  wire u2__abc_44228_n13103_1;
  wire u2__abc_44228_n13104;
  wire u2__abc_44228_n13105;
  wire u2__abc_44228_n13106;
  wire u2__abc_44228_n13107;
  wire u2__abc_44228_n13108;
  wire u2__abc_44228_n13109;
  wire u2__abc_44228_n13110_1;
  wire u2__abc_44228_n13111;
  wire u2__abc_44228_n13112;
  wire u2__abc_44228_n13113;
  wire u2__abc_44228_n13114;
  wire u2__abc_44228_n13115;
  wire u2__abc_44228_n13116;
  wire u2__abc_44228_n13118;
  wire u2__abc_44228_n13119_1;
  wire u2__abc_44228_n13120;
  wire u2__abc_44228_n13121;
  wire u2__abc_44228_n13122;
  wire u2__abc_44228_n13123;
  wire u2__abc_44228_n13124;
  wire u2__abc_44228_n13125;
  wire u2__abc_44228_n13126_1;
  wire u2__abc_44228_n13127;
  wire u2__abc_44228_n13128;
  wire u2__abc_44228_n13129;
  wire u2__abc_44228_n13130;
  wire u2__abc_44228_n13131;
  wire u2__abc_44228_n13132;
  wire u2__abc_44228_n13133;
  wire u2__abc_44228_n13134_1;
  wire u2__abc_44228_n13136;
  wire u2__abc_44228_n13137;
  wire u2__abc_44228_n13138;
  wire u2__abc_44228_n13139;
  wire u2__abc_44228_n13140;
  wire u2__abc_44228_n13141_1;
  wire u2__abc_44228_n13142;
  wire u2__abc_44228_n13143;
  wire u2__abc_44228_n13144;
  wire u2__abc_44228_n13145;
  wire u2__abc_44228_n13146;
  wire u2__abc_44228_n13147;
  wire u2__abc_44228_n13148;
  wire u2__abc_44228_n13149;
  wire u2__abc_44228_n13150;
  wire u2__abc_44228_n13151_1;
  wire u2__abc_44228_n13153;
  wire u2__abc_44228_n13154;
  wire u2__abc_44228_n13155;
  wire u2__abc_44228_n13156;
  wire u2__abc_44228_n13157;
  wire u2__abc_44228_n13158_1;
  wire u2__abc_44228_n13159;
  wire u2__abc_44228_n13160;
  wire u2__abc_44228_n13161;
  wire u2__abc_44228_n13162;
  wire u2__abc_44228_n13163;
  wire u2__abc_44228_n13164;
  wire u2__abc_44228_n13165;
  wire u2__abc_44228_n13166_1;
  wire u2__abc_44228_n13167;
  wire u2__abc_44228_n13168;
  wire u2__abc_44228_n13170;
  wire u2__abc_44228_n13171;
  wire u2__abc_44228_n13172;
  wire u2__abc_44228_n13173_1;
  wire u2__abc_44228_n13174;
  wire u2__abc_44228_n13175;
  wire u2__abc_44228_n13176;
  wire u2__abc_44228_n13177;
  wire u2__abc_44228_n13178;
  wire u2__abc_44228_n13179;
  wire u2__abc_44228_n13180;
  wire u2__abc_44228_n13181;
  wire u2__abc_44228_n13182_1;
  wire u2__abc_44228_n13183;
  wire u2__abc_44228_n13184;
  wire u2__abc_44228_n13185;
  wire u2__abc_44228_n13187;
  wire u2__abc_44228_n13188;
  wire u2__abc_44228_n13189_1;
  wire u2__abc_44228_n13190;
  wire u2__abc_44228_n13191;
  wire u2__abc_44228_n13192;
  wire u2__abc_44228_n13193;
  wire u2__abc_44228_n13194;
  wire u2__abc_44228_n13195;
  wire u2__abc_44228_n13196;
  wire u2__abc_44228_n13197_1;
  wire u2__abc_44228_n13198;
  wire u2__abc_44228_n13199;
  wire u2__abc_44228_n13200;
  wire u2__abc_44228_n13201;
  wire u2__abc_44228_n13202;
  wire u2__abc_44228_n13203;
  wire u2__abc_44228_n13205;
  wire u2__abc_44228_n13206;
  wire u2__abc_44228_n13207;
  wire u2__abc_44228_n13208;
  wire u2__abc_44228_n13209;
  wire u2__abc_44228_n13210;
  wire u2__abc_44228_n13211;
  wire u2__abc_44228_n13212;
  wire u2__abc_44228_n13213;
  wire u2__abc_44228_n13214;
  wire u2__abc_44228_n13215;
  wire u2__abc_44228_n13216;
  wire u2__abc_44228_n13217_1;
  wire u2__abc_44228_n13218;
  wire u2__abc_44228_n13219;
  wire u2__abc_44228_n13220;
  wire u2__abc_44228_n13222;
  wire u2__abc_44228_n13223;
  wire u2__abc_44228_n13224_1;
  wire u2__abc_44228_n13225;
  wire u2__abc_44228_n13226;
  wire u2__abc_44228_n13227;
  wire u2__abc_44228_n13228;
  wire u2__abc_44228_n13229;
  wire u2__abc_44228_n13230;
  wire u2__abc_44228_n13231;
  wire u2__abc_44228_n13232_1;
  wire u2__abc_44228_n13233;
  wire u2__abc_44228_n13234;
  wire u2__abc_44228_n13235;
  wire u2__abc_44228_n13236;
  wire u2__abc_44228_n13237;
  wire u2__abc_44228_n13239_1;
  wire u2__abc_44228_n13240;
  wire u2__abc_44228_n13241;
  wire u2__abc_44228_n13242;
  wire u2__abc_44228_n13243;
  wire u2__abc_44228_n13244;
  wire u2__abc_44228_n13245;
  wire u2__abc_44228_n13246;
  wire u2__abc_44228_n13247;
  wire u2__abc_44228_n13248_1;
  wire u2__abc_44228_n13249;
  wire u2__abc_44228_n13250;
  wire u2__abc_44228_n13251;
  wire u2__abc_44228_n13252;
  wire u2__abc_44228_n13253;
  wire u2__abc_44228_n13254;
  wire u2__abc_44228_n13256;
  wire u2__abc_44228_n13257;
  wire u2__abc_44228_n13258;
  wire u2__abc_44228_n13259;
  wire u2__abc_44228_n13260;
  wire u2__abc_44228_n13261;
  wire u2__abc_44228_n13262;
  wire u2__abc_44228_n13263_1;
  wire u2__abc_44228_n13264;
  wire u2__abc_44228_n13265;
  wire u2__abc_44228_n13266;
  wire u2__abc_44228_n13267;
  wire u2__abc_44228_n13268;
  wire u2__abc_44228_n13269;
  wire u2__abc_44228_n13270_1;
  wire u2__abc_44228_n13271;
  wire u2__abc_44228_n13272;
  wire u2__abc_44228_n13274;
  wire u2__abc_44228_n13275;
  wire u2__abc_44228_n13276;
  wire u2__abc_44228_n13277;
  wire u2__abc_44228_n13278;
  wire u2__abc_44228_n13279;
  wire u2__abc_44228_n13280_1;
  wire u2__abc_44228_n13281;
  wire u2__abc_44228_n13282;
  wire u2__abc_44228_n13283;
  wire u2__abc_44228_n13284;
  wire u2__abc_44228_n13285;
  wire u2__abc_44228_n13286;
  wire u2__abc_44228_n13287_1;
  wire u2__abc_44228_n13288;
  wire u2__abc_44228_n13289;
  wire u2__abc_44228_n13291;
  wire u2__abc_44228_n13292;
  wire u2__abc_44228_n13293;
  wire u2__abc_44228_n13294;
  wire u2__abc_44228_n13295_1;
  wire u2__abc_44228_n13296;
  wire u2__abc_44228_n13297;
  wire u2__abc_44228_n13298;
  wire u2__abc_44228_n13299;
  wire u2__abc_44228_n13300;
  wire u2__abc_44228_n13301;
  wire u2__abc_44228_n13302_1;
  wire u2__abc_44228_n13303;
  wire u2__abc_44228_n13304;
  wire u2__abc_44228_n13305;
  wire u2__abc_44228_n13306;
  wire u2__abc_44228_n13308;
  wire u2__abc_44228_n13309;
  wire u2__abc_44228_n13310;
  wire u2__abc_44228_n13311_1;
  wire u2__abc_44228_n13312;
  wire u2__abc_44228_n13313;
  wire u2__abc_44228_n13314;
  wire u2__abc_44228_n13315;
  wire u2__abc_44228_n13316;
  wire u2__abc_44228_n13317;
  wire u2__abc_44228_n13318_1;
  wire u2__abc_44228_n13319;
  wire u2__abc_44228_n13320;
  wire u2__abc_44228_n13321;
  wire u2__abc_44228_n13322;
  wire u2__abc_44228_n13323;
  wire u2__abc_44228_n13325;
  wire u2__abc_44228_n13326_1;
  wire u2__abc_44228_n13327;
  wire u2__abc_44228_n13328;
  wire u2__abc_44228_n13329;
  wire u2__abc_44228_n13330;
  wire u2__abc_44228_n13331;
  wire u2__abc_44228_n13332;
  wire u2__abc_44228_n13333_1;
  wire u2__abc_44228_n13334;
  wire u2__abc_44228_n13335;
  wire u2__abc_44228_n13336;
  wire u2__abc_44228_n13337;
  wire u2__abc_44228_n13338;
  wire u2__abc_44228_n13339;
  wire u2__abc_44228_n13340;
  wire u2__abc_44228_n13342;
  wire u2__abc_44228_n13343;
  wire u2__abc_44228_n13344_1;
  wire u2__abc_44228_n13345;
  wire u2__abc_44228_n13346;
  wire u2__abc_44228_n13347;
  wire u2__abc_44228_n13348;
  wire u2__abc_44228_n13349;
  wire u2__abc_44228_n13350;
  wire u2__abc_44228_n13351_1;
  wire u2__abc_44228_n13352;
  wire u2__abc_44228_n13353;
  wire u2__abc_44228_n13354;
  wire u2__abc_44228_n13355;
  wire u2__abc_44228_n13356;
  wire u2__abc_44228_n13357;
  wire u2__abc_44228_n13359_1;
  wire u2__abc_44228_n13360;
  wire u2__abc_44228_n13361;
  wire u2__abc_44228_n13362;
  wire u2__abc_44228_n13363;
  wire u2__abc_44228_n13364;
  wire u2__abc_44228_n13365;
  wire u2__abc_44228_n13366_1;
  wire u2__abc_44228_n13367;
  wire u2__abc_44228_n13368;
  wire u2__abc_44228_n13369;
  wire u2__abc_44228_n13370;
  wire u2__abc_44228_n13371;
  wire u2__abc_44228_n13372;
  wire u2__abc_44228_n13373;
  wire u2__abc_44228_n13374;
  wire u2__abc_44228_n13376;
  wire u2__abc_44228_n13377;
  wire u2__abc_44228_n13378;
  wire u2__abc_44228_n13379;
  wire u2__abc_44228_n13380;
  wire u2__abc_44228_n13381;
  wire u2__abc_44228_n13382_1;
  wire u2__abc_44228_n13383;
  wire u2__abc_44228_n13384;
  wire u2__abc_44228_n13385;
  wire u2__abc_44228_n13386;
  wire u2__abc_44228_n13387;
  wire u2__abc_44228_n13388;
  wire u2__abc_44228_n13389;
  wire u2__abc_44228_n13390_1;
  wire u2__abc_44228_n13391;
  wire u2__abc_44228_n13393;
  wire u2__abc_44228_n13394;
  wire u2__abc_44228_n13395;
  wire u2__abc_44228_n13396;
  wire u2__abc_44228_n13397_1;
  wire u2__abc_44228_n13398;
  wire u2__abc_44228_n13399;
  wire u2__abc_44228_n13400;
  wire u2__abc_44228_n13401;
  wire u2__abc_44228_n13402;
  wire u2__abc_44228_n13403;
  wire u2__abc_44228_n13404;
  wire u2__abc_44228_n13405;
  wire u2__abc_44228_n13406;
  wire u2__abc_44228_n13407_1;
  wire u2__abc_44228_n13408;
  wire u2__abc_44228_n13409;
  wire u2__abc_44228_n13411;
  wire u2__abc_44228_n13412;
  wire u2__abc_44228_n13413;
  wire u2__abc_44228_n13414_1;
  wire u2__abc_44228_n13415;
  wire u2__abc_44228_n13416;
  wire u2__abc_44228_n13417;
  wire u2__abc_44228_n13418;
  wire u2__abc_44228_n13419;
  wire u2__abc_44228_n13420;
  wire u2__abc_44228_n13421;
  wire u2__abc_44228_n13422_1;
  wire u2__abc_44228_n13423;
  wire u2__abc_44228_n13424;
  wire u2__abc_44228_n13425;
  wire u2__abc_44228_n13426;
  wire u2__abc_44228_n13428;
  wire u2__abc_44228_n13429_1;
  wire u2__abc_44228_n13430;
  wire u2__abc_44228_n13431;
  wire u2__abc_44228_n13432;
  wire u2__abc_44228_n13433;
  wire u2__abc_44228_n13434;
  wire u2__abc_44228_n13435;
  wire u2__abc_44228_n13436;
  wire u2__abc_44228_n13437;
  wire u2__abc_44228_n13438_1;
  wire u2__abc_44228_n13439;
  wire u2__abc_44228_n13440;
  wire u2__abc_44228_n13441;
  wire u2__abc_44228_n13442;
  wire u2__abc_44228_n13443;
  wire u2__abc_44228_n13445_1;
  wire u2__abc_44228_n13446;
  wire u2__abc_44228_n13447;
  wire u2__abc_44228_n13448;
  wire u2__abc_44228_n13449;
  wire u2__abc_44228_n13450;
  wire u2__abc_44228_n13451;
  wire u2__abc_44228_n13452;
  wire u2__abc_44228_n13453_1;
  wire u2__abc_44228_n13454;
  wire u2__abc_44228_n13455;
  wire u2__abc_44228_n13456;
  wire u2__abc_44228_n13457;
  wire u2__abc_44228_n13458;
  wire u2__abc_44228_n13459;
  wire u2__abc_44228_n13460_1;
  wire u2__abc_44228_n13462;
  wire u2__abc_44228_n13463;
  wire u2__abc_44228_n13464;
  wire u2__abc_44228_n13465;
  wire u2__abc_44228_n13466;
  wire u2__abc_44228_n13467;
  wire u2__abc_44228_n13468;
  wire u2__abc_44228_n13469;
  wire u2__abc_44228_n13470;
  wire u2__abc_44228_n13471;
  wire u2__abc_44228_n13472_1;
  wire u2__abc_44228_n13473;
  wire u2__abc_44228_n13474;
  wire u2__abc_44228_n13475;
  wire u2__abc_44228_n13476;
  wire u2__abc_44228_n13477;
  wire u2__abc_44228_n13479_1;
  wire u2__abc_44228_n13480;
  wire u2__abc_44228_n13481;
  wire u2__abc_44228_n13482;
  wire u2__abc_44228_n13483;
  wire u2__abc_44228_n13484;
  wire u2__abc_44228_n13485;
  wire u2__abc_44228_n13486;
  wire u2__abc_44228_n13487_1;
  wire u2__abc_44228_n13488;
  wire u2__abc_44228_n13489;
  wire u2__abc_44228_n13490;
  wire u2__abc_44228_n13491;
  wire u2__abc_44228_n13492;
  wire u2__abc_44228_n13493;
  wire u2__abc_44228_n13494_1;
  wire u2__abc_44228_n13496;
  wire u2__abc_44228_n13497;
  wire u2__abc_44228_n13498;
  wire u2__abc_44228_n13499;
  wire u2__abc_44228_n13500;
  wire u2__abc_44228_n13501;
  wire u2__abc_44228_n13502;
  wire u2__abc_44228_n13503_1;
  wire u2__abc_44228_n13504;
  wire u2__abc_44228_n13505;
  wire u2__abc_44228_n13506;
  wire u2__abc_44228_n13507;
  wire u2__abc_44228_n13508;
  wire u2__abc_44228_n13509;
  wire u2__abc_44228_n13510_1;
  wire u2__abc_44228_n13511;
  wire u2__abc_44228_n13512;
  wire u2__abc_44228_n13514;
  wire u2__abc_44228_n13515;
  wire u2__abc_44228_n13516;
  wire u2__abc_44228_n13517;
  wire u2__abc_44228_n13518_1;
  wire u2__abc_44228_n13519;
  wire u2__abc_44228_n13520;
  wire u2__abc_44228_n13521;
  wire u2__abc_44228_n13522;
  wire u2__abc_44228_n13523;
  wire u2__abc_44228_n13524;
  wire u2__abc_44228_n13525_1;
  wire u2__abc_44228_n13526;
  wire u2__abc_44228_n13527;
  wire u2__abc_44228_n13528;
  wire u2__abc_44228_n13529;
  wire u2__abc_44228_n13531;
  wire u2__abc_44228_n13532;
  wire u2__abc_44228_n13533;
  wire u2__abc_44228_n13534;
  wire u2__abc_44228_n13535_1;
  wire u2__abc_44228_n13536;
  wire u2__abc_44228_n13537;
  wire u2__abc_44228_n13538;
  wire u2__abc_44228_n13539;
  wire u2__abc_44228_n13540;
  wire u2__abc_44228_n13541;
  wire u2__abc_44228_n13542_1;
  wire u2__abc_44228_n13543;
  wire u2__abc_44228_n13544;
  wire u2__abc_44228_n13545;
  wire u2__abc_44228_n13546;
  wire u2__abc_44228_n13547;
  wire u2__abc_44228_n13549;
  wire u2__abc_44228_n13550_1;
  wire u2__abc_44228_n13551;
  wire u2__abc_44228_n13552;
  wire u2__abc_44228_n13553;
  wire u2__abc_44228_n13554;
  wire u2__abc_44228_n13555;
  wire u2__abc_44228_n13556;
  wire u2__abc_44228_n13557_1;
  wire u2__abc_44228_n13558;
  wire u2__abc_44228_n13559;
  wire u2__abc_44228_n13560;
  wire u2__abc_44228_n13561;
  wire u2__abc_44228_n13562;
  wire u2__abc_44228_n13563;
  wire u2__abc_44228_n13564;
  wire u2__abc_44228_n13566_1;
  wire u2__abc_44228_n13567;
  wire u2__abc_44228_n13568;
  wire u2__abc_44228_n13569;
  wire u2__abc_44228_n13570;
  wire u2__abc_44228_n13571;
  wire u2__abc_44228_n13572;
  wire u2__abc_44228_n13573_1;
  wire u2__abc_44228_n13574;
  wire u2__abc_44228_n13575;
  wire u2__abc_44228_n13576;
  wire u2__abc_44228_n13577;
  wire u2__abc_44228_n13578;
  wire u2__abc_44228_n13579;
  wire u2__abc_44228_n13580;
  wire u2__abc_44228_n13581_1;
  wire u2__abc_44228_n13583;
  wire u2__abc_44228_n13584;
  wire u2__abc_44228_n13585;
  wire u2__abc_44228_n13586;
  wire u2__abc_44228_n13587;
  wire u2__abc_44228_n13588_1;
  wire u2__abc_44228_n13589;
  wire u2__abc_44228_n13590;
  wire u2__abc_44228_n13591;
  wire u2__abc_44228_n13592;
  wire u2__abc_44228_n13593;
  wire u2__abc_44228_n13594;
  wire u2__abc_44228_n13595;
  wire u2__abc_44228_n13596;
  wire u2__abc_44228_n13597;
  wire u2__abc_44228_n13598;
  wire u2__abc_44228_n13600;
  wire u2__abc_44228_n13601;
  wire u2__abc_44228_n13602;
  wire u2__abc_44228_n13603;
  wire u2__abc_44228_n13604;
  wire u2__abc_44228_n13605;
  wire u2__abc_44228_n13606_1;
  wire u2__abc_44228_n13607;
  wire u2__abc_44228_n13608;
  wire u2__abc_44228_n13609;
  wire u2__abc_44228_n13610;
  wire u2__abc_44228_n13611;
  wire u2__abc_44228_n13612;
  wire u2__abc_44228_n13613;
  wire u2__abc_44228_n13614_1;
  wire u2__abc_44228_n13615;
  wire u2__abc_44228_n13617;
  wire u2__abc_44228_n13618;
  wire u2__abc_44228_n13619;
  wire u2__abc_44228_n13620;
  wire u2__abc_44228_n13621_1;
  wire u2__abc_44228_n13622;
  wire u2__abc_44228_n13623;
  wire u2__abc_44228_n13624;
  wire u2__abc_44228_n13625;
  wire u2__abc_44228_n13626;
  wire u2__abc_44228_n13627;
  wire u2__abc_44228_n13628;
  wire u2__abc_44228_n13629;
  wire u2__abc_44228_n13630_1;
  wire u2__abc_44228_n13631;
  wire u2__abc_44228_n13632;
  wire u2__abc_44228_n13634;
  wire u2__abc_44228_n13635;
  wire u2__abc_44228_n13636;
  wire u2__abc_44228_n13637_1;
  wire u2__abc_44228_n13638;
  wire u2__abc_44228_n13639;
  wire u2__abc_44228_n13640;
  wire u2__abc_44228_n13641;
  wire u2__abc_44228_n13642;
  wire u2__abc_44228_n13643;
  wire u2__abc_44228_n13644;
  wire u2__abc_44228_n13645_1;
  wire u2__abc_44228_n13646;
  wire u2__abc_44228_n13647;
  wire u2__abc_44228_n13648;
  wire u2__abc_44228_n13649;
  wire u2__abc_44228_n13651;
  wire u2__abc_44228_n13652_1;
  wire u2__abc_44228_n13653;
  wire u2__abc_44228_n13654;
  wire u2__abc_44228_n13655;
  wire u2__abc_44228_n13656;
  wire u2__abc_44228_n13657;
  wire u2__abc_44228_n13658;
  wire u2__abc_44228_n13659;
  wire u2__abc_44228_n13660;
  wire u2__abc_44228_n13661;
  wire u2__abc_44228_n13662_1;
  wire u2__abc_44228_n13663;
  wire u2__abc_44228_n13664;
  wire u2__abc_44228_n13665;
  wire u2__abc_44228_n13666;
  wire u2__abc_44228_n13668;
  wire u2__abc_44228_n13669_1;
  wire u2__abc_44228_n13670;
  wire u2__abc_44228_n13671;
  wire u2__abc_44228_n13672;
  wire u2__abc_44228_n13673;
  wire u2__abc_44228_n13674;
  wire u2__abc_44228_n13675;
  wire u2__abc_44228_n13676;
  wire u2__abc_44228_n13677_1;
  wire u2__abc_44228_n13678;
  wire u2__abc_44228_n13679;
  wire u2__abc_44228_n13680;
  wire u2__abc_44228_n13681;
  wire u2__abc_44228_n13682;
  wire u2__abc_44228_n13683;
  wire u2__abc_44228_n13684_1;
  wire u2__abc_44228_n13686;
  wire u2__abc_44228_n13687;
  wire u2__abc_44228_n13688;
  wire u2__abc_44228_n13689;
  wire u2__abc_44228_n13690;
  wire u2__abc_44228_n13691;
  wire u2__abc_44228_n13692;
  wire u2__abc_44228_n13693_1;
  wire u2__abc_44228_n13694;
  wire u2__abc_44228_n13695;
  wire u2__abc_44228_n13696;
  wire u2__abc_44228_n13697;
  wire u2__abc_44228_n13698;
  wire u2__abc_44228_n13699;
  wire u2__abc_44228_n13700_1;
  wire u2__abc_44228_n13701;
  wire u2__abc_44228_n13703;
  wire u2__abc_44228_n13704;
  wire u2__abc_44228_n13705;
  wire u2__abc_44228_n13706;
  wire u2__abc_44228_n13707;
  wire u2__abc_44228_n13708;
  wire u2__abc_44228_n13709_1;
  wire u2__abc_44228_n13710;
  wire u2__abc_44228_n13711;
  wire u2__abc_44228_n13712;
  wire u2__abc_44228_n13713;
  wire u2__abc_44228_n13714;
  wire u2__abc_44228_n13715;
  wire u2__abc_44228_n13716;
  wire u2__abc_44228_n13717_1;
  wire u2__abc_44228_n13718;
  wire u2__abc_44228_n13720;
  wire u2__abc_44228_n13721;
  wire u2__abc_44228_n13722;
  wire u2__abc_44228_n13723;
  wire u2__abc_44228_n13724;
  wire u2__abc_44228_n13725;
  wire u2__abc_44228_n13726;
  wire u2__abc_44228_n13727;
  wire u2__abc_44228_n13728;
  wire u2__abc_44228_n13729;
  wire u2__abc_44228_n13730;
  wire u2__abc_44228_n13731;
  wire u2__abc_44228_n13732_1;
  wire u2__abc_44228_n13733;
  wire u2__abc_44228_n13734;
  wire u2__abc_44228_n13735;
  wire u2__abc_44228_n13737;
  wire u2__abc_44228_n13738;
  wire u2__abc_44228_n13739;
  wire u2__abc_44228_n13740_1;
  wire u2__abc_44228_n13741;
  wire u2__abc_44228_n13742;
  wire u2__abc_44228_n13743;
  wire u2__abc_44228_n13744;
  wire u2__abc_44228_n13745;
  wire u2__abc_44228_n13746;
  wire u2__abc_44228_n13747;
  wire u2__abc_44228_n13748;
  wire u2__abc_44228_n13749_1;
  wire u2__abc_44228_n13750;
  wire u2__abc_44228_n13751;
  wire u2__abc_44228_n13752;
  wire u2__abc_44228_n13754;
  wire u2__abc_44228_n13755;
  wire u2__abc_44228_n13756;
  wire u2__abc_44228_n13757_1;
  wire u2__abc_44228_n13758;
  wire u2__abc_44228_n13759;
  wire u2__abc_44228_n13760;
  wire u2__abc_44228_n13761;
  wire u2__abc_44228_n13762;
  wire u2__abc_44228_n13763;
  wire u2__abc_44228_n13764;
  wire u2__abc_44228_n13765;
  wire u2__abc_44228_n13766;
  wire u2__abc_44228_n13767_1;
  wire u2__abc_44228_n13768;
  wire u2__abc_44228_n13769;
  wire u2__abc_44228_n13771;
  wire u2__abc_44228_n13772;
  wire u2__abc_44228_n13773;
  wire u2__abc_44228_n13774;
  wire u2__abc_44228_n13775_1;
  wire u2__abc_44228_n13776;
  wire u2__abc_44228_n13777;
  wire u2__abc_44228_n13778;
  wire u2__abc_44228_n13779;
  wire u2__abc_44228_n13780;
  wire u2__abc_44228_n13781;
  wire u2__abc_44228_n13782;
  wire u2__abc_44228_n13783;
  wire u2__abc_44228_n13784_1;
  wire u2__abc_44228_n13785;
  wire u2__abc_44228_n13786;
  wire u2__abc_44228_n13787;
  wire u2__abc_44228_n13789;
  wire u2__abc_44228_n13790;
  wire u2__abc_44228_n13791;
  wire u2__abc_44228_n13792_1;
  wire u2__abc_44228_n13793;
  wire u2__abc_44228_n13794;
  wire u2__abc_44228_n13795;
  wire u2__abc_44228_n13796;
  wire u2__abc_44228_n13797;
  wire u2__abc_44228_n13798;
  wire u2__abc_44228_n13799;
  wire u2__abc_44228_n13800;
  wire u2__abc_44228_n13801;
  wire u2__abc_44228_n13802;
  wire u2__abc_44228_n13803_1;
  wire u2__abc_44228_n13804;
  wire u2__abc_44228_n13806;
  wire u2__abc_44228_n13807;
  wire u2__abc_44228_n13808;
  wire u2__abc_44228_n13809;
  wire u2__abc_44228_n13810;
  wire u2__abc_44228_n13811_1;
  wire u2__abc_44228_n13812;
  wire u2__abc_44228_n13813;
  wire u2__abc_44228_n13814;
  wire u2__abc_44228_n13815;
  wire u2__abc_44228_n13816;
  wire u2__abc_44228_n13817;
  wire u2__abc_44228_n13818;
  wire u2__abc_44228_n13819;
  wire u2__abc_44228_n13820_1;
  wire u2__abc_44228_n13821;
  wire u2__abc_44228_n13823;
  wire u2__abc_44228_n13824;
  wire u2__abc_44228_n13825;
  wire u2__abc_44228_n13826;
  wire u2__abc_44228_n13827;
  wire u2__abc_44228_n13828_1;
  wire u2__abc_44228_n13829;
  wire u2__abc_44228_n13830;
  wire u2__abc_44228_n13831;
  wire u2__abc_44228_n13832;
  wire u2__abc_44228_n13833;
  wire u2__abc_44228_n13834;
  wire u2__abc_44228_n13835;
  wire u2__abc_44228_n13836;
  wire u2__abc_44228_n13837;
  wire u2__abc_44228_n13838_1;
  wire u2__abc_44228_n13840;
  wire u2__abc_44228_n13841;
  wire u2__abc_44228_n13842;
  wire u2__abc_44228_n13843;
  wire u2__abc_44228_n13844;
  wire u2__abc_44228_n13845;
  wire u2__abc_44228_n13846_1;
  wire u2__abc_44228_n13847;
  wire u2__abc_44228_n13848;
  wire u2__abc_44228_n13849;
  wire u2__abc_44228_n13850;
  wire u2__abc_44228_n13851;
  wire u2__abc_44228_n13852;
  wire u2__abc_44228_n13853;
  wire u2__abc_44228_n13854;
  wire u2__abc_44228_n13855_1;
  wire u2__abc_44228_n13857;
  wire u2__abc_44228_n13858;
  wire u2__abc_44228_n13859;
  wire u2__abc_44228_n13860;
  wire u2__abc_44228_n13861;
  wire u2__abc_44228_n13862;
  wire u2__abc_44228_n13863_1;
  wire u2__abc_44228_n13864;
  wire u2__abc_44228_n13865;
  wire u2__abc_44228_n13866;
  wire u2__abc_44228_n13867;
  wire u2__abc_44228_n13868;
  wire u2__abc_44228_n13869;
  wire u2__abc_44228_n13870;
  wire u2__abc_44228_n13871;
  wire u2__abc_44228_n13872;
  wire u2__abc_44228_n13874;
  wire u2__abc_44228_n13875_1;
  wire u2__abc_44228_n13876;
  wire u2__abc_44228_n13877;
  wire u2__abc_44228_n13878;
  wire u2__abc_44228_n13879;
  wire u2__abc_44228_n13880;
  wire u2__abc_44228_n13881;
  wire u2__abc_44228_n13882;
  wire u2__abc_44228_n13883_1;
  wire u2__abc_44228_n13884;
  wire u2__abc_44228_n13885;
  wire u2__abc_44228_n13886;
  wire u2__abc_44228_n13887;
  wire u2__abc_44228_n13888;
  wire u2__abc_44228_n13889;
  wire u2__abc_44228_n13891;
  wire u2__abc_44228_n13892_1;
  wire u2__abc_44228_n13893;
  wire u2__abc_44228_n13894;
  wire u2__abc_44228_n13895;
  wire u2__abc_44228_n13896;
  wire u2__abc_44228_n13897;
  wire u2__abc_44228_n13898;
  wire u2__abc_44228_n13899;
  wire u2__abc_44228_n13900_1;
  wire u2__abc_44228_n13901;
  wire u2__abc_44228_n13902;
  wire u2__abc_44228_n13903;
  wire u2__abc_44228_n13904;
  wire u2__abc_44228_n13905;
  wire u2__abc_44228_n13906;
  wire u2__abc_44228_n13908;
  wire u2__abc_44228_n13909;
  wire u2__abc_44228_n13910_1;
  wire u2__abc_44228_n13911;
  wire u2__abc_44228_n13912;
  wire u2__abc_44228_n13913;
  wire u2__abc_44228_n13914;
  wire u2__abc_44228_n13915;
  wire u2__abc_44228_n13916;
  wire u2__abc_44228_n13917;
  wire u2__abc_44228_n13918_1;
  wire u2__abc_44228_n13919;
  wire u2__abc_44228_n13920;
  wire u2__abc_44228_n13921;
  wire u2__abc_44228_n13922;
  wire u2__abc_44228_n13923;
  wire u2__abc_44228_n13924;
  wire u2__abc_44228_n13926;
  wire u2__abc_44228_n13927_1;
  wire u2__abc_44228_n13928;
  wire u2__abc_44228_n13929;
  wire u2__abc_44228_n13930;
  wire u2__abc_44228_n13931;
  wire u2__abc_44228_n13932;
  wire u2__abc_44228_n13933;
  wire u2__abc_44228_n13934;
  wire u2__abc_44228_n13935_1;
  wire u2__abc_44228_n13936;
  wire u2__abc_44228_n13937;
  wire u2__abc_44228_n13938;
  wire u2__abc_44228_n13939;
  wire u2__abc_44228_n13940;
  wire u2__abc_44228_n13941;
  wire u2__abc_44228_n13943;
  wire u2__abc_44228_n13944;
  wire u2__abc_44228_n13945;
  wire u2__abc_44228_n13946_1;
  wire u2__abc_44228_n13947;
  wire u2__abc_44228_n13948;
  wire u2__abc_44228_n13949;
  wire u2__abc_44228_n13950;
  wire u2__abc_44228_n13951;
  wire u2__abc_44228_n13952;
  wire u2__abc_44228_n13953;
  wire u2__abc_44228_n13954_1;
  wire u2__abc_44228_n13955;
  wire u2__abc_44228_n13956;
  wire u2__abc_44228_n13957;
  wire u2__abc_44228_n13958;
  wire u2__abc_44228_n13959;
  wire u2__abc_44228_n13961;
  wire u2__abc_44228_n13962;
  wire u2__abc_44228_n13963_1;
  wire u2__abc_44228_n13964;
  wire u2__abc_44228_n13965;
  wire u2__abc_44228_n13966;
  wire u2__abc_44228_n13967;
  wire u2__abc_44228_n13968;
  wire u2__abc_44228_n13969;
  wire u2__abc_44228_n13970;
  wire u2__abc_44228_n13971_1;
  wire u2__abc_44228_n13972;
  wire u2__abc_44228_n13973;
  wire u2__abc_44228_n13974;
  wire u2__abc_44228_n13975;
  wire u2__abc_44228_n13976;
  wire u2__abc_44228_n13978;
  wire u2__abc_44228_n13979;
  wire u2__abc_44228_n13980;
  wire u2__abc_44228_n13981_1;
  wire u2__abc_44228_n13982;
  wire u2__abc_44228_n13983;
  wire u2__abc_44228_n13984;
  wire u2__abc_44228_n13985;
  wire u2__abc_44228_n13986;
  wire u2__abc_44228_n13987;
  wire u2__abc_44228_n13988;
  wire u2__abc_44228_n13989_1;
  wire u2__abc_44228_n13990;
  wire u2__abc_44228_n13991;
  wire u2__abc_44228_n13992;
  wire u2__abc_44228_n13993;
  wire u2__abc_44228_n13995;
  wire u2__abc_44228_n13996;
  wire u2__abc_44228_n13997;
  wire u2__abc_44228_n13998_1;
  wire u2__abc_44228_n13999;
  wire u2__abc_44228_n14000;
  wire u2__abc_44228_n14001;
  wire u2__abc_44228_n14002;
  wire u2__abc_44228_n14003;
  wire u2__abc_44228_n14004;
  wire u2__abc_44228_n14005;
  wire u2__abc_44228_n14006_1;
  wire u2__abc_44228_n14007;
  wire u2__abc_44228_n14008;
  wire u2__abc_44228_n14009;
  wire u2__abc_44228_n14010;
  wire u2__abc_44228_n14012;
  wire u2__abc_44228_n14013;
  wire u2__abc_44228_n14014;
  wire u2__abc_44228_n14015;
  wire u2__abc_44228_n14016;
  wire u2__abc_44228_n14017;
  wire u2__abc_44228_n14018;
  wire u2__abc_44228_n14019_1;
  wire u2__abc_44228_n14020;
  wire u2__abc_44228_n14021;
  wire u2__abc_44228_n14022;
  wire u2__abc_44228_n14023;
  wire u2__abc_44228_n14024;
  wire u2__abc_44228_n14025;
  wire u2__abc_44228_n14026;
  wire u2__abc_44228_n14027_1;
  wire u2__abc_44228_n14029;
  wire u2__abc_44228_n14030;
  wire u2__abc_44228_n14031;
  wire u2__abc_44228_n14032;
  wire u2__abc_44228_n14033;
  wire u2__abc_44228_n14034;
  wire u2__abc_44228_n14035;
  wire u2__abc_44228_n14036_1;
  wire u2__abc_44228_n14037;
  wire u2__abc_44228_n14038;
  wire u2__abc_44228_n14039;
  wire u2__abc_44228_n14040;
  wire u2__abc_44228_n14041;
  wire u2__abc_44228_n14042;
  wire u2__abc_44228_n14043;
  wire u2__abc_44228_n14044_1;
  wire u2__abc_44228_n14046;
  wire u2__abc_44228_n14047;
  wire u2__abc_44228_n14048;
  wire u2__abc_44228_n14049;
  wire u2__abc_44228_n14050;
  wire u2__abc_44228_n14051;
  wire u2__abc_44228_n14052;
  wire u2__abc_44228_n14053;
  wire u2__abc_44228_n14054_1;
  wire u2__abc_44228_n14055;
  wire u2__abc_44228_n14056;
  wire u2__abc_44228_n14057;
  wire u2__abc_44228_n14058;
  wire u2__abc_44228_n14059;
  wire u2__abc_44228_n14060;
  wire u2__abc_44228_n14061;
  wire u2__abc_44228_n14062_1;
  wire u2__abc_44228_n14064;
  wire u2__abc_44228_n14065;
  wire u2__abc_44228_n14066;
  wire u2__abc_44228_n14067;
  wire u2__abc_44228_n14068;
  wire u2__abc_44228_n14069;
  wire u2__abc_44228_n14070;
  wire u2__abc_44228_n14071_1;
  wire u2__abc_44228_n14072;
  wire u2__abc_44228_n14073;
  wire u2__abc_44228_n14074;
  wire u2__abc_44228_n14075;
  wire u2__abc_44228_n14076;
  wire u2__abc_44228_n14077;
  wire u2__abc_44228_n14078;
  wire u2__abc_44228_n14079_1;
  wire u2__abc_44228_n14081;
  wire u2__abc_44228_n14082;
  wire u2__abc_44228_n14083;
  wire u2__abc_44228_n14084;
  wire u2__abc_44228_n14085;
  wire u2__abc_44228_n14086;
  wire u2__abc_44228_n14087;
  wire u2__abc_44228_n14088;
  wire u2__abc_44228_n14089;
  wire u2__abc_44228_n14090_1;
  wire u2__abc_44228_n14091;
  wire u2__abc_44228_n14092;
  wire u2__abc_44228_n14093;
  wire u2__abc_44228_n14094;
  wire u2__abc_44228_n14095;
  wire u2__abc_44228_n14096;
  wire u2__abc_44228_n14097;
  wire u2__abc_44228_n14099;
  wire u2__abc_44228_n14100;
  wire u2__abc_44228_n14101;
  wire u2__abc_44228_n14102;
  wire u2__abc_44228_n14103;
  wire u2__abc_44228_n14104;
  wire u2__abc_44228_n14105;
  wire u2__abc_44228_n14106;
  wire u2__abc_44228_n14107_1;
  wire u2__abc_44228_n14108;
  wire u2__abc_44228_n14109;
  wire u2__abc_44228_n14110;
  wire u2__abc_44228_n14111;
  wire u2__abc_44228_n14112;
  wire u2__abc_44228_n14113;
  wire u2__abc_44228_n14114;
  wire u2__abc_44228_n14116;
  wire u2__abc_44228_n14117;
  wire u2__abc_44228_n14118;
  wire u2__abc_44228_n14119;
  wire u2__abc_44228_n14120;
  wire u2__abc_44228_n14121;
  wire u2__abc_44228_n14122;
  wire u2__abc_44228_n14123;
  wire u2__abc_44228_n14124;
  wire u2__abc_44228_n14125_1;
  wire u2__abc_44228_n14126;
  wire u2__abc_44228_n14127;
  wire u2__abc_44228_n14128;
  wire u2__abc_44228_n14129;
  wire u2__abc_44228_n14131;
  wire u2__abc_44228_n14132;
  wire u2__abc_44228_n14133_1;
  wire u2__abc_44228_n14134;
  wire u2__abc_44228_n14135;
  wire u2__abc_44228_n14136;
  wire u2__abc_44228_n14137;
  wire u2__abc_44228_n14138;
  wire u2__abc_44228_n14139;
  wire u2__abc_44228_n14140;
  wire u2__abc_44228_n14141;
  wire u2__abc_44228_n14142_1;
  wire u2__abc_44228_n14143;
  wire u2__abc_44228_n14144;
  wire u2__abc_44228_n14145;
  wire u2__abc_44228_n14146;
  wire u2__abc_44228_n14148;
  wire u2__abc_44228_n14149;
  wire u2__abc_44228_n14150_1;
  wire u2__abc_44228_n14151;
  wire u2__abc_44228_n14152;
  wire u2__abc_44228_n14153;
  wire u2__abc_44228_n14154;
  wire u2__abc_44228_n14155;
  wire u2__abc_44228_n14156;
  wire u2__abc_44228_n14157;
  wire u2__abc_44228_n14158;
  wire u2__abc_44228_n14159;
  wire u2__abc_44228_n14160;
  wire u2__abc_44228_n14161;
  wire u2__abc_44228_n14162_1;
  wire u2__abc_44228_n14163;
  wire u2__abc_44228_n14165;
  wire u2__abc_44228_n14166;
  wire u2__abc_44228_n14167;
  wire u2__abc_44228_n14168;
  wire u2__abc_44228_n14169;
  wire u2__abc_44228_n14170_1;
  wire u2__abc_44228_n14171;
  wire u2__abc_44228_n14172;
  wire u2__abc_44228_n14173;
  wire u2__abc_44228_n14174;
  wire u2__abc_44228_n14175;
  wire u2__abc_44228_n14176;
  wire u2__abc_44228_n14177;
  wire u2__abc_44228_n14178;
  wire u2__abc_44228_n14179_1;
  wire u2__abc_44228_n14180;
  wire u2__abc_44228_n14182;
  wire u2__abc_44228_n14183;
  wire u2__abc_44228_n14184;
  wire u2__abc_44228_n14185;
  wire u2__abc_44228_n14186;
  wire u2__abc_44228_n14187_1;
  wire u2__abc_44228_n14188;
  wire u2__abc_44228_n14189;
  wire u2__abc_44228_n14190;
  wire u2__abc_44228_n14191;
  wire u2__abc_44228_n14192;
  wire u2__abc_44228_n14193;
  wire u2__abc_44228_n14194;
  wire u2__abc_44228_n14195;
  wire u2__abc_44228_n14196;
  wire u2__abc_44228_n14197_1;
  wire u2__abc_44228_n14199;
  wire u2__abc_44228_n14200;
  wire u2__abc_44228_n14201;
  wire u2__abc_44228_n14202;
  wire u2__abc_44228_n14203;
  wire u2__abc_44228_n14204;
  wire u2__abc_44228_n14205_1;
  wire u2__abc_44228_n14206;
  wire u2__abc_44228_n14207;
  wire u2__abc_44228_n14208;
  wire u2__abc_44228_n14209;
  wire u2__abc_44228_n14210;
  wire u2__abc_44228_n14211;
  wire u2__abc_44228_n14212;
  wire u2__abc_44228_n14213;
  wire u2__abc_44228_n14214_1;
  wire u2__abc_44228_n14216;
  wire u2__abc_44228_n14217;
  wire u2__abc_44228_n14218;
  wire u2__abc_44228_n14219;
  wire u2__abc_44228_n14220;
  wire u2__abc_44228_n14221;
  wire u2__abc_44228_n14222_1;
  wire u2__abc_44228_n14223;
  wire u2__abc_44228_n14224;
  wire u2__abc_44228_n14225;
  wire u2__abc_44228_n14226;
  wire u2__abc_44228_n14227;
  wire u2__abc_44228_n14228;
  wire u2__abc_44228_n14229;
  wire u2__abc_44228_n14230;
  wire u2__abc_44228_n14231;
  wire u2__abc_44228_n14232;
  wire u2__abc_44228_n14234;
  wire u2__abc_44228_n14235;
  wire u2__abc_44228_n14236;
  wire u2__abc_44228_n14237;
  wire u2__abc_44228_n14238;
  wire u2__abc_44228_n14239;
  wire u2__abc_44228_n14240;
  wire u2__abc_44228_n14241_1;
  wire u2__abc_44228_n14242;
  wire u2__abc_44228_n14243;
  wire u2__abc_44228_n14244;
  wire u2__abc_44228_n14245;
  wire u2__abc_44228_n14246;
  wire u2__abc_44228_n14247;
  wire u2__abc_44228_n14248;
  wire u2__abc_44228_n14249;
  wire u2__abc_44228_n14251;
  wire u2__abc_44228_n14252;
  wire u2__abc_44228_n14253;
  wire u2__abc_44228_n14254;
  wire u2__abc_44228_n14255;
  wire u2__abc_44228_n14256;
  wire u2__abc_44228_n14257;
  wire u2__abc_44228_n14258_1;
  wire u2__abc_44228_n14259;
  wire u2__abc_44228_n14260;
  wire u2__abc_44228_n14261;
  wire u2__abc_44228_n14262;
  wire u2__abc_44228_n14263;
  wire u2__abc_44228_n14264;
  wire u2__abc_44228_n14265;
  wire u2__abc_44228_n14266;
  wire u2__abc_44228_n14268_1;
  wire u2__abc_44228_n14269;
  wire u2__abc_44228_n14270;
  wire u2__abc_44228_n14271;
  wire u2__abc_44228_n14272;
  wire u2__abc_44228_n14273;
  wire u2__abc_44228_n14274;
  wire u2__abc_44228_n14275;
  wire u2__abc_44228_n14276_1;
  wire u2__abc_44228_n14277;
  wire u2__abc_44228_n14278;
  wire u2__abc_44228_n14279;
  wire u2__abc_44228_n14280;
  wire u2__abc_44228_n14281;
  wire u2__abc_44228_n14282;
  wire u2__abc_44228_n14283;
  wire u2__abc_44228_n14285_1;
  wire u2__abc_44228_n14286;
  wire u2__abc_44228_n14287;
  wire u2__abc_44228_n14288;
  wire u2__abc_44228_n14289;
  wire u2__abc_44228_n14290;
  wire u2__abc_44228_n14291;
  wire u2__abc_44228_n14292;
  wire u2__abc_44228_n14293_1;
  wire u2__abc_44228_n14294;
  wire u2__abc_44228_n14295;
  wire u2__abc_44228_n14296;
  wire u2__abc_44228_n14297;
  wire u2__abc_44228_n14298;
  wire u2__abc_44228_n14299;
  wire u2__abc_44228_n14300;
  wire u2__abc_44228_n14301;
  wire u2__abc_44228_n14303;
  wire u2__abc_44228_n14304;
  wire u2__abc_44228_n14305;
  wire u2__abc_44228_n14306;
  wire u2__abc_44228_n14307_1;
  wire u2__abc_44228_n14308;
  wire u2__abc_44228_n14309;
  wire u2__abc_44228_n14310;
  wire u2__abc_44228_n14311;
  wire u2__abc_44228_n14312;
  wire u2__abc_44228_n14313;
  wire u2__abc_44228_n14314;
  wire u2__abc_44228_n14315_1;
  wire u2__abc_44228_n14316;
  wire u2__abc_44228_n14317;
  wire u2__abc_44228_n14318;
  wire u2__abc_44228_n14320;
  wire u2__abc_44228_n14321;
  wire u2__abc_44228_n14322;
  wire u2__abc_44228_n14323;
  wire u2__abc_44228_n14324_1;
  wire u2__abc_44228_n14325;
  wire u2__abc_44228_n14326;
  wire u2__abc_44228_n14327;
  wire u2__abc_44228_n14328;
  wire u2__abc_44228_n14329;
  wire u2__abc_44228_n14330;
  wire u2__abc_44228_n14331;
  wire u2__abc_44228_n14332_1;
  wire u2__abc_44228_n14333;
  wire u2__abc_44228_n14334;
  wire u2__abc_44228_n14335;
  wire u2__abc_44228_n14337;
  wire u2__abc_44228_n14338;
  wire u2__abc_44228_n14339;
  wire u2__abc_44228_n14340;
  wire u2__abc_44228_n14341;
  wire u2__abc_44228_n14342_1;
  wire u2__abc_44228_n14343;
  wire u2__abc_44228_n14344;
  wire u2__abc_44228_n14345;
  wire u2__abc_44228_n14346;
  wire u2__abc_44228_n14347;
  wire u2__abc_44228_n14348;
  wire u2__abc_44228_n14349;
  wire u2__abc_44228_n14350_1;
  wire u2__abc_44228_n14351;
  wire u2__abc_44228_n14352;
  wire u2__abc_44228_n14354;
  wire u2__abc_44228_n14355;
  wire u2__abc_44228_n14356;
  wire u2__abc_44228_n14357;
  wire u2__abc_44228_n14358;
  wire u2__abc_44228_n14359_1;
  wire u2__abc_44228_n14360;
  wire u2__abc_44228_n14361;
  wire u2__abc_44228_n14362;
  wire u2__abc_44228_n14363;
  wire u2__abc_44228_n14364;
  wire u2__abc_44228_n14365;
  wire u2__abc_44228_n14366;
  wire u2__abc_44228_n14367_1;
  wire u2__abc_44228_n14368;
  wire u2__abc_44228_n14369;
  wire u2__abc_44228_n14370;
  wire u2__abc_44228_n14372;
  wire u2__abc_44228_n14373;
  wire u2__abc_44228_n14374;
  wire u2__abc_44228_n14375;
  wire u2__abc_44228_n14376;
  wire u2__abc_44228_n14377;
  wire u2__abc_44228_n14378_1;
  wire u2__abc_44228_n14379;
  wire u2__abc_44228_n14380;
  wire u2__abc_44228_n14381;
  wire u2__abc_44228_n14382;
  wire u2__abc_44228_n14383;
  wire u2__abc_44228_n14384;
  wire u2__abc_44228_n14385;
  wire u2__abc_44228_n14386_1;
  wire u2__abc_44228_n14387;
  wire u2__abc_44228_n14389;
  wire u2__abc_44228_n14390;
  wire u2__abc_44228_n14391;
  wire u2__abc_44228_n14392;
  wire u2__abc_44228_n14393;
  wire u2__abc_44228_n14394;
  wire u2__abc_44228_n14395_1;
  wire u2__abc_44228_n14396;
  wire u2__abc_44228_n14397;
  wire u2__abc_44228_n14398;
  wire u2__abc_44228_n14399;
  wire u2__abc_44228_n14400;
  wire u2__abc_44228_n14401;
  wire u2__abc_44228_n14402;
  wire u2__abc_44228_n14403_1;
  wire u2__abc_44228_n14404;
  wire u2__abc_44228_n14406;
  wire u2__abc_44228_n14407;
  wire u2__abc_44228_n14408;
  wire u2__abc_44228_n14409;
  wire u2__abc_44228_n14410;
  wire u2__abc_44228_n14411;
  wire u2__abc_44228_n14412;
  wire u2__abc_44228_n14413_1;
  wire u2__abc_44228_n14414;
  wire u2__abc_44228_n14415;
  wire u2__abc_44228_n14416;
  wire u2__abc_44228_n14417;
  wire u2__abc_44228_n14418;
  wire u2__abc_44228_n14419;
  wire u2__abc_44228_n14420;
  wire u2__abc_44228_n14421_1;
  wire u2__abc_44228_n14423;
  wire u2__abc_44228_n14424;
  wire u2__abc_44228_n14425;
  wire u2__abc_44228_n14426;
  wire u2__abc_44228_n14427;
  wire u2__abc_44228_n14428;
  wire u2__abc_44228_n14429;
  wire u2__abc_44228_n14430_1;
  wire u2__abc_44228_n14431;
  wire u2__abc_44228_n14432;
  wire u2__abc_44228_n14433;
  wire u2__abc_44228_n14434;
  wire u2__abc_44228_n14435;
  wire u2__abc_44228_n14436;
  wire u2__abc_44228_n14437;
  wire u2__abc_44228_n14438_1;
  wire u2__abc_44228_n14439;
  wire u2__abc_44228_n14441;
  wire u2__abc_44228_n14442;
  wire u2__abc_44228_n14443;
  wire u2__abc_44228_n14444;
  wire u2__abc_44228_n14445;
  wire u2__abc_44228_n14446;
  wire u2__abc_44228_n14447;
  wire u2__abc_44228_n14448;
  wire u2__abc_44228_n14449;
  wire u2__abc_44228_n14450_1;
  wire u2__abc_44228_n14451;
  wire u2__abc_44228_n14452;
  wire u2__abc_44228_n14453;
  wire u2__abc_44228_n14454;
  wire u2__abc_44228_n14455;
  wire u2__abc_44228_n14456;
  wire u2__abc_44228_n14458_1;
  wire u2__abc_44228_n14459;
  wire u2__abc_44228_n14460;
  wire u2__abc_44228_n14461;
  wire u2__abc_44228_n14462;
  wire u2__abc_44228_n14463;
  wire u2__abc_44228_n14464;
  wire u2__abc_44228_n14465;
  wire u2__abc_44228_n14466;
  wire u2__abc_44228_n14467_1;
  wire u2__abc_44228_n14468;
  wire u2__abc_44228_n14469;
  wire u2__abc_44228_n14470;
  wire u2__abc_44228_n14471;
  wire u2__abc_44228_n14472;
  wire u2__abc_44228_n14473;
  wire u2__abc_44228_n14475_1;
  wire u2__abc_44228_n14476;
  wire u2__abc_44228_n14477;
  wire u2__abc_44228_n14478;
  wire u2__abc_44228_n14479;
  wire u2__abc_44228_n14480;
  wire u2__abc_44228_n14481;
  wire u2__abc_44228_n14482;
  wire u2__abc_44228_n14483;
  wire u2__abc_44228_n14484;
  wire u2__abc_44228_n14485_1;
  wire u2__abc_44228_n14486;
  wire u2__abc_44228_n14487;
  wire u2__abc_44228_n14488;
  wire u2__abc_44228_n14489;
  wire u2__abc_44228_n14490;
  wire u2__abc_44228_n14492;
  wire u2__abc_44228_n14493_1;
  wire u2__abc_44228_n14494;
  wire u2__abc_44228_n14495;
  wire u2__abc_44228_n14496;
  wire u2__abc_44228_n14497;
  wire u2__abc_44228_n14498;
  wire u2__abc_44228_n14499;
  wire u2__abc_44228_n14500;
  wire u2__abc_44228_n14501;
  wire u2__abc_44228_n14502_1;
  wire u2__abc_44228_n14503;
  wire u2__abc_44228_n14504;
  wire u2__abc_44228_n14505;
  wire u2__abc_44228_n14506;
  wire u2__abc_44228_n14507;
  wire u2__abc_44228_n14509;
  wire u2__abc_44228_n14510_1;
  wire u2__abc_44228_n14511;
  wire u2__abc_44228_n14512;
  wire u2__abc_44228_n14513;
  wire u2__abc_44228_n14514;
  wire u2__abc_44228_n14515;
  wire u2__abc_44228_n14516;
  wire u2__abc_44228_n14517;
  wire u2__abc_44228_n14518;
  wire u2__abc_44228_n14519;
  wire u2__abc_44228_n14520;
  wire u2__abc_44228_n14521_1;
  wire u2__abc_44228_n14522;
  wire u2__abc_44228_n14523;
  wire u2__abc_44228_n14524;
  wire u2__abc_44228_n14526;
  wire u2__abc_44228_n14527;
  wire u2__abc_44228_n14528;
  wire u2__abc_44228_n14529_1;
  wire u2__abc_44228_n14530;
  wire u2__abc_44228_n14531;
  wire u2__abc_44228_n14532;
  wire u2__abc_44228_n14533;
  wire u2__abc_44228_n14534;
  wire u2__abc_44228_n14535;
  wire u2__abc_44228_n14536;
  wire u2__abc_44228_n14537;
  wire u2__abc_44228_n14538_1;
  wire u2__abc_44228_n14539;
  wire u2__abc_44228_n14540;
  wire u2__abc_44228_n14541;
  wire u2__abc_44228_n14543;
  wire u2__abc_44228_n14544;
  wire u2__abc_44228_n14545;
  wire u2__abc_44228_n14546_1;
  wire u2__abc_44228_n14547;
  wire u2__abc_44228_n14548;
  wire u2__abc_44228_n14549;
  wire u2__abc_44228_n14550;
  wire u2__abc_44228_n14551;
  wire u2__abc_44228_n14552;
  wire u2__abc_44228_n14553;
  wire u2__abc_44228_n14554;
  wire u2__abc_44228_n14555;
  wire u2__abc_44228_n14556_1;
  wire u2__abc_44228_n14557;
  wire u2__abc_44228_n14558;
  wire u2__abc_44228_n14560;
  wire u2__abc_44228_n14561;
  wire u2__abc_44228_n14562;
  wire u2__abc_44228_n14563;
  wire u2__abc_44228_n14564_1;
  wire u2__abc_44228_n14565;
  wire u2__abc_44228_n14566;
  wire u2__abc_44228_n14567;
  wire u2__abc_44228_n14568;
  wire u2__abc_44228_n14569;
  wire u2__abc_44228_n14570;
  wire u2__abc_44228_n14571;
  wire u2__abc_44228_n14572;
  wire u2__abc_44228_n14573_1;
  wire u2__abc_44228_n14574;
  wire u2__abc_44228_n14575;
  wire u2__abc_44228_n14576;
  wire u2__abc_44228_n14578;
  wire u2__abc_44228_n14579;
  wire u2__abc_44228_n14580;
  wire u2__abc_44228_n14581_1;
  wire u2__abc_44228_n14582;
  wire u2__abc_44228_n14583;
  wire u2__abc_44228_n14584;
  wire u2__abc_44228_n14585;
  wire u2__abc_44228_n14586;
  wire u2__abc_44228_n14587;
  wire u2__abc_44228_n14588;
  wire u2__abc_44228_n14589;
  wire u2__abc_44228_n14590;
  wire u2__abc_44228_n14591;
  wire u2__abc_44228_n14592;
  wire u2__abc_44228_n14593;
  wire u2__abc_44228_n14595;
  wire u2__abc_44228_n14596;
  wire u2__abc_44228_n14597;
  wire u2__abc_44228_n14598;
  wire u2__abc_44228_n14599;
  wire u2__abc_44228_n14600;
  wire u2__abc_44228_n14601;
  wire u2__abc_44228_n14602_1;
  wire u2__abc_44228_n14603;
  wire u2__abc_44228_n14604;
  wire u2__abc_44228_n14605;
  wire u2__abc_44228_n14606;
  wire u2__abc_44228_n14607;
  wire u2__abc_44228_n14608;
  wire u2__abc_44228_n14609;
  wire u2__abc_44228_n14610;
  wire u2__abc_44228_n14612;
  wire u2__abc_44228_n14613;
  wire u2__abc_44228_n14614;
  wire u2__abc_44228_n14615;
  wire u2__abc_44228_n14616;
  wire u2__abc_44228_n14617;
  wire u2__abc_44228_n14618;
  wire u2__abc_44228_n14619_1;
  wire u2__abc_44228_n14620;
  wire u2__abc_44228_n14621;
  wire u2__abc_44228_n14622;
  wire u2__abc_44228_n14623;
  wire u2__abc_44228_n14624;
  wire u2__abc_44228_n14625;
  wire u2__abc_44228_n14626;
  wire u2__abc_44228_n14627;
  wire u2__abc_44228_n14629_1;
  wire u2__abc_44228_n14630;
  wire u2__abc_44228_n14631;
  wire u2__abc_44228_n14632;
  wire u2__abc_44228_n14633;
  wire u2__abc_44228_n14634;
  wire u2__abc_44228_n14635;
  wire u2__abc_44228_n14636;
  wire u2__abc_44228_n14637_1;
  wire u2__abc_44228_n14638;
  wire u2__abc_44228_n14639;
  wire u2__abc_44228_n14640;
  wire u2__abc_44228_n14641;
  wire u2__abc_44228_n14642;
  wire u2__abc_44228_n14643;
  wire u2__abc_44228_n14644;
  wire u2__abc_44228_n14645;
  wire u2__abc_44228_n14647;
  wire u2__abc_44228_n14648;
  wire u2__abc_44228_n14649;
  wire u2__abc_44228_n14650;
  wire u2__abc_44228_n14651;
  wire u2__abc_44228_n14652;
  wire u2__abc_44228_n14653;
  wire u2__abc_44228_n14654_1;
  wire u2__abc_44228_n14655;
  wire u2__abc_44228_n14656;
  wire u2__abc_44228_n14657;
  wire u2__abc_44228_n14658;
  wire u2__abc_44228_n14659;
  wire u2__abc_44228_n14660;
  wire u2__abc_44228_n14661;
  wire u2__abc_44228_n14662;
  wire u2__abc_44228_n14664;
  wire u2__abc_44228_n14665_1;
  wire u2__abc_44228_n14666;
  wire u2__abc_44228_n14667;
  wire u2__abc_44228_n14668;
  wire u2__abc_44228_n14669;
  wire u2__abc_44228_n14670;
  wire u2__abc_44228_n14671;
  wire u2__abc_44228_n14672;
  wire u2__abc_44228_n14673_1;
  wire u2__abc_44228_n14674;
  wire u2__abc_44228_n14675;
  wire u2__abc_44228_n14676;
  wire u2__abc_44228_n14677;
  wire u2__abc_44228_n14678;
  wire u2__abc_44228_n14679;
  wire u2__abc_44228_n14681;
  wire u2__abc_44228_n14682_1;
  wire u2__abc_44228_n14683;
  wire u2__abc_44228_n14684;
  wire u2__abc_44228_n14685;
  wire u2__abc_44228_n14686;
  wire u2__abc_44228_n14687;
  wire u2__abc_44228_n14688;
  wire u2__abc_44228_n14689;
  wire u2__abc_44228_n14690_1;
  wire u2__abc_44228_n14691;
  wire u2__abc_44228_n14692;
  wire u2__abc_44228_n14693;
  wire u2__abc_44228_n14694;
  wire u2__abc_44228_n14695;
  wire u2__abc_44228_n14696;
  wire u2__abc_44228_n14698;
  wire u2__abc_44228_n14699;
  wire u2__abc_44228_n14700_1;
  wire u2__abc_44228_n14701;
  wire u2__abc_44228_n14702;
  wire u2__abc_44228_n14703;
  wire u2__abc_44228_n14704;
  wire u2__abc_44228_n14705;
  wire u2__abc_44228_n14706;
  wire u2__abc_44228_n14707;
  wire u2__abc_44228_n14708_1;
  wire u2__abc_44228_n14709;
  wire u2__abc_44228_n14710;
  wire u2__abc_44228_n14711;
  wire u2__abc_44228_n14712;
  wire u2__abc_44228_n14713;
  wire u2__abc_44228_n14714;
  wire u2__abc_44228_n14716;
  wire u2__abc_44228_n14717_1;
  wire u2__abc_44228_n14718;
  wire u2__abc_44228_n14719;
  wire u2__abc_44228_n14720;
  wire u2__abc_44228_n14721;
  wire u2__abc_44228_n14722;
  wire u2__abc_44228_n14723;
  wire u2__abc_44228_n14724;
  wire u2__abc_44228_n14725_1;
  wire u2__abc_44228_n14726;
  wire u2__abc_44228_n14727;
  wire u2__abc_44228_n14728;
  wire u2__abc_44228_n14729;
  wire u2__abc_44228_n14730;
  wire u2__abc_44228_n14731;
  wire u2__abc_44228_n14733;
  wire u2__abc_44228_n14734;
  wire u2__abc_44228_n14735;
  wire u2__abc_44228_n14736;
  wire u2__abc_44228_n14737_1;
  wire u2__abc_44228_n14738;
  wire u2__abc_44228_n14739;
  wire u2__abc_44228_n14740;
  wire u2__abc_44228_n14741;
  wire u2__abc_44228_n14742;
  wire u2__abc_44228_n14743;
  wire u2__abc_44228_n14744;
  wire u2__abc_44228_n14745_1;
  wire u2__abc_44228_n14746;
  wire u2__abc_44228_n14747;
  wire u2__abc_44228_n14748;
  wire u2__abc_44228_n14750;
  wire u2__abc_44228_n14751;
  wire u2__abc_44228_n14752;
  wire u2__abc_44228_n14753;
  wire u2__abc_44228_n14754_1;
  wire u2__abc_44228_n14755;
  wire u2__abc_44228_n14756;
  wire u2__abc_44228_n14757;
  wire u2__abc_44228_n14758;
  wire u2__abc_44228_n14759;
  wire u2__abc_44228_n14760;
  wire u2__abc_44228_n14761;
  wire u2__abc_44228_n14762_1;
  wire u2__abc_44228_n14763;
  wire u2__abc_44228_n14764;
  wire u2__abc_44228_n14765;
  wire u2__abc_44228_n14767;
  wire u2__abc_44228_n14768;
  wire u2__abc_44228_n14769;
  wire u2__abc_44228_n14770;
  wire u2__abc_44228_n14771;
  wire u2__abc_44228_n14772_1;
  wire u2__abc_44228_n14773;
  wire u2__abc_44228_n14774;
  wire u2__abc_44228_n14775;
  wire u2__abc_44228_n14776;
  wire u2__abc_44228_n14777;
  wire u2__abc_44228_n14778;
  wire u2__abc_44228_n14779;
  wire u2__abc_44228_n14780_1;
  wire u2__abc_44228_n14781;
  wire u2__abc_44228_n14782;
  wire u2__abc_44228_n14784;
  wire u2__abc_44228_n14785;
  wire u2__abc_44228_n14786;
  wire u2__abc_44228_n14787;
  wire u2__abc_44228_n14788;
  wire u2__abc_44228_n14789_1;
  wire u2__abc_44228_n14790;
  wire u2__abc_44228_n14791;
  wire u2__abc_44228_n14792;
  wire u2__abc_44228_n14793;
  wire u2__abc_44228_n14794;
  wire u2__abc_44228_n14795;
  wire u2__abc_44228_n14796;
  wire u2__abc_44228_n14797_1;
  wire u2__abc_44228_n14798;
  wire u2__abc_44228_n14799;
  wire u2__abc_44228_n14801;
  wire u2__abc_44228_n14802;
  wire u2__abc_44228_n14803;
  wire u2__abc_44228_n14804;
  wire u2__abc_44228_n14805;
  wire u2__abc_44228_n14806;
  wire u2__abc_44228_n14807;
  wire u2__abc_44228_n14808_1;
  wire u2__abc_44228_n14809;
  wire u2__abc_44228_n14810;
  wire u2__abc_44228_n14811;
  wire u2__abc_44228_n14812;
  wire u2__abc_44228_n14813;
  wire u2__abc_44228_n14814;
  wire u2__abc_44228_n14815;
  wire u2__abc_44228_n14816_1;
  wire u2__abc_44228_n14818;
  wire u2__abc_44228_n14819;
  wire u2__abc_44228_n14820;
  wire u2__abc_44228_n14821;
  wire u2__abc_44228_n14822;
  wire u2__abc_44228_n14823;
  wire u2__abc_44228_n14824;
  wire u2__abc_44228_n14825_1;
  wire u2__abc_44228_n14826;
  wire u2__abc_44228_n14827;
  wire u2__abc_44228_n14828;
  wire u2__abc_44228_n14829;
  wire u2__abc_44228_n14830;
  wire u2__abc_44228_n14831;
  wire u2__abc_44228_n14832;
  wire u2__abc_44228_n14833_1;
  wire u2__abc_44228_n14835;
  wire u2__abc_44228_n14836;
  wire u2__abc_44228_n14837;
  wire u2__abc_44228_n14838;
  wire u2__abc_44228_n14839;
  wire u2__abc_44228_n14840;
  wire u2__abc_44228_n14841;
  wire u2__abc_44228_n14842;
  wire u2__abc_44228_n14843_1;
  wire u2__abc_44228_n14844;
  wire u2__abc_44228_n14845;
  wire u2__abc_44228_n14846;
  wire u2__abc_44228_n14847;
  wire u2__abc_44228_n14848;
  wire u2__abc_44228_n14849;
  wire u2__abc_44228_n14850;
  wire u2__abc_44228_n14852;
  wire u2__abc_44228_n14853;
  wire u2__abc_44228_n14854;
  wire u2__abc_44228_n14855;
  wire u2__abc_44228_n14856;
  wire u2__abc_44228_n14857;
  wire u2__abc_44228_n14858;
  wire u2__abc_44228_n14859;
  wire u2__abc_44228_n14860_1;
  wire u2__abc_44228_n14861;
  wire u2__abc_44228_n14862;
  wire u2__abc_44228_n14863;
  wire u2__abc_44228_n14864;
  wire u2__abc_44228_n14865;
  wire u2__abc_44228_n14866;
  wire u2__abc_44228_n14867;
  wire u2__abc_44228_n14869;
  wire u2__abc_44228_n14870;
  wire u2__abc_44228_n14871;
  wire u2__abc_44228_n14872;
  wire u2__abc_44228_n14873;
  wire u2__abc_44228_n14874;
  wire u2__abc_44228_n14875;
  wire u2__abc_44228_n14876;
  wire u2__abc_44228_n14877;
  wire u2__abc_44228_n14878;
  wire u2__abc_44228_n14879;
  wire u2__abc_44228_n14880;
  wire u2__abc_44228_n14881;
  wire u2__abc_44228_n14882;
  wire u2__abc_44228_n14883_1;
  wire u2__abc_44228_n14884;
  wire u2__abc_44228_n14885;
  wire u2__abc_44228_n14887;
  wire u2__abc_44228_n14888;
  wire u2__abc_44228_n14889;
  wire u2__abc_44228_n14890;
  wire u2__abc_44228_n14891_1;
  wire u2__abc_44228_n14892;
  wire u2__abc_44228_n14893;
  wire u2__abc_44228_n14894;
  wire u2__abc_44228_n14895;
  wire u2__abc_44228_n14896;
  wire u2__abc_44228_n14897;
  wire u2__abc_44228_n14898;
  wire u2__abc_44228_n14899;
  wire u2__abc_44228_n14900_1;
  wire u2__abc_44228_n14901;
  wire u2__abc_44228_n14902;
  wire u2__abc_44228_n14904;
  wire u2__abc_44228_n14905;
  wire u2__abc_44228_n14906;
  wire u2__abc_44228_n14907;
  wire u2__abc_44228_n14908_1;
  wire u2__abc_44228_n14909;
  wire u2__abc_44228_n14910;
  wire u2__abc_44228_n14911;
  wire u2__abc_44228_n14912;
  wire u2__abc_44228_n14913;
  wire u2__abc_44228_n14914;
  wire u2__abc_44228_n14915;
  wire u2__abc_44228_n14916;
  wire u2__abc_44228_n14917;
  wire u2__abc_44228_n14918_1;
  wire u2__abc_44228_n14919;
  wire u2__abc_44228_n14920;
  wire u2__abc_44228_n14922;
  wire u2__abc_44228_n14923;
  wire u2__abc_44228_n14924;
  wire u2__abc_44228_n14925;
  wire u2__abc_44228_n14926_1;
  wire u2__abc_44228_n14927;
  wire u2__abc_44228_n14928;
  wire u2__abc_44228_n14929;
  wire u2__abc_44228_n14930;
  wire u2__abc_44228_n14931;
  wire u2__abc_44228_n14932;
  wire u2__abc_44228_n14933;
  wire u2__abc_44228_n14934;
  wire u2__abc_44228_n14935_1;
  wire u2__abc_44228_n14936;
  wire u2__abc_44228_n14937;
  wire u2__abc_44228_n14939;
  wire u2__abc_44228_n14940;
  wire u2__abc_44228_n14941;
  wire u2__abc_44228_n14942;
  wire u2__abc_44228_n14943_1;
  wire u2__abc_44228_n14944;
  wire u2__abc_44228_n14945;
  wire u2__abc_44228_n14946;
  wire u2__abc_44228_n14947;
  wire u2__abc_44228_n14948;
  wire u2__abc_44228_n14949;
  wire u2__abc_44228_n14950;
  wire u2__abc_44228_n14951;
  wire u2__abc_44228_n14952;
  wire u2__abc_44228_n14953;
  wire u2__abc_44228_n14954_1;
  wire u2__abc_44228_n14956;
  wire u2__abc_44228_n14957;
  wire u2__abc_44228_n14958;
  wire u2__abc_44228_n14959;
  wire u2__abc_44228_n14960;
  wire u2__abc_44228_n14961;
  wire u2__abc_44228_n14962_1;
  wire u2__abc_44228_n14963;
  wire u2__abc_44228_n14964;
  wire u2__abc_44228_n14965;
  wire u2__abc_44228_n14966;
  wire u2__abc_44228_n14967;
  wire u2__abc_44228_n14968;
  wire u2__abc_44228_n14969;
  wire u2__abc_44228_n14970;
  wire u2__abc_44228_n14971_1;
  wire u2__abc_44228_n14973;
  wire u2__abc_44228_n14974;
  wire u2__abc_44228_n14975;
  wire u2__abc_44228_n14976;
  wire u2__abc_44228_n14977;
  wire u2__abc_44228_n14978;
  wire u2__abc_44228_n14979_1;
  wire u2__abc_44228_n14980;
  wire u2__abc_44228_n14981;
  wire u2__abc_44228_n14982;
  wire u2__abc_44228_n14983;
  wire u2__abc_44228_n14984;
  wire u2__abc_44228_n14985;
  wire u2__abc_44228_n14986;
  wire u2__abc_44228_n14987;
  wire u2__abc_44228_n14988;
  wire u2__abc_44228_n14990;
  wire u2__abc_44228_n14991;
  wire u2__abc_44228_n14992;
  wire u2__abc_44228_n14993;
  wire u2__abc_44228_n14994;
  wire u2__abc_44228_n14995;
  wire u2__abc_44228_n14996;
  wire u2__abc_44228_n14997_1;
  wire u2__abc_44228_n14998;
  wire u2__abc_44228_n14999;
  wire u2__abc_44228_n15000;
  wire u2__abc_44228_n15001;
  wire u2__abc_44228_n15002;
  wire u2__abc_44228_n15003;
  wire u2__abc_44228_n15004;
  wire u2__abc_44228_n15005;
  wire u2__abc_44228_n15007;
  wire u2__abc_44228_n15008;
  wire u2__abc_44228_n15009;
  wire u2__abc_44228_n15010;
  wire u2__abc_44228_n15011;
  wire u2__abc_44228_n15012;
  wire u2__abc_44228_n15013;
  wire u2__abc_44228_n15014_1;
  wire u2__abc_44228_n15015;
  wire u2__abc_44228_n15016;
  wire u2__abc_44228_n15017;
  wire u2__abc_44228_n15018;
  wire u2__abc_44228_n15019;
  wire u2__abc_44228_n15020;
  wire u2__abc_44228_n15021;
  wire u2__abc_44228_n15022;
  wire u2__abc_44228_n15023;
  wire u2__abc_44228_n15025;
  wire u2__abc_44228_n15026_1;
  wire u2__abc_44228_n15027;
  wire u2__abc_44228_n15028;
  wire u2__abc_44228_n15029;
  wire u2__abc_44228_n15030;
  wire u2__abc_44228_n15031;
  wire u2__abc_44228_n15032;
  wire u2__abc_44228_n15033;
  wire u2__abc_44228_n15034_1;
  wire u2__abc_44228_n15035;
  wire u2__abc_44228_n15036;
  wire u2__abc_44228_n15037;
  wire u2__abc_44228_n15038;
  wire u2__abc_44228_n15039;
  wire u2__abc_44228_n15040;
  wire u2__abc_44228_n15042;
  wire u2__abc_44228_n15043_1;
  wire u2__abc_44228_n15044;
  wire u2__abc_44228_n15045;
  wire u2__abc_44228_n15046;
  wire u2__abc_44228_n15047;
  wire u2__abc_44228_n15048;
  wire u2__abc_44228_n15049;
  wire u2__abc_44228_n15050;
  wire u2__abc_44228_n15051_1;
  wire u2__abc_44228_n15052;
  wire u2__abc_44228_n15053;
  wire u2__abc_44228_n15054;
  wire u2__abc_44228_n15055;
  wire u2__abc_44228_n15056;
  wire u2__abc_44228_n15057;
  wire u2__abc_44228_n15058;
  wire u2__abc_44228_n15060;
  wire u2__abc_44228_n15061_1;
  wire u2__abc_44228_n15062;
  wire u2__abc_44228_n15063;
  wire u2__abc_44228_n15064;
  wire u2__abc_44228_n15065;
  wire u2__abc_44228_n15066;
  wire u2__abc_44228_n15067;
  wire u2__abc_44228_n15068;
  wire u2__abc_44228_n15069_1;
  wire u2__abc_44228_n15070;
  wire u2__abc_44228_n15071;
  wire u2__abc_44228_n15072;
  wire u2__abc_44228_n15073;
  wire u2__abc_44228_n15074;
  wire u2__abc_44228_n15075;
  wire u2__abc_44228_n15077;
  wire u2__abc_44228_n15078_1;
  wire u2__abc_44228_n15079;
  wire u2__abc_44228_n15080;
  wire u2__abc_44228_n15081;
  wire u2__abc_44228_n15082;
  wire u2__abc_44228_n15083;
  wire u2__abc_44228_n15084;
  wire u2__abc_44228_n15085;
  wire u2__abc_44228_n15086_1;
  wire u2__abc_44228_n15087;
  wire u2__abc_44228_n15088;
  wire u2__abc_44228_n15089;
  wire u2__abc_44228_n15090;
  wire u2__abc_44228_n15091;
  wire u2__abc_44228_n15092;
  wire u2__abc_44228_n15094;
  wire u2__abc_44228_n15095;
  wire u2__abc_44228_n15096;
  wire u2__abc_44228_n15097_1;
  wire u2__abc_44228_n15098;
  wire u2__abc_44228_n15099;
  wire u2__abc_44228_n15100;
  wire u2__abc_44228_n15101;
  wire u2__abc_44228_n15102;
  wire u2__abc_44228_n15103;
  wire u2__abc_44228_n15104;
  wire u2__abc_44228_n15105_1;
  wire u2__abc_44228_n15106;
  wire u2__abc_44228_n15107;
  wire u2__abc_44228_n15108;
  wire u2__abc_44228_n15109;
  wire u2__abc_44228_n15111;
  wire u2__abc_44228_n15112;
  wire u2__abc_44228_n15113;
  wire u2__abc_44228_n15114_1;
  wire u2__abc_44228_n15115;
  wire u2__abc_44228_n15116;
  wire u2__abc_44228_n15117;
  wire u2__abc_44228_n15118;
  wire u2__abc_44228_n15119;
  wire u2__abc_44228_n15120;
  wire u2__abc_44228_n15121;
  wire u2__abc_44228_n15122_1;
  wire u2__abc_44228_n15123;
  wire u2__abc_44228_n15124;
  wire u2__abc_44228_n15125;
  wire u2__abc_44228_n15126;
  wire u2__abc_44228_n15127;
  wire u2__abc_44228_n15129;
  wire u2__abc_44228_n15130;
  wire u2__abc_44228_n15131;
  wire u2__abc_44228_n15132_1;
  wire u2__abc_44228_n15133;
  wire u2__abc_44228_n15134;
  wire u2__abc_44228_n15135;
  wire u2__abc_44228_n15136;
  wire u2__abc_44228_n15137;
  wire u2__abc_44228_n15138;
  wire u2__abc_44228_n15139;
  wire u2__abc_44228_n15140_1;
  wire u2__abc_44228_n15141;
  wire u2__abc_44228_n15142;
  wire u2__abc_44228_n15143;
  wire u2__abc_44228_n15144;
  wire u2__abc_44228_n15146;
  wire u2__abc_44228_n15147;
  wire u2__abc_44228_n15148;
  wire u2__abc_44228_n15149_1;
  wire u2__abc_44228_n15150;
  wire u2__abc_44228_n15151;
  wire u2__abc_44228_n15152;
  wire u2__abc_44228_n15153;
  wire u2__abc_44228_n15154;
  wire u2__abc_44228_n15155;
  wire u2__abc_44228_n15156;
  wire u2__abc_44228_n15157_1;
  wire u2__abc_44228_n15158;
  wire u2__abc_44228_n15159;
  wire u2__abc_44228_n15160;
  wire u2__abc_44228_n15161;
  wire u2__abc_44228_n15163;
  wire u2__abc_44228_n15164;
  wire u2__abc_44228_n15165;
  wire u2__abc_44228_n15166;
  wire u2__abc_44228_n15167;
  wire u2__abc_44228_n15168;
  wire u2__abc_44228_n15169;
  wire u2__abc_44228_n15170_1;
  wire u2__abc_44228_n15171;
  wire u2__abc_44228_n15172;
  wire u2__abc_44228_n15173;
  wire u2__abc_44228_n15174;
  wire u2__abc_44228_n15175;
  wire u2__abc_44228_n15176;
  wire u2__abc_44228_n15177;
  wire u2__abc_44228_n15178_1;
  wire u2__abc_44228_n15180;
  wire u2__abc_44228_n15181;
  wire u2__abc_44228_n15182;
  wire u2__abc_44228_n15183;
  wire u2__abc_44228_n15184;
  wire u2__abc_44228_n15185;
  wire u2__abc_44228_n15186;
  wire u2__abc_44228_n15187_1;
  wire u2__abc_44228_n15188;
  wire u2__abc_44228_n15189;
  wire u2__abc_44228_n15190;
  wire u2__abc_44228_n15191;
  wire u2__abc_44228_n15192;
  wire u2__abc_44228_n15193;
  wire u2__abc_44228_n15194;
  wire u2__abc_44228_n15195_1;
  wire u2__abc_44228_n15197;
  wire u2__abc_44228_n15198;
  wire u2__abc_44228_n15199;
  wire u2__abc_44228_n15200;
  wire u2__abc_44228_n15201;
  wire u2__abc_44228_n15202;
  wire u2__abc_44228_n15203;
  wire u2__abc_44228_n15204;
  wire u2__abc_44228_n15205_1;
  wire u2__abc_44228_n15206;
  wire u2__abc_44228_n15207;
  wire u2__abc_44228_n15208;
  wire u2__abc_44228_n15209;
  wire u2__abc_44228_n15210;
  wire u2__abc_44228_n15211;
  wire u2__abc_44228_n15212;
  wire u2__abc_44228_n15214;
  wire u2__abc_44228_n15215;
  wire u2__abc_44228_n15216;
  wire u2__abc_44228_n15217;
  wire u2__abc_44228_n15218;
  wire u2__abc_44228_n15219;
  wire u2__abc_44228_n15220;
  wire u2__abc_44228_n15221;
  wire u2__abc_44228_n15222_1;
  wire u2__abc_44228_n15223;
  wire u2__abc_44228_n15224;
  wire u2__abc_44228_n15225;
  wire u2__abc_44228_n15226;
  wire u2__abc_44228_n15227;
  wire u2__abc_44228_n15229;
  wire u2__abc_44228_n15230_1;
  wire u2__abc_44228_n15231;
  wire u2__abc_44228_n15232;
  wire u2__abc_44228_n15233;
  wire u2__abc_44228_n15234;
  wire u2__abc_44228_n15235;
  wire u2__abc_44228_n15236;
  wire u2__abc_44228_n15237;
  wire u2__abc_44228_n15238;
  wire u2__abc_44228_n15239;
  wire u2__abc_44228_n15240;
  wire u2__abc_44228_n15241_1;
  wire u2__abc_44228_n15242;
  wire u2__abc_44228_n15243;
  wire u2__abc_44228_n15244;
  wire u2__abc_44228_n15246;
  wire u2__abc_44228_n15247;
  wire u2__abc_44228_n15247_bF_buf0;
  wire u2__abc_44228_n15247_bF_buf1;
  wire u2__abc_44228_n15247_bF_buf10;
  wire u2__abc_44228_n15247_bF_buf11;
  wire u2__abc_44228_n15247_bF_buf12;
  wire u2__abc_44228_n15247_bF_buf13;
  wire u2__abc_44228_n15247_bF_buf14;
  wire u2__abc_44228_n15247_bF_buf2;
  wire u2__abc_44228_n15247_bF_buf3;
  wire u2__abc_44228_n15247_bF_buf4;
  wire u2__abc_44228_n15247_bF_buf5;
  wire u2__abc_44228_n15247_bF_buf6;
  wire u2__abc_44228_n15247_bF_buf7;
  wire u2__abc_44228_n15247_bF_buf8;
  wire u2__abc_44228_n15247_bF_buf9;
  wire u2__abc_44228_n15248;
  wire u2__abc_44228_n15250;
  wire u2__abc_44228_n15252;
  wire u2__abc_44228_n15253;
  wire u2__abc_44228_n15254;
  wire u2__abc_44228_n15255;
  wire u2__abc_44228_n15257;
  wire u2__abc_44228_n15258_1;
  wire u2__abc_44228_n15259;
  wire u2__abc_44228_n15260;
  wire u2__abc_44228_n15262;
  wire u2__abc_44228_n15263;
  wire u2__abc_44228_n15264;
  wire u2__abc_44228_n15265;
  wire u2__abc_44228_n15267;
  wire u2__abc_44228_n15268;
  wire u2__abc_44228_n15269;
  wire u2__abc_44228_n15270;
  wire u2__abc_44228_n15272;
  wire u2__abc_44228_n15273;
  wire u2__abc_44228_n15274;
  wire u2__abc_44228_n15275;
  wire u2__abc_44228_n15277;
  wire u2__abc_44228_n15278;
  wire u2__abc_44228_n15279;
  wire u2__abc_44228_n15280;
  wire u2__abc_44228_n15282;
  wire u2__abc_44228_n15283;
  wire u2__abc_44228_n15284_1;
  wire u2__abc_44228_n15285;
  wire u2__abc_44228_n15287;
  wire u2__abc_44228_n15288;
  wire u2__abc_44228_n15289;
  wire u2__abc_44228_n15290;
  wire u2__abc_44228_n15292;
  wire u2__abc_44228_n15293_1;
  wire u2__abc_44228_n15294;
  wire u2__abc_44228_n15295;
  wire u2__abc_44228_n15297;
  wire u2__abc_44228_n15298;
  wire u2__abc_44228_n15299;
  wire u2__abc_44228_n15300;
  wire u2__abc_44228_n15302;
  wire u2__abc_44228_n15303;
  wire u2__abc_44228_n15304;
  wire u2__abc_44228_n15305;
  wire u2__abc_44228_n15307;
  wire u2__abc_44228_n15308;
  wire u2__abc_44228_n15309;
  wire u2__abc_44228_n15310;
  wire u2__abc_44228_n15312;
  wire u2__abc_44228_n15313_1;
  wire u2__abc_44228_n15314;
  wire u2__abc_44228_n15315;
  wire u2__abc_44228_n15317;
  wire u2__abc_44228_n15318;
  wire u2__abc_44228_n15319;
  wire u2__abc_44228_n15320;
  wire u2__abc_44228_n15322;
  wire u2__abc_44228_n15323;
  wire u2__abc_44228_n15324;
  wire u2__abc_44228_n15325;
  wire u2__abc_44228_n15327;
  wire u2__abc_44228_n15328;
  wire u2__abc_44228_n15329;
  wire u2__abc_44228_n15330_1;
  wire u2__abc_44228_n15332;
  wire u2__abc_44228_n15333;
  wire u2__abc_44228_n15334;
  wire u2__abc_44228_n15335;
  wire u2__abc_44228_n15337;
  wire u2__abc_44228_n15338_1;
  wire u2__abc_44228_n15339;
  wire u2__abc_44228_n15340;
  wire u2__abc_44228_n15342;
  wire u2__abc_44228_n15343;
  wire u2__abc_44228_n15344;
  wire u2__abc_44228_n15345;
  wire u2__abc_44228_n15347;
  wire u2__abc_44228_n15348_1;
  wire u2__abc_44228_n15349;
  wire u2__abc_44228_n15350;
  wire u2__abc_44228_n15352;
  wire u2__abc_44228_n15353;
  wire u2__abc_44228_n15354;
  wire u2__abc_44228_n15355;
  wire u2__abc_44228_n15357;
  wire u2__abc_44228_n15358;
  wire u2__abc_44228_n15359;
  wire u2__abc_44228_n15360;
  wire u2__abc_44228_n15362;
  wire u2__abc_44228_n15363;
  wire u2__abc_44228_n15364;
  wire u2__abc_44228_n15365_1;
  wire u2__abc_44228_n15367;
  wire u2__abc_44228_n15368;
  wire u2__abc_44228_n15369;
  wire u2__abc_44228_n15370;
  wire u2__abc_44228_n15372;
  wire u2__abc_44228_n15373_1;
  wire u2__abc_44228_n15374;
  wire u2__abc_44228_n15375;
  wire u2__abc_44228_n15377;
  wire u2__abc_44228_n15378;
  wire u2__abc_44228_n15379;
  wire u2__abc_44228_n15380;
  wire u2__abc_44228_n15382;
  wire u2__abc_44228_n15383;
  wire u2__abc_44228_n15384_1;
  wire u2__abc_44228_n15385;
  wire u2__abc_44228_n15387;
  wire u2__abc_44228_n15388;
  wire u2__abc_44228_n15389;
  wire u2__abc_44228_n15390;
  wire u2__abc_44228_n15392_1;
  wire u2__abc_44228_n15393;
  wire u2__abc_44228_n15394;
  wire u2__abc_44228_n15395;
  wire u2__abc_44228_n15397;
  wire u2__abc_44228_n15398;
  wire u2__abc_44228_n15399;
  wire u2__abc_44228_n15400;
  wire u2__abc_44228_n15402;
  wire u2__abc_44228_n15402_bF_buf0;
  wire u2__abc_44228_n15402_bF_buf1;
  wire u2__abc_44228_n15402_bF_buf2;
  wire u2__abc_44228_n15402_bF_buf3;
  wire u2__abc_44228_n15403;
  wire u2__abc_44228_n15403_bF_buf0;
  wire u2__abc_44228_n15403_bF_buf1;
  wire u2__abc_44228_n15403_bF_buf2;
  wire u2__abc_44228_n15403_bF_buf3;
  wire u2__abc_44228_n15404;
  wire u2__abc_44228_n15405;
  wire u2__abc_44228_n15405_bF_buf0;
  wire u2__abc_44228_n15405_bF_buf1;
  wire u2__abc_44228_n15405_bF_buf10;
  wire u2__abc_44228_n15405_bF_buf11;
  wire u2__abc_44228_n15405_bF_buf12;
  wire u2__abc_44228_n15405_bF_buf13;
  wire u2__abc_44228_n15405_bF_buf2;
  wire u2__abc_44228_n15405_bF_buf3;
  wire u2__abc_44228_n15405_bF_buf4;
  wire u2__abc_44228_n15405_bF_buf5;
  wire u2__abc_44228_n15405_bF_buf6;
  wire u2__abc_44228_n15405_bF_buf7;
  wire u2__abc_44228_n15405_bF_buf8;
  wire u2__abc_44228_n15405_bF_buf9;
  wire u2__abc_44228_n15406;
  wire u2__abc_44228_n15407;
  wire u2__abc_44228_n15408;
  wire u2__abc_44228_n15408_bF_buf0;
  wire u2__abc_44228_n15408_bF_buf1;
  wire u2__abc_44228_n15408_bF_buf10;
  wire u2__abc_44228_n15408_bF_buf11;
  wire u2__abc_44228_n15408_bF_buf12;
  wire u2__abc_44228_n15408_bF_buf13;
  wire u2__abc_44228_n15408_bF_buf14;
  wire u2__abc_44228_n15408_bF_buf2;
  wire u2__abc_44228_n15408_bF_buf3;
  wire u2__abc_44228_n15408_bF_buf4;
  wire u2__abc_44228_n15408_bF_buf5;
  wire u2__abc_44228_n15408_bF_buf6;
  wire u2__abc_44228_n15408_bF_buf7;
  wire u2__abc_44228_n15408_bF_buf8;
  wire u2__abc_44228_n15408_bF_buf9;
  wire u2__abc_44228_n15409_1;
  wire u2__abc_44228_n15410;
  wire u2__abc_44228_n15411;
  wire u2__abc_44228_n15413;
  wire u2__abc_44228_n15414;
  wire u2__abc_44228_n15415;
  wire u2__abc_44228_n15416;
  wire u2__abc_44228_n15417;
  wire u2__abc_44228_n15419_1;
  wire u2__abc_44228_n15420;
  wire u2__abc_44228_n15421;
  wire u2__abc_44228_n15422;
  wire u2__abc_44228_n15423;
  wire u2__abc_44228_n15425;
  wire u2__abc_44228_n15426;
  wire u2__abc_44228_n15427_1;
  wire u2__abc_44228_n15428;
  wire u2__abc_44228_n15429;
  wire u2__abc_44228_n15431;
  wire u2__abc_44228_n15432;
  wire u2__abc_44228_n15433;
  wire u2__abc_44228_n15434;
  wire u2__abc_44228_n15435_1;
  wire u2__abc_44228_n15436;
  wire u2__abc_44228_n15437;
  wire u2__abc_44228_n15439;
  wire u2__abc_44228_n15440;
  wire u2__abc_44228_n15441;
  wire u2__abc_44228_n15442_1;
  wire u2__abc_44228_n15443;
  wire u2__abc_44228_n15445;
  wire u2__abc_44228_n15446;
  wire u2__abc_44228_n15447;
  wire u2__abc_44228_n15448;
  wire u2__abc_44228_n15449;
  wire u2__abc_44228_n15451;
  wire u2__abc_44228_n15452;
  wire u2__abc_44228_n15453;
  wire u2__abc_44228_n15454;
  wire u2__abc_44228_n15455_1;
  wire u2__abc_44228_n15457;
  wire u2__abc_44228_n15458;
  wire u2__abc_44228_n15459;
  wire u2__abc_44228_n15460;
  wire u2__abc_44228_n15461;
  wire u2__abc_44228_n15463_1;
  wire u2__abc_44228_n15464;
  wire u2__abc_44228_n15465;
  wire u2__abc_44228_n15466;
  wire u2__abc_44228_n15467;
  wire u2__abc_44228_n15469;
  wire u2__abc_44228_n15470;
  wire u2__abc_44228_n15471;
  wire u2__abc_44228_n15472_1;
  wire u2__abc_44228_n15473_1;
  wire u2__abc_44228_n15475;
  wire u2__abc_44228_n15476;
  wire u2__abc_44228_n15477;
  wire u2__abc_44228_n15478;
  wire u2__abc_44228_n15479;
  wire u2__abc_44228_n15481_1;
  wire u2__abc_44228_n15482;
  wire u2__abc_44228_n15483;
  wire u2__abc_44228_n15484;
  wire u2__abc_44228_n15485;
  wire u2__abc_44228_n15487;
  wire u2__abc_44228_n15488;
  wire u2__abc_44228_n15489;
  wire u2__abc_44228_n15490;
  wire u2__abc_44228_n15491;
  wire u2__abc_44228_n15493;
  wire u2__abc_44228_n15494;
  wire u2__abc_44228_n15495;
  wire u2__abc_44228_n15496;
  wire u2__abc_44228_n15497;
  wire u2__abc_44228_n15499;
  wire u2__abc_44228_n15500;
  wire u2__abc_44228_n15501;
  wire u2__abc_44228_n15502;
  wire u2__abc_44228_n15503;
  wire u2__abc_44228_n15505;
  wire u2__abc_44228_n15506;
  wire u2__abc_44228_n15507;
  wire u2__abc_44228_n15508;
  wire u2__abc_44228_n15509;
  wire u2__abc_44228_n15511;
  wire u2__abc_44228_n15512;
  wire u2__abc_44228_n15513;
  wire u2__abc_44228_n15514;
  wire u2__abc_44228_n15515;
  wire u2__abc_44228_n15517;
  wire u2__abc_44228_n15518;
  wire u2__abc_44228_n15519;
  wire u2__abc_44228_n15520;
  wire u2__abc_44228_n15521;
  wire u2__abc_44228_n15523;
  wire u2__abc_44228_n15524;
  wire u2__abc_44228_n15525;
  wire u2__abc_44228_n15526;
  wire u2__abc_44228_n15527;
  wire u2__abc_44228_n15529;
  wire u2__abc_44228_n15530;
  wire u2__abc_44228_n15531;
  wire u2__abc_44228_n15532;
  wire u2__abc_44228_n15533;
  wire u2__abc_44228_n15535;
  wire u2__abc_44228_n15536;
  wire u2__abc_44228_n15537;
  wire u2__abc_44228_n15538;
  wire u2__abc_44228_n15539;
  wire u2__abc_44228_n15541;
  wire u2__abc_44228_n15542;
  wire u2__abc_44228_n15543;
  wire u2__abc_44228_n15544;
  wire u2__abc_44228_n15545;
  wire u2__abc_44228_n15546;
  wire u2__abc_44228_n15547;
  wire u2__abc_44228_n15549;
  wire u2__abc_44228_n15550;
  wire u2__abc_44228_n15551;
  wire u2__abc_44228_n15552;
  wire u2__abc_44228_n15553;
  wire u2__abc_44228_n15555;
  wire u2__abc_44228_n15556;
  wire u2__abc_44228_n15557;
  wire u2__abc_44228_n15558;
  wire u2__abc_44228_n15559;
  wire u2__abc_44228_n15561;
  wire u2__abc_44228_n15562;
  wire u2__abc_44228_n15563;
  wire u2__abc_44228_n15564;
  wire u2__abc_44228_n15565;
  wire u2__abc_44228_n15567;
  wire u2__abc_44228_n15568;
  wire u2__abc_44228_n15569;
  wire u2__abc_44228_n15570;
  wire u2__abc_44228_n15571;
  wire u2__abc_44228_n15573;
  wire u2__abc_44228_n15574;
  wire u2__abc_44228_n15575;
  wire u2__abc_44228_n15576;
  wire u2__abc_44228_n15577;
  wire u2__abc_44228_n15579;
  wire u2__abc_44228_n15580;
  wire u2__abc_44228_n15581;
  wire u2__abc_44228_n15582;
  wire u2__abc_44228_n15583;
  wire u2__abc_44228_n15585;
  wire u2__abc_44228_n15586;
  wire u2__abc_44228_n15587;
  wire u2__abc_44228_n15588;
  wire u2__abc_44228_n15589;
  wire u2__abc_44228_n15591;
  wire u2__abc_44228_n15592;
  wire u2__abc_44228_n15593;
  wire u2__abc_44228_n15594;
  wire u2__abc_44228_n15595;
  wire u2__abc_44228_n15597;
  wire u2__abc_44228_n15598;
  wire u2__abc_44228_n15599;
  wire u2__abc_44228_n15600;
  wire u2__abc_44228_n15601;
  wire u2__abc_44228_n15603;
  wire u2__abc_44228_n15604;
  wire u2__abc_44228_n15605;
  wire u2__abc_44228_n15606;
  wire u2__abc_44228_n15607;
  wire u2__abc_44228_n15609;
  wire u2__abc_44228_n15610;
  wire u2__abc_44228_n15611;
  wire u2__abc_44228_n15612;
  wire u2__abc_44228_n15613;
  wire u2__abc_44228_n15615;
  wire u2__abc_44228_n15616;
  wire u2__abc_44228_n15617;
  wire u2__abc_44228_n15618;
  wire u2__abc_44228_n15619;
  wire u2__abc_44228_n15621;
  wire u2__abc_44228_n15622;
  wire u2__abc_44228_n15623;
  wire u2__abc_44228_n15624;
  wire u2__abc_44228_n15625;
  wire u2__abc_44228_n15627;
  wire u2__abc_44228_n15628;
  wire u2__abc_44228_n15629;
  wire u2__abc_44228_n15630;
  wire u2__abc_44228_n15631;
  wire u2__abc_44228_n15633;
  wire u2__abc_44228_n15634;
  wire u2__abc_44228_n15635;
  wire u2__abc_44228_n15636;
  wire u2__abc_44228_n15637;
  wire u2__abc_44228_n15639;
  wire u2__abc_44228_n15640;
  wire u2__abc_44228_n15641;
  wire u2__abc_44228_n15642;
  wire u2__abc_44228_n15643;
  wire u2__abc_44228_n15645;
  wire u2__abc_44228_n15646;
  wire u2__abc_44228_n15647;
  wire u2__abc_44228_n15648;
  wire u2__abc_44228_n15649;
  wire u2__abc_44228_n15651;
  wire u2__abc_44228_n15652;
  wire u2__abc_44228_n15653;
  wire u2__abc_44228_n15654;
  wire u2__abc_44228_n15655;
  wire u2__abc_44228_n15657;
  wire u2__abc_44228_n15658;
  wire u2__abc_44228_n15659;
  wire u2__abc_44228_n15660;
  wire u2__abc_44228_n15661;
  wire u2__abc_44228_n15663;
  wire u2__abc_44228_n15664;
  wire u2__abc_44228_n15665;
  wire u2__abc_44228_n15666;
  wire u2__abc_44228_n15667;
  wire u2__abc_44228_n15669;
  wire u2__abc_44228_n15670;
  wire u2__abc_44228_n15671;
  wire u2__abc_44228_n15672;
  wire u2__abc_44228_n15673;
  wire u2__abc_44228_n15675;
  wire u2__abc_44228_n15676;
  wire u2__abc_44228_n15677;
  wire u2__abc_44228_n15678;
  wire u2__abc_44228_n15679;
  wire u2__abc_44228_n15681;
  wire u2__abc_44228_n15682;
  wire u2__abc_44228_n15683;
  wire u2__abc_44228_n15684;
  wire u2__abc_44228_n15685;
  wire u2__abc_44228_n15687;
  wire u2__abc_44228_n15688;
  wire u2__abc_44228_n15689;
  wire u2__abc_44228_n15690;
  wire u2__abc_44228_n15691;
  wire u2__abc_44228_n15693;
  wire u2__abc_44228_n15694;
  wire u2__abc_44228_n15695;
  wire u2__abc_44228_n15696;
  wire u2__abc_44228_n15697;
  wire u2__abc_44228_n15699;
  wire u2__abc_44228_n15700;
  wire u2__abc_44228_n15701;
  wire u2__abc_44228_n15702;
  wire u2__abc_44228_n15703;
  wire u2__abc_44228_n15705;
  wire u2__abc_44228_n15706;
  wire u2__abc_44228_n15707;
  wire u2__abc_44228_n15708;
  wire u2__abc_44228_n15709;
  wire u2__abc_44228_n15711;
  wire u2__abc_44228_n15712;
  wire u2__abc_44228_n15713;
  wire u2__abc_44228_n15714;
  wire u2__abc_44228_n15715;
  wire u2__abc_44228_n15717;
  wire u2__abc_44228_n15718;
  wire u2__abc_44228_n15719;
  wire u2__abc_44228_n15720;
  wire u2__abc_44228_n15721;
  wire u2__abc_44228_n15723;
  wire u2__abc_44228_n15724;
  wire u2__abc_44228_n15725;
  wire u2__abc_44228_n15726;
  wire u2__abc_44228_n15727;
  wire u2__abc_44228_n15729;
  wire u2__abc_44228_n15730;
  wire u2__abc_44228_n15731;
  wire u2__abc_44228_n15732;
  wire u2__abc_44228_n15733;
  wire u2__abc_44228_n15735;
  wire u2__abc_44228_n15736;
  wire u2__abc_44228_n15737;
  wire u2__abc_44228_n15738;
  wire u2__abc_44228_n15739;
  wire u2__abc_44228_n15740;
  wire u2__abc_44228_n15741;
  wire u2__abc_44228_n15743;
  wire u2__abc_44228_n15744;
  wire u2__abc_44228_n15745;
  wire u2__abc_44228_n15746;
  wire u2__abc_44228_n15747;
  wire u2__abc_44228_n15749;
  wire u2__abc_44228_n15750;
  wire u2__abc_44228_n15751;
  wire u2__abc_44228_n15752;
  wire u2__abc_44228_n15753;
  wire u2__abc_44228_n15755;
  wire u2__abc_44228_n15756;
  wire u2__abc_44228_n15757;
  wire u2__abc_44228_n15758;
  wire u2__abc_44228_n15759;
  wire u2__abc_44228_n15761;
  wire u2__abc_44228_n15762;
  wire u2__abc_44228_n15763;
  wire u2__abc_44228_n15764;
  wire u2__abc_44228_n15765;
  wire u2__abc_44228_n15766;
  wire u2__abc_44228_n15767;
  wire u2__abc_44228_n15769;
  wire u2__abc_44228_n15770;
  wire u2__abc_44228_n15771;
  wire u2__abc_44228_n15772;
  wire u2__abc_44228_n15773;
  wire u2__abc_44228_n15775;
  wire u2__abc_44228_n15776;
  wire u2__abc_44228_n15777;
  wire u2__abc_44228_n15778;
  wire u2__abc_44228_n15779;
  wire u2__abc_44228_n15781;
  wire u2__abc_44228_n15782;
  wire u2__abc_44228_n15783;
  wire u2__abc_44228_n15784;
  wire u2__abc_44228_n15785;
  wire u2__abc_44228_n15787;
  wire u2__abc_44228_n15788;
  wire u2__abc_44228_n15789;
  wire u2__abc_44228_n15790;
  wire u2__abc_44228_n15791;
  wire u2__abc_44228_n15793;
  wire u2__abc_44228_n15794;
  wire u2__abc_44228_n15795;
  wire u2__abc_44228_n15796;
  wire u2__abc_44228_n15797;
  wire u2__abc_44228_n15799;
  wire u2__abc_44228_n15800;
  wire u2__abc_44228_n15801;
  wire u2__abc_44228_n15802;
  wire u2__abc_44228_n15803;
  wire u2__abc_44228_n15805;
  wire u2__abc_44228_n15806;
  wire u2__abc_44228_n15807;
  wire u2__abc_44228_n15808;
  wire u2__abc_44228_n15809;
  wire u2__abc_44228_n15811;
  wire u2__abc_44228_n15812;
  wire u2__abc_44228_n15813;
  wire u2__abc_44228_n15814;
  wire u2__abc_44228_n15815;
  wire u2__abc_44228_n15817;
  wire u2__abc_44228_n15818;
  wire u2__abc_44228_n15819;
  wire u2__abc_44228_n15820;
  wire u2__abc_44228_n15821;
  wire u2__abc_44228_n15823;
  wire u2__abc_44228_n15824;
  wire u2__abc_44228_n15825;
  wire u2__abc_44228_n15826;
  wire u2__abc_44228_n15827;
  wire u2__abc_44228_n15829;
  wire u2__abc_44228_n15830;
  wire u2__abc_44228_n15831;
  wire u2__abc_44228_n15832;
  wire u2__abc_44228_n15833;
  wire u2__abc_44228_n15835;
  wire u2__abc_44228_n15836;
  wire u2__abc_44228_n15837;
  wire u2__abc_44228_n15838;
  wire u2__abc_44228_n15839;
  wire u2__abc_44228_n15841;
  wire u2__abc_44228_n15842;
  wire u2__abc_44228_n15843;
  wire u2__abc_44228_n15844;
  wire u2__abc_44228_n15845;
  wire u2__abc_44228_n15847;
  wire u2__abc_44228_n15848;
  wire u2__abc_44228_n15849;
  wire u2__abc_44228_n15850;
  wire u2__abc_44228_n15851;
  wire u2__abc_44228_n15853;
  wire u2__abc_44228_n15854;
  wire u2__abc_44228_n15855;
  wire u2__abc_44228_n15856;
  wire u2__abc_44228_n15857;
  wire u2__abc_44228_n15859;
  wire u2__abc_44228_n15860;
  wire u2__abc_44228_n15861;
  wire u2__abc_44228_n15862;
  wire u2__abc_44228_n15863;
  wire u2__abc_44228_n15865;
  wire u2__abc_44228_n15866;
  wire u2__abc_44228_n15867;
  wire u2__abc_44228_n15868;
  wire u2__abc_44228_n15869;
  wire u2__abc_44228_n15871;
  wire u2__abc_44228_n15872;
  wire u2__abc_44228_n15873;
  wire u2__abc_44228_n15874;
  wire u2__abc_44228_n15875;
  wire u2__abc_44228_n15877;
  wire u2__abc_44228_n15878;
  wire u2__abc_44228_n15879;
  wire u2__abc_44228_n15880;
  wire u2__abc_44228_n15881;
  wire u2__abc_44228_n15883;
  wire u2__abc_44228_n15884;
  wire u2__abc_44228_n15885;
  wire u2__abc_44228_n15886;
  wire u2__abc_44228_n15887;
  wire u2__abc_44228_n15889;
  wire u2__abc_44228_n15890;
  wire u2__abc_44228_n15891;
  wire u2__abc_44228_n15892;
  wire u2__abc_44228_n15893;
  wire u2__abc_44228_n15895;
  wire u2__abc_44228_n15896;
  wire u2__abc_44228_n15897;
  wire u2__abc_44228_n15898;
  wire u2__abc_44228_n15899;
  wire u2__abc_44228_n15901;
  wire u2__abc_44228_n15902;
  wire u2__abc_44228_n15903;
  wire u2__abc_44228_n15904;
  wire u2__abc_44228_n15905;
  wire u2__abc_44228_n15907;
  wire u2__abc_44228_n15908;
  wire u2__abc_44228_n15909;
  wire u2__abc_44228_n15910;
  wire u2__abc_44228_n15911;
  wire u2__abc_44228_n15913;
  wire u2__abc_44228_n15914;
  wire u2__abc_44228_n15915;
  wire u2__abc_44228_n15916;
  wire u2__abc_44228_n15917;
  wire u2__abc_44228_n15919;
  wire u2__abc_44228_n15920;
  wire u2__abc_44228_n15921;
  wire u2__abc_44228_n15922;
  wire u2__abc_44228_n15923;
  wire u2__abc_44228_n15925;
  wire u2__abc_44228_n15926;
  wire u2__abc_44228_n15927;
  wire u2__abc_44228_n15928;
  wire u2__abc_44228_n15929;
  wire u2__abc_44228_n15931;
  wire u2__abc_44228_n15932;
  wire u2__abc_44228_n15933;
  wire u2__abc_44228_n15934;
  wire u2__abc_44228_n15935;
  wire u2__abc_44228_n15936;
  wire u2__abc_44228_n15937;
  wire u2__abc_44228_n15939;
  wire u2__abc_44228_n15940;
  wire u2__abc_44228_n15941;
  wire u2__abc_44228_n15942;
  wire u2__abc_44228_n15943;
  wire u2__abc_44228_n15945;
  wire u2__abc_44228_n15946;
  wire u2__abc_44228_n15947;
  wire u2__abc_44228_n15948;
  wire u2__abc_44228_n15949;
  wire u2__abc_44228_n15951;
  wire u2__abc_44228_n15952;
  wire u2__abc_44228_n15953;
  wire u2__abc_44228_n15954;
  wire u2__abc_44228_n15955;
  wire u2__abc_44228_n15957;
  wire u2__abc_44228_n15958;
  wire u2__abc_44228_n15959;
  wire u2__abc_44228_n15960;
  wire u2__abc_44228_n15961;
  wire u2__abc_44228_n15963;
  wire u2__abc_44228_n15964;
  wire u2__abc_44228_n15965;
  wire u2__abc_44228_n15966;
  wire u2__abc_44228_n15967;
  wire u2__abc_44228_n15969;
  wire u2__abc_44228_n15970;
  wire u2__abc_44228_n15971;
  wire u2__abc_44228_n15972;
  wire u2__abc_44228_n15973;
  wire u2__abc_44228_n15975;
  wire u2__abc_44228_n15976;
  wire u2__abc_44228_n15977;
  wire u2__abc_44228_n15978;
  wire u2__abc_44228_n15979;
  wire u2__abc_44228_n15981;
  wire u2__abc_44228_n15982;
  wire u2__abc_44228_n15983;
  wire u2__abc_44228_n15984;
  wire u2__abc_44228_n15985;
  wire u2__abc_44228_n15987;
  wire u2__abc_44228_n15988;
  wire u2__abc_44228_n15989;
  wire u2__abc_44228_n15990;
  wire u2__abc_44228_n15991;
  wire u2__abc_44228_n15992;
  wire u2__abc_44228_n15993;
  wire u2__abc_44228_n15995;
  wire u2__abc_44228_n15996;
  wire u2__abc_44228_n15997;
  wire u2__abc_44228_n15998;
  wire u2__abc_44228_n15999;
  wire u2__abc_44228_n16001;
  wire u2__abc_44228_n16002;
  wire u2__abc_44228_n16003;
  wire u2__abc_44228_n16004;
  wire u2__abc_44228_n16005;
  wire u2__abc_44228_n16007;
  wire u2__abc_44228_n16008;
  wire u2__abc_44228_n16009;
  wire u2__abc_44228_n16010;
  wire u2__abc_44228_n16011;
  wire u2__abc_44228_n16013;
  wire u2__abc_44228_n16014;
  wire u2__abc_44228_n16015;
  wire u2__abc_44228_n16016;
  wire u2__abc_44228_n16017;
  wire u2__abc_44228_n16019;
  wire u2__abc_44228_n16020;
  wire u2__abc_44228_n16021;
  wire u2__abc_44228_n16022;
  wire u2__abc_44228_n16023;
  wire u2__abc_44228_n16025;
  wire u2__abc_44228_n16026;
  wire u2__abc_44228_n16027;
  wire u2__abc_44228_n16028;
  wire u2__abc_44228_n16029;
  wire u2__abc_44228_n16031;
  wire u2__abc_44228_n16032;
  wire u2__abc_44228_n16033;
  wire u2__abc_44228_n16034;
  wire u2__abc_44228_n16035;
  wire u2__abc_44228_n16037;
  wire u2__abc_44228_n16038;
  wire u2__abc_44228_n16039;
  wire u2__abc_44228_n16040;
  wire u2__abc_44228_n16041;
  wire u2__abc_44228_n16043;
  wire u2__abc_44228_n16044;
  wire u2__abc_44228_n16045;
  wire u2__abc_44228_n16046;
  wire u2__abc_44228_n16047;
  wire u2__abc_44228_n16049;
  wire u2__abc_44228_n16050;
  wire u2__abc_44228_n16051;
  wire u2__abc_44228_n16052;
  wire u2__abc_44228_n16053;
  wire u2__abc_44228_n16055;
  wire u2__abc_44228_n16056;
  wire u2__abc_44228_n16057;
  wire u2__abc_44228_n16058;
  wire u2__abc_44228_n16059;
  wire u2__abc_44228_n16061;
  wire u2__abc_44228_n16062;
  wire u2__abc_44228_n16063;
  wire u2__abc_44228_n16064;
  wire u2__abc_44228_n16065;
  wire u2__abc_44228_n16067;
  wire u2__abc_44228_n16068;
  wire u2__abc_44228_n16069;
  wire u2__abc_44228_n16070;
  wire u2__abc_44228_n16071;
  wire u2__abc_44228_n16073;
  wire u2__abc_44228_n16074;
  wire u2__abc_44228_n16075;
  wire u2__abc_44228_n16076;
  wire u2__abc_44228_n16077;
  wire u2__abc_44228_n16079;
  wire u2__abc_44228_n16080;
  wire u2__abc_44228_n16081;
  wire u2__abc_44228_n16082;
  wire u2__abc_44228_n16083;
  wire u2__abc_44228_n16085;
  wire u2__abc_44228_n16086;
  wire u2__abc_44228_n16087;
  wire u2__abc_44228_n16088;
  wire u2__abc_44228_n16089;
  wire u2__abc_44228_n16091;
  wire u2__abc_44228_n16092;
  wire u2__abc_44228_n16093;
  wire u2__abc_44228_n16094;
  wire u2__abc_44228_n16095;
  wire u2__abc_44228_n16097;
  wire u2__abc_44228_n16098;
  wire u2__abc_44228_n16099;
  wire u2__abc_44228_n16100;
  wire u2__abc_44228_n16101;
  wire u2__abc_44228_n16102;
  wire u2__abc_44228_n16103;
  wire u2__abc_44228_n16105;
  wire u2__abc_44228_n16106;
  wire u2__abc_44228_n16107;
  wire u2__abc_44228_n16108;
  wire u2__abc_44228_n16109;
  wire u2__abc_44228_n16110;
  wire u2__abc_44228_n16111;
  wire u2__abc_44228_n16113;
  wire u2__abc_44228_n16114;
  wire u2__abc_44228_n16115;
  wire u2__abc_44228_n16116;
  wire u2__abc_44228_n16117;
  wire u2__abc_44228_n16119;
  wire u2__abc_44228_n16120;
  wire u2__abc_44228_n16121;
  wire u2__abc_44228_n16122;
  wire u2__abc_44228_n16123;
  wire u2__abc_44228_n16125;
  wire u2__abc_44228_n16126;
  wire u2__abc_44228_n16127;
  wire u2__abc_44228_n16128;
  wire u2__abc_44228_n16129;
  wire u2__abc_44228_n16131;
  wire u2__abc_44228_n16132;
  wire u2__abc_44228_n16133;
  wire u2__abc_44228_n16134;
  wire u2__abc_44228_n16135;
  wire u2__abc_44228_n16136;
  wire u2__abc_44228_n16137;
  wire u2__abc_44228_n16139;
  wire u2__abc_44228_n16140;
  wire u2__abc_44228_n16141;
  wire u2__abc_44228_n16142;
  wire u2__abc_44228_n16143;
  wire u2__abc_44228_n16145;
  wire u2__abc_44228_n16146;
  wire u2__abc_44228_n16147;
  wire u2__abc_44228_n16148;
  wire u2__abc_44228_n16149;
  wire u2__abc_44228_n16151;
  wire u2__abc_44228_n16152;
  wire u2__abc_44228_n16153;
  wire u2__abc_44228_n16154;
  wire u2__abc_44228_n16155;
  wire u2__abc_44228_n16157;
  wire u2__abc_44228_n16158;
  wire u2__abc_44228_n16159;
  wire u2__abc_44228_n16160;
  wire u2__abc_44228_n16161;
  wire u2__abc_44228_n16163;
  wire u2__abc_44228_n16164;
  wire u2__abc_44228_n16165;
  wire u2__abc_44228_n16166;
  wire u2__abc_44228_n16167;
  wire u2__abc_44228_n16169;
  wire u2__abc_44228_n16170;
  wire u2__abc_44228_n16171;
  wire u2__abc_44228_n16172;
  wire u2__abc_44228_n16173;
  wire u2__abc_44228_n16175;
  wire u2__abc_44228_n16176;
  wire u2__abc_44228_n16177;
  wire u2__abc_44228_n16178;
  wire u2__abc_44228_n16179;
  wire u2__abc_44228_n16181;
  wire u2__abc_44228_n16182;
  wire u2__abc_44228_n16183;
  wire u2__abc_44228_n16184;
  wire u2__abc_44228_n16185;
  wire u2__abc_44228_n16187;
  wire u2__abc_44228_n16188;
  wire u2__abc_44228_n16189;
  wire u2__abc_44228_n16190;
  wire u2__abc_44228_n16191;
  wire u2__abc_44228_n16193;
  wire u2__abc_44228_n16194;
  wire u2__abc_44228_n16195;
  wire u2__abc_44228_n16196;
  wire u2__abc_44228_n16197;
  wire u2__abc_44228_n16199;
  wire u2__abc_44228_n16200;
  wire u2__abc_44228_n16201;
  wire u2__abc_44228_n16202;
  wire u2__abc_44228_n16203;
  wire u2__abc_44228_n16205;
  wire u2__abc_44228_n16206;
  wire u2__abc_44228_n16207;
  wire u2__abc_44228_n16208;
  wire u2__abc_44228_n16209;
  wire u2__abc_44228_n16211;
  wire u2__abc_44228_n16212;
  wire u2__abc_44228_n16213;
  wire u2__abc_44228_n16214;
  wire u2__abc_44228_n16215;
  wire u2__abc_44228_n16217;
  wire u2__abc_44228_n16218;
  wire u2__abc_44228_n16219;
  wire u2__abc_44228_n16220;
  wire u2__abc_44228_n16221;
  wire u2__abc_44228_n16223;
  wire u2__abc_44228_n16224;
  wire u2__abc_44228_n16225;
  wire u2__abc_44228_n16226;
  wire u2__abc_44228_n16227;
  wire u2__abc_44228_n16229;
  wire u2__abc_44228_n16230;
  wire u2__abc_44228_n16231;
  wire u2__abc_44228_n16232;
  wire u2__abc_44228_n16233;
  wire u2__abc_44228_n16235;
  wire u2__abc_44228_n16236;
  wire u2__abc_44228_n16237;
  wire u2__abc_44228_n16238;
  wire u2__abc_44228_n16239;
  wire u2__abc_44228_n16241;
  wire u2__abc_44228_n16242;
  wire u2__abc_44228_n16243;
  wire u2__abc_44228_n16244;
  wire u2__abc_44228_n16245;
  wire u2__abc_44228_n16247;
  wire u2__abc_44228_n16248;
  wire u2__abc_44228_n16249;
  wire u2__abc_44228_n16250;
  wire u2__abc_44228_n16251;
  wire u2__abc_44228_n16253;
  wire u2__abc_44228_n16254;
  wire u2__abc_44228_n16255;
  wire u2__abc_44228_n16256;
  wire u2__abc_44228_n16257;
  wire u2__abc_44228_n16259;
  wire u2__abc_44228_n16260;
  wire u2__abc_44228_n16261;
  wire u2__abc_44228_n16262;
  wire u2__abc_44228_n16263;
  wire u2__abc_44228_n16265;
  wire u2__abc_44228_n16266;
  wire u2__abc_44228_n16267;
  wire u2__abc_44228_n16268;
  wire u2__abc_44228_n16269;
  wire u2__abc_44228_n16271;
  wire u2__abc_44228_n16272;
  wire u2__abc_44228_n16273;
  wire u2__abc_44228_n16274;
  wire u2__abc_44228_n16275;
  wire u2__abc_44228_n16277;
  wire u2__abc_44228_n16278;
  wire u2__abc_44228_n16279;
  wire u2__abc_44228_n16280;
  wire u2__abc_44228_n16281;
  wire u2__abc_44228_n16283;
  wire u2__abc_44228_n16284;
  wire u2__abc_44228_n16285;
  wire u2__abc_44228_n16286;
  wire u2__abc_44228_n16287;
  wire u2__abc_44228_n16288;
  wire u2__abc_44228_n16289;
  wire u2__abc_44228_n16291;
  wire u2__abc_44228_n16292;
  wire u2__abc_44228_n16293;
  wire u2__abc_44228_n16294;
  wire u2__abc_44228_n16295;
  wire u2__abc_44228_n16297;
  wire u2__abc_44228_n16298;
  wire u2__abc_44228_n16299;
  wire u2__abc_44228_n16300;
  wire u2__abc_44228_n16301;
  wire u2__abc_44228_n16302;
  wire u2__abc_44228_n16303;
  wire u2__abc_44228_n16305;
  wire u2__abc_44228_n16306;
  wire u2__abc_44228_n16307;
  wire u2__abc_44228_n16308;
  wire u2__abc_44228_n16309;
  wire u2__abc_44228_n16310;
  wire u2__abc_44228_n16311;
  wire u2__abc_44228_n16313;
  wire u2__abc_44228_n16314;
  wire u2__abc_44228_n16315;
  wire u2__abc_44228_n16316;
  wire u2__abc_44228_n16317;
  wire u2__abc_44228_n16319;
  wire u2__abc_44228_n16320;
  wire u2__abc_44228_n16321;
  wire u2__abc_44228_n16322;
  wire u2__abc_44228_n16323;
  wire u2__abc_44228_n16325;
  wire u2__abc_44228_n16326;
  wire u2__abc_44228_n16327;
  wire u2__abc_44228_n16328;
  wire u2__abc_44228_n16329;
  wire u2__abc_44228_n16331;
  wire u2__abc_44228_n16332;
  wire u2__abc_44228_n16333;
  wire u2__abc_44228_n16334;
  wire u2__abc_44228_n16335;
  wire u2__abc_44228_n16336;
  wire u2__abc_44228_n16337;
  wire u2__abc_44228_n16339;
  wire u2__abc_44228_n16340;
  wire u2__abc_44228_n16341;
  wire u2__abc_44228_n16342;
  wire u2__abc_44228_n16343;
  wire u2__abc_44228_n16345;
  wire u2__abc_44228_n16346;
  wire u2__abc_44228_n16347;
  wire u2__abc_44228_n16348;
  wire u2__abc_44228_n16349;
  wire u2__abc_44228_n16351;
  wire u2__abc_44228_n16352;
  wire u2__abc_44228_n16353;
  wire u2__abc_44228_n16354;
  wire u2__abc_44228_n16355;
  wire u2__abc_44228_n16357;
  wire u2__abc_44228_n16358;
  wire u2__abc_44228_n16359;
  wire u2__abc_44228_n16360;
  wire u2__abc_44228_n16361;
  wire u2__abc_44228_n16363;
  wire u2__abc_44228_n16364;
  wire u2__abc_44228_n16365;
  wire u2__abc_44228_n16366;
  wire u2__abc_44228_n16367;
  wire u2__abc_44228_n16369;
  wire u2__abc_44228_n16370;
  wire u2__abc_44228_n16371;
  wire u2__abc_44228_n16372;
  wire u2__abc_44228_n16373;
  wire u2__abc_44228_n16375;
  wire u2__abc_44228_n16376;
  wire u2__abc_44228_n16377;
  wire u2__abc_44228_n16378;
  wire u2__abc_44228_n16379;
  wire u2__abc_44228_n16381;
  wire u2__abc_44228_n16382;
  wire u2__abc_44228_n16383;
  wire u2__abc_44228_n16384;
  wire u2__abc_44228_n16385;
  wire u2__abc_44228_n16387;
  wire u2__abc_44228_n16388;
  wire u2__abc_44228_n16389;
  wire u2__abc_44228_n16390;
  wire u2__abc_44228_n16391;
  wire u2__abc_44228_n16393;
  wire u2__abc_44228_n16394;
  wire u2__abc_44228_n16395;
  wire u2__abc_44228_n16396;
  wire u2__abc_44228_n16397;
  wire u2__abc_44228_n16399;
  wire u2__abc_44228_n16400;
  wire u2__abc_44228_n16401;
  wire u2__abc_44228_n16402;
  wire u2__abc_44228_n16403;
  wire u2__abc_44228_n16405;
  wire u2__abc_44228_n16406;
  wire u2__abc_44228_n16407;
  wire u2__abc_44228_n16408;
  wire u2__abc_44228_n16409;
  wire u2__abc_44228_n16411;
  wire u2__abc_44228_n16412;
  wire u2__abc_44228_n16413;
  wire u2__abc_44228_n16414;
  wire u2__abc_44228_n16415;
  wire u2__abc_44228_n16417;
  wire u2__abc_44228_n16418;
  wire u2__abc_44228_n16419;
  wire u2__abc_44228_n16420;
  wire u2__abc_44228_n16421;
  wire u2__abc_44228_n16423;
  wire u2__abc_44228_n16424;
  wire u2__abc_44228_n16425;
  wire u2__abc_44228_n16426;
  wire u2__abc_44228_n16427;
  wire u2__abc_44228_n16429;
  wire u2__abc_44228_n16430;
  wire u2__abc_44228_n16431;
  wire u2__abc_44228_n16432;
  wire u2__abc_44228_n16433;
  wire u2__abc_44228_n16435;
  wire u2__abc_44228_n16436;
  wire u2__abc_44228_n16437;
  wire u2__abc_44228_n16438;
  wire u2__abc_44228_n16439;
  wire u2__abc_44228_n16441;
  wire u2__abc_44228_n16442;
  wire u2__abc_44228_n16443;
  wire u2__abc_44228_n16444;
  wire u2__abc_44228_n16445;
  wire u2__abc_44228_n16447;
  wire u2__abc_44228_n16448;
  wire u2__abc_44228_n16449;
  wire u2__abc_44228_n16450;
  wire u2__abc_44228_n16451;
  wire u2__abc_44228_n16453;
  wire u2__abc_44228_n16454;
  wire u2__abc_44228_n16455;
  wire u2__abc_44228_n16456;
  wire u2__abc_44228_n16457;
  wire u2__abc_44228_n16459;
  wire u2__abc_44228_n16460;
  wire u2__abc_44228_n16461;
  wire u2__abc_44228_n16462;
  wire u2__abc_44228_n16463;
  wire u2__abc_44228_n16465;
  wire u2__abc_44228_n16466;
  wire u2__abc_44228_n16467;
  wire u2__abc_44228_n16468;
  wire u2__abc_44228_n16469;
  wire u2__abc_44228_n16471;
  wire u2__abc_44228_n16472;
  wire u2__abc_44228_n16473;
  wire u2__abc_44228_n16474;
  wire u2__abc_44228_n16475;
  wire u2__abc_44228_n16477;
  wire u2__abc_44228_n16478;
  wire u2__abc_44228_n16479;
  wire u2__abc_44228_n16480;
  wire u2__abc_44228_n16481;
  wire u2__abc_44228_n16483;
  wire u2__abc_44228_n16484;
  wire u2__abc_44228_n16485;
  wire u2__abc_44228_n16486;
  wire u2__abc_44228_n16487;
  wire u2__abc_44228_n16489;
  wire u2__abc_44228_n16490;
  wire u2__abc_44228_n16491;
  wire u2__abc_44228_n16492;
  wire u2__abc_44228_n16493;
  wire u2__abc_44228_n16495;
  wire u2__abc_44228_n16496;
  wire u2__abc_44228_n16497;
  wire u2__abc_44228_n16498;
  wire u2__abc_44228_n16499;
  wire u2__abc_44228_n16501;
  wire u2__abc_44228_n16502;
  wire u2__abc_44228_n16503;
  wire u2__abc_44228_n16504;
  wire u2__abc_44228_n16505;
  wire u2__abc_44228_n16506;
  wire u2__abc_44228_n16507;
  wire u2__abc_44228_n16509;
  wire u2__abc_44228_n16510;
  wire u2__abc_44228_n16511;
  wire u2__abc_44228_n16512;
  wire u2__abc_44228_n16513;
  wire u2__abc_44228_n16515;
  wire u2__abc_44228_n16516;
  wire u2__abc_44228_n16517;
  wire u2__abc_44228_n16518;
  wire u2__abc_44228_n16519;
  wire u2__abc_44228_n16521;
  wire u2__abc_44228_n16522;
  wire u2__abc_44228_n16523;
  wire u2__abc_44228_n16524;
  wire u2__abc_44228_n16525;
  wire u2__abc_44228_n16527;
  wire u2__abc_44228_n16528;
  wire u2__abc_44228_n16529;
  wire u2__abc_44228_n16530;
  wire u2__abc_44228_n16531;
  wire u2__abc_44228_n16532;
  wire u2__abc_44228_n16533;
  wire u2__abc_44228_n16535;
  wire u2__abc_44228_n16536;
  wire u2__abc_44228_n16537;
  wire u2__abc_44228_n16538;
  wire u2__abc_44228_n16539;
  wire u2__abc_44228_n16541;
  wire u2__abc_44228_n16542;
  wire u2__abc_44228_n16543;
  wire u2__abc_44228_n16544;
  wire u2__abc_44228_n16545;
  wire u2__abc_44228_n16547;
  wire u2__abc_44228_n16548;
  wire u2__abc_44228_n16549;
  wire u2__abc_44228_n16550;
  wire u2__abc_44228_n16551;
  wire u2__abc_44228_n16553;
  wire u2__abc_44228_n16554;
  wire u2__abc_44228_n16555;
  wire u2__abc_44228_n16556;
  wire u2__abc_44228_n16557;
  wire u2__abc_44228_n16558;
  wire u2__abc_44228_n16559;
  wire u2__abc_44228_n16561;
  wire u2__abc_44228_n16562;
  wire u2__abc_44228_n16563;
  wire u2__abc_44228_n16564;
  wire u2__abc_44228_n16565;
  wire u2__abc_44228_n16567;
  wire u2__abc_44228_n16568;
  wire u2__abc_44228_n16569;
  wire u2__abc_44228_n16570;
  wire u2__abc_44228_n16571;
  wire u2__abc_44228_n16573;
  wire u2__abc_44228_n16574;
  wire u2__abc_44228_n16575;
  wire u2__abc_44228_n16576;
  wire u2__abc_44228_n16577;
  wire u2__abc_44228_n16579;
  wire u2__abc_44228_n16580;
  wire u2__abc_44228_n16581;
  wire u2__abc_44228_n16582;
  wire u2__abc_44228_n16583;
  wire u2__abc_44228_n16584;
  wire u2__abc_44228_n16585;
  wire u2__abc_44228_n16587;
  wire u2__abc_44228_n16588;
  wire u2__abc_44228_n16589;
  wire u2__abc_44228_n16590;
  wire u2__abc_44228_n16591;
  wire u2__abc_44228_n16593;
  wire u2__abc_44228_n16594;
  wire u2__abc_44228_n16595;
  wire u2__abc_44228_n16596;
  wire u2__abc_44228_n16597;
  wire u2__abc_44228_n16599;
  wire u2__abc_44228_n16600;
  wire u2__abc_44228_n16601;
  wire u2__abc_44228_n16602;
  wire u2__abc_44228_n16603;
  wire u2__abc_44228_n16605;
  wire u2__abc_44228_n16606;
  wire u2__abc_44228_n16607;
  wire u2__abc_44228_n16608;
  wire u2__abc_44228_n16609;
  wire u2__abc_44228_n16611;
  wire u2__abc_44228_n16612;
  wire u2__abc_44228_n16613;
  wire u2__abc_44228_n16614;
  wire u2__abc_44228_n16615;
  wire u2__abc_44228_n16617;
  wire u2__abc_44228_n16618;
  wire u2__abc_44228_n16619;
  wire u2__abc_44228_n16620;
  wire u2__abc_44228_n16621;
  wire u2__abc_44228_n16623;
  wire u2__abc_44228_n16624;
  wire u2__abc_44228_n16625;
  wire u2__abc_44228_n16626;
  wire u2__abc_44228_n16627;
  wire u2__abc_44228_n16629;
  wire u2__abc_44228_n16630;
  wire u2__abc_44228_n16631;
  wire u2__abc_44228_n16632;
  wire u2__abc_44228_n16633;
  wire u2__abc_44228_n16635;
  wire u2__abc_44228_n16636;
  wire u2__abc_44228_n16637;
  wire u2__abc_44228_n16638;
  wire u2__abc_44228_n16639;
  wire u2__abc_44228_n16641;
  wire u2__abc_44228_n16642;
  wire u2__abc_44228_n16643;
  wire u2__abc_44228_n16644;
  wire u2__abc_44228_n16645;
  wire u2__abc_44228_n16647;
  wire u2__abc_44228_n16648;
  wire u2__abc_44228_n16649;
  wire u2__abc_44228_n16650;
  wire u2__abc_44228_n16651;
  wire u2__abc_44228_n16653;
  wire u2__abc_44228_n16654;
  wire u2__abc_44228_n16655;
  wire u2__abc_44228_n16656;
  wire u2__abc_44228_n16657;
  wire u2__abc_44228_n16659;
  wire u2__abc_44228_n16660;
  wire u2__abc_44228_n16661;
  wire u2__abc_44228_n16662;
  wire u2__abc_44228_n16663;
  wire u2__abc_44228_n16665;
  wire u2__abc_44228_n16666;
  wire u2__abc_44228_n16667;
  wire u2__abc_44228_n16668;
  wire u2__abc_44228_n16669;
  wire u2__abc_44228_n16671;
  wire u2__abc_44228_n16672;
  wire u2__abc_44228_n16673;
  wire u2__abc_44228_n16674;
  wire u2__abc_44228_n16675;
  wire u2__abc_44228_n16677;
  wire u2__abc_44228_n16678;
  wire u2__abc_44228_n16679;
  wire u2__abc_44228_n16680;
  wire u2__abc_44228_n16681;
  wire u2__abc_44228_n16683;
  wire u2__abc_44228_n16684;
  wire u2__abc_44228_n16685;
  wire u2__abc_44228_n16686;
  wire u2__abc_44228_n16687;
  wire u2__abc_44228_n16689;
  wire u2__abc_44228_n16690;
  wire u2__abc_44228_n16691;
  wire u2__abc_44228_n16692;
  wire u2__abc_44228_n16693;
  wire u2__abc_44228_n16695;
  wire u2__abc_44228_n16696;
  wire u2__abc_44228_n16697;
  wire u2__abc_44228_n16698;
  wire u2__abc_44228_n16699;
  wire u2__abc_44228_n16701;
  wire u2__abc_44228_n16702;
  wire u2__abc_44228_n16703;
  wire u2__abc_44228_n16704;
  wire u2__abc_44228_n16705;
  wire u2__abc_44228_n16706;
  wire u2__abc_44228_n16707;
  wire u2__abc_44228_n16709;
  wire u2__abc_44228_n16710;
  wire u2__abc_44228_n16711;
  wire u2__abc_44228_n16712;
  wire u2__abc_44228_n16713;
  wire u2__abc_44228_n16715;
  wire u2__abc_44228_n16716;
  wire u2__abc_44228_n16717;
  wire u2__abc_44228_n16718;
  wire u2__abc_44228_n16719;
  wire u2__abc_44228_n16721;
  wire u2__abc_44228_n16722;
  wire u2__abc_44228_n16723;
  wire u2__abc_44228_n16724;
  wire u2__abc_44228_n16725;
  wire u2__abc_44228_n16727;
  wire u2__abc_44228_n16728;
  wire u2__abc_44228_n16729;
  wire u2__abc_44228_n16730;
  wire u2__abc_44228_n16731;
  wire u2__abc_44228_n16732;
  wire u2__abc_44228_n16733;
  wire u2__abc_44228_n16735;
  wire u2__abc_44228_n16736;
  wire u2__abc_44228_n16737;
  wire u2__abc_44228_n16738;
  wire u2__abc_44228_n16739;
  wire u2__abc_44228_n16741;
  wire u2__abc_44228_n16742;
  wire u2__abc_44228_n16743;
  wire u2__abc_44228_n16744;
  wire u2__abc_44228_n16745;
  wire u2__abc_44228_n16747;
  wire u2__abc_44228_n16748;
  wire u2__abc_44228_n16749;
  wire u2__abc_44228_n16750;
  wire u2__abc_44228_n16751;
  wire u2__abc_44228_n16753;
  wire u2__abc_44228_n16754;
  wire u2__abc_44228_n16755;
  wire u2__abc_44228_n16756;
  wire u2__abc_44228_n16757;
  wire u2__abc_44228_n16759;
  wire u2__abc_44228_n16760;
  wire u2__abc_44228_n16761;
  wire u2__abc_44228_n16762;
  wire u2__abc_44228_n16763;
  wire u2__abc_44228_n16764;
  wire u2__abc_44228_n16765;
  wire u2__abc_44228_n16767;
  wire u2__abc_44228_n16768;
  wire u2__abc_44228_n16769;
  wire u2__abc_44228_n16770;
  wire u2__abc_44228_n16771;
  wire u2__abc_44228_n16773;
  wire u2__abc_44228_n16774;
  wire u2__abc_44228_n16775;
  wire u2__abc_44228_n16776;
  wire u2__abc_44228_n16777;
  wire u2__abc_44228_n16779;
  wire u2__abc_44228_n16780;
  wire u2__abc_44228_n16781;
  wire u2__abc_44228_n16782;
  wire u2__abc_44228_n16783;
  wire u2__abc_44228_n16785;
  wire u2__abc_44228_n16786;
  wire u2__abc_44228_n16787;
  wire u2__abc_44228_n16788;
  wire u2__abc_44228_n16789;
  wire u2__abc_44228_n16791;
  wire u2__abc_44228_n16792;
  wire u2__abc_44228_n16793;
  wire u2__abc_44228_n16794;
  wire u2__abc_44228_n16795;
  wire u2__abc_44228_n16797;
  wire u2__abc_44228_n16798;
  wire u2__abc_44228_n16799;
  wire u2__abc_44228_n16800;
  wire u2__abc_44228_n16801;
  wire u2__abc_44228_n16803;
  wire u2__abc_44228_n16804;
  wire u2__abc_44228_n16805;
  wire u2__abc_44228_n16806;
  wire u2__abc_44228_n16808;
  wire u2__abc_44228_n16809;
  wire u2__abc_44228_n16810;
  wire u2__abc_44228_n16811;
  wire u2__abc_44228_n16813;
  wire u2__abc_44228_n16814;
  wire u2__abc_44228_n16815;
  wire u2__abc_44228_n16816;
  wire u2__abc_44228_n16818;
  wire u2__abc_44228_n16819;
  wire u2__abc_44228_n16820;
  wire u2__abc_44228_n16821;
  wire u2__abc_44228_n16823;
  wire u2__abc_44228_n16824;
  wire u2__abc_44228_n16825;
  wire u2__abc_44228_n16826;
  wire u2__abc_44228_n16828;
  wire u2__abc_44228_n16829;
  wire u2__abc_44228_n16830;
  wire u2__abc_44228_n16831;
  wire u2__abc_44228_n16833;
  wire u2__abc_44228_n16834;
  wire u2__abc_44228_n16835;
  wire u2__abc_44228_n16836;
  wire u2__abc_44228_n16838;
  wire u2__abc_44228_n16839;
  wire u2__abc_44228_n16840;
  wire u2__abc_44228_n16841;
  wire u2__abc_44228_n16843;
  wire u2__abc_44228_n16844;
  wire u2__abc_44228_n16845;
  wire u2__abc_44228_n16846;
  wire u2__abc_44228_n16848;
  wire u2__abc_44228_n16849;
  wire u2__abc_44228_n16850;
  wire u2__abc_44228_n16851;
  wire u2__abc_44228_n16853;
  wire u2__abc_44228_n16854;
  wire u2__abc_44228_n16855;
  wire u2__abc_44228_n16856;
  wire u2__abc_44228_n16858;
  wire u2__abc_44228_n16859;
  wire u2__abc_44228_n16860;
  wire u2__abc_44228_n16861;
  wire u2__abc_44228_n16863;
  wire u2__abc_44228_n16864;
  wire u2__abc_44228_n16865;
  wire u2__abc_44228_n16866;
  wire u2__abc_44228_n16868;
  wire u2__abc_44228_n16869;
  wire u2__abc_44228_n16870;
  wire u2__abc_44228_n16871;
  wire u2__abc_44228_n16873;
  wire u2__abc_44228_n16874;
  wire u2__abc_44228_n16875;
  wire u2__abc_44228_n16876;
  wire u2__abc_44228_n16878;
  wire u2__abc_44228_n16879;
  wire u2__abc_44228_n16880;
  wire u2__abc_44228_n16881;
  wire u2__abc_44228_n16883;
  wire u2__abc_44228_n16884;
  wire u2__abc_44228_n16885;
  wire u2__abc_44228_n16886;
  wire u2__abc_44228_n16888;
  wire u2__abc_44228_n16889;
  wire u2__abc_44228_n16890;
  wire u2__abc_44228_n16891;
  wire u2__abc_44228_n16893;
  wire u2__abc_44228_n16894;
  wire u2__abc_44228_n16895;
  wire u2__abc_44228_n16896;
  wire u2__abc_44228_n16898;
  wire u2__abc_44228_n16899;
  wire u2__abc_44228_n16900;
  wire u2__abc_44228_n16901;
  wire u2__abc_44228_n16903;
  wire u2__abc_44228_n16904;
  wire u2__abc_44228_n16905;
  wire u2__abc_44228_n16906;
  wire u2__abc_44228_n16908;
  wire u2__abc_44228_n16909;
  wire u2__abc_44228_n16910;
  wire u2__abc_44228_n16911;
  wire u2__abc_44228_n16913;
  wire u2__abc_44228_n16914;
  wire u2__abc_44228_n16915;
  wire u2__abc_44228_n16916;
  wire u2__abc_44228_n16918;
  wire u2__abc_44228_n16919;
  wire u2__abc_44228_n16920;
  wire u2__abc_44228_n16921;
  wire u2__abc_44228_n16923;
  wire u2__abc_44228_n16924;
  wire u2__abc_44228_n16925;
  wire u2__abc_44228_n16926;
  wire u2__abc_44228_n16928;
  wire u2__abc_44228_n16929;
  wire u2__abc_44228_n16930;
  wire u2__abc_44228_n16931;
  wire u2__abc_44228_n16933;
  wire u2__abc_44228_n16934;
  wire u2__abc_44228_n16935;
  wire u2__abc_44228_n16936;
  wire u2__abc_44228_n16938;
  wire u2__abc_44228_n16939;
  wire u2__abc_44228_n16940;
  wire u2__abc_44228_n16941;
  wire u2__abc_44228_n16943;
  wire u2__abc_44228_n16944;
  wire u2__abc_44228_n16945;
  wire u2__abc_44228_n16946;
  wire u2__abc_44228_n16948;
  wire u2__abc_44228_n16949;
  wire u2__abc_44228_n16950;
  wire u2__abc_44228_n16951;
  wire u2__abc_44228_n16953;
  wire u2__abc_44228_n16954;
  wire u2__abc_44228_n16955;
  wire u2__abc_44228_n16956;
  wire u2__abc_44228_n16958;
  wire u2__abc_44228_n16959;
  wire u2__abc_44228_n16960;
  wire u2__abc_44228_n16961;
  wire u2__abc_44228_n16963;
  wire u2__abc_44228_n16964;
  wire u2__abc_44228_n16965;
  wire u2__abc_44228_n16966;
  wire u2__abc_44228_n16968;
  wire u2__abc_44228_n16969;
  wire u2__abc_44228_n16970;
  wire u2__abc_44228_n16971;
  wire u2__abc_44228_n16973;
  wire u2__abc_44228_n16974;
  wire u2__abc_44228_n16975;
  wire u2__abc_44228_n16976;
  wire u2__abc_44228_n16978;
  wire u2__abc_44228_n16979;
  wire u2__abc_44228_n16980;
  wire u2__abc_44228_n16981;
  wire u2__abc_44228_n16983;
  wire u2__abc_44228_n16984;
  wire u2__abc_44228_n16985;
  wire u2__abc_44228_n16986;
  wire u2__abc_44228_n16988;
  wire u2__abc_44228_n16989;
  wire u2__abc_44228_n16990;
  wire u2__abc_44228_n16991;
  wire u2__abc_44228_n16993;
  wire u2__abc_44228_n16994;
  wire u2__abc_44228_n16995;
  wire u2__abc_44228_n16996;
  wire u2__abc_44228_n16998;
  wire u2__abc_44228_n16999;
  wire u2__abc_44228_n17000;
  wire u2__abc_44228_n17001;
  wire u2__abc_44228_n17003;
  wire u2__abc_44228_n17004;
  wire u2__abc_44228_n17005;
  wire u2__abc_44228_n17006;
  wire u2__abc_44228_n17008;
  wire u2__abc_44228_n17009;
  wire u2__abc_44228_n17010;
  wire u2__abc_44228_n17011;
  wire u2__abc_44228_n17013;
  wire u2__abc_44228_n17014;
  wire u2__abc_44228_n17015;
  wire u2__abc_44228_n17016;
  wire u2__abc_44228_n17018;
  wire u2__abc_44228_n17019;
  wire u2__abc_44228_n17020;
  wire u2__abc_44228_n17021;
  wire u2__abc_44228_n17023;
  wire u2__abc_44228_n17024;
  wire u2__abc_44228_n17025;
  wire u2__abc_44228_n17026;
  wire u2__abc_44228_n17028;
  wire u2__abc_44228_n17029;
  wire u2__abc_44228_n17030;
  wire u2__abc_44228_n17031;
  wire u2__abc_44228_n17033;
  wire u2__abc_44228_n17034;
  wire u2__abc_44228_n17035;
  wire u2__abc_44228_n17036;
  wire u2__abc_44228_n17038;
  wire u2__abc_44228_n17039;
  wire u2__abc_44228_n17040;
  wire u2__abc_44228_n17041;
  wire u2__abc_44228_n17043;
  wire u2__abc_44228_n17044;
  wire u2__abc_44228_n17045;
  wire u2__abc_44228_n17046;
  wire u2__abc_44228_n17048;
  wire u2__abc_44228_n17049;
  wire u2__abc_44228_n17050;
  wire u2__abc_44228_n17051;
  wire u2__abc_44228_n17053;
  wire u2__abc_44228_n17054;
  wire u2__abc_44228_n17055;
  wire u2__abc_44228_n17056;
  wire u2__abc_44228_n17058;
  wire u2__abc_44228_n17059;
  wire u2__abc_44228_n17060;
  wire u2__abc_44228_n17061;
  wire u2__abc_44228_n17063;
  wire u2__abc_44228_n17064;
  wire u2__abc_44228_n17065;
  wire u2__abc_44228_n17066;
  wire u2__abc_44228_n17068;
  wire u2__abc_44228_n17069;
  wire u2__abc_44228_n17070;
  wire u2__abc_44228_n17071;
  wire u2__abc_44228_n17073;
  wire u2__abc_44228_n17074;
  wire u2__abc_44228_n17075;
  wire u2__abc_44228_n17076;
  wire u2__abc_44228_n17078;
  wire u2__abc_44228_n17079;
  wire u2__abc_44228_n17080;
  wire u2__abc_44228_n17081;
  wire u2__abc_44228_n17083;
  wire u2__abc_44228_n17084;
  wire u2__abc_44228_n17085;
  wire u2__abc_44228_n17086;
  wire u2__abc_44228_n17088;
  wire u2__abc_44228_n17089;
  wire u2__abc_44228_n17090;
  wire u2__abc_44228_n17091;
  wire u2__abc_44228_n17093;
  wire u2__abc_44228_n17094;
  wire u2__abc_44228_n17095;
  wire u2__abc_44228_n17096;
  wire u2__abc_44228_n17098;
  wire u2__abc_44228_n17099;
  wire u2__abc_44228_n17100;
  wire u2__abc_44228_n17101;
  wire u2__abc_44228_n17103;
  wire u2__abc_44228_n17104;
  wire u2__abc_44228_n17105;
  wire u2__abc_44228_n17106;
  wire u2__abc_44228_n17108;
  wire u2__abc_44228_n17109;
  wire u2__abc_44228_n17110;
  wire u2__abc_44228_n17111;
  wire u2__abc_44228_n17113;
  wire u2__abc_44228_n17114;
  wire u2__abc_44228_n17115;
  wire u2__abc_44228_n17116;
  wire u2__abc_44228_n17118;
  wire u2__abc_44228_n17119;
  wire u2__abc_44228_n17120;
  wire u2__abc_44228_n17121;
  wire u2__abc_44228_n17123;
  wire u2__abc_44228_n17124;
  wire u2__abc_44228_n17125;
  wire u2__abc_44228_n17126;
  wire u2__abc_44228_n17128;
  wire u2__abc_44228_n17129;
  wire u2__abc_44228_n17130;
  wire u2__abc_44228_n17131;
  wire u2__abc_44228_n17133;
  wire u2__abc_44228_n17134;
  wire u2__abc_44228_n17135;
  wire u2__abc_44228_n17136;
  wire u2__abc_44228_n17138;
  wire u2__abc_44228_n17139;
  wire u2__abc_44228_n17140;
  wire u2__abc_44228_n17141;
  wire u2__abc_44228_n17143;
  wire u2__abc_44228_n17144;
  wire u2__abc_44228_n17145;
  wire u2__abc_44228_n17146;
  wire u2__abc_44228_n17148;
  wire u2__abc_44228_n17149;
  wire u2__abc_44228_n17150;
  wire u2__abc_44228_n17151;
  wire u2__abc_44228_n17153;
  wire u2__abc_44228_n17154;
  wire u2__abc_44228_n17155;
  wire u2__abc_44228_n17156;
  wire u2__abc_44228_n17158;
  wire u2__abc_44228_n17159;
  wire u2__abc_44228_n17160;
  wire u2__abc_44228_n17161;
  wire u2__abc_44228_n17163;
  wire u2__abc_44228_n17164;
  wire u2__abc_44228_n17165;
  wire u2__abc_44228_n17166;
  wire u2__abc_44228_n17168;
  wire u2__abc_44228_n17169;
  wire u2__abc_44228_n17170;
  wire u2__abc_44228_n17171;
  wire u2__abc_44228_n17173;
  wire u2__abc_44228_n17174;
  wire u2__abc_44228_n17175;
  wire u2__abc_44228_n17176;
  wire u2__abc_44228_n17178;
  wire u2__abc_44228_n17179;
  wire u2__abc_44228_n17180;
  wire u2__abc_44228_n17181;
  wire u2__abc_44228_n17183;
  wire u2__abc_44228_n17184;
  wire u2__abc_44228_n17185;
  wire u2__abc_44228_n17186;
  wire u2__abc_44228_n17188;
  wire u2__abc_44228_n17189;
  wire u2__abc_44228_n17190;
  wire u2__abc_44228_n17191;
  wire u2__abc_44228_n17193;
  wire u2__abc_44228_n17194;
  wire u2__abc_44228_n17195;
  wire u2__abc_44228_n17196;
  wire u2__abc_44228_n17198;
  wire u2__abc_44228_n17199;
  wire u2__abc_44228_n17200;
  wire u2__abc_44228_n17201;
  wire u2__abc_44228_n17203;
  wire u2__abc_44228_n17204;
  wire u2__abc_44228_n17205;
  wire u2__abc_44228_n17206;
  wire u2__abc_44228_n17208;
  wire u2__abc_44228_n17209;
  wire u2__abc_44228_n17210;
  wire u2__abc_44228_n17211;
  wire u2__abc_44228_n17213;
  wire u2__abc_44228_n17214;
  wire u2__abc_44228_n17215;
  wire u2__abc_44228_n17216;
  wire u2__abc_44228_n17218;
  wire u2__abc_44228_n17219;
  wire u2__abc_44228_n17220;
  wire u2__abc_44228_n17221;
  wire u2__abc_44228_n17223;
  wire u2__abc_44228_n17224;
  wire u2__abc_44228_n17225;
  wire u2__abc_44228_n17226;
  wire u2__abc_44228_n17228;
  wire u2__abc_44228_n17229;
  wire u2__abc_44228_n17230;
  wire u2__abc_44228_n17231;
  wire u2__abc_44228_n17233;
  wire u2__abc_44228_n17234;
  wire u2__abc_44228_n17235;
  wire u2__abc_44228_n17236;
  wire u2__abc_44228_n17238;
  wire u2__abc_44228_n17239;
  wire u2__abc_44228_n17240;
  wire u2__abc_44228_n17241;
  wire u2__abc_44228_n17243;
  wire u2__abc_44228_n17244;
  wire u2__abc_44228_n17245;
  wire u2__abc_44228_n17246;
  wire u2__abc_44228_n17248;
  wire u2__abc_44228_n17249;
  wire u2__abc_44228_n17250;
  wire u2__abc_44228_n17251;
  wire u2__abc_44228_n17253;
  wire u2__abc_44228_n17254;
  wire u2__abc_44228_n17255;
  wire u2__abc_44228_n17256;
  wire u2__abc_44228_n17258;
  wire u2__abc_44228_n17259;
  wire u2__abc_44228_n17260;
  wire u2__abc_44228_n17261;
  wire u2__abc_44228_n17263;
  wire u2__abc_44228_n17264;
  wire u2__abc_44228_n17265;
  wire u2__abc_44228_n17266;
  wire u2__abc_44228_n17268;
  wire u2__abc_44228_n17269;
  wire u2__abc_44228_n17270;
  wire u2__abc_44228_n17271;
  wire u2__abc_44228_n17273;
  wire u2__abc_44228_n17274;
  wire u2__abc_44228_n17275;
  wire u2__abc_44228_n17276;
  wire u2__abc_44228_n17278;
  wire u2__abc_44228_n17279;
  wire u2__abc_44228_n17280;
  wire u2__abc_44228_n17281;
  wire u2__abc_44228_n17283;
  wire u2__abc_44228_n17284;
  wire u2__abc_44228_n17285;
  wire u2__abc_44228_n17286;
  wire u2__abc_44228_n17288;
  wire u2__abc_44228_n17289;
  wire u2__abc_44228_n17290;
  wire u2__abc_44228_n17291;
  wire u2__abc_44228_n17293;
  wire u2__abc_44228_n17294;
  wire u2__abc_44228_n17295;
  wire u2__abc_44228_n17296;
  wire u2__abc_44228_n17298;
  wire u2__abc_44228_n17299;
  wire u2__abc_44228_n17300;
  wire u2__abc_44228_n17301;
  wire u2__abc_44228_n17303;
  wire u2__abc_44228_n17304;
  wire u2__abc_44228_n17305;
  wire u2__abc_44228_n17306;
  wire u2__abc_44228_n17308;
  wire u2__abc_44228_n17309;
  wire u2__abc_44228_n17310;
  wire u2__abc_44228_n17311;
  wire u2__abc_44228_n17313;
  wire u2__abc_44228_n17314;
  wire u2__abc_44228_n17315;
  wire u2__abc_44228_n17316;
  wire u2__abc_44228_n17318;
  wire u2__abc_44228_n17319;
  wire u2__abc_44228_n17320;
  wire u2__abc_44228_n17321;
  wire u2__abc_44228_n17323;
  wire u2__abc_44228_n17324;
  wire u2__abc_44228_n17325;
  wire u2__abc_44228_n17326;
  wire u2__abc_44228_n17328;
  wire u2__abc_44228_n17329;
  wire u2__abc_44228_n17330;
  wire u2__abc_44228_n17331;
  wire u2__abc_44228_n17333;
  wire u2__abc_44228_n17334;
  wire u2__abc_44228_n17335;
  wire u2__abc_44228_n17336;
  wire u2__abc_44228_n17338;
  wire u2__abc_44228_n17339;
  wire u2__abc_44228_n17340;
  wire u2__abc_44228_n17341;
  wire u2__abc_44228_n17343;
  wire u2__abc_44228_n17344;
  wire u2__abc_44228_n17345;
  wire u2__abc_44228_n17346;
  wire u2__abc_44228_n17348;
  wire u2__abc_44228_n17349;
  wire u2__abc_44228_n17350;
  wire u2__abc_44228_n17351;
  wire u2__abc_44228_n17353;
  wire u2__abc_44228_n17354;
  wire u2__abc_44228_n17355;
  wire u2__abc_44228_n17356;
  wire u2__abc_44228_n17358;
  wire u2__abc_44228_n17359;
  wire u2__abc_44228_n17360;
  wire u2__abc_44228_n17361;
  wire u2__abc_44228_n17363;
  wire u2__abc_44228_n17364;
  wire u2__abc_44228_n17365;
  wire u2__abc_44228_n17366;
  wire u2__abc_44228_n17368;
  wire u2__abc_44228_n17369;
  wire u2__abc_44228_n17370;
  wire u2__abc_44228_n17371;
  wire u2__abc_44228_n17373;
  wire u2__abc_44228_n17374;
  wire u2__abc_44228_n17375;
  wire u2__abc_44228_n17376;
  wire u2__abc_44228_n17378;
  wire u2__abc_44228_n17379;
  wire u2__abc_44228_n17380;
  wire u2__abc_44228_n17381;
  wire u2__abc_44228_n17383;
  wire u2__abc_44228_n17384;
  wire u2__abc_44228_n17385;
  wire u2__abc_44228_n17386;
  wire u2__abc_44228_n17388;
  wire u2__abc_44228_n17389;
  wire u2__abc_44228_n17390;
  wire u2__abc_44228_n17391;
  wire u2__abc_44228_n17393;
  wire u2__abc_44228_n17394;
  wire u2__abc_44228_n17395;
  wire u2__abc_44228_n17396;
  wire u2__abc_44228_n17398;
  wire u2__abc_44228_n17399;
  wire u2__abc_44228_n17400;
  wire u2__abc_44228_n17401;
  wire u2__abc_44228_n17403;
  wire u2__abc_44228_n17404;
  wire u2__abc_44228_n17405;
  wire u2__abc_44228_n17406;
  wire u2__abc_44228_n17408;
  wire u2__abc_44228_n17409;
  wire u2__abc_44228_n17410;
  wire u2__abc_44228_n17411;
  wire u2__abc_44228_n17413;
  wire u2__abc_44228_n17414;
  wire u2__abc_44228_n17415;
  wire u2__abc_44228_n17416;
  wire u2__abc_44228_n17418;
  wire u2__abc_44228_n17419;
  wire u2__abc_44228_n17420;
  wire u2__abc_44228_n17421;
  wire u2__abc_44228_n17423;
  wire u2__abc_44228_n17424;
  wire u2__abc_44228_n17425;
  wire u2__abc_44228_n17426;
  wire u2__abc_44228_n17428;
  wire u2__abc_44228_n17429;
  wire u2__abc_44228_n17430;
  wire u2__abc_44228_n17431;
  wire u2__abc_44228_n17433;
  wire u2__abc_44228_n17434;
  wire u2__abc_44228_n17435;
  wire u2__abc_44228_n17436;
  wire u2__abc_44228_n17438;
  wire u2__abc_44228_n17439;
  wire u2__abc_44228_n17440;
  wire u2__abc_44228_n17441;
  wire u2__abc_44228_n17443;
  wire u2__abc_44228_n17444;
  wire u2__abc_44228_n17445;
  wire u2__abc_44228_n17446;
  wire u2__abc_44228_n17448;
  wire u2__abc_44228_n17449;
  wire u2__abc_44228_n17450;
  wire u2__abc_44228_n17451;
  wire u2__abc_44228_n17453;
  wire u2__abc_44228_n17454;
  wire u2__abc_44228_n17455;
  wire u2__abc_44228_n17456;
  wire u2__abc_44228_n17458;
  wire u2__abc_44228_n17459;
  wire u2__abc_44228_n17460;
  wire u2__abc_44228_n17461;
  wire u2__abc_44228_n17463;
  wire u2__abc_44228_n17464;
  wire u2__abc_44228_n17465;
  wire u2__abc_44228_n17466;
  wire u2__abc_44228_n17468;
  wire u2__abc_44228_n17469;
  wire u2__abc_44228_n17470;
  wire u2__abc_44228_n17471;
  wire u2__abc_44228_n17473;
  wire u2__abc_44228_n17474;
  wire u2__abc_44228_n17475;
  wire u2__abc_44228_n17476;
  wire u2__abc_44228_n17478;
  wire u2__abc_44228_n17479;
  wire u2__abc_44228_n17480;
  wire u2__abc_44228_n17481;
  wire u2__abc_44228_n17483;
  wire u2__abc_44228_n17484;
  wire u2__abc_44228_n17485;
  wire u2__abc_44228_n17486;
  wire u2__abc_44228_n17488;
  wire u2__abc_44228_n17489;
  wire u2__abc_44228_n17490;
  wire u2__abc_44228_n17491;
  wire u2__abc_44228_n17493;
  wire u2__abc_44228_n17494;
  wire u2__abc_44228_n17495;
  wire u2__abc_44228_n17496;
  wire u2__abc_44228_n17498;
  wire u2__abc_44228_n17499;
  wire u2__abc_44228_n17500;
  wire u2__abc_44228_n17501;
  wire u2__abc_44228_n17503;
  wire u2__abc_44228_n17504;
  wire u2__abc_44228_n17505;
  wire u2__abc_44228_n17506;
  wire u2__abc_44228_n17508;
  wire u2__abc_44228_n17509;
  wire u2__abc_44228_n17510;
  wire u2__abc_44228_n17511;
  wire u2__abc_44228_n17513;
  wire u2__abc_44228_n17514;
  wire u2__abc_44228_n17515;
  wire u2__abc_44228_n17516;
  wire u2__abc_44228_n17518;
  wire u2__abc_44228_n17519;
  wire u2__abc_44228_n17520;
  wire u2__abc_44228_n17521;
  wire u2__abc_44228_n17523;
  wire u2__abc_44228_n17524;
  wire u2__abc_44228_n17525;
  wire u2__abc_44228_n17526;
  wire u2__abc_44228_n17528;
  wire u2__abc_44228_n17529;
  wire u2__abc_44228_n17530;
  wire u2__abc_44228_n17531;
  wire u2__abc_44228_n17533;
  wire u2__abc_44228_n17534;
  wire u2__abc_44228_n17535;
  wire u2__abc_44228_n17536;
  wire u2__abc_44228_n17538;
  wire u2__abc_44228_n17539;
  wire u2__abc_44228_n17540;
  wire u2__abc_44228_n17541;
  wire u2__abc_44228_n17543;
  wire u2__abc_44228_n17544;
  wire u2__abc_44228_n17545;
  wire u2__abc_44228_n17546;
  wire u2__abc_44228_n17548;
  wire u2__abc_44228_n17549;
  wire u2__abc_44228_n17550;
  wire u2__abc_44228_n17551;
  wire u2__abc_44228_n17553;
  wire u2__abc_44228_n17554;
  wire u2__abc_44228_n17555;
  wire u2__abc_44228_n17556;
  wire u2__abc_44228_n17558;
  wire u2__abc_44228_n17559;
  wire u2__abc_44228_n17560;
  wire u2__abc_44228_n17561;
  wire u2__abc_44228_n17563;
  wire u2__abc_44228_n17564;
  wire u2__abc_44228_n17565;
  wire u2__abc_44228_n17566;
  wire u2__abc_44228_n17568;
  wire u2__abc_44228_n17569;
  wire u2__abc_44228_n17570;
  wire u2__abc_44228_n17571;
  wire u2__abc_44228_n17573;
  wire u2__abc_44228_n17574;
  wire u2__abc_44228_n17575;
  wire u2__abc_44228_n17576;
  wire u2__abc_44228_n17578;
  wire u2__abc_44228_n17579;
  wire u2__abc_44228_n17580;
  wire u2__abc_44228_n17581;
  wire u2__abc_44228_n17583;
  wire u2__abc_44228_n17584;
  wire u2__abc_44228_n17585;
  wire u2__abc_44228_n17586;
  wire u2__abc_44228_n17588;
  wire u2__abc_44228_n17589;
  wire u2__abc_44228_n17590;
  wire u2__abc_44228_n17591;
  wire u2__abc_44228_n17593;
  wire u2__abc_44228_n17594;
  wire u2__abc_44228_n17595;
  wire u2__abc_44228_n17596;
  wire u2__abc_44228_n17598;
  wire u2__abc_44228_n17599;
  wire u2__abc_44228_n17600;
  wire u2__abc_44228_n17601;
  wire u2__abc_44228_n17603;
  wire u2__abc_44228_n17604;
  wire u2__abc_44228_n17605;
  wire u2__abc_44228_n17606;
  wire u2__abc_44228_n17608;
  wire u2__abc_44228_n17609;
  wire u2__abc_44228_n17610;
  wire u2__abc_44228_n17611;
  wire u2__abc_44228_n17613;
  wire u2__abc_44228_n17614;
  wire u2__abc_44228_n17615;
  wire u2__abc_44228_n17616;
  wire u2__abc_44228_n17618;
  wire u2__abc_44228_n17619;
  wire u2__abc_44228_n17620;
  wire u2__abc_44228_n17621;
  wire u2__abc_44228_n17623;
  wire u2__abc_44228_n17624;
  wire u2__abc_44228_n17625;
  wire u2__abc_44228_n17626;
  wire u2__abc_44228_n17628;
  wire u2__abc_44228_n17629;
  wire u2__abc_44228_n17630;
  wire u2__abc_44228_n17631;
  wire u2__abc_44228_n17633;
  wire u2__abc_44228_n17634;
  wire u2__abc_44228_n17635;
  wire u2__abc_44228_n17636;
  wire u2__abc_44228_n17638;
  wire u2__abc_44228_n17639;
  wire u2__abc_44228_n17640;
  wire u2__abc_44228_n17641;
  wire u2__abc_44228_n17643;
  wire u2__abc_44228_n17644;
  wire u2__abc_44228_n17645;
  wire u2__abc_44228_n17646;
  wire u2__abc_44228_n17648;
  wire u2__abc_44228_n17649;
  wire u2__abc_44228_n17650;
  wire u2__abc_44228_n17651;
  wire u2__abc_44228_n17653;
  wire u2__abc_44228_n17654;
  wire u2__abc_44228_n17655;
  wire u2__abc_44228_n17656;
  wire u2__abc_44228_n17658;
  wire u2__abc_44228_n17659;
  wire u2__abc_44228_n17660;
  wire u2__abc_44228_n17661;
  wire u2__abc_44228_n17663;
  wire u2__abc_44228_n17664;
  wire u2__abc_44228_n17665;
  wire u2__abc_44228_n17666;
  wire u2__abc_44228_n17668;
  wire u2__abc_44228_n17669;
  wire u2__abc_44228_n17670;
  wire u2__abc_44228_n17671;
  wire u2__abc_44228_n17673;
  wire u2__abc_44228_n17674;
  wire u2__abc_44228_n17675;
  wire u2__abc_44228_n17676;
  wire u2__abc_44228_n17678;
  wire u2__abc_44228_n17679;
  wire u2__abc_44228_n17680;
  wire u2__abc_44228_n17681;
  wire u2__abc_44228_n17683;
  wire u2__abc_44228_n17684;
  wire u2__abc_44228_n17685;
  wire u2__abc_44228_n17686;
  wire u2__abc_44228_n17688;
  wire u2__abc_44228_n17689;
  wire u2__abc_44228_n17690;
  wire u2__abc_44228_n17691;
  wire u2__abc_44228_n17693;
  wire u2__abc_44228_n17694;
  wire u2__abc_44228_n17695;
  wire u2__abc_44228_n17696;
  wire u2__abc_44228_n17698;
  wire u2__abc_44228_n17699;
  wire u2__abc_44228_n17700;
  wire u2__abc_44228_n17701;
  wire u2__abc_44228_n17703;
  wire u2__abc_44228_n17704;
  wire u2__abc_44228_n17705;
  wire u2__abc_44228_n17706;
  wire u2__abc_44228_n17708;
  wire u2__abc_44228_n17709;
  wire u2__abc_44228_n17710;
  wire u2__abc_44228_n17711;
  wire u2__abc_44228_n17713;
  wire u2__abc_44228_n17714;
  wire u2__abc_44228_n17715;
  wire u2__abc_44228_n17716;
  wire u2__abc_44228_n17718;
  wire u2__abc_44228_n17719;
  wire u2__abc_44228_n17720;
  wire u2__abc_44228_n17721;
  wire u2__abc_44228_n17723;
  wire u2__abc_44228_n17724;
  wire u2__abc_44228_n17725;
  wire u2__abc_44228_n17726;
  wire u2__abc_44228_n17728;
  wire u2__abc_44228_n17729;
  wire u2__abc_44228_n17730;
  wire u2__abc_44228_n17731;
  wire u2__abc_44228_n17733;
  wire u2__abc_44228_n17734;
  wire u2__abc_44228_n17735;
  wire u2__abc_44228_n17736;
  wire u2__abc_44228_n17738;
  wire u2__abc_44228_n17739;
  wire u2__abc_44228_n17740;
  wire u2__abc_44228_n17741;
  wire u2__abc_44228_n17743;
  wire u2__abc_44228_n17744;
  wire u2__abc_44228_n17745;
  wire u2__abc_44228_n17746;
  wire u2__abc_44228_n17748;
  wire u2__abc_44228_n17749;
  wire u2__abc_44228_n17750;
  wire u2__abc_44228_n17751;
  wire u2__abc_44228_n17753;
  wire u2__abc_44228_n17754;
  wire u2__abc_44228_n17755;
  wire u2__abc_44228_n17756;
  wire u2__abc_44228_n17758;
  wire u2__abc_44228_n17759;
  wire u2__abc_44228_n17760;
  wire u2__abc_44228_n17761;
  wire u2__abc_44228_n17763;
  wire u2__abc_44228_n17764;
  wire u2__abc_44228_n17765;
  wire u2__abc_44228_n17766;
  wire u2__abc_44228_n17768;
  wire u2__abc_44228_n17769;
  wire u2__abc_44228_n17770;
  wire u2__abc_44228_n17771;
  wire u2__abc_44228_n17773;
  wire u2__abc_44228_n17775;
  wire u2__abc_44228_n17776;
  wire u2__abc_44228_n17777;
  wire u2__abc_44228_n17778;
  wire u2__abc_44228_n17779;
  wire u2__abc_44228_n17780;
  wire u2__abc_44228_n17781;
  wire u2__abc_44228_n17782;
  wire u2__abc_44228_n17783;
  wire u2__abc_44228_n17784;
  wire u2__abc_44228_n17785;
  wire u2__abc_44228_n17787;
  wire u2__abc_44228_n17788;
  wire u2__abc_44228_n17789;
  wire u2__abc_44228_n17790;
  wire u2__abc_44228_n17791;
  wire u2__abc_44228_n17792;
  wire u2__abc_44228_n17793;
  wire u2__abc_44228_n17794;
  wire u2__abc_44228_n17795;
  wire u2__abc_44228_n17796;
  wire u2__abc_44228_n17797;
  wire u2__abc_44228_n17799;
  wire u2__abc_44228_n17800;
  wire u2__abc_44228_n17801;
  wire u2__abc_44228_n17802;
  wire u2__abc_44228_n17803;
  wire u2__abc_44228_n17804;
  wire u2__abc_44228_n17805;
  wire u2__abc_44228_n17806;
  wire u2__abc_44228_n17807;
  wire u2__abc_44228_n17808;
  wire u2__abc_44228_n17809;
  wire u2__abc_44228_n17811;
  wire u2__abc_44228_n17812;
  wire u2__abc_44228_n17813;
  wire u2__abc_44228_n17814;
  wire u2__abc_44228_n17815;
  wire u2__abc_44228_n17816;
  wire u2__abc_44228_n17817;
  wire u2__abc_44228_n17818;
  wire u2__abc_44228_n17819;
  wire u2__abc_44228_n17820;
  wire u2__abc_44228_n17821;
  wire u2__abc_44228_n17823;
  wire u2__abc_44228_n17824;
  wire u2__abc_44228_n17825;
  wire u2__abc_44228_n17826;
  wire u2__abc_44228_n17827;
  wire u2__abc_44228_n17828;
  wire u2__abc_44228_n17829;
  wire u2__abc_44228_n17830;
  wire u2__abc_44228_n17831;
  wire u2__abc_44228_n17832;
  wire u2__abc_44228_n17833;
  wire u2__abc_44228_n17835;
  wire u2__abc_44228_n17836;
  wire u2__abc_44228_n17837;
  wire u2__abc_44228_n17838;
  wire u2__abc_44228_n17839;
  wire u2__abc_44228_n17840;
  wire u2__abc_44228_n17841;
  wire u2__abc_44228_n17842;
  wire u2__abc_44228_n17843;
  wire u2__abc_44228_n17844;
  wire u2__abc_44228_n17845;
  wire u2__abc_44228_n17847;
  wire u2__abc_44228_n17848;
  wire u2__abc_44228_n17849;
  wire u2__abc_44228_n17850;
  wire u2__abc_44228_n17851;
  wire u2__abc_44228_n17852;
  wire u2__abc_44228_n17853;
  wire u2__abc_44228_n17854;
  wire u2__abc_44228_n17855;
  wire u2__abc_44228_n17856;
  wire u2__abc_44228_n17857;
  wire u2__abc_44228_n17859;
  wire u2__abc_44228_n17860;
  wire u2__abc_44228_n17861;
  wire u2__abc_44228_n17862;
  wire u2__abc_44228_n17863;
  wire u2__abc_44228_n17864;
  wire u2__abc_44228_n17865;
  wire u2__abc_44228_n17866;
  wire u2__abc_44228_n17867;
  wire u2__abc_44228_n17868;
  wire u2__abc_44228_n17869;
  wire u2__abc_44228_n17871;
  wire u2__abc_44228_n17872;
  wire u2__abc_44228_n17873;
  wire u2__abc_44228_n17874;
  wire u2__abc_44228_n17875;
  wire u2__abc_44228_n17876;
  wire u2__abc_44228_n17877;
  wire u2__abc_44228_n17878;
  wire u2__abc_44228_n17879;
  wire u2__abc_44228_n17880;
  wire u2__abc_44228_n17881;
  wire u2__abc_44228_n17883;
  wire u2__abc_44228_n17884;
  wire u2__abc_44228_n17885;
  wire u2__abc_44228_n17886;
  wire u2__abc_44228_n17887;
  wire u2__abc_44228_n17888;
  wire u2__abc_44228_n17889;
  wire u2__abc_44228_n17890;
  wire u2__abc_44228_n17891;
  wire u2__abc_44228_n17892;
  wire u2__abc_44228_n17893;
  wire u2__abc_44228_n17895;
  wire u2__abc_44228_n17896;
  wire u2__abc_44228_n17897;
  wire u2__abc_44228_n17898;
  wire u2__abc_44228_n17899;
  wire u2__abc_44228_n17900;
  wire u2__abc_44228_n17901;
  wire u2__abc_44228_n17902;
  wire u2__abc_44228_n17903;
  wire u2__abc_44228_n17904;
  wire u2__abc_44228_n17905;
  wire u2__abc_44228_n17907;
  wire u2__abc_44228_n17908;
  wire u2__abc_44228_n17909;
  wire u2__abc_44228_n17910;
  wire u2__abc_44228_n17911;
  wire u2__abc_44228_n17912;
  wire u2__abc_44228_n17913;
  wire u2__abc_44228_n17914;
  wire u2__abc_44228_n17915;
  wire u2__abc_44228_n17916;
  wire u2__abc_44228_n17917;
  wire u2__abc_44228_n17919;
  wire u2__abc_44228_n17920;
  wire u2__abc_44228_n17921;
  wire u2__abc_44228_n17922;
  wire u2__abc_44228_n17923;
  wire u2__abc_44228_n17924;
  wire u2__abc_44228_n17925;
  wire u2__abc_44228_n17926;
  wire u2__abc_44228_n17927;
  wire u2__abc_44228_n17928;
  wire u2__abc_44228_n17929;
  wire u2__abc_44228_n17931;
  wire u2__abc_44228_n17932;
  wire u2__abc_44228_n17933;
  wire u2__abc_44228_n17934;
  wire u2__abc_44228_n17935;
  wire u2__abc_44228_n17936;
  wire u2__abc_44228_n17937;
  wire u2__abc_44228_n17938;
  wire u2__abc_44228_n17939;
  wire u2__abc_44228_n17940;
  wire u2__abc_44228_n17941;
  wire u2__abc_44228_n17943;
  wire u2__abc_44228_n17944;
  wire u2__abc_44228_n17945;
  wire u2__abc_44228_n17946;
  wire u2__abc_44228_n17947;
  wire u2__abc_44228_n17948;
  wire u2__abc_44228_n17949;
  wire u2__abc_44228_n17950;
  wire u2__abc_44228_n17951;
  wire u2__abc_44228_n17952;
  wire u2__abc_44228_n17953;
  wire u2__abc_44228_n17955;
  wire u2__abc_44228_n17956;
  wire u2__abc_44228_n17957;
  wire u2__abc_44228_n17958;
  wire u2__abc_44228_n17959;
  wire u2__abc_44228_n17960;
  wire u2__abc_44228_n17961;
  wire u2__abc_44228_n17962;
  wire u2__abc_44228_n17963;
  wire u2__abc_44228_n17964;
  wire u2__abc_44228_n17965;
  wire u2__abc_44228_n17967;
  wire u2__abc_44228_n17968;
  wire u2__abc_44228_n17969;
  wire u2__abc_44228_n17970;
  wire u2__abc_44228_n17971;
  wire u2__abc_44228_n17972;
  wire u2__abc_44228_n17973;
  wire u2__abc_44228_n17974;
  wire u2__abc_44228_n17975;
  wire u2__abc_44228_n17976;
  wire u2__abc_44228_n17977;
  wire u2__abc_44228_n17979;
  wire u2__abc_44228_n17980;
  wire u2__abc_44228_n17981;
  wire u2__abc_44228_n17982;
  wire u2__abc_44228_n17983;
  wire u2__abc_44228_n17984;
  wire u2__abc_44228_n17985;
  wire u2__abc_44228_n17986;
  wire u2__abc_44228_n17987;
  wire u2__abc_44228_n17988;
  wire u2__abc_44228_n17989;
  wire u2__abc_44228_n17991;
  wire u2__abc_44228_n17992;
  wire u2__abc_44228_n17993;
  wire u2__abc_44228_n17994;
  wire u2__abc_44228_n17995;
  wire u2__abc_44228_n17996;
  wire u2__abc_44228_n17997;
  wire u2__abc_44228_n17998;
  wire u2__abc_44228_n17999;
  wire u2__abc_44228_n18000;
  wire u2__abc_44228_n18001;
  wire u2__abc_44228_n18003;
  wire u2__abc_44228_n18004;
  wire u2__abc_44228_n18005;
  wire u2__abc_44228_n18006;
  wire u2__abc_44228_n18007;
  wire u2__abc_44228_n18008;
  wire u2__abc_44228_n18009;
  wire u2__abc_44228_n18010;
  wire u2__abc_44228_n18011;
  wire u2__abc_44228_n18012;
  wire u2__abc_44228_n18013;
  wire u2__abc_44228_n18015;
  wire u2__abc_44228_n18016;
  wire u2__abc_44228_n18017;
  wire u2__abc_44228_n18018;
  wire u2__abc_44228_n18019;
  wire u2__abc_44228_n18020;
  wire u2__abc_44228_n18021;
  wire u2__abc_44228_n18022;
  wire u2__abc_44228_n18023;
  wire u2__abc_44228_n18024;
  wire u2__abc_44228_n18025;
  wire u2__abc_44228_n18027;
  wire u2__abc_44228_n18028;
  wire u2__abc_44228_n18029;
  wire u2__abc_44228_n18030;
  wire u2__abc_44228_n18031;
  wire u2__abc_44228_n18032;
  wire u2__abc_44228_n18033;
  wire u2__abc_44228_n18034;
  wire u2__abc_44228_n18035;
  wire u2__abc_44228_n18036;
  wire u2__abc_44228_n18037;
  wire u2__abc_44228_n18039;
  wire u2__abc_44228_n18040;
  wire u2__abc_44228_n18041;
  wire u2__abc_44228_n18042;
  wire u2__abc_44228_n18043;
  wire u2__abc_44228_n18044;
  wire u2__abc_44228_n18045;
  wire u2__abc_44228_n18046;
  wire u2__abc_44228_n18047;
  wire u2__abc_44228_n18048;
  wire u2__abc_44228_n18049;
  wire u2__abc_44228_n18051;
  wire u2__abc_44228_n18052;
  wire u2__abc_44228_n18053;
  wire u2__abc_44228_n18054;
  wire u2__abc_44228_n18055;
  wire u2__abc_44228_n18056;
  wire u2__abc_44228_n18057;
  wire u2__abc_44228_n18058;
  wire u2__abc_44228_n18059;
  wire u2__abc_44228_n18060;
  wire u2__abc_44228_n18061;
  wire u2__abc_44228_n18063;
  wire u2__abc_44228_n18064;
  wire u2__abc_44228_n18065;
  wire u2__abc_44228_n18066;
  wire u2__abc_44228_n18067;
  wire u2__abc_44228_n18068;
  wire u2__abc_44228_n18069;
  wire u2__abc_44228_n18070;
  wire u2__abc_44228_n18071;
  wire u2__abc_44228_n18072;
  wire u2__abc_44228_n18073;
  wire u2__abc_44228_n18075;
  wire u2__abc_44228_n18076;
  wire u2__abc_44228_n18077;
  wire u2__abc_44228_n18078;
  wire u2__abc_44228_n18079;
  wire u2__abc_44228_n18080;
  wire u2__abc_44228_n18081;
  wire u2__abc_44228_n18082;
  wire u2__abc_44228_n18083;
  wire u2__abc_44228_n18084;
  wire u2__abc_44228_n18085;
  wire u2__abc_44228_n18087;
  wire u2__abc_44228_n18088;
  wire u2__abc_44228_n18089;
  wire u2__abc_44228_n18090;
  wire u2__abc_44228_n18091;
  wire u2__abc_44228_n18092;
  wire u2__abc_44228_n18093;
  wire u2__abc_44228_n18094;
  wire u2__abc_44228_n18095;
  wire u2__abc_44228_n18096;
  wire u2__abc_44228_n18097;
  wire u2__abc_44228_n18099;
  wire u2__abc_44228_n18100;
  wire u2__abc_44228_n18101;
  wire u2__abc_44228_n18102;
  wire u2__abc_44228_n18103;
  wire u2__abc_44228_n18104;
  wire u2__abc_44228_n18105;
  wire u2__abc_44228_n18106;
  wire u2__abc_44228_n18107;
  wire u2__abc_44228_n18108;
  wire u2__abc_44228_n18109;
  wire u2__abc_44228_n18111;
  wire u2__abc_44228_n18112;
  wire u2__abc_44228_n18113;
  wire u2__abc_44228_n18114;
  wire u2__abc_44228_n18115;
  wire u2__abc_44228_n18116;
  wire u2__abc_44228_n18117;
  wire u2__abc_44228_n18118;
  wire u2__abc_44228_n18119;
  wire u2__abc_44228_n18120;
  wire u2__abc_44228_n18121;
  wire u2__abc_44228_n18123;
  wire u2__abc_44228_n18124;
  wire u2__abc_44228_n18125;
  wire u2__abc_44228_n18126;
  wire u2__abc_44228_n18127;
  wire u2__abc_44228_n18128;
  wire u2__abc_44228_n18129;
  wire u2__abc_44228_n18130;
  wire u2__abc_44228_n18131;
  wire u2__abc_44228_n18132;
  wire u2__abc_44228_n18133;
  wire u2__abc_44228_n18135;
  wire u2__abc_44228_n18136;
  wire u2__abc_44228_n18137;
  wire u2__abc_44228_n18138;
  wire u2__abc_44228_n18139;
  wire u2__abc_44228_n18140;
  wire u2__abc_44228_n18141;
  wire u2__abc_44228_n18142;
  wire u2__abc_44228_n18143;
  wire u2__abc_44228_n18144;
  wire u2__abc_44228_n18145;
  wire u2__abc_44228_n18147;
  wire u2__abc_44228_n18148;
  wire u2__abc_44228_n18149;
  wire u2__abc_44228_n18150;
  wire u2__abc_44228_n18151;
  wire u2__abc_44228_n18152;
  wire u2__abc_44228_n18153;
  wire u2__abc_44228_n18154;
  wire u2__abc_44228_n18155;
  wire u2__abc_44228_n18156;
  wire u2__abc_44228_n18157;
  wire u2__abc_44228_n18159;
  wire u2__abc_44228_n18160;
  wire u2__abc_44228_n18161;
  wire u2__abc_44228_n18162;
  wire u2__abc_44228_n18163;
  wire u2__abc_44228_n18164;
  wire u2__abc_44228_n18165;
  wire u2__abc_44228_n18166;
  wire u2__abc_44228_n18167;
  wire u2__abc_44228_n18168;
  wire u2__abc_44228_n18169;
  wire u2__abc_44228_n18171;
  wire u2__abc_44228_n18172;
  wire u2__abc_44228_n18173;
  wire u2__abc_44228_n18174;
  wire u2__abc_44228_n18175;
  wire u2__abc_44228_n18176;
  wire u2__abc_44228_n18177;
  wire u2__abc_44228_n18178;
  wire u2__abc_44228_n18179;
  wire u2__abc_44228_n18180;
  wire u2__abc_44228_n18181;
  wire u2__abc_44228_n18183;
  wire u2__abc_44228_n18184;
  wire u2__abc_44228_n18185;
  wire u2__abc_44228_n18186;
  wire u2__abc_44228_n18187;
  wire u2__abc_44228_n18188;
  wire u2__abc_44228_n18189;
  wire u2__abc_44228_n18190;
  wire u2__abc_44228_n18191;
  wire u2__abc_44228_n18192;
  wire u2__abc_44228_n18193;
  wire u2__abc_44228_n18195;
  wire u2__abc_44228_n18196;
  wire u2__abc_44228_n18197;
  wire u2__abc_44228_n18198;
  wire u2__abc_44228_n18199;
  wire u2__abc_44228_n18200;
  wire u2__abc_44228_n18201;
  wire u2__abc_44228_n18202;
  wire u2__abc_44228_n18203;
  wire u2__abc_44228_n18204;
  wire u2__abc_44228_n18205;
  wire u2__abc_44228_n18207;
  wire u2__abc_44228_n18208;
  wire u2__abc_44228_n18209;
  wire u2__abc_44228_n18210;
  wire u2__abc_44228_n18211;
  wire u2__abc_44228_n18212;
  wire u2__abc_44228_n18213;
  wire u2__abc_44228_n18214;
  wire u2__abc_44228_n18215;
  wire u2__abc_44228_n18216;
  wire u2__abc_44228_n18217;
  wire u2__abc_44228_n18219;
  wire u2__abc_44228_n18220;
  wire u2__abc_44228_n18221;
  wire u2__abc_44228_n18222;
  wire u2__abc_44228_n18223;
  wire u2__abc_44228_n18224;
  wire u2__abc_44228_n18225;
  wire u2__abc_44228_n18226;
  wire u2__abc_44228_n18227;
  wire u2__abc_44228_n18228;
  wire u2__abc_44228_n18229;
  wire u2__abc_44228_n18231;
  wire u2__abc_44228_n18232;
  wire u2__abc_44228_n18233;
  wire u2__abc_44228_n18234;
  wire u2__abc_44228_n18235;
  wire u2__abc_44228_n18236;
  wire u2__abc_44228_n18237;
  wire u2__abc_44228_n18238;
  wire u2__abc_44228_n18239;
  wire u2__abc_44228_n18240;
  wire u2__abc_44228_n18241;
  wire u2__abc_44228_n18243;
  wire u2__abc_44228_n18244;
  wire u2__abc_44228_n18245;
  wire u2__abc_44228_n18246;
  wire u2__abc_44228_n18247;
  wire u2__abc_44228_n18248;
  wire u2__abc_44228_n18249;
  wire u2__abc_44228_n18250;
  wire u2__abc_44228_n18251;
  wire u2__abc_44228_n18252;
  wire u2__abc_44228_n18253;
  wire u2__abc_44228_n18255;
  wire u2__abc_44228_n18256;
  wire u2__abc_44228_n18257;
  wire u2__abc_44228_n18258;
  wire u2__abc_44228_n18259;
  wire u2__abc_44228_n18260;
  wire u2__abc_44228_n18261;
  wire u2__abc_44228_n18262;
  wire u2__abc_44228_n18263;
  wire u2__abc_44228_n18264;
  wire u2__abc_44228_n18265;
  wire u2__abc_44228_n18267;
  wire u2__abc_44228_n18268;
  wire u2__abc_44228_n18269;
  wire u2__abc_44228_n18270;
  wire u2__abc_44228_n18271;
  wire u2__abc_44228_n18272;
  wire u2__abc_44228_n18273;
  wire u2__abc_44228_n18274;
  wire u2__abc_44228_n18275;
  wire u2__abc_44228_n18276;
  wire u2__abc_44228_n18277;
  wire u2__abc_44228_n18279;
  wire u2__abc_44228_n18280;
  wire u2__abc_44228_n18281;
  wire u2__abc_44228_n18282;
  wire u2__abc_44228_n18283;
  wire u2__abc_44228_n18284;
  wire u2__abc_44228_n18285;
  wire u2__abc_44228_n18286;
  wire u2__abc_44228_n18287;
  wire u2__abc_44228_n18288;
  wire u2__abc_44228_n18289;
  wire u2__abc_44228_n18291;
  wire u2__abc_44228_n18292;
  wire u2__abc_44228_n18293;
  wire u2__abc_44228_n18294;
  wire u2__abc_44228_n18295;
  wire u2__abc_44228_n18296;
  wire u2__abc_44228_n18297;
  wire u2__abc_44228_n18298;
  wire u2__abc_44228_n18299;
  wire u2__abc_44228_n18300;
  wire u2__abc_44228_n18301;
  wire u2__abc_44228_n18303;
  wire u2__abc_44228_n18304;
  wire u2__abc_44228_n18305;
  wire u2__abc_44228_n18306;
  wire u2__abc_44228_n18307;
  wire u2__abc_44228_n18308;
  wire u2__abc_44228_n18309;
  wire u2__abc_44228_n18310;
  wire u2__abc_44228_n18311;
  wire u2__abc_44228_n18312;
  wire u2__abc_44228_n18313;
  wire u2__abc_44228_n18315;
  wire u2__abc_44228_n18316;
  wire u2__abc_44228_n18317;
  wire u2__abc_44228_n18318;
  wire u2__abc_44228_n18319;
  wire u2__abc_44228_n18320;
  wire u2__abc_44228_n18321;
  wire u2__abc_44228_n18322;
  wire u2__abc_44228_n18323;
  wire u2__abc_44228_n18324;
  wire u2__abc_44228_n18325;
  wire u2__abc_44228_n18327;
  wire u2__abc_44228_n18328;
  wire u2__abc_44228_n18329;
  wire u2__abc_44228_n18330;
  wire u2__abc_44228_n18331;
  wire u2__abc_44228_n18332;
  wire u2__abc_44228_n18333;
  wire u2__abc_44228_n18334;
  wire u2__abc_44228_n18335;
  wire u2__abc_44228_n18336;
  wire u2__abc_44228_n18337;
  wire u2__abc_44228_n18339;
  wire u2__abc_44228_n18340;
  wire u2__abc_44228_n18341;
  wire u2__abc_44228_n18342;
  wire u2__abc_44228_n18343;
  wire u2__abc_44228_n18344;
  wire u2__abc_44228_n18345;
  wire u2__abc_44228_n18346;
  wire u2__abc_44228_n18347;
  wire u2__abc_44228_n18348;
  wire u2__abc_44228_n18349;
  wire u2__abc_44228_n18351;
  wire u2__abc_44228_n18352;
  wire u2__abc_44228_n18353;
  wire u2__abc_44228_n18354;
  wire u2__abc_44228_n18355;
  wire u2__abc_44228_n18356;
  wire u2__abc_44228_n18357;
  wire u2__abc_44228_n18358;
  wire u2__abc_44228_n18359;
  wire u2__abc_44228_n18360;
  wire u2__abc_44228_n18361;
  wire u2__abc_44228_n18363;
  wire u2__abc_44228_n18364;
  wire u2__abc_44228_n18365;
  wire u2__abc_44228_n18366;
  wire u2__abc_44228_n18367;
  wire u2__abc_44228_n18368;
  wire u2__abc_44228_n18369;
  wire u2__abc_44228_n18370;
  wire u2__abc_44228_n18371;
  wire u2__abc_44228_n18372;
  wire u2__abc_44228_n18373;
  wire u2__abc_44228_n18375;
  wire u2__abc_44228_n18376;
  wire u2__abc_44228_n18377;
  wire u2__abc_44228_n18378;
  wire u2__abc_44228_n18379;
  wire u2__abc_44228_n18380;
  wire u2__abc_44228_n18381;
  wire u2__abc_44228_n18382;
  wire u2__abc_44228_n18383;
  wire u2__abc_44228_n18384;
  wire u2__abc_44228_n18385;
  wire u2__abc_44228_n18387;
  wire u2__abc_44228_n18388;
  wire u2__abc_44228_n18389;
  wire u2__abc_44228_n18390;
  wire u2__abc_44228_n18391;
  wire u2__abc_44228_n18392;
  wire u2__abc_44228_n18393;
  wire u2__abc_44228_n18394;
  wire u2__abc_44228_n18395;
  wire u2__abc_44228_n18396;
  wire u2__abc_44228_n18397;
  wire u2__abc_44228_n18399;
  wire u2__abc_44228_n18400;
  wire u2__abc_44228_n18401;
  wire u2__abc_44228_n18402;
  wire u2__abc_44228_n18403;
  wire u2__abc_44228_n18404;
  wire u2__abc_44228_n18405;
  wire u2__abc_44228_n18406;
  wire u2__abc_44228_n18407;
  wire u2__abc_44228_n18408;
  wire u2__abc_44228_n18409;
  wire u2__abc_44228_n18411;
  wire u2__abc_44228_n18412;
  wire u2__abc_44228_n18413;
  wire u2__abc_44228_n18414;
  wire u2__abc_44228_n18415;
  wire u2__abc_44228_n18416;
  wire u2__abc_44228_n18417;
  wire u2__abc_44228_n18418;
  wire u2__abc_44228_n18419;
  wire u2__abc_44228_n18420;
  wire u2__abc_44228_n18421;
  wire u2__abc_44228_n18423;
  wire u2__abc_44228_n18424;
  wire u2__abc_44228_n18425;
  wire u2__abc_44228_n18426;
  wire u2__abc_44228_n18427;
  wire u2__abc_44228_n18428;
  wire u2__abc_44228_n18429;
  wire u2__abc_44228_n18430;
  wire u2__abc_44228_n18431;
  wire u2__abc_44228_n18432;
  wire u2__abc_44228_n18433;
  wire u2__abc_44228_n18435;
  wire u2__abc_44228_n18436;
  wire u2__abc_44228_n18437;
  wire u2__abc_44228_n18438;
  wire u2__abc_44228_n18439;
  wire u2__abc_44228_n18440;
  wire u2__abc_44228_n18441;
  wire u2__abc_44228_n18442;
  wire u2__abc_44228_n18443;
  wire u2__abc_44228_n18444;
  wire u2__abc_44228_n18445;
  wire u2__abc_44228_n18447;
  wire u2__abc_44228_n18448;
  wire u2__abc_44228_n18449;
  wire u2__abc_44228_n18450;
  wire u2__abc_44228_n18451;
  wire u2__abc_44228_n18452;
  wire u2__abc_44228_n18453;
  wire u2__abc_44228_n18454;
  wire u2__abc_44228_n18455;
  wire u2__abc_44228_n18456;
  wire u2__abc_44228_n18457;
  wire u2__abc_44228_n18459;
  wire u2__abc_44228_n18460;
  wire u2__abc_44228_n18461;
  wire u2__abc_44228_n18462;
  wire u2__abc_44228_n18463;
  wire u2__abc_44228_n18464;
  wire u2__abc_44228_n18465;
  wire u2__abc_44228_n18466;
  wire u2__abc_44228_n18467;
  wire u2__abc_44228_n18468;
  wire u2__abc_44228_n18469;
  wire u2__abc_44228_n18471;
  wire u2__abc_44228_n18472;
  wire u2__abc_44228_n18473;
  wire u2__abc_44228_n18474;
  wire u2__abc_44228_n18475;
  wire u2__abc_44228_n18476;
  wire u2__abc_44228_n18477;
  wire u2__abc_44228_n18478;
  wire u2__abc_44228_n18479;
  wire u2__abc_44228_n18480;
  wire u2__abc_44228_n18481;
  wire u2__abc_44228_n18483;
  wire u2__abc_44228_n18484;
  wire u2__abc_44228_n18485;
  wire u2__abc_44228_n18486;
  wire u2__abc_44228_n18487;
  wire u2__abc_44228_n18488;
  wire u2__abc_44228_n18489;
  wire u2__abc_44228_n18490;
  wire u2__abc_44228_n18491;
  wire u2__abc_44228_n18492;
  wire u2__abc_44228_n18493;
  wire u2__abc_44228_n18495;
  wire u2__abc_44228_n18496;
  wire u2__abc_44228_n18497;
  wire u2__abc_44228_n18498;
  wire u2__abc_44228_n18499;
  wire u2__abc_44228_n18500;
  wire u2__abc_44228_n18501;
  wire u2__abc_44228_n18502;
  wire u2__abc_44228_n18503;
  wire u2__abc_44228_n18504;
  wire u2__abc_44228_n18505;
  wire u2__abc_44228_n18507;
  wire u2__abc_44228_n18508;
  wire u2__abc_44228_n18509;
  wire u2__abc_44228_n18510;
  wire u2__abc_44228_n18511;
  wire u2__abc_44228_n18512;
  wire u2__abc_44228_n18513;
  wire u2__abc_44228_n18514;
  wire u2__abc_44228_n18515;
  wire u2__abc_44228_n18516;
  wire u2__abc_44228_n18517;
  wire u2__abc_44228_n18519;
  wire u2__abc_44228_n18520;
  wire u2__abc_44228_n18521;
  wire u2__abc_44228_n18522;
  wire u2__abc_44228_n18523;
  wire u2__abc_44228_n18524;
  wire u2__abc_44228_n18525;
  wire u2__abc_44228_n18526;
  wire u2__abc_44228_n18527;
  wire u2__abc_44228_n18528;
  wire u2__abc_44228_n18529;
  wire u2__abc_44228_n18531;
  wire u2__abc_44228_n18532;
  wire u2__abc_44228_n18533;
  wire u2__abc_44228_n18534;
  wire u2__abc_44228_n18535;
  wire u2__abc_44228_n18536;
  wire u2__abc_44228_n18537;
  wire u2__abc_44228_n18538;
  wire u2__abc_44228_n18539;
  wire u2__abc_44228_n18540;
  wire u2__abc_44228_n18541;
  wire u2__abc_44228_n18543;
  wire u2__abc_44228_n18544;
  wire u2__abc_44228_n18545;
  wire u2__abc_44228_n18546;
  wire u2__abc_44228_n18547;
  wire u2__abc_44228_n18548;
  wire u2__abc_44228_n18549;
  wire u2__abc_44228_n18550;
  wire u2__abc_44228_n18551;
  wire u2__abc_44228_n18552;
  wire u2__abc_44228_n18553;
  wire u2__abc_44228_n18555;
  wire u2__abc_44228_n18556;
  wire u2__abc_44228_n18557;
  wire u2__abc_44228_n18558;
  wire u2__abc_44228_n18559;
  wire u2__abc_44228_n18560;
  wire u2__abc_44228_n18561;
  wire u2__abc_44228_n18562;
  wire u2__abc_44228_n18563;
  wire u2__abc_44228_n18564;
  wire u2__abc_44228_n18565;
  wire u2__abc_44228_n18567;
  wire u2__abc_44228_n18568;
  wire u2__abc_44228_n18569;
  wire u2__abc_44228_n18570;
  wire u2__abc_44228_n18571;
  wire u2__abc_44228_n18572;
  wire u2__abc_44228_n18573;
  wire u2__abc_44228_n18574;
  wire u2__abc_44228_n18575;
  wire u2__abc_44228_n18576;
  wire u2__abc_44228_n18577;
  wire u2__abc_44228_n18579;
  wire u2__abc_44228_n18580;
  wire u2__abc_44228_n18581;
  wire u2__abc_44228_n18582;
  wire u2__abc_44228_n18583;
  wire u2__abc_44228_n18584;
  wire u2__abc_44228_n18585;
  wire u2__abc_44228_n18586;
  wire u2__abc_44228_n18587;
  wire u2__abc_44228_n18588;
  wire u2__abc_44228_n18589;
  wire u2__abc_44228_n18591;
  wire u2__abc_44228_n18592;
  wire u2__abc_44228_n18593;
  wire u2__abc_44228_n18594;
  wire u2__abc_44228_n18595;
  wire u2__abc_44228_n18596;
  wire u2__abc_44228_n18597;
  wire u2__abc_44228_n18598;
  wire u2__abc_44228_n18599;
  wire u2__abc_44228_n18600;
  wire u2__abc_44228_n18601;
  wire u2__abc_44228_n18603;
  wire u2__abc_44228_n18604;
  wire u2__abc_44228_n18605;
  wire u2__abc_44228_n18606;
  wire u2__abc_44228_n18607;
  wire u2__abc_44228_n18608;
  wire u2__abc_44228_n18609;
  wire u2__abc_44228_n18610;
  wire u2__abc_44228_n18611;
  wire u2__abc_44228_n18612;
  wire u2__abc_44228_n18613;
  wire u2__abc_44228_n18615;
  wire u2__abc_44228_n18616;
  wire u2__abc_44228_n18617;
  wire u2__abc_44228_n18618;
  wire u2__abc_44228_n18619;
  wire u2__abc_44228_n18620;
  wire u2__abc_44228_n18621;
  wire u2__abc_44228_n18622;
  wire u2__abc_44228_n18623;
  wire u2__abc_44228_n18624;
  wire u2__abc_44228_n18625;
  wire u2__abc_44228_n18627;
  wire u2__abc_44228_n18628;
  wire u2__abc_44228_n18629;
  wire u2__abc_44228_n18630;
  wire u2__abc_44228_n18631;
  wire u2__abc_44228_n18632;
  wire u2__abc_44228_n18633;
  wire u2__abc_44228_n18634;
  wire u2__abc_44228_n18635;
  wire u2__abc_44228_n18636;
  wire u2__abc_44228_n18637;
  wire u2__abc_44228_n18639;
  wire u2__abc_44228_n18640;
  wire u2__abc_44228_n18641;
  wire u2__abc_44228_n18642;
  wire u2__abc_44228_n18643;
  wire u2__abc_44228_n18644;
  wire u2__abc_44228_n18645;
  wire u2__abc_44228_n18646;
  wire u2__abc_44228_n18647;
  wire u2__abc_44228_n18648;
  wire u2__abc_44228_n18649;
  wire u2__abc_44228_n18651;
  wire u2__abc_44228_n18652;
  wire u2__abc_44228_n18653;
  wire u2__abc_44228_n18654;
  wire u2__abc_44228_n18655;
  wire u2__abc_44228_n18656;
  wire u2__abc_44228_n18657;
  wire u2__abc_44228_n18658;
  wire u2__abc_44228_n18659;
  wire u2__abc_44228_n18660;
  wire u2__abc_44228_n18661;
  wire u2__abc_44228_n18663;
  wire u2__abc_44228_n18664;
  wire u2__abc_44228_n18665;
  wire u2__abc_44228_n18666;
  wire u2__abc_44228_n18667;
  wire u2__abc_44228_n18668;
  wire u2__abc_44228_n18669;
  wire u2__abc_44228_n18670;
  wire u2__abc_44228_n18671;
  wire u2__abc_44228_n18672;
  wire u2__abc_44228_n18673;
  wire u2__abc_44228_n18675;
  wire u2__abc_44228_n18676;
  wire u2__abc_44228_n18677;
  wire u2__abc_44228_n18678;
  wire u2__abc_44228_n18679;
  wire u2__abc_44228_n18680;
  wire u2__abc_44228_n18681;
  wire u2__abc_44228_n18682;
  wire u2__abc_44228_n18683;
  wire u2__abc_44228_n18684;
  wire u2__abc_44228_n18685;
  wire u2__abc_44228_n18687;
  wire u2__abc_44228_n18688;
  wire u2__abc_44228_n18689;
  wire u2__abc_44228_n18690;
  wire u2__abc_44228_n18691;
  wire u2__abc_44228_n18692;
  wire u2__abc_44228_n18693;
  wire u2__abc_44228_n18694;
  wire u2__abc_44228_n18695;
  wire u2__abc_44228_n18696;
  wire u2__abc_44228_n18697;
  wire u2__abc_44228_n18699;
  wire u2__abc_44228_n18700;
  wire u2__abc_44228_n18701;
  wire u2__abc_44228_n18702;
  wire u2__abc_44228_n18703;
  wire u2__abc_44228_n18704;
  wire u2__abc_44228_n18705;
  wire u2__abc_44228_n18706;
  wire u2__abc_44228_n18707;
  wire u2__abc_44228_n18708;
  wire u2__abc_44228_n18709;
  wire u2__abc_44228_n18711;
  wire u2__abc_44228_n18712;
  wire u2__abc_44228_n18713;
  wire u2__abc_44228_n18714;
  wire u2__abc_44228_n18715;
  wire u2__abc_44228_n18716;
  wire u2__abc_44228_n18717;
  wire u2__abc_44228_n18718;
  wire u2__abc_44228_n18719;
  wire u2__abc_44228_n18720;
  wire u2__abc_44228_n18721;
  wire u2__abc_44228_n18723;
  wire u2__abc_44228_n18724;
  wire u2__abc_44228_n18725;
  wire u2__abc_44228_n18726;
  wire u2__abc_44228_n18727;
  wire u2__abc_44228_n18728;
  wire u2__abc_44228_n18729;
  wire u2__abc_44228_n18730;
  wire u2__abc_44228_n18731;
  wire u2__abc_44228_n18732;
  wire u2__abc_44228_n18733;
  wire u2__abc_44228_n18735;
  wire u2__abc_44228_n18736;
  wire u2__abc_44228_n18737;
  wire u2__abc_44228_n18738;
  wire u2__abc_44228_n18739;
  wire u2__abc_44228_n18740;
  wire u2__abc_44228_n18741;
  wire u2__abc_44228_n18742;
  wire u2__abc_44228_n18743;
  wire u2__abc_44228_n18744;
  wire u2__abc_44228_n18745;
  wire u2__abc_44228_n18747;
  wire u2__abc_44228_n18748;
  wire u2__abc_44228_n18749;
  wire u2__abc_44228_n18750;
  wire u2__abc_44228_n18751;
  wire u2__abc_44228_n18752;
  wire u2__abc_44228_n18753;
  wire u2__abc_44228_n18754;
  wire u2__abc_44228_n18755;
  wire u2__abc_44228_n18756;
  wire u2__abc_44228_n18757;
  wire u2__abc_44228_n18759;
  wire u2__abc_44228_n18760;
  wire u2__abc_44228_n18761;
  wire u2__abc_44228_n18762;
  wire u2__abc_44228_n18763;
  wire u2__abc_44228_n18764;
  wire u2__abc_44228_n18765;
  wire u2__abc_44228_n18766;
  wire u2__abc_44228_n18767;
  wire u2__abc_44228_n18768;
  wire u2__abc_44228_n18769;
  wire u2__abc_44228_n18771;
  wire u2__abc_44228_n18772;
  wire u2__abc_44228_n18773;
  wire u2__abc_44228_n18774;
  wire u2__abc_44228_n18775;
  wire u2__abc_44228_n18776;
  wire u2__abc_44228_n18777;
  wire u2__abc_44228_n18778;
  wire u2__abc_44228_n18779;
  wire u2__abc_44228_n18780;
  wire u2__abc_44228_n18781;
  wire u2__abc_44228_n18783;
  wire u2__abc_44228_n18784;
  wire u2__abc_44228_n18785;
  wire u2__abc_44228_n18786;
  wire u2__abc_44228_n18787;
  wire u2__abc_44228_n18788;
  wire u2__abc_44228_n18789;
  wire u2__abc_44228_n18790;
  wire u2__abc_44228_n18791;
  wire u2__abc_44228_n18792;
  wire u2__abc_44228_n18793;
  wire u2__abc_44228_n18795;
  wire u2__abc_44228_n18796;
  wire u2__abc_44228_n18797;
  wire u2__abc_44228_n18798;
  wire u2__abc_44228_n18799;
  wire u2__abc_44228_n18800;
  wire u2__abc_44228_n18801;
  wire u2__abc_44228_n18802;
  wire u2__abc_44228_n18803;
  wire u2__abc_44228_n18804;
  wire u2__abc_44228_n18805;
  wire u2__abc_44228_n18807;
  wire u2__abc_44228_n18808;
  wire u2__abc_44228_n18809;
  wire u2__abc_44228_n18810;
  wire u2__abc_44228_n18811;
  wire u2__abc_44228_n18812;
  wire u2__abc_44228_n18813;
  wire u2__abc_44228_n18814;
  wire u2__abc_44228_n18815;
  wire u2__abc_44228_n18816;
  wire u2__abc_44228_n18817;
  wire u2__abc_44228_n18819;
  wire u2__abc_44228_n18820;
  wire u2__abc_44228_n18821;
  wire u2__abc_44228_n18822;
  wire u2__abc_44228_n18823;
  wire u2__abc_44228_n18824;
  wire u2__abc_44228_n18825;
  wire u2__abc_44228_n18826;
  wire u2__abc_44228_n18827;
  wire u2__abc_44228_n18828;
  wire u2__abc_44228_n18829;
  wire u2__abc_44228_n18831;
  wire u2__abc_44228_n18832;
  wire u2__abc_44228_n18833;
  wire u2__abc_44228_n18834;
  wire u2__abc_44228_n18835;
  wire u2__abc_44228_n18836;
  wire u2__abc_44228_n18837;
  wire u2__abc_44228_n18838;
  wire u2__abc_44228_n18839;
  wire u2__abc_44228_n18840;
  wire u2__abc_44228_n18841;
  wire u2__abc_44228_n18843;
  wire u2__abc_44228_n18844;
  wire u2__abc_44228_n18845;
  wire u2__abc_44228_n18846;
  wire u2__abc_44228_n18847;
  wire u2__abc_44228_n18848;
  wire u2__abc_44228_n18849;
  wire u2__abc_44228_n18850;
  wire u2__abc_44228_n18851;
  wire u2__abc_44228_n18852;
  wire u2__abc_44228_n18853;
  wire u2__abc_44228_n18855;
  wire u2__abc_44228_n18856;
  wire u2__abc_44228_n18857;
  wire u2__abc_44228_n18858;
  wire u2__abc_44228_n18859;
  wire u2__abc_44228_n18860;
  wire u2__abc_44228_n18861;
  wire u2__abc_44228_n18862;
  wire u2__abc_44228_n18863;
  wire u2__abc_44228_n18864;
  wire u2__abc_44228_n18865;
  wire u2__abc_44228_n18867;
  wire u2__abc_44228_n18868;
  wire u2__abc_44228_n18869;
  wire u2__abc_44228_n18870;
  wire u2__abc_44228_n18871;
  wire u2__abc_44228_n18872;
  wire u2__abc_44228_n18873;
  wire u2__abc_44228_n18874;
  wire u2__abc_44228_n18875;
  wire u2__abc_44228_n18876;
  wire u2__abc_44228_n18877;
  wire u2__abc_44228_n18879;
  wire u2__abc_44228_n18880;
  wire u2__abc_44228_n18881;
  wire u2__abc_44228_n18882;
  wire u2__abc_44228_n18883;
  wire u2__abc_44228_n18884;
  wire u2__abc_44228_n18885;
  wire u2__abc_44228_n18886;
  wire u2__abc_44228_n18887;
  wire u2__abc_44228_n18888;
  wire u2__abc_44228_n18889;
  wire u2__abc_44228_n18891;
  wire u2__abc_44228_n18892;
  wire u2__abc_44228_n18893;
  wire u2__abc_44228_n18894;
  wire u2__abc_44228_n18895;
  wire u2__abc_44228_n18896;
  wire u2__abc_44228_n18897;
  wire u2__abc_44228_n18898;
  wire u2__abc_44228_n18899;
  wire u2__abc_44228_n18900;
  wire u2__abc_44228_n18901;
  wire u2__abc_44228_n18903;
  wire u2__abc_44228_n18904;
  wire u2__abc_44228_n18905;
  wire u2__abc_44228_n18906;
  wire u2__abc_44228_n18907;
  wire u2__abc_44228_n18908;
  wire u2__abc_44228_n18909;
  wire u2__abc_44228_n18910;
  wire u2__abc_44228_n18911;
  wire u2__abc_44228_n18912;
  wire u2__abc_44228_n18913;
  wire u2__abc_44228_n18915;
  wire u2__abc_44228_n18916;
  wire u2__abc_44228_n18917;
  wire u2__abc_44228_n18918;
  wire u2__abc_44228_n18919;
  wire u2__abc_44228_n18920;
  wire u2__abc_44228_n18921;
  wire u2__abc_44228_n18922;
  wire u2__abc_44228_n18923;
  wire u2__abc_44228_n18924;
  wire u2__abc_44228_n18925;
  wire u2__abc_44228_n18927;
  wire u2__abc_44228_n18928;
  wire u2__abc_44228_n18929;
  wire u2__abc_44228_n18930;
  wire u2__abc_44228_n18931;
  wire u2__abc_44228_n18932;
  wire u2__abc_44228_n18933;
  wire u2__abc_44228_n18934;
  wire u2__abc_44228_n18935;
  wire u2__abc_44228_n18936;
  wire u2__abc_44228_n18937;
  wire u2__abc_44228_n18939;
  wire u2__abc_44228_n18940;
  wire u2__abc_44228_n18941;
  wire u2__abc_44228_n18942;
  wire u2__abc_44228_n18943;
  wire u2__abc_44228_n18944;
  wire u2__abc_44228_n18945;
  wire u2__abc_44228_n18946;
  wire u2__abc_44228_n18947;
  wire u2__abc_44228_n18948;
  wire u2__abc_44228_n18949;
  wire u2__abc_44228_n18951;
  wire u2__abc_44228_n18952;
  wire u2__abc_44228_n18953;
  wire u2__abc_44228_n18954;
  wire u2__abc_44228_n18955;
  wire u2__abc_44228_n18956;
  wire u2__abc_44228_n18957;
  wire u2__abc_44228_n18958;
  wire u2__abc_44228_n18959;
  wire u2__abc_44228_n18960;
  wire u2__abc_44228_n18961;
  wire u2__abc_44228_n18963;
  wire u2__abc_44228_n18964;
  wire u2__abc_44228_n18965;
  wire u2__abc_44228_n18966;
  wire u2__abc_44228_n18967;
  wire u2__abc_44228_n18968;
  wire u2__abc_44228_n18969;
  wire u2__abc_44228_n18970;
  wire u2__abc_44228_n18971;
  wire u2__abc_44228_n18972;
  wire u2__abc_44228_n18973;
  wire u2__abc_44228_n18975;
  wire u2__abc_44228_n18976;
  wire u2__abc_44228_n18977;
  wire u2__abc_44228_n18978;
  wire u2__abc_44228_n18979;
  wire u2__abc_44228_n18980;
  wire u2__abc_44228_n18981;
  wire u2__abc_44228_n18982;
  wire u2__abc_44228_n18983;
  wire u2__abc_44228_n18984;
  wire u2__abc_44228_n18985;
  wire u2__abc_44228_n18987;
  wire u2__abc_44228_n18988;
  wire u2__abc_44228_n18989;
  wire u2__abc_44228_n18990;
  wire u2__abc_44228_n18991;
  wire u2__abc_44228_n18992;
  wire u2__abc_44228_n18993;
  wire u2__abc_44228_n18994;
  wire u2__abc_44228_n18995;
  wire u2__abc_44228_n18996;
  wire u2__abc_44228_n18997;
  wire u2__abc_44228_n18999;
  wire u2__abc_44228_n19000;
  wire u2__abc_44228_n19001;
  wire u2__abc_44228_n19002;
  wire u2__abc_44228_n19003;
  wire u2__abc_44228_n19004;
  wire u2__abc_44228_n19005;
  wire u2__abc_44228_n19006;
  wire u2__abc_44228_n19007;
  wire u2__abc_44228_n19008;
  wire u2__abc_44228_n19009;
  wire u2__abc_44228_n19011;
  wire u2__abc_44228_n19012;
  wire u2__abc_44228_n19013;
  wire u2__abc_44228_n19014;
  wire u2__abc_44228_n19015;
  wire u2__abc_44228_n19016;
  wire u2__abc_44228_n19017;
  wire u2__abc_44228_n19018;
  wire u2__abc_44228_n19019;
  wire u2__abc_44228_n19020;
  wire u2__abc_44228_n19021;
  wire u2__abc_44228_n19023;
  wire u2__abc_44228_n19024;
  wire u2__abc_44228_n19025;
  wire u2__abc_44228_n19026;
  wire u2__abc_44228_n19027;
  wire u2__abc_44228_n19028;
  wire u2__abc_44228_n19029;
  wire u2__abc_44228_n19030;
  wire u2__abc_44228_n19031;
  wire u2__abc_44228_n19032;
  wire u2__abc_44228_n19033;
  wire u2__abc_44228_n19035;
  wire u2__abc_44228_n19036;
  wire u2__abc_44228_n19037;
  wire u2__abc_44228_n19038;
  wire u2__abc_44228_n19039;
  wire u2__abc_44228_n19040;
  wire u2__abc_44228_n19041;
  wire u2__abc_44228_n19042;
  wire u2__abc_44228_n19043;
  wire u2__abc_44228_n19044;
  wire u2__abc_44228_n19045;
  wire u2__abc_44228_n19047;
  wire u2__abc_44228_n19048;
  wire u2__abc_44228_n19049;
  wire u2__abc_44228_n19050;
  wire u2__abc_44228_n19051;
  wire u2__abc_44228_n19052;
  wire u2__abc_44228_n19053;
  wire u2__abc_44228_n19054;
  wire u2__abc_44228_n19055;
  wire u2__abc_44228_n19056;
  wire u2__abc_44228_n19057;
  wire u2__abc_44228_n19059;
  wire u2__abc_44228_n19060;
  wire u2__abc_44228_n19061;
  wire u2__abc_44228_n19062;
  wire u2__abc_44228_n19063;
  wire u2__abc_44228_n19064;
  wire u2__abc_44228_n19065;
  wire u2__abc_44228_n19066;
  wire u2__abc_44228_n19067;
  wire u2__abc_44228_n19068;
  wire u2__abc_44228_n19069;
  wire u2__abc_44228_n19071;
  wire u2__abc_44228_n19072;
  wire u2__abc_44228_n19073;
  wire u2__abc_44228_n19074;
  wire u2__abc_44228_n19075;
  wire u2__abc_44228_n19076;
  wire u2__abc_44228_n19077;
  wire u2__abc_44228_n19078;
  wire u2__abc_44228_n19079;
  wire u2__abc_44228_n19080;
  wire u2__abc_44228_n19081;
  wire u2__abc_44228_n19083;
  wire u2__abc_44228_n19084;
  wire u2__abc_44228_n19085;
  wire u2__abc_44228_n19086;
  wire u2__abc_44228_n19087;
  wire u2__abc_44228_n19088;
  wire u2__abc_44228_n19089;
  wire u2__abc_44228_n19090;
  wire u2__abc_44228_n19091;
  wire u2__abc_44228_n19092;
  wire u2__abc_44228_n19093;
  wire u2__abc_44228_n19095;
  wire u2__abc_44228_n19096;
  wire u2__abc_44228_n19097;
  wire u2__abc_44228_n19098;
  wire u2__abc_44228_n19099;
  wire u2__abc_44228_n19100;
  wire u2__abc_44228_n19101;
  wire u2__abc_44228_n19102;
  wire u2__abc_44228_n19103;
  wire u2__abc_44228_n19104;
  wire u2__abc_44228_n19105;
  wire u2__abc_44228_n19107;
  wire u2__abc_44228_n19108;
  wire u2__abc_44228_n19109;
  wire u2__abc_44228_n19110;
  wire u2__abc_44228_n19111;
  wire u2__abc_44228_n19112;
  wire u2__abc_44228_n19113;
  wire u2__abc_44228_n19114;
  wire u2__abc_44228_n19115;
  wire u2__abc_44228_n19116;
  wire u2__abc_44228_n19117;
  wire u2__abc_44228_n19119;
  wire u2__abc_44228_n19120;
  wire u2__abc_44228_n19121;
  wire u2__abc_44228_n19122;
  wire u2__abc_44228_n19123;
  wire u2__abc_44228_n19124;
  wire u2__abc_44228_n19125;
  wire u2__abc_44228_n19126;
  wire u2__abc_44228_n19127;
  wire u2__abc_44228_n19128;
  wire u2__abc_44228_n19129;
  wire u2__abc_44228_n19131;
  wire u2__abc_44228_n19132;
  wire u2__abc_44228_n19133;
  wire u2__abc_44228_n19134;
  wire u2__abc_44228_n19135;
  wire u2__abc_44228_n19136;
  wire u2__abc_44228_n19137;
  wire u2__abc_44228_n19138;
  wire u2__abc_44228_n19139;
  wire u2__abc_44228_n19140;
  wire u2__abc_44228_n19141;
  wire u2__abc_44228_n19143;
  wire u2__abc_44228_n19144;
  wire u2__abc_44228_n19145;
  wire u2__abc_44228_n19146;
  wire u2__abc_44228_n19147;
  wire u2__abc_44228_n19148;
  wire u2__abc_44228_n19149;
  wire u2__abc_44228_n19150;
  wire u2__abc_44228_n19151;
  wire u2__abc_44228_n19152;
  wire u2__abc_44228_n19153;
  wire u2__abc_44228_n19155;
  wire u2__abc_44228_n19156;
  wire u2__abc_44228_n19157;
  wire u2__abc_44228_n19158;
  wire u2__abc_44228_n19159;
  wire u2__abc_44228_n19160;
  wire u2__abc_44228_n19161;
  wire u2__abc_44228_n19162;
  wire u2__abc_44228_n19163;
  wire u2__abc_44228_n19164;
  wire u2__abc_44228_n19165;
  wire u2__abc_44228_n19167;
  wire u2__abc_44228_n19168;
  wire u2__abc_44228_n19169;
  wire u2__abc_44228_n19170;
  wire u2__abc_44228_n19171;
  wire u2__abc_44228_n19172;
  wire u2__abc_44228_n19173;
  wire u2__abc_44228_n19174;
  wire u2__abc_44228_n19175;
  wire u2__abc_44228_n19176;
  wire u2__abc_44228_n19177;
  wire u2__abc_44228_n19179;
  wire u2__abc_44228_n19180;
  wire u2__abc_44228_n19181;
  wire u2__abc_44228_n19182;
  wire u2__abc_44228_n19183;
  wire u2__abc_44228_n19184;
  wire u2__abc_44228_n19185;
  wire u2__abc_44228_n19186;
  wire u2__abc_44228_n19187;
  wire u2__abc_44228_n19188;
  wire u2__abc_44228_n19189;
  wire u2__abc_44228_n19191;
  wire u2__abc_44228_n19192;
  wire u2__abc_44228_n19193;
  wire u2__abc_44228_n19194;
  wire u2__abc_44228_n19195;
  wire u2__abc_44228_n19196;
  wire u2__abc_44228_n19197;
  wire u2__abc_44228_n19198;
  wire u2__abc_44228_n19199;
  wire u2__abc_44228_n19200;
  wire u2__abc_44228_n19201;
  wire u2__abc_44228_n19203;
  wire u2__abc_44228_n19204;
  wire u2__abc_44228_n19205;
  wire u2__abc_44228_n19206;
  wire u2__abc_44228_n19207;
  wire u2__abc_44228_n19208;
  wire u2__abc_44228_n19209;
  wire u2__abc_44228_n19210;
  wire u2__abc_44228_n19211;
  wire u2__abc_44228_n19212;
  wire u2__abc_44228_n19213;
  wire u2__abc_44228_n19215;
  wire u2__abc_44228_n19216;
  wire u2__abc_44228_n19217;
  wire u2__abc_44228_n19218;
  wire u2__abc_44228_n19219;
  wire u2__abc_44228_n19220;
  wire u2__abc_44228_n19221;
  wire u2__abc_44228_n19222;
  wire u2__abc_44228_n19223;
  wire u2__abc_44228_n19224;
  wire u2__abc_44228_n19225;
  wire u2__abc_44228_n19227;
  wire u2__abc_44228_n19228;
  wire u2__abc_44228_n19229;
  wire u2__abc_44228_n19230;
  wire u2__abc_44228_n19231;
  wire u2__abc_44228_n19232;
  wire u2__abc_44228_n19233;
  wire u2__abc_44228_n19234;
  wire u2__abc_44228_n19235;
  wire u2__abc_44228_n19236;
  wire u2__abc_44228_n19237;
  wire u2__abc_44228_n19239;
  wire u2__abc_44228_n19240;
  wire u2__abc_44228_n19241;
  wire u2__abc_44228_n19242;
  wire u2__abc_44228_n19243;
  wire u2__abc_44228_n19244;
  wire u2__abc_44228_n19245;
  wire u2__abc_44228_n19246;
  wire u2__abc_44228_n19247;
  wire u2__abc_44228_n19248;
  wire u2__abc_44228_n19249;
  wire u2__abc_44228_n19251;
  wire u2__abc_44228_n19252;
  wire u2__abc_44228_n19253;
  wire u2__abc_44228_n19254;
  wire u2__abc_44228_n19255;
  wire u2__abc_44228_n19256;
  wire u2__abc_44228_n19257;
  wire u2__abc_44228_n19258;
  wire u2__abc_44228_n19259;
  wire u2__abc_44228_n19260;
  wire u2__abc_44228_n19261;
  wire u2__abc_44228_n19263;
  wire u2__abc_44228_n19264;
  wire u2__abc_44228_n19265;
  wire u2__abc_44228_n19266;
  wire u2__abc_44228_n19267;
  wire u2__abc_44228_n19268;
  wire u2__abc_44228_n19269;
  wire u2__abc_44228_n19270;
  wire u2__abc_44228_n19271;
  wire u2__abc_44228_n19272;
  wire u2__abc_44228_n19273;
  wire u2__abc_44228_n19275;
  wire u2__abc_44228_n19276;
  wire u2__abc_44228_n19277;
  wire u2__abc_44228_n19278;
  wire u2__abc_44228_n19279;
  wire u2__abc_44228_n19280;
  wire u2__abc_44228_n19281;
  wire u2__abc_44228_n19282;
  wire u2__abc_44228_n19283;
  wire u2__abc_44228_n19284;
  wire u2__abc_44228_n19285;
  wire u2__abc_44228_n19287;
  wire u2__abc_44228_n19288;
  wire u2__abc_44228_n19289;
  wire u2__abc_44228_n19290;
  wire u2__abc_44228_n19291;
  wire u2__abc_44228_n19292;
  wire u2__abc_44228_n19293;
  wire u2__abc_44228_n19294;
  wire u2__abc_44228_n19295;
  wire u2__abc_44228_n19296;
  wire u2__abc_44228_n19297;
  wire u2__abc_44228_n19299;
  wire u2__abc_44228_n19300;
  wire u2__abc_44228_n19301;
  wire u2__abc_44228_n19302;
  wire u2__abc_44228_n19303;
  wire u2__abc_44228_n19304;
  wire u2__abc_44228_n19305;
  wire u2__abc_44228_n19306;
  wire u2__abc_44228_n19307;
  wire u2__abc_44228_n19308;
  wire u2__abc_44228_n19309;
  wire u2__abc_44228_n19311;
  wire u2__abc_44228_n19312;
  wire u2__abc_44228_n19313;
  wire u2__abc_44228_n19314;
  wire u2__abc_44228_n19315;
  wire u2__abc_44228_n19316;
  wire u2__abc_44228_n19317;
  wire u2__abc_44228_n19318;
  wire u2__abc_44228_n19319;
  wire u2__abc_44228_n19320;
  wire u2__abc_44228_n19321;
  wire u2__abc_44228_n19323;
  wire u2__abc_44228_n19324;
  wire u2__abc_44228_n19325;
  wire u2__abc_44228_n19326;
  wire u2__abc_44228_n19327;
  wire u2__abc_44228_n19328;
  wire u2__abc_44228_n19329;
  wire u2__abc_44228_n19330;
  wire u2__abc_44228_n19331;
  wire u2__abc_44228_n19332;
  wire u2__abc_44228_n19333;
  wire u2__abc_44228_n19335;
  wire u2__abc_44228_n19336;
  wire u2__abc_44228_n19337;
  wire u2__abc_44228_n19338;
  wire u2__abc_44228_n19339;
  wire u2__abc_44228_n19340;
  wire u2__abc_44228_n19341;
  wire u2__abc_44228_n19342;
  wire u2__abc_44228_n19343;
  wire u2__abc_44228_n19344;
  wire u2__abc_44228_n19345;
  wire u2__abc_44228_n19347;
  wire u2__abc_44228_n19348;
  wire u2__abc_44228_n19349;
  wire u2__abc_44228_n19350;
  wire u2__abc_44228_n19351;
  wire u2__abc_44228_n19352;
  wire u2__abc_44228_n19353;
  wire u2__abc_44228_n19354;
  wire u2__abc_44228_n19355;
  wire u2__abc_44228_n19356;
  wire u2__abc_44228_n19357;
  wire u2__abc_44228_n19359;
  wire u2__abc_44228_n19360;
  wire u2__abc_44228_n19361;
  wire u2__abc_44228_n19362;
  wire u2__abc_44228_n19363;
  wire u2__abc_44228_n19364;
  wire u2__abc_44228_n19365;
  wire u2__abc_44228_n19366;
  wire u2__abc_44228_n19367;
  wire u2__abc_44228_n19368;
  wire u2__abc_44228_n19369;
  wire u2__abc_44228_n19371;
  wire u2__abc_44228_n19372;
  wire u2__abc_44228_n19373;
  wire u2__abc_44228_n19374;
  wire u2__abc_44228_n19375;
  wire u2__abc_44228_n19376;
  wire u2__abc_44228_n19377;
  wire u2__abc_44228_n19378;
  wire u2__abc_44228_n19379;
  wire u2__abc_44228_n19380;
  wire u2__abc_44228_n19381;
  wire u2__abc_44228_n19383;
  wire u2__abc_44228_n19384;
  wire u2__abc_44228_n19385;
  wire u2__abc_44228_n19386;
  wire u2__abc_44228_n19387;
  wire u2__abc_44228_n19388;
  wire u2__abc_44228_n19389;
  wire u2__abc_44228_n19390;
  wire u2__abc_44228_n19391;
  wire u2__abc_44228_n19392;
  wire u2__abc_44228_n19393;
  wire u2__abc_44228_n19395;
  wire u2__abc_44228_n19396;
  wire u2__abc_44228_n19397;
  wire u2__abc_44228_n19398;
  wire u2__abc_44228_n19399;
  wire u2__abc_44228_n19400;
  wire u2__abc_44228_n19401;
  wire u2__abc_44228_n19402;
  wire u2__abc_44228_n19403;
  wire u2__abc_44228_n19404;
  wire u2__abc_44228_n19405;
  wire u2__abc_44228_n19407;
  wire u2__abc_44228_n19408;
  wire u2__abc_44228_n19409;
  wire u2__abc_44228_n19410;
  wire u2__abc_44228_n19411;
  wire u2__abc_44228_n19412;
  wire u2__abc_44228_n19413;
  wire u2__abc_44228_n19414;
  wire u2__abc_44228_n19415;
  wire u2__abc_44228_n19416;
  wire u2__abc_44228_n19417;
  wire u2__abc_44228_n19419;
  wire u2__abc_44228_n19420;
  wire u2__abc_44228_n19421;
  wire u2__abc_44228_n19422;
  wire u2__abc_44228_n19423;
  wire u2__abc_44228_n19424;
  wire u2__abc_44228_n19425;
  wire u2__abc_44228_n19426;
  wire u2__abc_44228_n19427;
  wire u2__abc_44228_n19428;
  wire u2__abc_44228_n19429;
  wire u2__abc_44228_n19431;
  wire u2__abc_44228_n19432;
  wire u2__abc_44228_n19433;
  wire u2__abc_44228_n19434;
  wire u2__abc_44228_n19435;
  wire u2__abc_44228_n19436;
  wire u2__abc_44228_n19437;
  wire u2__abc_44228_n19438;
  wire u2__abc_44228_n19439;
  wire u2__abc_44228_n19440;
  wire u2__abc_44228_n19441;
  wire u2__abc_44228_n19443;
  wire u2__abc_44228_n19444;
  wire u2__abc_44228_n19445;
  wire u2__abc_44228_n19446;
  wire u2__abc_44228_n19447;
  wire u2__abc_44228_n19448;
  wire u2__abc_44228_n19449;
  wire u2__abc_44228_n19450;
  wire u2__abc_44228_n19451;
  wire u2__abc_44228_n19452;
  wire u2__abc_44228_n19453;
  wire u2__abc_44228_n19455;
  wire u2__abc_44228_n19456;
  wire u2__abc_44228_n19457;
  wire u2__abc_44228_n19458;
  wire u2__abc_44228_n19459;
  wire u2__abc_44228_n19460;
  wire u2__abc_44228_n19461;
  wire u2__abc_44228_n19462;
  wire u2__abc_44228_n19463;
  wire u2__abc_44228_n19464;
  wire u2__abc_44228_n19465;
  wire u2__abc_44228_n19467;
  wire u2__abc_44228_n19468;
  wire u2__abc_44228_n19469;
  wire u2__abc_44228_n19470;
  wire u2__abc_44228_n19471;
  wire u2__abc_44228_n19472;
  wire u2__abc_44228_n19473;
  wire u2__abc_44228_n19474;
  wire u2__abc_44228_n19475;
  wire u2__abc_44228_n19476;
  wire u2__abc_44228_n19477;
  wire u2__abc_44228_n19479;
  wire u2__abc_44228_n19480;
  wire u2__abc_44228_n19481;
  wire u2__abc_44228_n19482;
  wire u2__abc_44228_n19483;
  wire u2__abc_44228_n19484;
  wire u2__abc_44228_n19485;
  wire u2__abc_44228_n19486;
  wire u2__abc_44228_n19487;
  wire u2__abc_44228_n19488;
  wire u2__abc_44228_n19489;
  wire u2__abc_44228_n19491;
  wire u2__abc_44228_n19492;
  wire u2__abc_44228_n19493;
  wire u2__abc_44228_n19494;
  wire u2__abc_44228_n19495;
  wire u2__abc_44228_n19496;
  wire u2__abc_44228_n19497;
  wire u2__abc_44228_n19498;
  wire u2__abc_44228_n19499;
  wire u2__abc_44228_n19500;
  wire u2__abc_44228_n19501;
  wire u2__abc_44228_n19503;
  wire u2__abc_44228_n19504;
  wire u2__abc_44228_n19505;
  wire u2__abc_44228_n19506;
  wire u2__abc_44228_n19507;
  wire u2__abc_44228_n19508;
  wire u2__abc_44228_n19509;
  wire u2__abc_44228_n19510;
  wire u2__abc_44228_n19511;
  wire u2__abc_44228_n19512;
  wire u2__abc_44228_n19513;
  wire u2__abc_44228_n19515;
  wire u2__abc_44228_n19516;
  wire u2__abc_44228_n19517;
  wire u2__abc_44228_n19518;
  wire u2__abc_44228_n19519;
  wire u2__abc_44228_n19520;
  wire u2__abc_44228_n19521;
  wire u2__abc_44228_n19522;
  wire u2__abc_44228_n19523;
  wire u2__abc_44228_n19524;
  wire u2__abc_44228_n19525;
  wire u2__abc_44228_n19527;
  wire u2__abc_44228_n19528;
  wire u2__abc_44228_n19529;
  wire u2__abc_44228_n19530;
  wire u2__abc_44228_n19531;
  wire u2__abc_44228_n19532;
  wire u2__abc_44228_n19533;
  wire u2__abc_44228_n19534;
  wire u2__abc_44228_n19535;
  wire u2__abc_44228_n19536;
  wire u2__abc_44228_n19537;
  wire u2__abc_44228_n19539;
  wire u2__abc_44228_n19540;
  wire u2__abc_44228_n19541;
  wire u2__abc_44228_n19542;
  wire u2__abc_44228_n19543;
  wire u2__abc_44228_n19544;
  wire u2__abc_44228_n19545;
  wire u2__abc_44228_n19546;
  wire u2__abc_44228_n19547;
  wire u2__abc_44228_n19548;
  wire u2__abc_44228_n19549;
  wire u2__abc_44228_n19551;
  wire u2__abc_44228_n19552;
  wire u2__abc_44228_n19553;
  wire u2__abc_44228_n19554;
  wire u2__abc_44228_n19555;
  wire u2__abc_44228_n19556;
  wire u2__abc_44228_n19557;
  wire u2__abc_44228_n19558;
  wire u2__abc_44228_n19559;
  wire u2__abc_44228_n19560;
  wire u2__abc_44228_n19561;
  wire u2__abc_44228_n19563;
  wire u2__abc_44228_n19564;
  wire u2__abc_44228_n19565;
  wire u2__abc_44228_n19566;
  wire u2__abc_44228_n19567;
  wire u2__abc_44228_n19568;
  wire u2__abc_44228_n19569;
  wire u2__abc_44228_n19570;
  wire u2__abc_44228_n19571;
  wire u2__abc_44228_n19572;
  wire u2__abc_44228_n19573;
  wire u2__abc_44228_n19575;
  wire u2__abc_44228_n19576;
  wire u2__abc_44228_n19577;
  wire u2__abc_44228_n19578;
  wire u2__abc_44228_n19579;
  wire u2__abc_44228_n19580;
  wire u2__abc_44228_n19581;
  wire u2__abc_44228_n19582;
  wire u2__abc_44228_n19583;
  wire u2__abc_44228_n19584;
  wire u2__abc_44228_n19585;
  wire u2__abc_44228_n19587;
  wire u2__abc_44228_n19588;
  wire u2__abc_44228_n19589;
  wire u2__abc_44228_n19590;
  wire u2__abc_44228_n19591;
  wire u2__abc_44228_n19592;
  wire u2__abc_44228_n19593;
  wire u2__abc_44228_n19594;
  wire u2__abc_44228_n19595;
  wire u2__abc_44228_n19596;
  wire u2__abc_44228_n19597;
  wire u2__abc_44228_n19599;
  wire u2__abc_44228_n19600;
  wire u2__abc_44228_n19601;
  wire u2__abc_44228_n19602;
  wire u2__abc_44228_n19603;
  wire u2__abc_44228_n19604;
  wire u2__abc_44228_n19605;
  wire u2__abc_44228_n19606;
  wire u2__abc_44228_n19607;
  wire u2__abc_44228_n19608;
  wire u2__abc_44228_n19609;
  wire u2__abc_44228_n19611;
  wire u2__abc_44228_n19612;
  wire u2__abc_44228_n19613;
  wire u2__abc_44228_n19614;
  wire u2__abc_44228_n19615;
  wire u2__abc_44228_n19616;
  wire u2__abc_44228_n19617;
  wire u2__abc_44228_n19618;
  wire u2__abc_44228_n19619;
  wire u2__abc_44228_n19620;
  wire u2__abc_44228_n19621;
  wire u2__abc_44228_n19623;
  wire u2__abc_44228_n19624;
  wire u2__abc_44228_n19625;
  wire u2__abc_44228_n19626;
  wire u2__abc_44228_n19627;
  wire u2__abc_44228_n19628;
  wire u2__abc_44228_n19629;
  wire u2__abc_44228_n19630;
  wire u2__abc_44228_n19631;
  wire u2__abc_44228_n19632;
  wire u2__abc_44228_n19633;
  wire u2__abc_44228_n19635;
  wire u2__abc_44228_n19636;
  wire u2__abc_44228_n19637;
  wire u2__abc_44228_n19638;
  wire u2__abc_44228_n19639;
  wire u2__abc_44228_n19640;
  wire u2__abc_44228_n19641;
  wire u2__abc_44228_n19642;
  wire u2__abc_44228_n19643;
  wire u2__abc_44228_n19644;
  wire u2__abc_44228_n19645;
  wire u2__abc_44228_n19647;
  wire u2__abc_44228_n19648;
  wire u2__abc_44228_n19649;
  wire u2__abc_44228_n19650;
  wire u2__abc_44228_n19651;
  wire u2__abc_44228_n19652;
  wire u2__abc_44228_n19653;
  wire u2__abc_44228_n19654;
  wire u2__abc_44228_n19655;
  wire u2__abc_44228_n19656;
  wire u2__abc_44228_n19657;
  wire u2__abc_44228_n19659;
  wire u2__abc_44228_n19660;
  wire u2__abc_44228_n19661;
  wire u2__abc_44228_n19662;
  wire u2__abc_44228_n19663;
  wire u2__abc_44228_n19664;
  wire u2__abc_44228_n19665;
  wire u2__abc_44228_n19666;
  wire u2__abc_44228_n19667;
  wire u2__abc_44228_n19668;
  wire u2__abc_44228_n19669;
  wire u2__abc_44228_n19671;
  wire u2__abc_44228_n19672;
  wire u2__abc_44228_n19673;
  wire u2__abc_44228_n19674;
  wire u2__abc_44228_n19675;
  wire u2__abc_44228_n19676;
  wire u2__abc_44228_n19677;
  wire u2__abc_44228_n19678;
  wire u2__abc_44228_n19679;
  wire u2__abc_44228_n19680;
  wire u2__abc_44228_n19681;
  wire u2__abc_44228_n19683;
  wire u2__abc_44228_n19684;
  wire u2__abc_44228_n19685;
  wire u2__abc_44228_n19686;
  wire u2__abc_44228_n19687;
  wire u2__abc_44228_n19688;
  wire u2__abc_44228_n19689;
  wire u2__abc_44228_n19690;
  wire u2__abc_44228_n19691;
  wire u2__abc_44228_n19692;
  wire u2__abc_44228_n19693;
  wire u2__abc_44228_n19695;
  wire u2__abc_44228_n19696;
  wire u2__abc_44228_n19697;
  wire u2__abc_44228_n19698;
  wire u2__abc_44228_n19699;
  wire u2__abc_44228_n19700;
  wire u2__abc_44228_n19701;
  wire u2__abc_44228_n19702;
  wire u2__abc_44228_n19703;
  wire u2__abc_44228_n19704;
  wire u2__abc_44228_n19705;
  wire u2__abc_44228_n19707;
  wire u2__abc_44228_n19708;
  wire u2__abc_44228_n19709;
  wire u2__abc_44228_n19710;
  wire u2__abc_44228_n19711;
  wire u2__abc_44228_n19712;
  wire u2__abc_44228_n19713;
  wire u2__abc_44228_n19714;
  wire u2__abc_44228_n19715;
  wire u2__abc_44228_n19716;
  wire u2__abc_44228_n19717;
  wire u2__abc_44228_n19719;
  wire u2__abc_44228_n19720;
  wire u2__abc_44228_n19721;
  wire u2__abc_44228_n19722;
  wire u2__abc_44228_n19723;
  wire u2__abc_44228_n19724;
  wire u2__abc_44228_n19725;
  wire u2__abc_44228_n19726;
  wire u2__abc_44228_n19727;
  wire u2__abc_44228_n19728;
  wire u2__abc_44228_n19729;
  wire u2__abc_44228_n19731;
  wire u2__abc_44228_n19732;
  wire u2__abc_44228_n19733;
  wire u2__abc_44228_n19734;
  wire u2__abc_44228_n19735;
  wire u2__abc_44228_n19736;
  wire u2__abc_44228_n19737;
  wire u2__abc_44228_n19738;
  wire u2__abc_44228_n19739;
  wire u2__abc_44228_n19740;
  wire u2__abc_44228_n19741;
  wire u2__abc_44228_n19743;
  wire u2__abc_44228_n19744;
  wire u2__abc_44228_n19745;
  wire u2__abc_44228_n19746;
  wire u2__abc_44228_n19747;
  wire u2__abc_44228_n19748;
  wire u2__abc_44228_n19749;
  wire u2__abc_44228_n19750;
  wire u2__abc_44228_n19751;
  wire u2__abc_44228_n19752;
  wire u2__abc_44228_n19753;
  wire u2__abc_44228_n19755;
  wire u2__abc_44228_n19756;
  wire u2__abc_44228_n19757;
  wire u2__abc_44228_n19758;
  wire u2__abc_44228_n19759;
  wire u2__abc_44228_n19760;
  wire u2__abc_44228_n19761;
  wire u2__abc_44228_n19762;
  wire u2__abc_44228_n19763;
  wire u2__abc_44228_n19764;
  wire u2__abc_44228_n19765;
  wire u2__abc_44228_n19767;
  wire u2__abc_44228_n19768;
  wire u2__abc_44228_n19769;
  wire u2__abc_44228_n19770;
  wire u2__abc_44228_n19771;
  wire u2__abc_44228_n19772;
  wire u2__abc_44228_n19773;
  wire u2__abc_44228_n19774;
  wire u2__abc_44228_n19775;
  wire u2__abc_44228_n19776;
  wire u2__abc_44228_n19777;
  wire u2__abc_44228_n19779;
  wire u2__abc_44228_n19780;
  wire u2__abc_44228_n19781;
  wire u2__abc_44228_n19782;
  wire u2__abc_44228_n19783;
  wire u2__abc_44228_n19784;
  wire u2__abc_44228_n19785;
  wire u2__abc_44228_n19786;
  wire u2__abc_44228_n19787;
  wire u2__abc_44228_n19788;
  wire u2__abc_44228_n19789;
  wire u2__abc_44228_n19791;
  wire u2__abc_44228_n19792;
  wire u2__abc_44228_n19793;
  wire u2__abc_44228_n19794;
  wire u2__abc_44228_n19795;
  wire u2__abc_44228_n19796;
  wire u2__abc_44228_n19797;
  wire u2__abc_44228_n19798;
  wire u2__abc_44228_n19799;
  wire u2__abc_44228_n19800;
  wire u2__abc_44228_n19801;
  wire u2__abc_44228_n19803;
  wire u2__abc_44228_n19804;
  wire u2__abc_44228_n19805;
  wire u2__abc_44228_n19806;
  wire u2__abc_44228_n19807;
  wire u2__abc_44228_n19808;
  wire u2__abc_44228_n19809;
  wire u2__abc_44228_n19810;
  wire u2__abc_44228_n19811;
  wire u2__abc_44228_n19812;
  wire u2__abc_44228_n19813;
  wire u2__abc_44228_n19815;
  wire u2__abc_44228_n19816;
  wire u2__abc_44228_n19817;
  wire u2__abc_44228_n19818;
  wire u2__abc_44228_n19819;
  wire u2__abc_44228_n19820;
  wire u2__abc_44228_n19821;
  wire u2__abc_44228_n19822;
  wire u2__abc_44228_n19823;
  wire u2__abc_44228_n19824;
  wire u2__abc_44228_n19825;
  wire u2__abc_44228_n19827;
  wire u2__abc_44228_n19828;
  wire u2__abc_44228_n19829;
  wire u2__abc_44228_n19830;
  wire u2__abc_44228_n19831;
  wire u2__abc_44228_n19832;
  wire u2__abc_44228_n19833;
  wire u2__abc_44228_n19834;
  wire u2__abc_44228_n19835;
  wire u2__abc_44228_n19836;
  wire u2__abc_44228_n19837;
  wire u2__abc_44228_n19839;
  wire u2__abc_44228_n19840;
  wire u2__abc_44228_n19841;
  wire u2__abc_44228_n19842;
  wire u2__abc_44228_n19843;
  wire u2__abc_44228_n19844;
  wire u2__abc_44228_n19845;
  wire u2__abc_44228_n19846;
  wire u2__abc_44228_n19847;
  wire u2__abc_44228_n19848;
  wire u2__abc_44228_n19849;
  wire u2__abc_44228_n19851;
  wire u2__abc_44228_n19852;
  wire u2__abc_44228_n19853;
  wire u2__abc_44228_n19854;
  wire u2__abc_44228_n19855;
  wire u2__abc_44228_n19856;
  wire u2__abc_44228_n19857;
  wire u2__abc_44228_n19858;
  wire u2__abc_44228_n19859;
  wire u2__abc_44228_n19860;
  wire u2__abc_44228_n19861;
  wire u2__abc_44228_n19863;
  wire u2__abc_44228_n19864;
  wire u2__abc_44228_n19865;
  wire u2__abc_44228_n19866;
  wire u2__abc_44228_n19867;
  wire u2__abc_44228_n19868;
  wire u2__abc_44228_n19869;
  wire u2__abc_44228_n19870;
  wire u2__abc_44228_n19871;
  wire u2__abc_44228_n19872;
  wire u2__abc_44228_n19873;
  wire u2__abc_44228_n19875;
  wire u2__abc_44228_n19876;
  wire u2__abc_44228_n19877;
  wire u2__abc_44228_n19878;
  wire u2__abc_44228_n19879;
  wire u2__abc_44228_n19880;
  wire u2__abc_44228_n19881;
  wire u2__abc_44228_n19882;
  wire u2__abc_44228_n19883;
  wire u2__abc_44228_n19884;
  wire u2__abc_44228_n19885;
  wire u2__abc_44228_n19887;
  wire u2__abc_44228_n19888;
  wire u2__abc_44228_n19889;
  wire u2__abc_44228_n19890;
  wire u2__abc_44228_n19891;
  wire u2__abc_44228_n19892;
  wire u2__abc_44228_n19893;
  wire u2__abc_44228_n19894;
  wire u2__abc_44228_n19895;
  wire u2__abc_44228_n19896;
  wire u2__abc_44228_n19897;
  wire u2__abc_44228_n19899;
  wire u2__abc_44228_n19900;
  wire u2__abc_44228_n19901;
  wire u2__abc_44228_n19902;
  wire u2__abc_44228_n19903;
  wire u2__abc_44228_n19904;
  wire u2__abc_44228_n19905;
  wire u2__abc_44228_n19906;
  wire u2__abc_44228_n19907;
  wire u2__abc_44228_n19908;
  wire u2__abc_44228_n19909;
  wire u2__abc_44228_n19911;
  wire u2__abc_44228_n19912;
  wire u2__abc_44228_n19913;
  wire u2__abc_44228_n19914;
  wire u2__abc_44228_n19915;
  wire u2__abc_44228_n19916;
  wire u2__abc_44228_n19917;
  wire u2__abc_44228_n19918;
  wire u2__abc_44228_n19919;
  wire u2__abc_44228_n19920;
  wire u2__abc_44228_n19921;
  wire u2__abc_44228_n19923;
  wire u2__abc_44228_n19924;
  wire u2__abc_44228_n19925;
  wire u2__abc_44228_n19926;
  wire u2__abc_44228_n19927;
  wire u2__abc_44228_n19928;
  wire u2__abc_44228_n19929;
  wire u2__abc_44228_n19930;
  wire u2__abc_44228_n19931;
  wire u2__abc_44228_n19932;
  wire u2__abc_44228_n19933;
  wire u2__abc_44228_n19935;
  wire u2__abc_44228_n19936;
  wire u2__abc_44228_n19937;
  wire u2__abc_44228_n19938;
  wire u2__abc_44228_n19939;
  wire u2__abc_44228_n19940;
  wire u2__abc_44228_n19941;
  wire u2__abc_44228_n19942;
  wire u2__abc_44228_n19943;
  wire u2__abc_44228_n19944;
  wire u2__abc_44228_n19945;
  wire u2__abc_44228_n19947;
  wire u2__abc_44228_n19948;
  wire u2__abc_44228_n19949;
  wire u2__abc_44228_n19950;
  wire u2__abc_44228_n19951;
  wire u2__abc_44228_n19952;
  wire u2__abc_44228_n19953;
  wire u2__abc_44228_n19954;
  wire u2__abc_44228_n19955;
  wire u2__abc_44228_n19956;
  wire u2__abc_44228_n19957;
  wire u2__abc_44228_n19959;
  wire u2__abc_44228_n19960;
  wire u2__abc_44228_n19961;
  wire u2__abc_44228_n19962;
  wire u2__abc_44228_n19963;
  wire u2__abc_44228_n19964;
  wire u2__abc_44228_n19965;
  wire u2__abc_44228_n19966;
  wire u2__abc_44228_n19967;
  wire u2__abc_44228_n19968;
  wire u2__abc_44228_n19969;
  wire u2__abc_44228_n19971;
  wire u2__abc_44228_n19972;
  wire u2__abc_44228_n19973;
  wire u2__abc_44228_n19974;
  wire u2__abc_44228_n19975;
  wire u2__abc_44228_n19976;
  wire u2__abc_44228_n19977;
  wire u2__abc_44228_n19978;
  wire u2__abc_44228_n19979;
  wire u2__abc_44228_n19980;
  wire u2__abc_44228_n19981;
  wire u2__abc_44228_n19983;
  wire u2__abc_44228_n19984;
  wire u2__abc_44228_n19985;
  wire u2__abc_44228_n19986;
  wire u2__abc_44228_n19987;
  wire u2__abc_44228_n19988;
  wire u2__abc_44228_n19989;
  wire u2__abc_44228_n19990;
  wire u2__abc_44228_n19991;
  wire u2__abc_44228_n19992;
  wire u2__abc_44228_n19993;
  wire u2__abc_44228_n19995;
  wire u2__abc_44228_n19996;
  wire u2__abc_44228_n19997;
  wire u2__abc_44228_n19998;
  wire u2__abc_44228_n19999;
  wire u2__abc_44228_n20000;
  wire u2__abc_44228_n20001;
  wire u2__abc_44228_n20002;
  wire u2__abc_44228_n20003;
  wire u2__abc_44228_n20004;
  wire u2__abc_44228_n20005;
  wire u2__abc_44228_n20007;
  wire u2__abc_44228_n20008;
  wire u2__abc_44228_n20009;
  wire u2__abc_44228_n20010;
  wire u2__abc_44228_n20011;
  wire u2__abc_44228_n20012;
  wire u2__abc_44228_n20013;
  wire u2__abc_44228_n20014;
  wire u2__abc_44228_n20015;
  wire u2__abc_44228_n20016;
  wire u2__abc_44228_n20017;
  wire u2__abc_44228_n20019;
  wire u2__abc_44228_n20020;
  wire u2__abc_44228_n20021;
  wire u2__abc_44228_n20022;
  wire u2__abc_44228_n20023;
  wire u2__abc_44228_n20024;
  wire u2__abc_44228_n20025;
  wire u2__abc_44228_n20026;
  wire u2__abc_44228_n20027;
  wire u2__abc_44228_n20028;
  wire u2__abc_44228_n20029;
  wire u2__abc_44228_n20031;
  wire u2__abc_44228_n20032;
  wire u2__abc_44228_n20033;
  wire u2__abc_44228_n20034;
  wire u2__abc_44228_n20035;
  wire u2__abc_44228_n20036;
  wire u2__abc_44228_n20037;
  wire u2__abc_44228_n20038;
  wire u2__abc_44228_n20039;
  wire u2__abc_44228_n20040;
  wire u2__abc_44228_n20041;
  wire u2__abc_44228_n20043;
  wire u2__abc_44228_n20044;
  wire u2__abc_44228_n20045;
  wire u2__abc_44228_n20046;
  wire u2__abc_44228_n20047;
  wire u2__abc_44228_n20048;
  wire u2__abc_44228_n20049;
  wire u2__abc_44228_n20050;
  wire u2__abc_44228_n20051;
  wire u2__abc_44228_n20052;
  wire u2__abc_44228_n20053;
  wire u2__abc_44228_n20055;
  wire u2__abc_44228_n20056;
  wire u2__abc_44228_n20057;
  wire u2__abc_44228_n20058;
  wire u2__abc_44228_n20059;
  wire u2__abc_44228_n20060;
  wire u2__abc_44228_n20061;
  wire u2__abc_44228_n20062;
  wire u2__abc_44228_n20063;
  wire u2__abc_44228_n20064;
  wire u2__abc_44228_n20065;
  wire u2__abc_44228_n20067;
  wire u2__abc_44228_n20068;
  wire u2__abc_44228_n20069;
  wire u2__abc_44228_n20070;
  wire u2__abc_44228_n20071;
  wire u2__abc_44228_n20072;
  wire u2__abc_44228_n20073;
  wire u2__abc_44228_n20074;
  wire u2__abc_44228_n20075;
  wire u2__abc_44228_n20076;
  wire u2__abc_44228_n20077;
  wire u2__abc_44228_n20079;
  wire u2__abc_44228_n20080;
  wire u2__abc_44228_n20081;
  wire u2__abc_44228_n20082;
  wire u2__abc_44228_n20083;
  wire u2__abc_44228_n20084;
  wire u2__abc_44228_n20085;
  wire u2__abc_44228_n20086;
  wire u2__abc_44228_n20087;
  wire u2__abc_44228_n20088;
  wire u2__abc_44228_n20089;
  wire u2__abc_44228_n20091;
  wire u2__abc_44228_n20092;
  wire u2__abc_44228_n20093;
  wire u2__abc_44228_n20094;
  wire u2__abc_44228_n20095;
  wire u2__abc_44228_n20096;
  wire u2__abc_44228_n20097;
  wire u2__abc_44228_n20098;
  wire u2__abc_44228_n20099;
  wire u2__abc_44228_n20100;
  wire u2__abc_44228_n20101;
  wire u2__abc_44228_n20103;
  wire u2__abc_44228_n20104;
  wire u2__abc_44228_n20105;
  wire u2__abc_44228_n20106;
  wire u2__abc_44228_n20107;
  wire u2__abc_44228_n20108;
  wire u2__abc_44228_n20109;
  wire u2__abc_44228_n20110;
  wire u2__abc_44228_n20111;
  wire u2__abc_44228_n20112;
  wire u2__abc_44228_n20113;
  wire u2__abc_44228_n20115;
  wire u2__abc_44228_n20116;
  wire u2__abc_44228_n20117;
  wire u2__abc_44228_n20118;
  wire u2__abc_44228_n20119;
  wire u2__abc_44228_n20120;
  wire u2__abc_44228_n20121;
  wire u2__abc_44228_n20122;
  wire u2__abc_44228_n20123;
  wire u2__abc_44228_n20124;
  wire u2__abc_44228_n20125;
  wire u2__abc_44228_n20127;
  wire u2__abc_44228_n20128;
  wire u2__abc_44228_n20129;
  wire u2__abc_44228_n20130;
  wire u2__abc_44228_n20131;
  wire u2__abc_44228_n20132;
  wire u2__abc_44228_n20133;
  wire u2__abc_44228_n20134;
  wire u2__abc_44228_n20135;
  wire u2__abc_44228_n20136;
  wire u2__abc_44228_n20137;
  wire u2__abc_44228_n20139;
  wire u2__abc_44228_n20140;
  wire u2__abc_44228_n20141;
  wire u2__abc_44228_n20142;
  wire u2__abc_44228_n20143;
  wire u2__abc_44228_n20144;
  wire u2__abc_44228_n20145;
  wire u2__abc_44228_n20146;
  wire u2__abc_44228_n20147;
  wire u2__abc_44228_n20148;
  wire u2__abc_44228_n20149;
  wire u2__abc_44228_n20151;
  wire u2__abc_44228_n20152;
  wire u2__abc_44228_n20153;
  wire u2__abc_44228_n20154;
  wire u2__abc_44228_n20155;
  wire u2__abc_44228_n20156;
  wire u2__abc_44228_n20157;
  wire u2__abc_44228_n20158;
  wire u2__abc_44228_n20159;
  wire u2__abc_44228_n20160;
  wire u2__abc_44228_n20161;
  wire u2__abc_44228_n20163;
  wire u2__abc_44228_n20164;
  wire u2__abc_44228_n20165;
  wire u2__abc_44228_n20166;
  wire u2__abc_44228_n20167;
  wire u2__abc_44228_n20168;
  wire u2__abc_44228_n20169;
  wire u2__abc_44228_n20170;
  wire u2__abc_44228_n20171;
  wire u2__abc_44228_n20172;
  wire u2__abc_44228_n20173;
  wire u2__abc_44228_n20175;
  wire u2__abc_44228_n20176;
  wire u2__abc_44228_n20177;
  wire u2__abc_44228_n20178;
  wire u2__abc_44228_n20179;
  wire u2__abc_44228_n20180;
  wire u2__abc_44228_n20181;
  wire u2__abc_44228_n20182;
  wire u2__abc_44228_n20183;
  wire u2__abc_44228_n20184;
  wire u2__abc_44228_n20185;
  wire u2__abc_44228_n20187;
  wire u2__abc_44228_n20188;
  wire u2__abc_44228_n20189;
  wire u2__abc_44228_n20190;
  wire u2__abc_44228_n20191;
  wire u2__abc_44228_n20192;
  wire u2__abc_44228_n20193;
  wire u2__abc_44228_n20194;
  wire u2__abc_44228_n20195;
  wire u2__abc_44228_n20196;
  wire u2__abc_44228_n20197;
  wire u2__abc_44228_n20199;
  wire u2__abc_44228_n20200;
  wire u2__abc_44228_n20201;
  wire u2__abc_44228_n20202;
  wire u2__abc_44228_n20203;
  wire u2__abc_44228_n20204;
  wire u2__abc_44228_n20205;
  wire u2__abc_44228_n20206;
  wire u2__abc_44228_n20207;
  wire u2__abc_44228_n20208;
  wire u2__abc_44228_n20209;
  wire u2__abc_44228_n20211;
  wire u2__abc_44228_n20212;
  wire u2__abc_44228_n20213;
  wire u2__abc_44228_n20214;
  wire u2__abc_44228_n20215;
  wire u2__abc_44228_n20216;
  wire u2__abc_44228_n20217;
  wire u2__abc_44228_n20218;
  wire u2__abc_44228_n20219;
  wire u2__abc_44228_n20220;
  wire u2__abc_44228_n20221;
  wire u2__abc_44228_n20223;
  wire u2__abc_44228_n20224;
  wire u2__abc_44228_n20225;
  wire u2__abc_44228_n20226;
  wire u2__abc_44228_n20227;
  wire u2__abc_44228_n20228;
  wire u2__abc_44228_n20229;
  wire u2__abc_44228_n20230;
  wire u2__abc_44228_n20231;
  wire u2__abc_44228_n20232;
  wire u2__abc_44228_n20233;
  wire u2__abc_44228_n20235;
  wire u2__abc_44228_n20236;
  wire u2__abc_44228_n20237;
  wire u2__abc_44228_n20238;
  wire u2__abc_44228_n20239;
  wire u2__abc_44228_n20240;
  wire u2__abc_44228_n20241;
  wire u2__abc_44228_n20242;
  wire u2__abc_44228_n20243;
  wire u2__abc_44228_n20244;
  wire u2__abc_44228_n20245;
  wire u2__abc_44228_n20247;
  wire u2__abc_44228_n20248;
  wire u2__abc_44228_n20249;
  wire u2__abc_44228_n20250;
  wire u2__abc_44228_n20251;
  wire u2__abc_44228_n20252;
  wire u2__abc_44228_n20253;
  wire u2__abc_44228_n20254;
  wire u2__abc_44228_n20255;
  wire u2__abc_44228_n20256;
  wire u2__abc_44228_n20257;
  wire u2__abc_44228_n20259;
  wire u2__abc_44228_n20260;
  wire u2__abc_44228_n20261;
  wire u2__abc_44228_n20262;
  wire u2__abc_44228_n20263;
  wire u2__abc_44228_n20264;
  wire u2__abc_44228_n20265;
  wire u2__abc_44228_n20266;
  wire u2__abc_44228_n20267;
  wire u2__abc_44228_n20268;
  wire u2__abc_44228_n20269;
  wire u2__abc_44228_n20271;
  wire u2__abc_44228_n20272;
  wire u2__abc_44228_n20273;
  wire u2__abc_44228_n20274;
  wire u2__abc_44228_n20275;
  wire u2__abc_44228_n20276;
  wire u2__abc_44228_n20277;
  wire u2__abc_44228_n20278;
  wire u2__abc_44228_n20279;
  wire u2__abc_44228_n20280;
  wire u2__abc_44228_n20281;
  wire u2__abc_44228_n20283;
  wire u2__abc_44228_n20284;
  wire u2__abc_44228_n20285;
  wire u2__abc_44228_n20286;
  wire u2__abc_44228_n20287;
  wire u2__abc_44228_n20288;
  wire u2__abc_44228_n20289;
  wire u2__abc_44228_n20290;
  wire u2__abc_44228_n20291;
  wire u2__abc_44228_n20292;
  wire u2__abc_44228_n20293;
  wire u2__abc_44228_n20295;
  wire u2__abc_44228_n20296;
  wire u2__abc_44228_n20297;
  wire u2__abc_44228_n20298;
  wire u2__abc_44228_n20299;
  wire u2__abc_44228_n20300;
  wire u2__abc_44228_n20301;
  wire u2__abc_44228_n20302;
  wire u2__abc_44228_n20303;
  wire u2__abc_44228_n20304;
  wire u2__abc_44228_n20305;
  wire u2__abc_44228_n20307;
  wire u2__abc_44228_n20308;
  wire u2__abc_44228_n20309;
  wire u2__abc_44228_n20310;
  wire u2__abc_44228_n20311;
  wire u2__abc_44228_n20312;
  wire u2__abc_44228_n20313;
  wire u2__abc_44228_n20314;
  wire u2__abc_44228_n20315;
  wire u2__abc_44228_n20316;
  wire u2__abc_44228_n20317;
  wire u2__abc_44228_n20319;
  wire u2__abc_44228_n20320;
  wire u2__abc_44228_n20321;
  wire u2__abc_44228_n20322;
  wire u2__abc_44228_n20323;
  wire u2__abc_44228_n20324;
  wire u2__abc_44228_n20325;
  wire u2__abc_44228_n20326;
  wire u2__abc_44228_n20327;
  wire u2__abc_44228_n20328;
  wire u2__abc_44228_n20329;
  wire u2__abc_44228_n20331;
  wire u2__abc_44228_n20332;
  wire u2__abc_44228_n20333;
  wire u2__abc_44228_n20334;
  wire u2__abc_44228_n20335;
  wire u2__abc_44228_n20336;
  wire u2__abc_44228_n20337;
  wire u2__abc_44228_n20338;
  wire u2__abc_44228_n20339;
  wire u2__abc_44228_n20340;
  wire u2__abc_44228_n20341;
  wire u2__abc_44228_n20343;
  wire u2__abc_44228_n20344;
  wire u2__abc_44228_n20345;
  wire u2__abc_44228_n20346;
  wire u2__abc_44228_n20347;
  wire u2__abc_44228_n20348;
  wire u2__abc_44228_n20349;
  wire u2__abc_44228_n20350;
  wire u2__abc_44228_n20351;
  wire u2__abc_44228_n20352;
  wire u2__abc_44228_n20353;
  wire u2__abc_44228_n20355;
  wire u2__abc_44228_n20356;
  wire u2__abc_44228_n20357;
  wire u2__abc_44228_n20358;
  wire u2__abc_44228_n20359;
  wire u2__abc_44228_n20360;
  wire u2__abc_44228_n20361;
  wire u2__abc_44228_n20362;
  wire u2__abc_44228_n20363;
  wire u2__abc_44228_n20364;
  wire u2__abc_44228_n20365;
  wire u2__abc_44228_n20367;
  wire u2__abc_44228_n20368;
  wire u2__abc_44228_n20369;
  wire u2__abc_44228_n20370;
  wire u2__abc_44228_n20371;
  wire u2__abc_44228_n20372;
  wire u2__abc_44228_n20373;
  wire u2__abc_44228_n20374;
  wire u2__abc_44228_n20375;
  wire u2__abc_44228_n20376;
  wire u2__abc_44228_n20377;
  wire u2__abc_44228_n20379;
  wire u2__abc_44228_n20380;
  wire u2__abc_44228_n20381;
  wire u2__abc_44228_n20382;
  wire u2__abc_44228_n20383;
  wire u2__abc_44228_n20384;
  wire u2__abc_44228_n20385;
  wire u2__abc_44228_n20386;
  wire u2__abc_44228_n20387;
  wire u2__abc_44228_n20388;
  wire u2__abc_44228_n20389;
  wire u2__abc_44228_n20391;
  wire u2__abc_44228_n20392;
  wire u2__abc_44228_n20393;
  wire u2__abc_44228_n20394;
  wire u2__abc_44228_n20395;
  wire u2__abc_44228_n20396;
  wire u2__abc_44228_n20397;
  wire u2__abc_44228_n20398;
  wire u2__abc_44228_n20399;
  wire u2__abc_44228_n20400;
  wire u2__abc_44228_n20401;
  wire u2__abc_44228_n20403;
  wire u2__abc_44228_n20404;
  wire u2__abc_44228_n20405;
  wire u2__abc_44228_n20406;
  wire u2__abc_44228_n20407;
  wire u2__abc_44228_n20408;
  wire u2__abc_44228_n20409;
  wire u2__abc_44228_n20410;
  wire u2__abc_44228_n20411;
  wire u2__abc_44228_n20412;
  wire u2__abc_44228_n20413;
  wire u2__abc_44228_n20415;
  wire u2__abc_44228_n20416;
  wire u2__abc_44228_n20417;
  wire u2__abc_44228_n20418;
  wire u2__abc_44228_n20419;
  wire u2__abc_44228_n20420;
  wire u2__abc_44228_n20421;
  wire u2__abc_44228_n20422;
  wire u2__abc_44228_n20423;
  wire u2__abc_44228_n20424;
  wire u2__abc_44228_n20425;
  wire u2__abc_44228_n20427;
  wire u2__abc_44228_n20428;
  wire u2__abc_44228_n20429;
  wire u2__abc_44228_n20430;
  wire u2__abc_44228_n20431;
  wire u2__abc_44228_n20432;
  wire u2__abc_44228_n20433;
  wire u2__abc_44228_n20434;
  wire u2__abc_44228_n20435;
  wire u2__abc_44228_n20436;
  wire u2__abc_44228_n20437;
  wire u2__abc_44228_n20439;
  wire u2__abc_44228_n20440;
  wire u2__abc_44228_n20441;
  wire u2__abc_44228_n20442;
  wire u2__abc_44228_n20443;
  wire u2__abc_44228_n20444;
  wire u2__abc_44228_n20445;
  wire u2__abc_44228_n20446;
  wire u2__abc_44228_n20447;
  wire u2__abc_44228_n20448;
  wire u2__abc_44228_n20449;
  wire u2__abc_44228_n20451;
  wire u2__abc_44228_n20452;
  wire u2__abc_44228_n20453;
  wire u2__abc_44228_n20454;
  wire u2__abc_44228_n20455;
  wire u2__abc_44228_n20456;
  wire u2__abc_44228_n20457;
  wire u2__abc_44228_n20458;
  wire u2__abc_44228_n20459;
  wire u2__abc_44228_n20460;
  wire u2__abc_44228_n20461;
  wire u2__abc_44228_n20463;
  wire u2__abc_44228_n20464;
  wire u2__abc_44228_n20465;
  wire u2__abc_44228_n20466;
  wire u2__abc_44228_n20467;
  wire u2__abc_44228_n20468;
  wire u2__abc_44228_n20469;
  wire u2__abc_44228_n20470;
  wire u2__abc_44228_n20471;
  wire u2__abc_44228_n20472;
  wire u2__abc_44228_n20473;
  wire u2__abc_44228_n20475;
  wire u2__abc_44228_n20476;
  wire u2__abc_44228_n20477;
  wire u2__abc_44228_n20478;
  wire u2__abc_44228_n20479;
  wire u2__abc_44228_n20480;
  wire u2__abc_44228_n20481;
  wire u2__abc_44228_n20482;
  wire u2__abc_44228_n20483;
  wire u2__abc_44228_n20484;
  wire u2__abc_44228_n20485;
  wire u2__abc_44228_n20487;
  wire u2__abc_44228_n20488;
  wire u2__abc_44228_n20489;
  wire u2__abc_44228_n20490;
  wire u2__abc_44228_n20491;
  wire u2__abc_44228_n20492;
  wire u2__abc_44228_n20493;
  wire u2__abc_44228_n20494;
  wire u2__abc_44228_n20495;
  wire u2__abc_44228_n20496;
  wire u2__abc_44228_n20497;
  wire u2__abc_44228_n20499;
  wire u2__abc_44228_n20500;
  wire u2__abc_44228_n20501;
  wire u2__abc_44228_n20502;
  wire u2__abc_44228_n20503;
  wire u2__abc_44228_n20504;
  wire u2__abc_44228_n20505;
  wire u2__abc_44228_n20506;
  wire u2__abc_44228_n20507;
  wire u2__abc_44228_n20508;
  wire u2__abc_44228_n20509;
  wire u2__abc_44228_n20511;
  wire u2__abc_44228_n20512;
  wire u2__abc_44228_n20513;
  wire u2__abc_44228_n20514;
  wire u2__abc_44228_n20515;
  wire u2__abc_44228_n20516;
  wire u2__abc_44228_n20517;
  wire u2__abc_44228_n20518;
  wire u2__abc_44228_n20519;
  wire u2__abc_44228_n20520;
  wire u2__abc_44228_n20521;
  wire u2__abc_44228_n20523;
  wire u2__abc_44228_n20524;
  wire u2__abc_44228_n20525;
  wire u2__abc_44228_n20526;
  wire u2__abc_44228_n20527;
  wire u2__abc_44228_n20528;
  wire u2__abc_44228_n20529;
  wire u2__abc_44228_n20530;
  wire u2__abc_44228_n20531;
  wire u2__abc_44228_n20532;
  wire u2__abc_44228_n20533;
  wire u2__abc_44228_n20535;
  wire u2__abc_44228_n20536;
  wire u2__abc_44228_n20537;
  wire u2__abc_44228_n20538;
  wire u2__abc_44228_n20539;
  wire u2__abc_44228_n20540;
  wire u2__abc_44228_n20541;
  wire u2__abc_44228_n20542;
  wire u2__abc_44228_n20543;
  wire u2__abc_44228_n20544;
  wire u2__abc_44228_n20545;
  wire u2__abc_44228_n20547;
  wire u2__abc_44228_n20548;
  wire u2__abc_44228_n20549;
  wire u2__abc_44228_n20550;
  wire u2__abc_44228_n20551;
  wire u2__abc_44228_n20552;
  wire u2__abc_44228_n20553;
  wire u2__abc_44228_n20554;
  wire u2__abc_44228_n20555;
  wire u2__abc_44228_n20556;
  wire u2__abc_44228_n20557;
  wire u2__abc_44228_n20559;
  wire u2__abc_44228_n20560;
  wire u2__abc_44228_n20561;
  wire u2__abc_44228_n20562;
  wire u2__abc_44228_n20563;
  wire u2__abc_44228_n20564;
  wire u2__abc_44228_n20565;
  wire u2__abc_44228_n20566;
  wire u2__abc_44228_n20567;
  wire u2__abc_44228_n20568;
  wire u2__abc_44228_n20569;
  wire u2__abc_44228_n20571;
  wire u2__abc_44228_n20572;
  wire u2__abc_44228_n20573;
  wire u2__abc_44228_n20574;
  wire u2__abc_44228_n20575;
  wire u2__abc_44228_n20576;
  wire u2__abc_44228_n20577;
  wire u2__abc_44228_n20578;
  wire u2__abc_44228_n20579;
  wire u2__abc_44228_n20580;
  wire u2__abc_44228_n20581;
  wire u2__abc_44228_n20583;
  wire u2__abc_44228_n20584;
  wire u2__abc_44228_n20585;
  wire u2__abc_44228_n20586;
  wire u2__abc_44228_n20587;
  wire u2__abc_44228_n20588;
  wire u2__abc_44228_n20589;
  wire u2__abc_44228_n20590;
  wire u2__abc_44228_n20591;
  wire u2__abc_44228_n20592;
  wire u2__abc_44228_n20593;
  wire u2__abc_44228_n20595;
  wire u2__abc_44228_n20596;
  wire u2__abc_44228_n20597;
  wire u2__abc_44228_n20598;
  wire u2__abc_44228_n20599;
  wire u2__abc_44228_n20600;
  wire u2__abc_44228_n20601;
  wire u2__abc_44228_n20602;
  wire u2__abc_44228_n20603;
  wire u2__abc_44228_n20604;
  wire u2__abc_44228_n20605;
  wire u2__abc_44228_n20607;
  wire u2__abc_44228_n20608;
  wire u2__abc_44228_n20609;
  wire u2__abc_44228_n20610;
  wire u2__abc_44228_n20611;
  wire u2__abc_44228_n20612;
  wire u2__abc_44228_n20613;
  wire u2__abc_44228_n20614;
  wire u2__abc_44228_n20615;
  wire u2__abc_44228_n20616;
  wire u2__abc_44228_n20617;
  wire u2__abc_44228_n20619;
  wire u2__abc_44228_n20620;
  wire u2__abc_44228_n20621;
  wire u2__abc_44228_n20622;
  wire u2__abc_44228_n20623;
  wire u2__abc_44228_n20624;
  wire u2__abc_44228_n20625;
  wire u2__abc_44228_n20626;
  wire u2__abc_44228_n20627;
  wire u2__abc_44228_n20628;
  wire u2__abc_44228_n20629;
  wire u2__abc_44228_n20631;
  wire u2__abc_44228_n20632;
  wire u2__abc_44228_n20633;
  wire u2__abc_44228_n20634;
  wire u2__abc_44228_n20635;
  wire u2__abc_44228_n20636;
  wire u2__abc_44228_n20637;
  wire u2__abc_44228_n20638;
  wire u2__abc_44228_n20639;
  wire u2__abc_44228_n20640;
  wire u2__abc_44228_n20641;
  wire u2__abc_44228_n20643;
  wire u2__abc_44228_n20644;
  wire u2__abc_44228_n20645;
  wire u2__abc_44228_n20646;
  wire u2__abc_44228_n20647;
  wire u2__abc_44228_n20648;
  wire u2__abc_44228_n20649;
  wire u2__abc_44228_n20650;
  wire u2__abc_44228_n20651;
  wire u2__abc_44228_n20652;
  wire u2__abc_44228_n20653;
  wire u2__abc_44228_n20655;
  wire u2__abc_44228_n20656;
  wire u2__abc_44228_n20657;
  wire u2__abc_44228_n20658;
  wire u2__abc_44228_n20659;
  wire u2__abc_44228_n20660;
  wire u2__abc_44228_n20661;
  wire u2__abc_44228_n20662;
  wire u2__abc_44228_n20663;
  wire u2__abc_44228_n20664;
  wire u2__abc_44228_n20665;
  wire u2__abc_44228_n20667;
  wire u2__abc_44228_n20668;
  wire u2__abc_44228_n20669;
  wire u2__abc_44228_n20670;
  wire u2__abc_44228_n20671;
  wire u2__abc_44228_n20672;
  wire u2__abc_44228_n20673;
  wire u2__abc_44228_n20674;
  wire u2__abc_44228_n20675;
  wire u2__abc_44228_n20676;
  wire u2__abc_44228_n20677;
  wire u2__abc_44228_n20679;
  wire u2__abc_44228_n20680;
  wire u2__abc_44228_n20681;
  wire u2__abc_44228_n20682;
  wire u2__abc_44228_n20683;
  wire u2__abc_44228_n20684;
  wire u2__abc_44228_n20685;
  wire u2__abc_44228_n20686;
  wire u2__abc_44228_n20687;
  wire u2__abc_44228_n20688;
  wire u2__abc_44228_n20689;
  wire u2__abc_44228_n20691;
  wire u2__abc_44228_n20692;
  wire u2__abc_44228_n20693;
  wire u2__abc_44228_n20694;
  wire u2__abc_44228_n20695;
  wire u2__abc_44228_n20696;
  wire u2__abc_44228_n20697;
  wire u2__abc_44228_n20698;
  wire u2__abc_44228_n20699;
  wire u2__abc_44228_n20700;
  wire u2__abc_44228_n20701;
  wire u2__abc_44228_n20703;
  wire u2__abc_44228_n20704;
  wire u2__abc_44228_n20705;
  wire u2__abc_44228_n20706;
  wire u2__abc_44228_n20707;
  wire u2__abc_44228_n20708;
  wire u2__abc_44228_n20709;
  wire u2__abc_44228_n20710;
  wire u2__abc_44228_n20711;
  wire u2__abc_44228_n20712;
  wire u2__abc_44228_n20713;
  wire u2__abc_44228_n20715;
  wire u2__abc_44228_n20716;
  wire u2__abc_44228_n20717;
  wire u2__abc_44228_n20718;
  wire u2__abc_44228_n20719;
  wire u2__abc_44228_n20720;
  wire u2__abc_44228_n20721;
  wire u2__abc_44228_n20722;
  wire u2__abc_44228_n20723;
  wire u2__abc_44228_n20724;
  wire u2__abc_44228_n20725;
  wire u2__abc_44228_n20727;
  wire u2__abc_44228_n20728;
  wire u2__abc_44228_n20729;
  wire u2__abc_44228_n20730;
  wire u2__abc_44228_n20731;
  wire u2__abc_44228_n20732;
  wire u2__abc_44228_n20733;
  wire u2__abc_44228_n20734;
  wire u2__abc_44228_n20735;
  wire u2__abc_44228_n20736;
  wire u2__abc_44228_n20737;
  wire u2__abc_44228_n20739;
  wire u2__abc_44228_n20740;
  wire u2__abc_44228_n20741;
  wire u2__abc_44228_n20742;
  wire u2__abc_44228_n20743;
  wire u2__abc_44228_n20744;
  wire u2__abc_44228_n20745;
  wire u2__abc_44228_n20746;
  wire u2__abc_44228_n20747;
  wire u2__abc_44228_n20748;
  wire u2__abc_44228_n20749;
  wire u2__abc_44228_n20751;
  wire u2__abc_44228_n20752;
  wire u2__abc_44228_n20753;
  wire u2__abc_44228_n20754;
  wire u2__abc_44228_n20755;
  wire u2__abc_44228_n20756;
  wire u2__abc_44228_n20757;
  wire u2__abc_44228_n20758;
  wire u2__abc_44228_n20759;
  wire u2__abc_44228_n20760;
  wire u2__abc_44228_n20761;
  wire u2__abc_44228_n20763;
  wire u2__abc_44228_n20764;
  wire u2__abc_44228_n20765;
  wire u2__abc_44228_n20766;
  wire u2__abc_44228_n20767;
  wire u2__abc_44228_n20768;
  wire u2__abc_44228_n20769;
  wire u2__abc_44228_n20770;
  wire u2__abc_44228_n20771;
  wire u2__abc_44228_n20772;
  wire u2__abc_44228_n20773;
  wire u2__abc_44228_n20775;
  wire u2__abc_44228_n20776;
  wire u2__abc_44228_n20777;
  wire u2__abc_44228_n20778;
  wire u2__abc_44228_n20779;
  wire u2__abc_44228_n20780;
  wire u2__abc_44228_n20781;
  wire u2__abc_44228_n20782;
  wire u2__abc_44228_n20783;
  wire u2__abc_44228_n20784;
  wire u2__abc_44228_n20785;
  wire u2__abc_44228_n20787;
  wire u2__abc_44228_n20788;
  wire u2__abc_44228_n20789;
  wire u2__abc_44228_n20790;
  wire u2__abc_44228_n20791;
  wire u2__abc_44228_n20792;
  wire u2__abc_44228_n20793;
  wire u2__abc_44228_n20794;
  wire u2__abc_44228_n20795;
  wire u2__abc_44228_n20796;
  wire u2__abc_44228_n20797;
  wire u2__abc_44228_n20799;
  wire u2__abc_44228_n20800;
  wire u2__abc_44228_n20801;
  wire u2__abc_44228_n20802;
  wire u2__abc_44228_n20803;
  wire u2__abc_44228_n20804;
  wire u2__abc_44228_n20805;
  wire u2__abc_44228_n20806;
  wire u2__abc_44228_n20807;
  wire u2__abc_44228_n20808;
  wire u2__abc_44228_n20809;
  wire u2__abc_44228_n20811;
  wire u2__abc_44228_n20812;
  wire u2__abc_44228_n20813;
  wire u2__abc_44228_n20814;
  wire u2__abc_44228_n20815;
  wire u2__abc_44228_n20816;
  wire u2__abc_44228_n20817;
  wire u2__abc_44228_n20818;
  wire u2__abc_44228_n20819;
  wire u2__abc_44228_n20820;
  wire u2__abc_44228_n20821;
  wire u2__abc_44228_n20823;
  wire u2__abc_44228_n20824;
  wire u2__abc_44228_n20825;
  wire u2__abc_44228_n20826;
  wire u2__abc_44228_n20827;
  wire u2__abc_44228_n20828;
  wire u2__abc_44228_n20829;
  wire u2__abc_44228_n20830;
  wire u2__abc_44228_n20831;
  wire u2__abc_44228_n20832;
  wire u2__abc_44228_n20833;
  wire u2__abc_44228_n20835;
  wire u2__abc_44228_n20836;
  wire u2__abc_44228_n20837;
  wire u2__abc_44228_n20838;
  wire u2__abc_44228_n20839;
  wire u2__abc_44228_n20840;
  wire u2__abc_44228_n20841;
  wire u2__abc_44228_n20842;
  wire u2__abc_44228_n20843;
  wire u2__abc_44228_n20844;
  wire u2__abc_44228_n20845;
  wire u2__abc_44228_n20847;
  wire u2__abc_44228_n20848;
  wire u2__abc_44228_n20849;
  wire u2__abc_44228_n20850;
  wire u2__abc_44228_n20851;
  wire u2__abc_44228_n20852;
  wire u2__abc_44228_n20853;
  wire u2__abc_44228_n20854;
  wire u2__abc_44228_n20855;
  wire u2__abc_44228_n20856;
  wire u2__abc_44228_n20857;
  wire u2__abc_44228_n20859;
  wire u2__abc_44228_n20860;
  wire u2__abc_44228_n20861;
  wire u2__abc_44228_n20862;
  wire u2__abc_44228_n20863;
  wire u2__abc_44228_n20864;
  wire u2__abc_44228_n20865;
  wire u2__abc_44228_n20866;
  wire u2__abc_44228_n20867;
  wire u2__abc_44228_n20868;
  wire u2__abc_44228_n20869;
  wire u2__abc_44228_n20871;
  wire u2__abc_44228_n20872;
  wire u2__abc_44228_n20873;
  wire u2__abc_44228_n20874;
  wire u2__abc_44228_n20875;
  wire u2__abc_44228_n20876;
  wire u2__abc_44228_n20877;
  wire u2__abc_44228_n20878;
  wire u2__abc_44228_n20879;
  wire u2__abc_44228_n20880;
  wire u2__abc_44228_n20881;
  wire u2__abc_44228_n20883;
  wire u2__abc_44228_n20884;
  wire u2__abc_44228_n20885;
  wire u2__abc_44228_n20886;
  wire u2__abc_44228_n20887;
  wire u2__abc_44228_n20888;
  wire u2__abc_44228_n20889;
  wire u2__abc_44228_n20890;
  wire u2__abc_44228_n20891;
  wire u2__abc_44228_n20892;
  wire u2__abc_44228_n20893;
  wire u2__abc_44228_n20895;
  wire u2__abc_44228_n20896;
  wire u2__abc_44228_n20897;
  wire u2__abc_44228_n20898;
  wire u2__abc_44228_n20899;
  wire u2__abc_44228_n20900;
  wire u2__abc_44228_n20901;
  wire u2__abc_44228_n20902;
  wire u2__abc_44228_n20903;
  wire u2__abc_44228_n20904;
  wire u2__abc_44228_n20905;
  wire u2__abc_44228_n20907;
  wire u2__abc_44228_n20908;
  wire u2__abc_44228_n20909;
  wire u2__abc_44228_n20910;
  wire u2__abc_44228_n20911;
  wire u2__abc_44228_n20912;
  wire u2__abc_44228_n20913;
  wire u2__abc_44228_n20914;
  wire u2__abc_44228_n20915;
  wire u2__abc_44228_n20916;
  wire u2__abc_44228_n20917;
  wire u2__abc_44228_n20919;
  wire u2__abc_44228_n20920;
  wire u2__abc_44228_n20921;
  wire u2__abc_44228_n20922;
  wire u2__abc_44228_n20923;
  wire u2__abc_44228_n20924;
  wire u2__abc_44228_n20925;
  wire u2__abc_44228_n20926;
  wire u2__abc_44228_n20927;
  wire u2__abc_44228_n20928;
  wire u2__abc_44228_n20929;
  wire u2__abc_44228_n20931;
  wire u2__abc_44228_n20932;
  wire u2__abc_44228_n20933;
  wire u2__abc_44228_n20934;
  wire u2__abc_44228_n20935;
  wire u2__abc_44228_n20936;
  wire u2__abc_44228_n20937;
  wire u2__abc_44228_n20938;
  wire u2__abc_44228_n20939;
  wire u2__abc_44228_n20940;
  wire u2__abc_44228_n20941;
  wire u2__abc_44228_n20943;
  wire u2__abc_44228_n20944;
  wire u2__abc_44228_n20945;
  wire u2__abc_44228_n20946;
  wire u2__abc_44228_n20947;
  wire u2__abc_44228_n20948;
  wire u2__abc_44228_n20949;
  wire u2__abc_44228_n20950;
  wire u2__abc_44228_n20951;
  wire u2__abc_44228_n20952;
  wire u2__abc_44228_n20953;
  wire u2__abc_44228_n20955;
  wire u2__abc_44228_n20956;
  wire u2__abc_44228_n20957;
  wire u2__abc_44228_n20958;
  wire u2__abc_44228_n20959;
  wire u2__abc_44228_n20960;
  wire u2__abc_44228_n20961;
  wire u2__abc_44228_n20962;
  wire u2__abc_44228_n20963;
  wire u2__abc_44228_n20964;
  wire u2__abc_44228_n20965;
  wire u2__abc_44228_n20967;
  wire u2__abc_44228_n20968;
  wire u2__abc_44228_n20969;
  wire u2__abc_44228_n20970;
  wire u2__abc_44228_n20971;
  wire u2__abc_44228_n20972;
  wire u2__abc_44228_n20973;
  wire u2__abc_44228_n20974;
  wire u2__abc_44228_n20975;
  wire u2__abc_44228_n20976;
  wire u2__abc_44228_n20977;
  wire u2__abc_44228_n20979;
  wire u2__abc_44228_n20980;
  wire u2__abc_44228_n20981;
  wire u2__abc_44228_n20982;
  wire u2__abc_44228_n20983;
  wire u2__abc_44228_n20984;
  wire u2__abc_44228_n20985;
  wire u2__abc_44228_n20986;
  wire u2__abc_44228_n20987;
  wire u2__abc_44228_n20988;
  wire u2__abc_44228_n20989;
  wire u2__abc_44228_n20991;
  wire u2__abc_44228_n20992;
  wire u2__abc_44228_n20993;
  wire u2__abc_44228_n20994;
  wire u2__abc_44228_n20995;
  wire u2__abc_44228_n20996;
  wire u2__abc_44228_n20997;
  wire u2__abc_44228_n20998;
  wire u2__abc_44228_n20999;
  wire u2__abc_44228_n21000;
  wire u2__abc_44228_n21001;
  wire u2__abc_44228_n21003;
  wire u2__abc_44228_n21004;
  wire u2__abc_44228_n21005;
  wire u2__abc_44228_n21006;
  wire u2__abc_44228_n21007;
  wire u2__abc_44228_n21008;
  wire u2__abc_44228_n21009;
  wire u2__abc_44228_n21010;
  wire u2__abc_44228_n21011;
  wire u2__abc_44228_n21012;
  wire u2__abc_44228_n21013;
  wire u2__abc_44228_n21015;
  wire u2__abc_44228_n21016;
  wire u2__abc_44228_n21017;
  wire u2__abc_44228_n21018;
  wire u2__abc_44228_n21019;
  wire u2__abc_44228_n21020;
  wire u2__abc_44228_n21021;
  wire u2__abc_44228_n21022;
  wire u2__abc_44228_n21023;
  wire u2__abc_44228_n21024;
  wire u2__abc_44228_n21025;
  wire u2__abc_44228_n21027;
  wire u2__abc_44228_n21028;
  wire u2__abc_44228_n21029;
  wire u2__abc_44228_n21030;
  wire u2__abc_44228_n21031;
  wire u2__abc_44228_n21032;
  wire u2__abc_44228_n21033;
  wire u2__abc_44228_n21034;
  wire u2__abc_44228_n21035;
  wire u2__abc_44228_n21036;
  wire u2__abc_44228_n21037;
  wire u2__abc_44228_n21039;
  wire u2__abc_44228_n21040;
  wire u2__abc_44228_n21041;
  wire u2__abc_44228_n21042;
  wire u2__abc_44228_n21043;
  wire u2__abc_44228_n21044;
  wire u2__abc_44228_n21045;
  wire u2__abc_44228_n21046;
  wire u2__abc_44228_n21047;
  wire u2__abc_44228_n21048;
  wire u2__abc_44228_n21049;
  wire u2__abc_44228_n21051;
  wire u2__abc_44228_n21052;
  wire u2__abc_44228_n21053;
  wire u2__abc_44228_n21054;
  wire u2__abc_44228_n21055;
  wire u2__abc_44228_n21056;
  wire u2__abc_44228_n21057;
  wire u2__abc_44228_n21058;
  wire u2__abc_44228_n21059;
  wire u2__abc_44228_n21060;
  wire u2__abc_44228_n21061;
  wire u2__abc_44228_n21063;
  wire u2__abc_44228_n21064;
  wire u2__abc_44228_n21065;
  wire u2__abc_44228_n21066;
  wire u2__abc_44228_n21067;
  wire u2__abc_44228_n21068;
  wire u2__abc_44228_n21069;
  wire u2__abc_44228_n21070;
  wire u2__abc_44228_n21071;
  wire u2__abc_44228_n21072;
  wire u2__abc_44228_n21073;
  wire u2__abc_44228_n21075;
  wire u2__abc_44228_n21076;
  wire u2__abc_44228_n21077;
  wire u2__abc_44228_n21078;
  wire u2__abc_44228_n21079;
  wire u2__abc_44228_n21080;
  wire u2__abc_44228_n21081;
  wire u2__abc_44228_n21082;
  wire u2__abc_44228_n21083;
  wire u2__abc_44228_n21084;
  wire u2__abc_44228_n21085;
  wire u2__abc_44228_n21087;
  wire u2__abc_44228_n21088;
  wire u2__abc_44228_n21089;
  wire u2__abc_44228_n21090;
  wire u2__abc_44228_n21091;
  wire u2__abc_44228_n21092;
  wire u2__abc_44228_n21093;
  wire u2__abc_44228_n21094;
  wire u2__abc_44228_n21095;
  wire u2__abc_44228_n21096;
  wire u2__abc_44228_n21097;
  wire u2__abc_44228_n21099;
  wire u2__abc_44228_n21100;
  wire u2__abc_44228_n21101;
  wire u2__abc_44228_n21102;
  wire u2__abc_44228_n21103;
  wire u2__abc_44228_n21104;
  wire u2__abc_44228_n21105;
  wire u2__abc_44228_n21106;
  wire u2__abc_44228_n21107;
  wire u2__abc_44228_n21108;
  wire u2__abc_44228_n21109;
  wire u2__abc_44228_n21111;
  wire u2__abc_44228_n21112;
  wire u2__abc_44228_n21113;
  wire u2__abc_44228_n21114;
  wire u2__abc_44228_n21115;
  wire u2__abc_44228_n21116;
  wire u2__abc_44228_n21117;
  wire u2__abc_44228_n21118;
  wire u2__abc_44228_n21119;
  wire u2__abc_44228_n21120;
  wire u2__abc_44228_n21121;
  wire u2__abc_44228_n21123;
  wire u2__abc_44228_n21124;
  wire u2__abc_44228_n21125;
  wire u2__abc_44228_n21126;
  wire u2__abc_44228_n21127;
  wire u2__abc_44228_n21128;
  wire u2__abc_44228_n21129;
  wire u2__abc_44228_n21130;
  wire u2__abc_44228_n21131;
  wire u2__abc_44228_n21132;
  wire u2__abc_44228_n21133;
  wire u2__abc_44228_n21135;
  wire u2__abc_44228_n21136;
  wire u2__abc_44228_n21137;
  wire u2__abc_44228_n21138;
  wire u2__abc_44228_n21139;
  wire u2__abc_44228_n21140;
  wire u2__abc_44228_n21141;
  wire u2__abc_44228_n21142;
  wire u2__abc_44228_n21143;
  wire u2__abc_44228_n21144;
  wire u2__abc_44228_n21145;
  wire u2__abc_44228_n21147;
  wire u2__abc_44228_n21148;
  wire u2__abc_44228_n21149;
  wire u2__abc_44228_n21150;
  wire u2__abc_44228_n21151;
  wire u2__abc_44228_n21152;
  wire u2__abc_44228_n21153;
  wire u2__abc_44228_n21154;
  wire u2__abc_44228_n21155;
  wire u2__abc_44228_n21156;
  wire u2__abc_44228_n21157;
  wire u2__abc_44228_n21159;
  wire u2__abc_44228_n21160;
  wire u2__abc_44228_n21161;
  wire u2__abc_44228_n21162;
  wire u2__abc_44228_n21163;
  wire u2__abc_44228_n21164;
  wire u2__abc_44228_n21165;
  wire u2__abc_44228_n21166;
  wire u2__abc_44228_n21167;
  wire u2__abc_44228_n21168;
  wire u2__abc_44228_n21169;
  wire u2__abc_44228_n21171;
  wire u2__abc_44228_n21172;
  wire u2__abc_44228_n21173;
  wire u2__abc_44228_n21174;
  wire u2__abc_44228_n21175;
  wire u2__abc_44228_n21176;
  wire u2__abc_44228_n21177;
  wire u2__abc_44228_n21178;
  wire u2__abc_44228_n21179;
  wire u2__abc_44228_n21180;
  wire u2__abc_44228_n21181;
  wire u2__abc_44228_n21183;
  wire u2__abc_44228_n21184;
  wire u2__abc_44228_n21185;
  wire u2__abc_44228_n21186;
  wire u2__abc_44228_n21187;
  wire u2__abc_44228_n21188;
  wire u2__abc_44228_n21189;
  wire u2__abc_44228_n21190;
  wire u2__abc_44228_n21191;
  wire u2__abc_44228_n21192;
  wire u2__abc_44228_n21193;
  wire u2__abc_44228_n21195;
  wire u2__abc_44228_n21196;
  wire u2__abc_44228_n21197;
  wire u2__abc_44228_n21198;
  wire u2__abc_44228_n21199;
  wire u2__abc_44228_n21200;
  wire u2__abc_44228_n21201;
  wire u2__abc_44228_n21202;
  wire u2__abc_44228_n21203;
  wire u2__abc_44228_n21204;
  wire u2__abc_44228_n21205;
  wire u2__abc_44228_n21207;
  wire u2__abc_44228_n21208;
  wire u2__abc_44228_n21209;
  wire u2__abc_44228_n21210;
  wire u2__abc_44228_n21211;
  wire u2__abc_44228_n21212;
  wire u2__abc_44228_n21213;
  wire u2__abc_44228_n21214;
  wire u2__abc_44228_n21215;
  wire u2__abc_44228_n21216;
  wire u2__abc_44228_n21217;
  wire u2__abc_44228_n21219;
  wire u2__abc_44228_n21220;
  wire u2__abc_44228_n21221;
  wire u2__abc_44228_n21222;
  wire u2__abc_44228_n21223;
  wire u2__abc_44228_n21224;
  wire u2__abc_44228_n21225;
  wire u2__abc_44228_n21226;
  wire u2__abc_44228_n21227;
  wire u2__abc_44228_n21228;
  wire u2__abc_44228_n21229;
  wire u2__abc_44228_n21231;
  wire u2__abc_44228_n21232;
  wire u2__abc_44228_n21233;
  wire u2__abc_44228_n21234;
  wire u2__abc_44228_n21235;
  wire u2__abc_44228_n21236;
  wire u2__abc_44228_n21237;
  wire u2__abc_44228_n21238;
  wire u2__abc_44228_n21239;
  wire u2__abc_44228_n21240;
  wire u2__abc_44228_n21241;
  wire u2__abc_44228_n21243;
  wire u2__abc_44228_n21244;
  wire u2__abc_44228_n21245;
  wire u2__abc_44228_n21246;
  wire u2__abc_44228_n21247;
  wire u2__abc_44228_n21248;
  wire u2__abc_44228_n21249;
  wire u2__abc_44228_n21250;
  wire u2__abc_44228_n21251;
  wire u2__abc_44228_n21252;
  wire u2__abc_44228_n21253;
  wire u2__abc_44228_n21255;
  wire u2__abc_44228_n21256;
  wire u2__abc_44228_n21257;
  wire u2__abc_44228_n21258;
  wire u2__abc_44228_n21259;
  wire u2__abc_44228_n21260;
  wire u2__abc_44228_n21261;
  wire u2__abc_44228_n21262;
  wire u2__abc_44228_n21263;
  wire u2__abc_44228_n21264;
  wire u2__abc_44228_n21265;
  wire u2__abc_44228_n21267;
  wire u2__abc_44228_n21268;
  wire u2__abc_44228_n21269;
  wire u2__abc_44228_n21270;
  wire u2__abc_44228_n21271;
  wire u2__abc_44228_n21272;
  wire u2__abc_44228_n21273;
  wire u2__abc_44228_n21274;
  wire u2__abc_44228_n21275;
  wire u2__abc_44228_n21276;
  wire u2__abc_44228_n21277;
  wire u2__abc_44228_n21279;
  wire u2__abc_44228_n21280;
  wire u2__abc_44228_n21281;
  wire u2__abc_44228_n21282;
  wire u2__abc_44228_n21283;
  wire u2__abc_44228_n21284;
  wire u2__abc_44228_n21285;
  wire u2__abc_44228_n21286;
  wire u2__abc_44228_n21287;
  wire u2__abc_44228_n21288;
  wire u2__abc_44228_n21289;
  wire u2__abc_44228_n21291;
  wire u2__abc_44228_n21292;
  wire u2__abc_44228_n21293;
  wire u2__abc_44228_n21294;
  wire u2__abc_44228_n21295;
  wire u2__abc_44228_n21296;
  wire u2__abc_44228_n21297;
  wire u2__abc_44228_n21298;
  wire u2__abc_44228_n21299;
  wire u2__abc_44228_n21300;
  wire u2__abc_44228_n21301;
  wire u2__abc_44228_n21303;
  wire u2__abc_44228_n21304;
  wire u2__abc_44228_n21305;
  wire u2__abc_44228_n21306;
  wire u2__abc_44228_n21307;
  wire u2__abc_44228_n21308;
  wire u2__abc_44228_n21309;
  wire u2__abc_44228_n21310;
  wire u2__abc_44228_n21311;
  wire u2__abc_44228_n21312;
  wire u2__abc_44228_n21313;
  wire u2__abc_44228_n21315;
  wire u2__abc_44228_n21316;
  wire u2__abc_44228_n21317;
  wire u2__abc_44228_n21318;
  wire u2__abc_44228_n21319;
  wire u2__abc_44228_n21320;
  wire u2__abc_44228_n21321;
  wire u2__abc_44228_n21322;
  wire u2__abc_44228_n21323;
  wire u2__abc_44228_n21324;
  wire u2__abc_44228_n21325;
  wire u2__abc_44228_n21327;
  wire u2__abc_44228_n21328;
  wire u2__abc_44228_n21329;
  wire u2__abc_44228_n21330;
  wire u2__abc_44228_n21331;
  wire u2__abc_44228_n21332;
  wire u2__abc_44228_n21333;
  wire u2__abc_44228_n21334;
  wire u2__abc_44228_n21335;
  wire u2__abc_44228_n21336;
  wire u2__abc_44228_n21337;
  wire u2__abc_44228_n21339;
  wire u2__abc_44228_n21340;
  wire u2__abc_44228_n21341;
  wire u2__abc_44228_n21342;
  wire u2__abc_44228_n21343;
  wire u2__abc_44228_n21344;
  wire u2__abc_44228_n21345;
  wire u2__abc_44228_n21346;
  wire u2__abc_44228_n21347;
  wire u2__abc_44228_n21348;
  wire u2__abc_44228_n21349;
  wire u2__abc_44228_n21351;
  wire u2__abc_44228_n21352;
  wire u2__abc_44228_n21353;
  wire u2__abc_44228_n21354;
  wire u2__abc_44228_n21355;
  wire u2__abc_44228_n21356;
  wire u2__abc_44228_n21357;
  wire u2__abc_44228_n21358;
  wire u2__abc_44228_n21359;
  wire u2__abc_44228_n21360;
  wire u2__abc_44228_n21361;
  wire u2__abc_44228_n21363;
  wire u2__abc_44228_n21364;
  wire u2__abc_44228_n21365;
  wire u2__abc_44228_n21366;
  wire u2__abc_44228_n21367;
  wire u2__abc_44228_n21368;
  wire u2__abc_44228_n21369;
  wire u2__abc_44228_n21370;
  wire u2__abc_44228_n21371;
  wire u2__abc_44228_n21372;
  wire u2__abc_44228_n21373;
  wire u2__abc_44228_n21375;
  wire u2__abc_44228_n21376;
  wire u2__abc_44228_n21377;
  wire u2__abc_44228_n21378;
  wire u2__abc_44228_n21379;
  wire u2__abc_44228_n21380;
  wire u2__abc_44228_n21381;
  wire u2__abc_44228_n21382;
  wire u2__abc_44228_n21383;
  wire u2__abc_44228_n21384;
  wire u2__abc_44228_n21385;
  wire u2__abc_44228_n21387;
  wire u2__abc_44228_n21388;
  wire u2__abc_44228_n21389;
  wire u2__abc_44228_n21390;
  wire u2__abc_44228_n21391;
  wire u2__abc_44228_n21392;
  wire u2__abc_44228_n21393;
  wire u2__abc_44228_n21394;
  wire u2__abc_44228_n21395;
  wire u2__abc_44228_n21396;
  wire u2__abc_44228_n21397;
  wire u2__abc_44228_n21399;
  wire u2__abc_44228_n21400;
  wire u2__abc_44228_n21401;
  wire u2__abc_44228_n21402;
  wire u2__abc_44228_n21403;
  wire u2__abc_44228_n21404;
  wire u2__abc_44228_n21405;
  wire u2__abc_44228_n21406;
  wire u2__abc_44228_n21407;
  wire u2__abc_44228_n21408;
  wire u2__abc_44228_n21409;
  wire u2__abc_44228_n21411;
  wire u2__abc_44228_n21412;
  wire u2__abc_44228_n21413;
  wire u2__abc_44228_n21414;
  wire u2__abc_44228_n21415;
  wire u2__abc_44228_n21416;
  wire u2__abc_44228_n21417;
  wire u2__abc_44228_n21418;
  wire u2__abc_44228_n21419;
  wire u2__abc_44228_n21420;
  wire u2__abc_44228_n21421;
  wire u2__abc_44228_n21423;
  wire u2__abc_44228_n21424;
  wire u2__abc_44228_n21425;
  wire u2__abc_44228_n21426;
  wire u2__abc_44228_n21427;
  wire u2__abc_44228_n21428;
  wire u2__abc_44228_n21429;
  wire u2__abc_44228_n21430;
  wire u2__abc_44228_n21431;
  wire u2__abc_44228_n21432;
  wire u2__abc_44228_n21433;
  wire u2__abc_44228_n21435;
  wire u2__abc_44228_n21436;
  wire u2__abc_44228_n21437;
  wire u2__abc_44228_n21438;
  wire u2__abc_44228_n21439;
  wire u2__abc_44228_n21440;
  wire u2__abc_44228_n21441;
  wire u2__abc_44228_n21442;
  wire u2__abc_44228_n21443;
  wire u2__abc_44228_n21444;
  wire u2__abc_44228_n21445;
  wire u2__abc_44228_n21447;
  wire u2__abc_44228_n21448;
  wire u2__abc_44228_n21449;
  wire u2__abc_44228_n21450;
  wire u2__abc_44228_n21451;
  wire u2__abc_44228_n21452;
  wire u2__abc_44228_n21453;
  wire u2__abc_44228_n21454;
  wire u2__abc_44228_n21455;
  wire u2__abc_44228_n21456;
  wire u2__abc_44228_n21457;
  wire u2__abc_44228_n21459;
  wire u2__abc_44228_n21460;
  wire u2__abc_44228_n21461;
  wire u2__abc_44228_n21462;
  wire u2__abc_44228_n21463;
  wire u2__abc_44228_n21464;
  wire u2__abc_44228_n21465;
  wire u2__abc_44228_n21466;
  wire u2__abc_44228_n21467;
  wire u2__abc_44228_n21468;
  wire u2__abc_44228_n21469;
  wire u2__abc_44228_n21471;
  wire u2__abc_44228_n21472;
  wire u2__abc_44228_n21473;
  wire u2__abc_44228_n21474;
  wire u2__abc_44228_n21475;
  wire u2__abc_44228_n21476;
  wire u2__abc_44228_n21477;
  wire u2__abc_44228_n21478;
  wire u2__abc_44228_n21479;
  wire u2__abc_44228_n21480;
  wire u2__abc_44228_n21481;
  wire u2__abc_44228_n21483;
  wire u2__abc_44228_n21484;
  wire u2__abc_44228_n21485;
  wire u2__abc_44228_n21486;
  wire u2__abc_44228_n21487;
  wire u2__abc_44228_n21488;
  wire u2__abc_44228_n21489;
  wire u2__abc_44228_n21490;
  wire u2__abc_44228_n21491;
  wire u2__abc_44228_n21492;
  wire u2__abc_44228_n21493;
  wire u2__abc_44228_n21495;
  wire u2__abc_44228_n21496;
  wire u2__abc_44228_n21497;
  wire u2__abc_44228_n21498;
  wire u2__abc_44228_n21499;
  wire u2__abc_44228_n21500;
  wire u2__abc_44228_n21501;
  wire u2__abc_44228_n21502;
  wire u2__abc_44228_n21503;
  wire u2__abc_44228_n21504;
  wire u2__abc_44228_n21505;
  wire u2__abc_44228_n21507;
  wire u2__abc_44228_n21508;
  wire u2__abc_44228_n21509;
  wire u2__abc_44228_n21510;
  wire u2__abc_44228_n21511;
  wire u2__abc_44228_n21512;
  wire u2__abc_44228_n21513;
  wire u2__abc_44228_n21514;
  wire u2__abc_44228_n21515;
  wire u2__abc_44228_n21516;
  wire u2__abc_44228_n21517;
  wire u2__abc_44228_n21519;
  wire u2__abc_44228_n21520;
  wire u2__abc_44228_n21521;
  wire u2__abc_44228_n21522;
  wire u2__abc_44228_n21523;
  wire u2__abc_44228_n21524;
  wire u2__abc_44228_n21525;
  wire u2__abc_44228_n21526;
  wire u2__abc_44228_n21527;
  wire u2__abc_44228_n21528;
  wire u2__abc_44228_n21529;
  wire u2__abc_44228_n21531;
  wire u2__abc_44228_n21532;
  wire u2__abc_44228_n21533;
  wire u2__abc_44228_n21534;
  wire u2__abc_44228_n21535;
  wire u2__abc_44228_n21536;
  wire u2__abc_44228_n21537;
  wire u2__abc_44228_n21538;
  wire u2__abc_44228_n21539;
  wire u2__abc_44228_n21540;
  wire u2__abc_44228_n21541;
  wire u2__abc_44228_n21543;
  wire u2__abc_44228_n21544;
  wire u2__abc_44228_n21545;
  wire u2__abc_44228_n21546;
  wire u2__abc_44228_n21547;
  wire u2__abc_44228_n21548;
  wire u2__abc_44228_n21549;
  wire u2__abc_44228_n21550;
  wire u2__abc_44228_n21551;
  wire u2__abc_44228_n21552;
  wire u2__abc_44228_n21553;
  wire u2__abc_44228_n21555;
  wire u2__abc_44228_n21556;
  wire u2__abc_44228_n21557;
  wire u2__abc_44228_n21558;
  wire u2__abc_44228_n21559;
  wire u2__abc_44228_n21560;
  wire u2__abc_44228_n21561;
  wire u2__abc_44228_n21562;
  wire u2__abc_44228_n21563;
  wire u2__abc_44228_n21564;
  wire u2__abc_44228_n21565;
  wire u2__abc_44228_n21567;
  wire u2__abc_44228_n21568;
  wire u2__abc_44228_n21569;
  wire u2__abc_44228_n21570;
  wire u2__abc_44228_n21571;
  wire u2__abc_44228_n21572;
  wire u2__abc_44228_n21573;
  wire u2__abc_44228_n21574;
  wire u2__abc_44228_n21575;
  wire u2__abc_44228_n21576;
  wire u2__abc_44228_n21577;
  wire u2__abc_44228_n21579;
  wire u2__abc_44228_n21580;
  wire u2__abc_44228_n21581;
  wire u2__abc_44228_n21582;
  wire u2__abc_44228_n21583;
  wire u2__abc_44228_n21584;
  wire u2__abc_44228_n21585;
  wire u2__abc_44228_n21586;
  wire u2__abc_44228_n21587;
  wire u2__abc_44228_n21588;
  wire u2__abc_44228_n21589;
  wire u2__abc_44228_n21591;
  wire u2__abc_44228_n21592;
  wire u2__abc_44228_n21593;
  wire u2__abc_44228_n21594;
  wire u2__abc_44228_n21595;
  wire u2__abc_44228_n21596;
  wire u2__abc_44228_n21597;
  wire u2__abc_44228_n21598;
  wire u2__abc_44228_n21599;
  wire u2__abc_44228_n21600;
  wire u2__abc_44228_n21601;
  wire u2__abc_44228_n21603;
  wire u2__abc_44228_n21604;
  wire u2__abc_44228_n21605;
  wire u2__abc_44228_n21606;
  wire u2__abc_44228_n21607;
  wire u2__abc_44228_n21608;
  wire u2__abc_44228_n21609;
  wire u2__abc_44228_n21610;
  wire u2__abc_44228_n21611;
  wire u2__abc_44228_n21612;
  wire u2__abc_44228_n21613;
  wire u2__abc_44228_n21615;
  wire u2__abc_44228_n21616;
  wire u2__abc_44228_n21617;
  wire u2__abc_44228_n21618;
  wire u2__abc_44228_n21619;
  wire u2__abc_44228_n21620;
  wire u2__abc_44228_n21621;
  wire u2__abc_44228_n21622;
  wire u2__abc_44228_n21623;
  wire u2__abc_44228_n21624;
  wire u2__abc_44228_n21625;
  wire u2__abc_44228_n21627;
  wire u2__abc_44228_n21628;
  wire u2__abc_44228_n21629;
  wire u2__abc_44228_n21630;
  wire u2__abc_44228_n21631;
  wire u2__abc_44228_n21632;
  wire u2__abc_44228_n21633;
  wire u2__abc_44228_n21634;
  wire u2__abc_44228_n21635;
  wire u2__abc_44228_n21636;
  wire u2__abc_44228_n21637;
  wire u2__abc_44228_n21639;
  wire u2__abc_44228_n21640;
  wire u2__abc_44228_n21641;
  wire u2__abc_44228_n21642;
  wire u2__abc_44228_n21643;
  wire u2__abc_44228_n21644;
  wire u2__abc_44228_n21645;
  wire u2__abc_44228_n21646;
  wire u2__abc_44228_n21647;
  wire u2__abc_44228_n21648;
  wire u2__abc_44228_n21649;
  wire u2__abc_44228_n21651;
  wire u2__abc_44228_n21652;
  wire u2__abc_44228_n21653;
  wire u2__abc_44228_n21654;
  wire u2__abc_44228_n21655;
  wire u2__abc_44228_n21656;
  wire u2__abc_44228_n21657;
  wire u2__abc_44228_n21658;
  wire u2__abc_44228_n21659;
  wire u2__abc_44228_n21660;
  wire u2__abc_44228_n21661;
  wire u2__abc_44228_n21663;
  wire u2__abc_44228_n21664;
  wire u2__abc_44228_n21665;
  wire u2__abc_44228_n21666;
  wire u2__abc_44228_n21667;
  wire u2__abc_44228_n21668;
  wire u2__abc_44228_n21669;
  wire u2__abc_44228_n21670;
  wire u2__abc_44228_n21671;
  wire u2__abc_44228_n21672;
  wire u2__abc_44228_n21673;
  wire u2__abc_44228_n21675;
  wire u2__abc_44228_n21676;
  wire u2__abc_44228_n21677;
  wire u2__abc_44228_n21678;
  wire u2__abc_44228_n21679;
  wire u2__abc_44228_n21680;
  wire u2__abc_44228_n21681;
  wire u2__abc_44228_n21682;
  wire u2__abc_44228_n21683;
  wire u2__abc_44228_n21684;
  wire u2__abc_44228_n21685;
  wire u2__abc_44228_n21687;
  wire u2__abc_44228_n21688;
  wire u2__abc_44228_n21689;
  wire u2__abc_44228_n21690;
  wire u2__abc_44228_n21691;
  wire u2__abc_44228_n21692;
  wire u2__abc_44228_n21693;
  wire u2__abc_44228_n21694;
  wire u2__abc_44228_n21695;
  wire u2__abc_44228_n21696;
  wire u2__abc_44228_n21697;
  wire u2__abc_44228_n21699;
  wire u2__abc_44228_n21700;
  wire u2__abc_44228_n21701;
  wire u2__abc_44228_n21702;
  wire u2__abc_44228_n21703;
  wire u2__abc_44228_n21704;
  wire u2__abc_44228_n21705;
  wire u2__abc_44228_n21706;
  wire u2__abc_44228_n21707;
  wire u2__abc_44228_n21708;
  wire u2__abc_44228_n21709;
  wire u2__abc_44228_n21711;
  wire u2__abc_44228_n21712;
  wire u2__abc_44228_n21713;
  wire u2__abc_44228_n21714;
  wire u2__abc_44228_n21715;
  wire u2__abc_44228_n21716;
  wire u2__abc_44228_n21717;
  wire u2__abc_44228_n21718;
  wire u2__abc_44228_n21719;
  wire u2__abc_44228_n21720;
  wire u2__abc_44228_n21721;
  wire u2__abc_44228_n21723;
  wire u2__abc_44228_n21724;
  wire u2__abc_44228_n21725;
  wire u2__abc_44228_n21726;
  wire u2__abc_44228_n21727;
  wire u2__abc_44228_n21728;
  wire u2__abc_44228_n21729;
  wire u2__abc_44228_n21730;
  wire u2__abc_44228_n21731;
  wire u2__abc_44228_n21732;
  wire u2__abc_44228_n21733;
  wire u2__abc_44228_n21735;
  wire u2__abc_44228_n21736;
  wire u2__abc_44228_n21737;
  wire u2__abc_44228_n21738;
  wire u2__abc_44228_n21739;
  wire u2__abc_44228_n21740;
  wire u2__abc_44228_n21741;
  wire u2__abc_44228_n21742;
  wire u2__abc_44228_n21743;
  wire u2__abc_44228_n21744;
  wire u2__abc_44228_n21745;
  wire u2__abc_44228_n21747;
  wire u2__abc_44228_n21748;
  wire u2__abc_44228_n21749;
  wire u2__abc_44228_n21750;
  wire u2__abc_44228_n21751;
  wire u2__abc_44228_n21752;
  wire u2__abc_44228_n21753;
  wire u2__abc_44228_n21754;
  wire u2__abc_44228_n21755;
  wire u2__abc_44228_n21756;
  wire u2__abc_44228_n21757;
  wire u2__abc_44228_n21759;
  wire u2__abc_44228_n21760;
  wire u2__abc_44228_n21761;
  wire u2__abc_44228_n21762;
  wire u2__abc_44228_n21763;
  wire u2__abc_44228_n21764;
  wire u2__abc_44228_n21765;
  wire u2__abc_44228_n21766;
  wire u2__abc_44228_n21767;
  wire u2__abc_44228_n21768;
  wire u2__abc_44228_n21769;
  wire u2__abc_44228_n21771;
  wire u2__abc_44228_n21772;
  wire u2__abc_44228_n21773;
  wire u2__abc_44228_n21774;
  wire u2__abc_44228_n21775;
  wire u2__abc_44228_n21776;
  wire u2__abc_44228_n21777;
  wire u2__abc_44228_n21778;
  wire u2__abc_44228_n21779;
  wire u2__abc_44228_n21780;
  wire u2__abc_44228_n21781;
  wire u2__abc_44228_n21783;
  wire u2__abc_44228_n21784;
  wire u2__abc_44228_n21785;
  wire u2__abc_44228_n21786;
  wire u2__abc_44228_n21787;
  wire u2__abc_44228_n21788;
  wire u2__abc_44228_n21789;
  wire u2__abc_44228_n21790;
  wire u2__abc_44228_n21791;
  wire u2__abc_44228_n21792;
  wire u2__abc_44228_n21793;
  wire u2__abc_44228_n21795;
  wire u2__abc_44228_n21796;
  wire u2__abc_44228_n21797;
  wire u2__abc_44228_n21798;
  wire u2__abc_44228_n21799;
  wire u2__abc_44228_n21800;
  wire u2__abc_44228_n21801;
  wire u2__abc_44228_n21802;
  wire u2__abc_44228_n21803;
  wire u2__abc_44228_n21804;
  wire u2__abc_44228_n21805;
  wire u2__abc_44228_n21807;
  wire u2__abc_44228_n21808;
  wire u2__abc_44228_n21809;
  wire u2__abc_44228_n21810;
  wire u2__abc_44228_n21811;
  wire u2__abc_44228_n21812;
  wire u2__abc_44228_n21813;
  wire u2__abc_44228_n21814;
  wire u2__abc_44228_n21815;
  wire u2__abc_44228_n21816;
  wire u2__abc_44228_n21817;
  wire u2__abc_44228_n21819;
  wire u2__abc_44228_n21820;
  wire u2__abc_44228_n21821;
  wire u2__abc_44228_n21822;
  wire u2__abc_44228_n21823;
  wire u2__abc_44228_n21824;
  wire u2__abc_44228_n21825;
  wire u2__abc_44228_n21826;
  wire u2__abc_44228_n21827;
  wire u2__abc_44228_n21828;
  wire u2__abc_44228_n21829;
  wire u2__abc_44228_n21831;
  wire u2__abc_44228_n21832;
  wire u2__abc_44228_n21833;
  wire u2__abc_44228_n21834;
  wire u2__abc_44228_n21835;
  wire u2__abc_44228_n21836;
  wire u2__abc_44228_n21837;
  wire u2__abc_44228_n21838;
  wire u2__abc_44228_n21839;
  wire u2__abc_44228_n21840;
  wire u2__abc_44228_n21841;
  wire u2__abc_44228_n21843;
  wire u2__abc_44228_n21844;
  wire u2__abc_44228_n21845;
  wire u2__abc_44228_n21846;
  wire u2__abc_44228_n21847;
  wire u2__abc_44228_n21848;
  wire u2__abc_44228_n21849;
  wire u2__abc_44228_n21850;
  wire u2__abc_44228_n21851;
  wire u2__abc_44228_n21852;
  wire u2__abc_44228_n21853;
  wire u2__abc_44228_n21855;
  wire u2__abc_44228_n21856;
  wire u2__abc_44228_n21857;
  wire u2__abc_44228_n21858;
  wire u2__abc_44228_n21859;
  wire u2__abc_44228_n21860;
  wire u2__abc_44228_n21861;
  wire u2__abc_44228_n21862;
  wire u2__abc_44228_n21863;
  wire u2__abc_44228_n21864;
  wire u2__abc_44228_n21865;
  wire u2__abc_44228_n21867;
  wire u2__abc_44228_n21868;
  wire u2__abc_44228_n21869;
  wire u2__abc_44228_n21870;
  wire u2__abc_44228_n21871;
  wire u2__abc_44228_n21872;
  wire u2__abc_44228_n21873;
  wire u2__abc_44228_n21874;
  wire u2__abc_44228_n21875;
  wire u2__abc_44228_n21876;
  wire u2__abc_44228_n21877;
  wire u2__abc_44228_n21879;
  wire u2__abc_44228_n21880;
  wire u2__abc_44228_n21881;
  wire u2__abc_44228_n21882;
  wire u2__abc_44228_n21883;
  wire u2__abc_44228_n21884;
  wire u2__abc_44228_n21885;
  wire u2__abc_44228_n21886;
  wire u2__abc_44228_n21887;
  wire u2__abc_44228_n21888;
  wire u2__abc_44228_n21889;
  wire u2__abc_44228_n21891;
  wire u2__abc_44228_n21892;
  wire u2__abc_44228_n21893;
  wire u2__abc_44228_n21894;
  wire u2__abc_44228_n21895;
  wire u2__abc_44228_n21896;
  wire u2__abc_44228_n21897;
  wire u2__abc_44228_n21898;
  wire u2__abc_44228_n21899;
  wire u2__abc_44228_n21900;
  wire u2__abc_44228_n21901;
  wire u2__abc_44228_n21903;
  wire u2__abc_44228_n21904;
  wire u2__abc_44228_n21905;
  wire u2__abc_44228_n21906;
  wire u2__abc_44228_n21907;
  wire u2__abc_44228_n21908;
  wire u2__abc_44228_n21909;
  wire u2__abc_44228_n21910;
  wire u2__abc_44228_n21911;
  wire u2__abc_44228_n21912;
  wire u2__abc_44228_n21913;
  wire u2__abc_44228_n21915;
  wire u2__abc_44228_n21916;
  wire u2__abc_44228_n21917;
  wire u2__abc_44228_n21918;
  wire u2__abc_44228_n21919;
  wire u2__abc_44228_n21920;
  wire u2__abc_44228_n21921;
  wire u2__abc_44228_n21922;
  wire u2__abc_44228_n21923;
  wire u2__abc_44228_n21924;
  wire u2__abc_44228_n21925;
  wire u2__abc_44228_n21927;
  wire u2__abc_44228_n21928;
  wire u2__abc_44228_n21929;
  wire u2__abc_44228_n21930;
  wire u2__abc_44228_n21931;
  wire u2__abc_44228_n21932;
  wire u2__abc_44228_n21933;
  wire u2__abc_44228_n21934;
  wire u2__abc_44228_n21935;
  wire u2__abc_44228_n21936;
  wire u2__abc_44228_n21937;
  wire u2__abc_44228_n21939;
  wire u2__abc_44228_n21940;
  wire u2__abc_44228_n21941;
  wire u2__abc_44228_n21942;
  wire u2__abc_44228_n21943;
  wire u2__abc_44228_n21944;
  wire u2__abc_44228_n21945;
  wire u2__abc_44228_n21946;
  wire u2__abc_44228_n21947;
  wire u2__abc_44228_n21948;
  wire u2__abc_44228_n21949;
  wire u2__abc_44228_n21951;
  wire u2__abc_44228_n21952;
  wire u2__abc_44228_n21953;
  wire u2__abc_44228_n21954;
  wire u2__abc_44228_n21955;
  wire u2__abc_44228_n21956;
  wire u2__abc_44228_n21957;
  wire u2__abc_44228_n21958;
  wire u2__abc_44228_n21959;
  wire u2__abc_44228_n21960;
  wire u2__abc_44228_n21961;
  wire u2__abc_44228_n21963;
  wire u2__abc_44228_n21964;
  wire u2__abc_44228_n21965;
  wire u2__abc_44228_n21966;
  wire u2__abc_44228_n21967;
  wire u2__abc_44228_n21968;
  wire u2__abc_44228_n21969;
  wire u2__abc_44228_n21970;
  wire u2__abc_44228_n21971;
  wire u2__abc_44228_n21972;
  wire u2__abc_44228_n21973;
  wire u2__abc_44228_n21975;
  wire u2__abc_44228_n21976;
  wire u2__abc_44228_n21977;
  wire u2__abc_44228_n21978;
  wire u2__abc_44228_n21979;
  wire u2__abc_44228_n21980;
  wire u2__abc_44228_n21981;
  wire u2__abc_44228_n21982;
  wire u2__abc_44228_n21983;
  wire u2__abc_44228_n21984;
  wire u2__abc_44228_n21985;
  wire u2__abc_44228_n21987;
  wire u2__abc_44228_n21988;
  wire u2__abc_44228_n21989;
  wire u2__abc_44228_n21990;
  wire u2__abc_44228_n21991;
  wire u2__abc_44228_n21992;
  wire u2__abc_44228_n21993;
  wire u2__abc_44228_n21994;
  wire u2__abc_44228_n21995;
  wire u2__abc_44228_n21996;
  wire u2__abc_44228_n21997;
  wire u2__abc_44228_n21999;
  wire u2__abc_44228_n22000;
  wire u2__abc_44228_n22001;
  wire u2__abc_44228_n22002;
  wire u2__abc_44228_n22003;
  wire u2__abc_44228_n22004;
  wire u2__abc_44228_n22005;
  wire u2__abc_44228_n22006;
  wire u2__abc_44228_n22007;
  wire u2__abc_44228_n22008;
  wire u2__abc_44228_n22009;
  wire u2__abc_44228_n22011;
  wire u2__abc_44228_n22012;
  wire u2__abc_44228_n22013;
  wire u2__abc_44228_n22014;
  wire u2__abc_44228_n22015;
  wire u2__abc_44228_n22016;
  wire u2__abc_44228_n22017;
  wire u2__abc_44228_n22018;
  wire u2__abc_44228_n22019;
  wire u2__abc_44228_n22020;
  wire u2__abc_44228_n22021;
  wire u2__abc_44228_n22023;
  wire u2__abc_44228_n22024;
  wire u2__abc_44228_n22025;
  wire u2__abc_44228_n22026;
  wire u2__abc_44228_n22027;
  wire u2__abc_44228_n22028;
  wire u2__abc_44228_n22029;
  wire u2__abc_44228_n22030;
  wire u2__abc_44228_n22031;
  wire u2__abc_44228_n22032;
  wire u2__abc_44228_n22033;
  wire u2__abc_44228_n22035;
  wire u2__abc_44228_n22036;
  wire u2__abc_44228_n22037;
  wire u2__abc_44228_n22038;
  wire u2__abc_44228_n22039;
  wire u2__abc_44228_n22040;
  wire u2__abc_44228_n22041;
  wire u2__abc_44228_n22042;
  wire u2__abc_44228_n22043;
  wire u2__abc_44228_n22044;
  wire u2__abc_44228_n22045;
  wire u2__abc_44228_n22047;
  wire u2__abc_44228_n22048;
  wire u2__abc_44228_n22049;
  wire u2__abc_44228_n22050;
  wire u2__abc_44228_n22051;
  wire u2__abc_44228_n22052;
  wire u2__abc_44228_n22053;
  wire u2__abc_44228_n22054;
  wire u2__abc_44228_n22055;
  wire u2__abc_44228_n22056;
  wire u2__abc_44228_n22057;
  wire u2__abc_44228_n22059;
  wire u2__abc_44228_n22060;
  wire u2__abc_44228_n22061;
  wire u2__abc_44228_n22062;
  wire u2__abc_44228_n22063;
  wire u2__abc_44228_n22064;
  wire u2__abc_44228_n22065;
  wire u2__abc_44228_n22066;
  wire u2__abc_44228_n22067;
  wire u2__abc_44228_n22068;
  wire u2__abc_44228_n22069;
  wire u2__abc_44228_n22071;
  wire u2__abc_44228_n22072;
  wire u2__abc_44228_n22073;
  wire u2__abc_44228_n22074;
  wire u2__abc_44228_n22075;
  wire u2__abc_44228_n22076;
  wire u2__abc_44228_n22077;
  wire u2__abc_44228_n22078;
  wire u2__abc_44228_n22079;
  wire u2__abc_44228_n22080;
  wire u2__abc_44228_n22081;
  wire u2__abc_44228_n22083;
  wire u2__abc_44228_n22084;
  wire u2__abc_44228_n22085;
  wire u2__abc_44228_n22086;
  wire u2__abc_44228_n22087;
  wire u2__abc_44228_n22088;
  wire u2__abc_44228_n22089;
  wire u2__abc_44228_n22090;
  wire u2__abc_44228_n22091;
  wire u2__abc_44228_n22092;
  wire u2__abc_44228_n22093;
  wire u2__abc_44228_n22095;
  wire u2__abc_44228_n22096;
  wire u2__abc_44228_n22097;
  wire u2__abc_44228_n22098;
  wire u2__abc_44228_n22099;
  wire u2__abc_44228_n22100;
  wire u2__abc_44228_n22101;
  wire u2__abc_44228_n22102;
  wire u2__abc_44228_n22103;
  wire u2__abc_44228_n22104;
  wire u2__abc_44228_n22105;
  wire u2__abc_44228_n22107;
  wire u2__abc_44228_n22108;
  wire u2__abc_44228_n22109;
  wire u2__abc_44228_n22110;
  wire u2__abc_44228_n22111;
  wire u2__abc_44228_n22112;
  wire u2__abc_44228_n22113;
  wire u2__abc_44228_n22114;
  wire u2__abc_44228_n22115;
  wire u2__abc_44228_n22116;
  wire u2__abc_44228_n22117;
  wire u2__abc_44228_n22119;
  wire u2__abc_44228_n22120;
  wire u2__abc_44228_n22121;
  wire u2__abc_44228_n22122;
  wire u2__abc_44228_n22123;
  wire u2__abc_44228_n22124;
  wire u2__abc_44228_n22125;
  wire u2__abc_44228_n22126;
  wire u2__abc_44228_n22127;
  wire u2__abc_44228_n22128;
  wire u2__abc_44228_n22129;
  wire u2__abc_44228_n22131;
  wire u2__abc_44228_n22132;
  wire u2__abc_44228_n22133;
  wire u2__abc_44228_n22134;
  wire u2__abc_44228_n22135;
  wire u2__abc_44228_n22136;
  wire u2__abc_44228_n22137;
  wire u2__abc_44228_n22138;
  wire u2__abc_44228_n22139;
  wire u2__abc_44228_n22140;
  wire u2__abc_44228_n22141;
  wire u2__abc_44228_n22143;
  wire u2__abc_44228_n22144;
  wire u2__abc_44228_n22145;
  wire u2__abc_44228_n22146;
  wire u2__abc_44228_n22147;
  wire u2__abc_44228_n22148;
  wire u2__abc_44228_n22149;
  wire u2__abc_44228_n22150;
  wire u2__abc_44228_n22151;
  wire u2__abc_44228_n22152;
  wire u2__abc_44228_n22153;
  wire u2__abc_44228_n22155;
  wire u2__abc_44228_n22156;
  wire u2__abc_44228_n22157;
  wire u2__abc_44228_n22158;
  wire u2__abc_44228_n22159;
  wire u2__abc_44228_n22160;
  wire u2__abc_44228_n22161;
  wire u2__abc_44228_n22162;
  wire u2__abc_44228_n22163;
  wire u2__abc_44228_n22164;
  wire u2__abc_44228_n22165;
  wire u2__abc_44228_n22167;
  wire u2__abc_44228_n22168;
  wire u2__abc_44228_n22169;
  wire u2__abc_44228_n22170;
  wire u2__abc_44228_n22171;
  wire u2__abc_44228_n22172;
  wire u2__abc_44228_n22173;
  wire u2__abc_44228_n22174;
  wire u2__abc_44228_n22175;
  wire u2__abc_44228_n22176;
  wire u2__abc_44228_n22177;
  wire u2__abc_44228_n22179;
  wire u2__abc_44228_n22180;
  wire u2__abc_44228_n22181;
  wire u2__abc_44228_n22182;
  wire u2__abc_44228_n22183;
  wire u2__abc_44228_n22184;
  wire u2__abc_44228_n22185;
  wire u2__abc_44228_n22186;
  wire u2__abc_44228_n22187;
  wire u2__abc_44228_n22188;
  wire u2__abc_44228_n22189;
  wire u2__abc_44228_n22191;
  wire u2__abc_44228_n22192;
  wire u2__abc_44228_n22193;
  wire u2__abc_44228_n22194;
  wire u2__abc_44228_n22195;
  wire u2__abc_44228_n22196;
  wire u2__abc_44228_n22197;
  wire u2__abc_44228_n22198;
  wire u2__abc_44228_n22199;
  wire u2__abc_44228_n22200;
  wire u2__abc_44228_n22201;
  wire u2__abc_44228_n22203;
  wire u2__abc_44228_n22204;
  wire u2__abc_44228_n22205;
  wire u2__abc_44228_n22206;
  wire u2__abc_44228_n22207;
  wire u2__abc_44228_n22208;
  wire u2__abc_44228_n22209;
  wire u2__abc_44228_n22210;
  wire u2__abc_44228_n22211;
  wire u2__abc_44228_n22212;
  wire u2__abc_44228_n22213;
  wire u2__abc_44228_n22215;
  wire u2__abc_44228_n22216;
  wire u2__abc_44228_n22217;
  wire u2__abc_44228_n22218;
  wire u2__abc_44228_n22219;
  wire u2__abc_44228_n22220;
  wire u2__abc_44228_n22221;
  wire u2__abc_44228_n22222;
  wire u2__abc_44228_n22223;
  wire u2__abc_44228_n22224;
  wire u2__abc_44228_n22225;
  wire u2__abc_44228_n22227;
  wire u2__abc_44228_n22228;
  wire u2__abc_44228_n22229;
  wire u2__abc_44228_n22230;
  wire u2__abc_44228_n22231;
  wire u2__abc_44228_n22232;
  wire u2__abc_44228_n22233;
  wire u2__abc_44228_n22234;
  wire u2__abc_44228_n22235;
  wire u2__abc_44228_n22236;
  wire u2__abc_44228_n22237;
  wire u2__abc_44228_n22239;
  wire u2__abc_44228_n22240;
  wire u2__abc_44228_n22241;
  wire u2__abc_44228_n22242;
  wire u2__abc_44228_n22243;
  wire u2__abc_44228_n22244;
  wire u2__abc_44228_n22245;
  wire u2__abc_44228_n22246;
  wire u2__abc_44228_n22247;
  wire u2__abc_44228_n22248;
  wire u2__abc_44228_n22249;
  wire u2__abc_44228_n22251;
  wire u2__abc_44228_n22252;
  wire u2__abc_44228_n22253;
  wire u2__abc_44228_n22254;
  wire u2__abc_44228_n22255;
  wire u2__abc_44228_n22256;
  wire u2__abc_44228_n22257;
  wire u2__abc_44228_n22258;
  wire u2__abc_44228_n22259;
  wire u2__abc_44228_n22260;
  wire u2__abc_44228_n22261;
  wire u2__abc_44228_n22263;
  wire u2__abc_44228_n22264;
  wire u2__abc_44228_n22265;
  wire u2__abc_44228_n22266;
  wire u2__abc_44228_n22267;
  wire u2__abc_44228_n22268;
  wire u2__abc_44228_n22269;
  wire u2__abc_44228_n22270;
  wire u2__abc_44228_n22271;
  wire u2__abc_44228_n22272;
  wire u2__abc_44228_n22273;
  wire u2__abc_44228_n22275;
  wire u2__abc_44228_n22276;
  wire u2__abc_44228_n22277;
  wire u2__abc_44228_n22278;
  wire u2__abc_44228_n22279;
  wire u2__abc_44228_n22280;
  wire u2__abc_44228_n22281;
  wire u2__abc_44228_n22282;
  wire u2__abc_44228_n22283;
  wire u2__abc_44228_n22284;
  wire u2__abc_44228_n22285;
  wire u2__abc_44228_n22287;
  wire u2__abc_44228_n22288;
  wire u2__abc_44228_n22289;
  wire u2__abc_44228_n22290;
  wire u2__abc_44228_n22291;
  wire u2__abc_44228_n22292;
  wire u2__abc_44228_n22293;
  wire u2__abc_44228_n22294;
  wire u2__abc_44228_n22295;
  wire u2__abc_44228_n22296;
  wire u2__abc_44228_n22297;
  wire u2__abc_44228_n22299;
  wire u2__abc_44228_n22300;
  wire u2__abc_44228_n22301;
  wire u2__abc_44228_n22302;
  wire u2__abc_44228_n22303;
  wire u2__abc_44228_n22304;
  wire u2__abc_44228_n22305;
  wire u2__abc_44228_n22306;
  wire u2__abc_44228_n22307;
  wire u2__abc_44228_n22308;
  wire u2__abc_44228_n22309;
  wire u2__abc_44228_n22311;
  wire u2__abc_44228_n22312;
  wire u2__abc_44228_n22313;
  wire u2__abc_44228_n22314;
  wire u2__abc_44228_n22315;
  wire u2__abc_44228_n22316;
  wire u2__abc_44228_n22317;
  wire u2__abc_44228_n22318;
  wire u2__abc_44228_n22319;
  wire u2__abc_44228_n22320;
  wire u2__abc_44228_n22321;
  wire u2__abc_44228_n22323;
  wire u2__abc_44228_n22324;
  wire u2__abc_44228_n22325;
  wire u2__abc_44228_n22326;
  wire u2__abc_44228_n22327;
  wire u2__abc_44228_n22328;
  wire u2__abc_44228_n22329;
  wire u2__abc_44228_n22330;
  wire u2__abc_44228_n22331;
  wire u2__abc_44228_n22332;
  wire u2__abc_44228_n22333;
  wire u2__abc_44228_n22335;
  wire u2__abc_44228_n22336;
  wire u2__abc_44228_n22337;
  wire u2__abc_44228_n22338;
  wire u2__abc_44228_n22339;
  wire u2__abc_44228_n22340;
  wire u2__abc_44228_n22341;
  wire u2__abc_44228_n22342;
  wire u2__abc_44228_n22343;
  wire u2__abc_44228_n22344;
  wire u2__abc_44228_n22345;
  wire u2__abc_44228_n22347;
  wire u2__abc_44228_n22348;
  wire u2__abc_44228_n22349;
  wire u2__abc_44228_n22350;
  wire u2__abc_44228_n22351;
  wire u2__abc_44228_n22352;
  wire u2__abc_44228_n22353;
  wire u2__abc_44228_n22354;
  wire u2__abc_44228_n22355;
  wire u2__abc_44228_n22356;
  wire u2__abc_44228_n22357;
  wire u2__abc_44228_n22359;
  wire u2__abc_44228_n22360;
  wire u2__abc_44228_n22361;
  wire u2__abc_44228_n22362;
  wire u2__abc_44228_n22363;
  wire u2__abc_44228_n22364;
  wire u2__abc_44228_n22365;
  wire u2__abc_44228_n22366;
  wire u2__abc_44228_n22367;
  wire u2__abc_44228_n22368;
  wire u2__abc_44228_n22369;
  wire u2__abc_44228_n22371;
  wire u2__abc_44228_n22372;
  wire u2__abc_44228_n22373;
  wire u2__abc_44228_n22374;
  wire u2__abc_44228_n22375;
  wire u2__abc_44228_n22376;
  wire u2__abc_44228_n22377;
  wire u2__abc_44228_n22378;
  wire u2__abc_44228_n22379;
  wire u2__abc_44228_n22380;
  wire u2__abc_44228_n22381;
  wire u2__abc_44228_n22383;
  wire u2__abc_44228_n22384;
  wire u2__abc_44228_n22385;
  wire u2__abc_44228_n22386;
  wire u2__abc_44228_n22387;
  wire u2__abc_44228_n22388;
  wire u2__abc_44228_n22389;
  wire u2__abc_44228_n22390;
  wire u2__abc_44228_n22391;
  wire u2__abc_44228_n22392;
  wire u2__abc_44228_n22393;
  wire u2__abc_44228_n22395;
  wire u2__abc_44228_n22396;
  wire u2__abc_44228_n22397;
  wire u2__abc_44228_n22398;
  wire u2__abc_44228_n22399;
  wire u2__abc_44228_n22400;
  wire u2__abc_44228_n22401;
  wire u2__abc_44228_n22402;
  wire u2__abc_44228_n22403;
  wire u2__abc_44228_n22404;
  wire u2__abc_44228_n22405;
  wire u2__abc_44228_n22407;
  wire u2__abc_44228_n22408;
  wire u2__abc_44228_n22409;
  wire u2__abc_44228_n22410;
  wire u2__abc_44228_n22411;
  wire u2__abc_44228_n22412;
  wire u2__abc_44228_n22413;
  wire u2__abc_44228_n22414;
  wire u2__abc_44228_n22415;
  wire u2__abc_44228_n22416;
  wire u2__abc_44228_n22417;
  wire u2__abc_44228_n22419;
  wire u2__abc_44228_n22420;
  wire u2__abc_44228_n22421;
  wire u2__abc_44228_n22422;
  wire u2__abc_44228_n22423;
  wire u2__abc_44228_n22424;
  wire u2__abc_44228_n22425;
  wire u2__abc_44228_n22426;
  wire u2__abc_44228_n22427;
  wire u2__abc_44228_n22428;
  wire u2__abc_44228_n22429;
  wire u2__abc_44228_n22431;
  wire u2__abc_44228_n22432;
  wire u2__abc_44228_n22433;
  wire u2__abc_44228_n22434;
  wire u2__abc_44228_n22435;
  wire u2__abc_44228_n22436;
  wire u2__abc_44228_n22437;
  wire u2__abc_44228_n22438;
  wire u2__abc_44228_n22439;
  wire u2__abc_44228_n22440;
  wire u2__abc_44228_n22441;
  wire u2__abc_44228_n22443;
  wire u2__abc_44228_n22444;
  wire u2__abc_44228_n22445;
  wire u2__abc_44228_n22446;
  wire u2__abc_44228_n22447;
  wire u2__abc_44228_n22448;
  wire u2__abc_44228_n22449;
  wire u2__abc_44228_n22450;
  wire u2__abc_44228_n22451;
  wire u2__abc_44228_n22452;
  wire u2__abc_44228_n22453;
  wire u2__abc_44228_n22455;
  wire u2__abc_44228_n22456;
  wire u2__abc_44228_n22457;
  wire u2__abc_44228_n22458;
  wire u2__abc_44228_n22459;
  wire u2__abc_44228_n22460;
  wire u2__abc_44228_n22461;
  wire u2__abc_44228_n22462;
  wire u2__abc_44228_n22463;
  wire u2__abc_44228_n22464;
  wire u2__abc_44228_n22465;
  wire u2__abc_44228_n22467;
  wire u2__abc_44228_n22468;
  wire u2__abc_44228_n22469;
  wire u2__abc_44228_n22470;
  wire u2__abc_44228_n22471;
  wire u2__abc_44228_n22472;
  wire u2__abc_44228_n22473;
  wire u2__abc_44228_n22474;
  wire u2__abc_44228_n22475;
  wire u2__abc_44228_n22476;
  wire u2__abc_44228_n22477;
  wire u2__abc_44228_n22479;
  wire u2__abc_44228_n22480;
  wire u2__abc_44228_n22481;
  wire u2__abc_44228_n22482;
  wire u2__abc_44228_n22483;
  wire u2__abc_44228_n22484;
  wire u2__abc_44228_n22485;
  wire u2__abc_44228_n22486;
  wire u2__abc_44228_n22487;
  wire u2__abc_44228_n22488;
  wire u2__abc_44228_n22489;
  wire u2__abc_44228_n22491;
  wire u2__abc_44228_n22492;
  wire u2__abc_44228_n22493;
  wire u2__abc_44228_n22494;
  wire u2__abc_44228_n22495;
  wire u2__abc_44228_n22496;
  wire u2__abc_44228_n22497;
  wire u2__abc_44228_n22498;
  wire u2__abc_44228_n22499;
  wire u2__abc_44228_n22500;
  wire u2__abc_44228_n22501;
  wire u2__abc_44228_n22503;
  wire u2__abc_44228_n22504;
  wire u2__abc_44228_n22505;
  wire u2__abc_44228_n22506;
  wire u2__abc_44228_n22507;
  wire u2__abc_44228_n22508;
  wire u2__abc_44228_n22509;
  wire u2__abc_44228_n22510;
  wire u2__abc_44228_n22511;
  wire u2__abc_44228_n22512;
  wire u2__abc_44228_n22513;
  wire u2__abc_44228_n22515;
  wire u2__abc_44228_n22516;
  wire u2__abc_44228_n22517;
  wire u2__abc_44228_n22518;
  wire u2__abc_44228_n22519;
  wire u2__abc_44228_n22520;
  wire u2__abc_44228_n22521;
  wire u2__abc_44228_n22522;
  wire u2__abc_44228_n22523;
  wire u2__abc_44228_n22524;
  wire u2__abc_44228_n22525;
  wire u2__abc_44228_n22527;
  wire u2__abc_44228_n22528;
  wire u2__abc_44228_n22529;
  wire u2__abc_44228_n22530;
  wire u2__abc_44228_n22531;
  wire u2__abc_44228_n22532;
  wire u2__abc_44228_n22533;
  wire u2__abc_44228_n22534;
  wire u2__abc_44228_n22535;
  wire u2__abc_44228_n22536;
  wire u2__abc_44228_n22537;
  wire u2__abc_44228_n22539;
  wire u2__abc_44228_n22540;
  wire u2__abc_44228_n22541;
  wire u2__abc_44228_n22542;
  wire u2__abc_44228_n22543;
  wire u2__abc_44228_n22544;
  wire u2__abc_44228_n22545;
  wire u2__abc_44228_n22546;
  wire u2__abc_44228_n22547;
  wire u2__abc_44228_n22548;
  wire u2__abc_44228_n22549;
  wire u2__abc_44228_n22551;
  wire u2__abc_44228_n22552;
  wire u2__abc_44228_n22553;
  wire u2__abc_44228_n22554;
  wire u2__abc_44228_n22555;
  wire u2__abc_44228_n22556;
  wire u2__abc_44228_n22557;
  wire u2__abc_44228_n22558;
  wire u2__abc_44228_n22559;
  wire u2__abc_44228_n22560;
  wire u2__abc_44228_n22561;
  wire u2__abc_44228_n22563;
  wire u2__abc_44228_n22564;
  wire u2__abc_44228_n22565;
  wire u2__abc_44228_n22566;
  wire u2__abc_44228_n22567;
  wire u2__abc_44228_n22568;
  wire u2__abc_44228_n22569;
  wire u2__abc_44228_n22570;
  wire u2__abc_44228_n22571;
  wire u2__abc_44228_n22572;
  wire u2__abc_44228_n22573;
  wire u2__abc_44228_n22575;
  wire u2__abc_44228_n22576;
  wire u2__abc_44228_n22577;
  wire u2__abc_44228_n22578;
  wire u2__abc_44228_n22579;
  wire u2__abc_44228_n22580;
  wire u2__abc_44228_n22581;
  wire u2__abc_44228_n22582;
  wire u2__abc_44228_n22583;
  wire u2__abc_44228_n22584;
  wire u2__abc_44228_n22585;
  wire u2__abc_44228_n22587;
  wire u2__abc_44228_n22588;
  wire u2__abc_44228_n22589;
  wire u2__abc_44228_n22590;
  wire u2__abc_44228_n22591;
  wire u2__abc_44228_n22592;
  wire u2__abc_44228_n22593;
  wire u2__abc_44228_n22594;
  wire u2__abc_44228_n22595;
  wire u2__abc_44228_n22596;
  wire u2__abc_44228_n22597;
  wire u2__abc_44228_n22599;
  wire u2__abc_44228_n22600;
  wire u2__abc_44228_n22601;
  wire u2__abc_44228_n22602;
  wire u2__abc_44228_n22603;
  wire u2__abc_44228_n22604;
  wire u2__abc_44228_n22605;
  wire u2__abc_44228_n22606;
  wire u2__abc_44228_n22607;
  wire u2__abc_44228_n22608;
  wire u2__abc_44228_n22609;
  wire u2__abc_44228_n22611;
  wire u2__abc_44228_n22612;
  wire u2__abc_44228_n22613;
  wire u2__abc_44228_n22614;
  wire u2__abc_44228_n22615;
  wire u2__abc_44228_n22616;
  wire u2__abc_44228_n22617;
  wire u2__abc_44228_n22618;
  wire u2__abc_44228_n22619;
  wire u2__abc_44228_n22620;
  wire u2__abc_44228_n22621;
  wire u2__abc_44228_n22623;
  wire u2__abc_44228_n22624;
  wire u2__abc_44228_n22625;
  wire u2__abc_44228_n22626;
  wire u2__abc_44228_n22627;
  wire u2__abc_44228_n22628;
  wire u2__abc_44228_n22629;
  wire u2__abc_44228_n22630;
  wire u2__abc_44228_n22631;
  wire u2__abc_44228_n22632;
  wire u2__abc_44228_n22633;
  wire u2__abc_44228_n22635;
  wire u2__abc_44228_n22636;
  wire u2__abc_44228_n22637;
  wire u2__abc_44228_n22638;
  wire u2__abc_44228_n22639;
  wire u2__abc_44228_n22640;
  wire u2__abc_44228_n22641;
  wire u2__abc_44228_n22642;
  wire u2__abc_44228_n22643;
  wire u2__abc_44228_n22644;
  wire u2__abc_44228_n22645;
  wire u2__abc_44228_n22647;
  wire u2__abc_44228_n22648;
  wire u2__abc_44228_n22649;
  wire u2__abc_44228_n22650;
  wire u2__abc_44228_n22651;
  wire u2__abc_44228_n22652;
  wire u2__abc_44228_n22653;
  wire u2__abc_44228_n22654;
  wire u2__abc_44228_n22655;
  wire u2__abc_44228_n22656;
  wire u2__abc_44228_n22657;
  wire u2__abc_44228_n22659;
  wire u2__abc_44228_n22660;
  wire u2__abc_44228_n22661;
  wire u2__abc_44228_n22662;
  wire u2__abc_44228_n22663;
  wire u2__abc_44228_n22664;
  wire u2__abc_44228_n22665;
  wire u2__abc_44228_n22666;
  wire u2__abc_44228_n22667;
  wire u2__abc_44228_n22668;
  wire u2__abc_44228_n22669;
  wire u2__abc_44228_n22671;
  wire u2__abc_44228_n22672;
  wire u2__abc_44228_n22673;
  wire u2__abc_44228_n22674;
  wire u2__abc_44228_n22675;
  wire u2__abc_44228_n22676;
  wire u2__abc_44228_n22677;
  wire u2__abc_44228_n22678;
  wire u2__abc_44228_n22679;
  wire u2__abc_44228_n22680;
  wire u2__abc_44228_n22681;
  wire u2__abc_44228_n22683;
  wire u2__abc_44228_n22684;
  wire u2__abc_44228_n22685;
  wire u2__abc_44228_n22686;
  wire u2__abc_44228_n22687;
  wire u2__abc_44228_n22688;
  wire u2__abc_44228_n22689;
  wire u2__abc_44228_n22690;
  wire u2__abc_44228_n22691;
  wire u2__abc_44228_n22692;
  wire u2__abc_44228_n22693;
  wire u2__abc_44228_n22695;
  wire u2__abc_44228_n22696;
  wire u2__abc_44228_n22697;
  wire u2__abc_44228_n22698;
  wire u2__abc_44228_n22699;
  wire u2__abc_44228_n22700;
  wire u2__abc_44228_n22701;
  wire u2__abc_44228_n22702;
  wire u2__abc_44228_n22703;
  wire u2__abc_44228_n22704;
  wire u2__abc_44228_n22705;
  wire u2__abc_44228_n22707;
  wire u2__abc_44228_n22708;
  wire u2__abc_44228_n22709;
  wire u2__abc_44228_n22710;
  wire u2__abc_44228_n22711;
  wire u2__abc_44228_n22712;
  wire u2__abc_44228_n22713;
  wire u2__abc_44228_n22714;
  wire u2__abc_44228_n22715;
  wire u2__abc_44228_n22716;
  wire u2__abc_44228_n22717;
  wire u2__abc_44228_n22719;
  wire u2__abc_44228_n22720;
  wire u2__abc_44228_n22721;
  wire u2__abc_44228_n22722;
  wire u2__abc_44228_n22723;
  wire u2__abc_44228_n22724;
  wire u2__abc_44228_n22725;
  wire u2__abc_44228_n22726;
  wire u2__abc_44228_n22727;
  wire u2__abc_44228_n22728;
  wire u2__abc_44228_n22729;
  wire u2__abc_44228_n22731;
  wire u2__abc_44228_n22732;
  wire u2__abc_44228_n22733;
  wire u2__abc_44228_n22734;
  wire u2__abc_44228_n22735;
  wire u2__abc_44228_n22736;
  wire u2__abc_44228_n22737;
  wire u2__abc_44228_n22738;
  wire u2__abc_44228_n22739;
  wire u2__abc_44228_n22740;
  wire u2__abc_44228_n22741;
  wire u2__abc_44228_n22743;
  wire u2__abc_44228_n22744;
  wire u2__abc_44228_n22745;
  wire u2__abc_44228_n22746;
  wire u2__abc_44228_n22747;
  wire u2__abc_44228_n22748;
  wire u2__abc_44228_n22749;
  wire u2__abc_44228_n22750;
  wire u2__abc_44228_n22751;
  wire u2__abc_44228_n22752;
  wire u2__abc_44228_n22753;
  wire u2__abc_44228_n22755;
  wire u2__abc_44228_n22756;
  wire u2__abc_44228_n22757;
  wire u2__abc_44228_n22758;
  wire u2__abc_44228_n22759;
  wire u2__abc_44228_n22760;
  wire u2__abc_44228_n22761;
  wire u2__abc_44228_n22762;
  wire u2__abc_44228_n22763;
  wire u2__abc_44228_n22764;
  wire u2__abc_44228_n22765;
  wire u2__abc_44228_n22767;
  wire u2__abc_44228_n22768;
  wire u2__abc_44228_n22769;
  wire u2__abc_44228_n22770;
  wire u2__abc_44228_n22771;
  wire u2__abc_44228_n22772;
  wire u2__abc_44228_n22773;
  wire u2__abc_44228_n22774;
  wire u2__abc_44228_n22775;
  wire u2__abc_44228_n22776;
  wire u2__abc_44228_n22777;
  wire u2__abc_44228_n22779;
  wire u2__abc_44228_n22780;
  wire u2__abc_44228_n22781;
  wire u2__abc_44228_n22782;
  wire u2__abc_44228_n22783;
  wire u2__abc_44228_n22784;
  wire u2__abc_44228_n22785;
  wire u2__abc_44228_n22786;
  wire u2__abc_44228_n22787;
  wire u2__abc_44228_n22788;
  wire u2__abc_44228_n22789;
  wire u2__abc_44228_n22791;
  wire u2__abc_44228_n22792;
  wire u2__abc_44228_n22793;
  wire u2__abc_44228_n22794;
  wire u2__abc_44228_n22795;
  wire u2__abc_44228_n22796;
  wire u2__abc_44228_n22797;
  wire u2__abc_44228_n22798;
  wire u2__abc_44228_n22799;
  wire u2__abc_44228_n22800;
  wire u2__abc_44228_n22801;
  wire u2__abc_44228_n22803;
  wire u2__abc_44228_n22804;
  wire u2__abc_44228_n22805;
  wire u2__abc_44228_n22806;
  wire u2__abc_44228_n22807;
  wire u2__abc_44228_n22808;
  wire u2__abc_44228_n22809;
  wire u2__abc_44228_n22810;
  wire u2__abc_44228_n22811;
  wire u2__abc_44228_n22812;
  wire u2__abc_44228_n22813;
  wire u2__abc_44228_n22815;
  wire u2__abc_44228_n22816;
  wire u2__abc_44228_n22817;
  wire u2__abc_44228_n22818;
  wire u2__abc_44228_n22819;
  wire u2__abc_44228_n22820;
  wire u2__abc_44228_n22821;
  wire u2__abc_44228_n22822;
  wire u2__abc_44228_n22823;
  wire u2__abc_44228_n22824;
  wire u2__abc_44228_n22825;
  wire u2__abc_44228_n22827;
  wire u2__abc_44228_n22828;
  wire u2__abc_44228_n22829;
  wire u2__abc_44228_n22830;
  wire u2__abc_44228_n22831;
  wire u2__abc_44228_n22832;
  wire u2__abc_44228_n22833;
  wire u2__abc_44228_n22834;
  wire u2__abc_44228_n22835;
  wire u2__abc_44228_n22836;
  wire u2__abc_44228_n22837;
  wire u2__abc_44228_n22839;
  wire u2__abc_44228_n22840;
  wire u2__abc_44228_n22841;
  wire u2__abc_44228_n22842;
  wire u2__abc_44228_n22843;
  wire u2__abc_44228_n22844;
  wire u2__abc_44228_n22845;
  wire u2__abc_44228_n22846;
  wire u2__abc_44228_n22847;
  wire u2__abc_44228_n22848;
  wire u2__abc_44228_n22849;
  wire u2__abc_44228_n22851;
  wire u2__abc_44228_n22852;
  wire u2__abc_44228_n22853;
  wire u2__abc_44228_n22854;
  wire u2__abc_44228_n22855;
  wire u2__abc_44228_n22856;
  wire u2__abc_44228_n22857;
  wire u2__abc_44228_n22858;
  wire u2__abc_44228_n22859;
  wire u2__abc_44228_n22860;
  wire u2__abc_44228_n22861;
  wire u2__abc_44228_n22863;
  wire u2__abc_44228_n22864;
  wire u2__abc_44228_n22865;
  wire u2__abc_44228_n22866;
  wire u2__abc_44228_n22867;
  wire u2__abc_44228_n22868;
  wire u2__abc_44228_n22869;
  wire u2__abc_44228_n22870;
  wire u2__abc_44228_n22871;
  wire u2__abc_44228_n22872;
  wire u2__abc_44228_n22873;
  wire u2__abc_44228_n22875;
  wire u2__abc_44228_n22876;
  wire u2__abc_44228_n22877;
  wire u2__abc_44228_n22878;
  wire u2__abc_44228_n22879;
  wire u2__abc_44228_n22880;
  wire u2__abc_44228_n22881;
  wire u2__abc_44228_n22882;
  wire u2__abc_44228_n22883;
  wire u2__abc_44228_n22884;
  wire u2__abc_44228_n22885;
  wire u2__abc_44228_n22887;
  wire u2__abc_44228_n22888;
  wire u2__abc_44228_n22889;
  wire u2__abc_44228_n22890;
  wire u2__abc_44228_n22891;
  wire u2__abc_44228_n22892;
  wire u2__abc_44228_n22893;
  wire u2__abc_44228_n22894;
  wire u2__abc_44228_n22895;
  wire u2__abc_44228_n22896;
  wire u2__abc_44228_n22897;
  wire u2__abc_44228_n22899;
  wire u2__abc_44228_n22900;
  wire u2__abc_44228_n22901;
  wire u2__abc_44228_n22902;
  wire u2__abc_44228_n22903;
  wire u2__abc_44228_n22904;
  wire u2__abc_44228_n22905;
  wire u2__abc_44228_n22906;
  wire u2__abc_44228_n22907;
  wire u2__abc_44228_n22908;
  wire u2__abc_44228_n22909;
  wire u2__abc_44228_n22911;
  wire u2__abc_44228_n22912;
  wire u2__abc_44228_n22913;
  wire u2__abc_44228_n22914;
  wire u2__abc_44228_n22915;
  wire u2__abc_44228_n22916;
  wire u2__abc_44228_n22917;
  wire u2__abc_44228_n22918;
  wire u2__abc_44228_n22919;
  wire u2__abc_44228_n22920;
  wire u2__abc_44228_n22921;
  wire u2__abc_44228_n22923;
  wire u2__abc_44228_n22924;
  wire u2__abc_44228_n22925;
  wire u2__abc_44228_n22926;
  wire u2__abc_44228_n22927;
  wire u2__abc_44228_n22928;
  wire u2__abc_44228_n22929;
  wire u2__abc_44228_n22930;
  wire u2__abc_44228_n22931;
  wire u2__abc_44228_n22932;
  wire u2__abc_44228_n22933;
  wire u2__abc_44228_n22935;
  wire u2__abc_44228_n22936;
  wire u2__abc_44228_n22937;
  wire u2__abc_44228_n22938;
  wire u2__abc_44228_n22939;
  wire u2__abc_44228_n22940;
  wire u2__abc_44228_n22941;
  wire u2__abc_44228_n22942;
  wire u2__abc_44228_n22943;
  wire u2__abc_44228_n22944;
  wire u2__abc_44228_n22945;
  wire u2__abc_44228_n22947;
  wire u2__abc_44228_n22948;
  wire u2__abc_44228_n22949;
  wire u2__abc_44228_n22950;
  wire u2__abc_44228_n22951;
  wire u2__abc_44228_n22952;
  wire u2__abc_44228_n22953;
  wire u2__abc_44228_n22954;
  wire u2__abc_44228_n22955;
  wire u2__abc_44228_n22956;
  wire u2__abc_44228_n22957;
  wire u2__abc_44228_n22959;
  wire u2__abc_44228_n22960;
  wire u2__abc_44228_n22961;
  wire u2__abc_44228_n22962;
  wire u2__abc_44228_n22963;
  wire u2__abc_44228_n22964;
  wire u2__abc_44228_n22965;
  wire u2__abc_44228_n22966;
  wire u2__abc_44228_n22967;
  wire u2__abc_44228_n22968;
  wire u2__abc_44228_n22969;
  wire u2__abc_44228_n22971;
  wire u2__abc_44228_n22972;
  wire u2__abc_44228_n22973;
  wire u2__abc_44228_n22974;
  wire u2__abc_44228_n22975;
  wire u2__abc_44228_n22976;
  wire u2__abc_44228_n22977;
  wire u2__abc_44228_n22978;
  wire u2__abc_44228_n22979;
  wire u2__abc_44228_n22980;
  wire u2__abc_44228_n22981;
  wire u2__abc_44228_n22983;
  wire u2__abc_44228_n22984;
  wire u2__abc_44228_n22985;
  wire u2__abc_44228_n22986;
  wire u2__abc_44228_n22987;
  wire u2__abc_44228_n22988;
  wire u2__abc_44228_n22989;
  wire u2__abc_44228_n22990;
  wire u2__abc_44228_n22991;
  wire u2__abc_44228_n22992;
  wire u2__abc_44228_n22993;
  wire u2__abc_44228_n22995;
  wire u2__abc_44228_n22996;
  wire u2__abc_44228_n22997;
  wire u2__abc_44228_n22998;
  wire u2__abc_44228_n22999;
  wire u2__abc_44228_n23000;
  wire u2__abc_44228_n23001;
  wire u2__abc_44228_n23002;
  wire u2__abc_44228_n23003;
  wire u2__abc_44228_n23004;
  wire u2__abc_44228_n23005;
  wire u2__abc_44228_n23007;
  wire u2__abc_44228_n23008;
  wire u2__abc_44228_n23009;
  wire u2__abc_44228_n23010;
  wire u2__abc_44228_n23011;
  wire u2__abc_44228_n23012;
  wire u2__abc_44228_n23013;
  wire u2__abc_44228_n23014;
  wire u2__abc_44228_n23015;
  wire u2__abc_44228_n23016;
  wire u2__abc_44228_n23017;
  wire u2__abc_44228_n23019;
  wire u2__abc_44228_n23020;
  wire u2__abc_44228_n23021;
  wire u2__abc_44228_n23022;
  wire u2__abc_44228_n23023;
  wire u2__abc_44228_n23024;
  wire u2__abc_44228_n23025;
  wire u2__abc_44228_n23026;
  wire u2__abc_44228_n23027;
  wire u2__abc_44228_n23028;
  wire u2__abc_44228_n23029;
  wire u2__abc_44228_n23031;
  wire u2__abc_44228_n23032;
  wire u2__abc_44228_n23033;
  wire u2__abc_44228_n23034;
  wire u2__abc_44228_n23035;
  wire u2__abc_44228_n23036;
  wire u2__abc_44228_n23037;
  wire u2__abc_44228_n23038;
  wire u2__abc_44228_n23039;
  wire u2__abc_44228_n23040;
  wire u2__abc_44228_n23041;
  wire u2__abc_44228_n23043;
  wire u2__abc_44228_n23044;
  wire u2__abc_44228_n23045;
  wire u2__abc_44228_n23046;
  wire u2__abc_44228_n23047;
  wire u2__abc_44228_n23048;
  wire u2__abc_44228_n23049;
  wire u2__abc_44228_n23050;
  wire u2__abc_44228_n23051;
  wire u2__abc_44228_n23052;
  wire u2__abc_44228_n23053;
  wire u2__abc_44228_n23055;
  wire u2__abc_44228_n23056;
  wire u2__abc_44228_n23057;
  wire u2__abc_44228_n23058;
  wire u2__abc_44228_n23059;
  wire u2__abc_44228_n23060;
  wire u2__abc_44228_n23061;
  wire u2__abc_44228_n23062;
  wire u2__abc_44228_n23063;
  wire u2__abc_44228_n23064;
  wire u2__abc_44228_n23065;
  wire u2__abc_44228_n23067;
  wire u2__abc_44228_n23068;
  wire u2__abc_44228_n23069;
  wire u2__abc_44228_n23070;
  wire u2__abc_44228_n23071;
  wire u2__abc_44228_n23072;
  wire u2__abc_44228_n23073;
  wire u2__abc_44228_n23074;
  wire u2__abc_44228_n23075;
  wire u2__abc_44228_n23076;
  wire u2__abc_44228_n23077;
  wire u2__abc_44228_n23079;
  wire u2__abc_44228_n23080;
  wire u2__abc_44228_n23081;
  wire u2__abc_44228_n23082;
  wire u2__abc_44228_n23083;
  wire u2__abc_44228_n23084;
  wire u2__abc_44228_n23085;
  wire u2__abc_44228_n23086;
  wire u2__abc_44228_n23087;
  wire u2__abc_44228_n23088;
  wire u2__abc_44228_n23089;
  wire u2__abc_44228_n23091;
  wire u2__abc_44228_n23092;
  wire u2__abc_44228_n23093;
  wire u2__abc_44228_n23094;
  wire u2__abc_44228_n23095;
  wire u2__abc_44228_n23096;
  wire u2__abc_44228_n23097;
  wire u2__abc_44228_n23098;
  wire u2__abc_44228_n23099;
  wire u2__abc_44228_n23100;
  wire u2__abc_44228_n23101;
  wire u2__abc_44228_n23103;
  wire u2__abc_44228_n23104;
  wire u2__abc_44228_n23105;
  wire u2__abc_44228_n23106;
  wire u2__abc_44228_n23107;
  wire u2__abc_44228_n23108;
  wire u2__abc_44228_n23109;
  wire u2__abc_44228_n23110;
  wire u2__abc_44228_n23111;
  wire u2__abc_44228_n23112;
  wire u2__abc_44228_n23113;
  wire u2__abc_44228_n23115;
  wire u2__abc_44228_n23116;
  wire u2__abc_44228_n23117;
  wire u2__abc_44228_n23118;
  wire u2__abc_44228_n23119;
  wire u2__abc_44228_n23120;
  wire u2__abc_44228_n23121;
  wire u2__abc_44228_n23122;
  wire u2__abc_44228_n23123;
  wire u2__abc_44228_n23124;
  wire u2__abc_44228_n23125;
  wire u2__abc_44228_n23127;
  wire u2__abc_44228_n23128;
  wire u2__abc_44228_n23129;
  wire u2__abc_44228_n23130;
  wire u2__abc_44228_n23131;
  wire u2__abc_44228_n23132;
  wire u2__abc_44228_n23133;
  wire u2__abc_44228_n23134;
  wire u2__abc_44228_n23135;
  wire u2__abc_44228_n23136;
  wire u2__abc_44228_n23137;
  wire u2__abc_44228_n23139;
  wire u2__abc_44228_n23140;
  wire u2__abc_44228_n23141;
  wire u2__abc_44228_n23142;
  wire u2__abc_44228_n23143;
  wire u2__abc_44228_n23144;
  wire u2__abc_44228_n23145;
  wire u2__abc_44228_n23146;
  wire u2__abc_44228_n23147;
  wire u2__abc_44228_n23148;
  wire u2__abc_44228_n23149;
  wire u2__abc_44228_n23151;
  wire u2__abc_44228_n23152;
  wire u2__abc_44228_n23153;
  wire u2__abc_44228_n23154;
  wire u2__abc_44228_n23155;
  wire u2__abc_44228_n23156;
  wire u2__abc_44228_n23157;
  wire u2__abc_44228_n23158;
  wire u2__abc_44228_n23159;
  wire u2__abc_44228_n23160;
  wire u2__abc_44228_n23161;
  wire u2__abc_44228_n23163;
  wire u2__abc_44228_n23164;
  wire u2__abc_44228_n23165;
  wire u2__abc_44228_n23166;
  wire u2__abc_44228_n23167;
  wire u2__abc_44228_n23168;
  wire u2__abc_44228_n23169;
  wire u2__abc_44228_n23170;
  wire u2__abc_44228_n23171;
  wire u2__abc_44228_n23172;
  wire u2__abc_44228_n23173;
  wire u2__abc_44228_n2962;
  wire u2__abc_44228_n2963;
  wire u2__abc_44228_n2964;
  wire u2__abc_44228_n2965;
  wire u2__abc_44228_n2966;
  wire u2__abc_44228_n2966_bF_buf0;
  wire u2__abc_44228_n2966_bF_buf1;
  wire u2__abc_44228_n2966_bF_buf10;
  wire u2__abc_44228_n2966_bF_buf100;
  wire u2__abc_44228_n2966_bF_buf101;
  wire u2__abc_44228_n2966_bF_buf102;
  wire u2__abc_44228_n2966_bF_buf103;
  wire u2__abc_44228_n2966_bF_buf104;
  wire u2__abc_44228_n2966_bF_buf105;
  wire u2__abc_44228_n2966_bF_buf106;
  wire u2__abc_44228_n2966_bF_buf107;
  wire u2__abc_44228_n2966_bF_buf11;
  wire u2__abc_44228_n2966_bF_buf12;
  wire u2__abc_44228_n2966_bF_buf13;
  wire u2__abc_44228_n2966_bF_buf14;
  wire u2__abc_44228_n2966_bF_buf15;
  wire u2__abc_44228_n2966_bF_buf16;
  wire u2__abc_44228_n2966_bF_buf17;
  wire u2__abc_44228_n2966_bF_buf18;
  wire u2__abc_44228_n2966_bF_buf19;
  wire u2__abc_44228_n2966_bF_buf2;
  wire u2__abc_44228_n2966_bF_buf20;
  wire u2__abc_44228_n2966_bF_buf21;
  wire u2__abc_44228_n2966_bF_buf22;
  wire u2__abc_44228_n2966_bF_buf23;
  wire u2__abc_44228_n2966_bF_buf24;
  wire u2__abc_44228_n2966_bF_buf25;
  wire u2__abc_44228_n2966_bF_buf26;
  wire u2__abc_44228_n2966_bF_buf27;
  wire u2__abc_44228_n2966_bF_buf28;
  wire u2__abc_44228_n2966_bF_buf29;
  wire u2__abc_44228_n2966_bF_buf3;
  wire u2__abc_44228_n2966_bF_buf30;
  wire u2__abc_44228_n2966_bF_buf31;
  wire u2__abc_44228_n2966_bF_buf32;
  wire u2__abc_44228_n2966_bF_buf33;
  wire u2__abc_44228_n2966_bF_buf34;
  wire u2__abc_44228_n2966_bF_buf35;
  wire u2__abc_44228_n2966_bF_buf36;
  wire u2__abc_44228_n2966_bF_buf37;
  wire u2__abc_44228_n2966_bF_buf38;
  wire u2__abc_44228_n2966_bF_buf39;
  wire u2__abc_44228_n2966_bF_buf4;
  wire u2__abc_44228_n2966_bF_buf40;
  wire u2__abc_44228_n2966_bF_buf41;
  wire u2__abc_44228_n2966_bF_buf42;
  wire u2__abc_44228_n2966_bF_buf43;
  wire u2__abc_44228_n2966_bF_buf44;
  wire u2__abc_44228_n2966_bF_buf45;
  wire u2__abc_44228_n2966_bF_buf46;
  wire u2__abc_44228_n2966_bF_buf47;
  wire u2__abc_44228_n2966_bF_buf48;
  wire u2__abc_44228_n2966_bF_buf49;
  wire u2__abc_44228_n2966_bF_buf5;
  wire u2__abc_44228_n2966_bF_buf50;
  wire u2__abc_44228_n2966_bF_buf51;
  wire u2__abc_44228_n2966_bF_buf52;
  wire u2__abc_44228_n2966_bF_buf53;
  wire u2__abc_44228_n2966_bF_buf54;
  wire u2__abc_44228_n2966_bF_buf55;
  wire u2__abc_44228_n2966_bF_buf56;
  wire u2__abc_44228_n2966_bF_buf57;
  wire u2__abc_44228_n2966_bF_buf58;
  wire u2__abc_44228_n2966_bF_buf59;
  wire u2__abc_44228_n2966_bF_buf6;
  wire u2__abc_44228_n2966_bF_buf60;
  wire u2__abc_44228_n2966_bF_buf61;
  wire u2__abc_44228_n2966_bF_buf62;
  wire u2__abc_44228_n2966_bF_buf63;
  wire u2__abc_44228_n2966_bF_buf64;
  wire u2__abc_44228_n2966_bF_buf65;
  wire u2__abc_44228_n2966_bF_buf66;
  wire u2__abc_44228_n2966_bF_buf67;
  wire u2__abc_44228_n2966_bF_buf68;
  wire u2__abc_44228_n2966_bF_buf69;
  wire u2__abc_44228_n2966_bF_buf7;
  wire u2__abc_44228_n2966_bF_buf70;
  wire u2__abc_44228_n2966_bF_buf71;
  wire u2__abc_44228_n2966_bF_buf72;
  wire u2__abc_44228_n2966_bF_buf73;
  wire u2__abc_44228_n2966_bF_buf74;
  wire u2__abc_44228_n2966_bF_buf75;
  wire u2__abc_44228_n2966_bF_buf76;
  wire u2__abc_44228_n2966_bF_buf77;
  wire u2__abc_44228_n2966_bF_buf78;
  wire u2__abc_44228_n2966_bF_buf79;
  wire u2__abc_44228_n2966_bF_buf8;
  wire u2__abc_44228_n2966_bF_buf80;
  wire u2__abc_44228_n2966_bF_buf81;
  wire u2__abc_44228_n2966_bF_buf82;
  wire u2__abc_44228_n2966_bF_buf83;
  wire u2__abc_44228_n2966_bF_buf84;
  wire u2__abc_44228_n2966_bF_buf85;
  wire u2__abc_44228_n2966_bF_buf86;
  wire u2__abc_44228_n2966_bF_buf87;
  wire u2__abc_44228_n2966_bF_buf88;
  wire u2__abc_44228_n2966_bF_buf89;
  wire u2__abc_44228_n2966_bF_buf9;
  wire u2__abc_44228_n2966_bF_buf90;
  wire u2__abc_44228_n2966_bF_buf91;
  wire u2__abc_44228_n2966_bF_buf92;
  wire u2__abc_44228_n2966_bF_buf93;
  wire u2__abc_44228_n2966_bF_buf94;
  wire u2__abc_44228_n2966_bF_buf95;
  wire u2__abc_44228_n2966_bF_buf96;
  wire u2__abc_44228_n2966_bF_buf97;
  wire u2__abc_44228_n2966_bF_buf98;
  wire u2__abc_44228_n2966_bF_buf99;
  wire u2__abc_44228_n2966_hier0_bF_buf0;
  wire u2__abc_44228_n2966_hier0_bF_buf1;
  wire u2__abc_44228_n2966_hier0_bF_buf2;
  wire u2__abc_44228_n2966_hier0_bF_buf3;
  wire u2__abc_44228_n2966_hier0_bF_buf4;
  wire u2__abc_44228_n2966_hier0_bF_buf5;
  wire u2__abc_44228_n2966_hier0_bF_buf6;
  wire u2__abc_44228_n2966_hier0_bF_buf7;
  wire u2__abc_44228_n2966_hier0_bF_buf8;
  wire u2__abc_44228_n2966_hier0_bF_buf9;
  wire u2__abc_44228_n2967;
  wire u2__abc_44228_n2968;
  wire u2__abc_44228_n2969;
  wire u2__abc_44228_n2970;
  wire u2__abc_44228_n2972;
  wire u2__abc_44228_n2972_bF_buf0;
  wire u2__abc_44228_n2972_bF_buf1;
  wire u2__abc_44228_n2972_bF_buf10;
  wire u2__abc_44228_n2972_bF_buf100;
  wire u2__abc_44228_n2972_bF_buf101;
  wire u2__abc_44228_n2972_bF_buf102;
  wire u2__abc_44228_n2972_bF_buf103;
  wire u2__abc_44228_n2972_bF_buf104;
  wire u2__abc_44228_n2972_bF_buf105;
  wire u2__abc_44228_n2972_bF_buf106;
  wire u2__abc_44228_n2972_bF_buf107;
  wire u2__abc_44228_n2972_bF_buf11;
  wire u2__abc_44228_n2972_bF_buf12;
  wire u2__abc_44228_n2972_bF_buf13;
  wire u2__abc_44228_n2972_bF_buf14;
  wire u2__abc_44228_n2972_bF_buf15;
  wire u2__abc_44228_n2972_bF_buf16;
  wire u2__abc_44228_n2972_bF_buf17;
  wire u2__abc_44228_n2972_bF_buf18;
  wire u2__abc_44228_n2972_bF_buf19;
  wire u2__abc_44228_n2972_bF_buf2;
  wire u2__abc_44228_n2972_bF_buf20;
  wire u2__abc_44228_n2972_bF_buf21;
  wire u2__abc_44228_n2972_bF_buf22;
  wire u2__abc_44228_n2972_bF_buf23;
  wire u2__abc_44228_n2972_bF_buf24;
  wire u2__abc_44228_n2972_bF_buf25;
  wire u2__abc_44228_n2972_bF_buf26;
  wire u2__abc_44228_n2972_bF_buf27;
  wire u2__abc_44228_n2972_bF_buf28;
  wire u2__abc_44228_n2972_bF_buf29;
  wire u2__abc_44228_n2972_bF_buf3;
  wire u2__abc_44228_n2972_bF_buf30;
  wire u2__abc_44228_n2972_bF_buf31;
  wire u2__abc_44228_n2972_bF_buf32;
  wire u2__abc_44228_n2972_bF_buf33;
  wire u2__abc_44228_n2972_bF_buf34;
  wire u2__abc_44228_n2972_bF_buf35;
  wire u2__abc_44228_n2972_bF_buf36;
  wire u2__abc_44228_n2972_bF_buf37;
  wire u2__abc_44228_n2972_bF_buf38;
  wire u2__abc_44228_n2972_bF_buf39;
  wire u2__abc_44228_n2972_bF_buf4;
  wire u2__abc_44228_n2972_bF_buf40;
  wire u2__abc_44228_n2972_bF_buf41;
  wire u2__abc_44228_n2972_bF_buf42;
  wire u2__abc_44228_n2972_bF_buf43;
  wire u2__abc_44228_n2972_bF_buf44;
  wire u2__abc_44228_n2972_bF_buf45;
  wire u2__abc_44228_n2972_bF_buf46;
  wire u2__abc_44228_n2972_bF_buf47;
  wire u2__abc_44228_n2972_bF_buf48;
  wire u2__abc_44228_n2972_bF_buf49;
  wire u2__abc_44228_n2972_bF_buf5;
  wire u2__abc_44228_n2972_bF_buf50;
  wire u2__abc_44228_n2972_bF_buf51;
  wire u2__abc_44228_n2972_bF_buf52;
  wire u2__abc_44228_n2972_bF_buf53;
  wire u2__abc_44228_n2972_bF_buf54;
  wire u2__abc_44228_n2972_bF_buf55;
  wire u2__abc_44228_n2972_bF_buf56;
  wire u2__abc_44228_n2972_bF_buf57;
  wire u2__abc_44228_n2972_bF_buf58;
  wire u2__abc_44228_n2972_bF_buf59;
  wire u2__abc_44228_n2972_bF_buf6;
  wire u2__abc_44228_n2972_bF_buf60;
  wire u2__abc_44228_n2972_bF_buf61;
  wire u2__abc_44228_n2972_bF_buf62;
  wire u2__abc_44228_n2972_bF_buf63;
  wire u2__abc_44228_n2972_bF_buf64;
  wire u2__abc_44228_n2972_bF_buf65;
  wire u2__abc_44228_n2972_bF_buf66;
  wire u2__abc_44228_n2972_bF_buf67;
  wire u2__abc_44228_n2972_bF_buf68;
  wire u2__abc_44228_n2972_bF_buf69;
  wire u2__abc_44228_n2972_bF_buf7;
  wire u2__abc_44228_n2972_bF_buf70;
  wire u2__abc_44228_n2972_bF_buf71;
  wire u2__abc_44228_n2972_bF_buf72;
  wire u2__abc_44228_n2972_bF_buf73;
  wire u2__abc_44228_n2972_bF_buf74;
  wire u2__abc_44228_n2972_bF_buf75;
  wire u2__abc_44228_n2972_bF_buf76;
  wire u2__abc_44228_n2972_bF_buf77;
  wire u2__abc_44228_n2972_bF_buf78;
  wire u2__abc_44228_n2972_bF_buf79;
  wire u2__abc_44228_n2972_bF_buf8;
  wire u2__abc_44228_n2972_bF_buf80;
  wire u2__abc_44228_n2972_bF_buf81;
  wire u2__abc_44228_n2972_bF_buf82;
  wire u2__abc_44228_n2972_bF_buf83;
  wire u2__abc_44228_n2972_bF_buf84;
  wire u2__abc_44228_n2972_bF_buf85;
  wire u2__abc_44228_n2972_bF_buf86;
  wire u2__abc_44228_n2972_bF_buf87;
  wire u2__abc_44228_n2972_bF_buf88;
  wire u2__abc_44228_n2972_bF_buf89;
  wire u2__abc_44228_n2972_bF_buf9;
  wire u2__abc_44228_n2972_bF_buf90;
  wire u2__abc_44228_n2972_bF_buf91;
  wire u2__abc_44228_n2972_bF_buf92;
  wire u2__abc_44228_n2972_bF_buf93;
  wire u2__abc_44228_n2972_bF_buf94;
  wire u2__abc_44228_n2972_bF_buf95;
  wire u2__abc_44228_n2972_bF_buf96;
  wire u2__abc_44228_n2972_bF_buf97;
  wire u2__abc_44228_n2972_bF_buf98;
  wire u2__abc_44228_n2972_bF_buf99;
  wire u2__abc_44228_n2972_hier0_bF_buf0;
  wire u2__abc_44228_n2972_hier0_bF_buf1;
  wire u2__abc_44228_n2972_hier0_bF_buf2;
  wire u2__abc_44228_n2972_hier0_bF_buf3;
  wire u2__abc_44228_n2972_hier0_bF_buf4;
  wire u2__abc_44228_n2972_hier0_bF_buf5;
  wire u2__abc_44228_n2972_hier0_bF_buf6;
  wire u2__abc_44228_n2972_hier0_bF_buf7;
  wire u2__abc_44228_n2972_hier0_bF_buf8;
  wire u2__abc_44228_n2972_hier0_bF_buf9;
  wire u2__abc_44228_n2973;
  wire u2__abc_44228_n2974;
  wire u2__abc_44228_n2975;
  wire u2__abc_44228_n2976;
  wire u2__abc_44228_n2977;
  wire u2__abc_44228_n2978;
  wire u2__abc_44228_n2979;
  wire u2__abc_44228_n2980;
  wire u2__abc_44228_n2981;
  wire u2__abc_44228_n2982;
  wire u2__abc_44228_n2983;
  wire u2__abc_44228_n2983_bF_buf0;
  wire u2__abc_44228_n2983_bF_buf1;
  wire u2__abc_44228_n2983_bF_buf10;
  wire u2__abc_44228_n2983_bF_buf100;
  wire u2__abc_44228_n2983_bF_buf101;
  wire u2__abc_44228_n2983_bF_buf102;
  wire u2__abc_44228_n2983_bF_buf103;
  wire u2__abc_44228_n2983_bF_buf104;
  wire u2__abc_44228_n2983_bF_buf105;
  wire u2__abc_44228_n2983_bF_buf106;
  wire u2__abc_44228_n2983_bF_buf107;
  wire u2__abc_44228_n2983_bF_buf108;
  wire u2__abc_44228_n2983_bF_buf109;
  wire u2__abc_44228_n2983_bF_buf11;
  wire u2__abc_44228_n2983_bF_buf110;
  wire u2__abc_44228_n2983_bF_buf111;
  wire u2__abc_44228_n2983_bF_buf112;
  wire u2__abc_44228_n2983_bF_buf113;
  wire u2__abc_44228_n2983_bF_buf114;
  wire u2__abc_44228_n2983_bF_buf115;
  wire u2__abc_44228_n2983_bF_buf116;
  wire u2__abc_44228_n2983_bF_buf117;
  wire u2__abc_44228_n2983_bF_buf118;
  wire u2__abc_44228_n2983_bF_buf119;
  wire u2__abc_44228_n2983_bF_buf12;
  wire u2__abc_44228_n2983_bF_buf120;
  wire u2__abc_44228_n2983_bF_buf121;
  wire u2__abc_44228_n2983_bF_buf122;
  wire u2__abc_44228_n2983_bF_buf123;
  wire u2__abc_44228_n2983_bF_buf124;
  wire u2__abc_44228_n2983_bF_buf125;
  wire u2__abc_44228_n2983_bF_buf126;
  wire u2__abc_44228_n2983_bF_buf127;
  wire u2__abc_44228_n2983_bF_buf128;
  wire u2__abc_44228_n2983_bF_buf129;
  wire u2__abc_44228_n2983_bF_buf13;
  wire u2__abc_44228_n2983_bF_buf130;
  wire u2__abc_44228_n2983_bF_buf131;
  wire u2__abc_44228_n2983_bF_buf132;
  wire u2__abc_44228_n2983_bF_buf133;
  wire u2__abc_44228_n2983_bF_buf134;
  wire u2__abc_44228_n2983_bF_buf135;
  wire u2__abc_44228_n2983_bF_buf136;
  wire u2__abc_44228_n2983_bF_buf137;
  wire u2__abc_44228_n2983_bF_buf138;
  wire u2__abc_44228_n2983_bF_buf139;
  wire u2__abc_44228_n2983_bF_buf14;
  wire u2__abc_44228_n2983_bF_buf140;
  wire u2__abc_44228_n2983_bF_buf141;
  wire u2__abc_44228_n2983_bF_buf15;
  wire u2__abc_44228_n2983_bF_buf16;
  wire u2__abc_44228_n2983_bF_buf17;
  wire u2__abc_44228_n2983_bF_buf18;
  wire u2__abc_44228_n2983_bF_buf19;
  wire u2__abc_44228_n2983_bF_buf2;
  wire u2__abc_44228_n2983_bF_buf20;
  wire u2__abc_44228_n2983_bF_buf21;
  wire u2__abc_44228_n2983_bF_buf22;
  wire u2__abc_44228_n2983_bF_buf23;
  wire u2__abc_44228_n2983_bF_buf24;
  wire u2__abc_44228_n2983_bF_buf25;
  wire u2__abc_44228_n2983_bF_buf26;
  wire u2__abc_44228_n2983_bF_buf27;
  wire u2__abc_44228_n2983_bF_buf28;
  wire u2__abc_44228_n2983_bF_buf29;
  wire u2__abc_44228_n2983_bF_buf3;
  wire u2__abc_44228_n2983_bF_buf30;
  wire u2__abc_44228_n2983_bF_buf31;
  wire u2__abc_44228_n2983_bF_buf32;
  wire u2__abc_44228_n2983_bF_buf33;
  wire u2__abc_44228_n2983_bF_buf34;
  wire u2__abc_44228_n2983_bF_buf35;
  wire u2__abc_44228_n2983_bF_buf36;
  wire u2__abc_44228_n2983_bF_buf37;
  wire u2__abc_44228_n2983_bF_buf38;
  wire u2__abc_44228_n2983_bF_buf39;
  wire u2__abc_44228_n2983_bF_buf4;
  wire u2__abc_44228_n2983_bF_buf40;
  wire u2__abc_44228_n2983_bF_buf41;
  wire u2__abc_44228_n2983_bF_buf42;
  wire u2__abc_44228_n2983_bF_buf43;
  wire u2__abc_44228_n2983_bF_buf44;
  wire u2__abc_44228_n2983_bF_buf45;
  wire u2__abc_44228_n2983_bF_buf46;
  wire u2__abc_44228_n2983_bF_buf47;
  wire u2__abc_44228_n2983_bF_buf48;
  wire u2__abc_44228_n2983_bF_buf49;
  wire u2__abc_44228_n2983_bF_buf5;
  wire u2__abc_44228_n2983_bF_buf50;
  wire u2__abc_44228_n2983_bF_buf51;
  wire u2__abc_44228_n2983_bF_buf52;
  wire u2__abc_44228_n2983_bF_buf53;
  wire u2__abc_44228_n2983_bF_buf54;
  wire u2__abc_44228_n2983_bF_buf55;
  wire u2__abc_44228_n2983_bF_buf56;
  wire u2__abc_44228_n2983_bF_buf57;
  wire u2__abc_44228_n2983_bF_buf58;
  wire u2__abc_44228_n2983_bF_buf59;
  wire u2__abc_44228_n2983_bF_buf6;
  wire u2__abc_44228_n2983_bF_buf60;
  wire u2__abc_44228_n2983_bF_buf61;
  wire u2__abc_44228_n2983_bF_buf62;
  wire u2__abc_44228_n2983_bF_buf63;
  wire u2__abc_44228_n2983_bF_buf64;
  wire u2__abc_44228_n2983_bF_buf65;
  wire u2__abc_44228_n2983_bF_buf66;
  wire u2__abc_44228_n2983_bF_buf67;
  wire u2__abc_44228_n2983_bF_buf68;
  wire u2__abc_44228_n2983_bF_buf69;
  wire u2__abc_44228_n2983_bF_buf7;
  wire u2__abc_44228_n2983_bF_buf70;
  wire u2__abc_44228_n2983_bF_buf71;
  wire u2__abc_44228_n2983_bF_buf72;
  wire u2__abc_44228_n2983_bF_buf73;
  wire u2__abc_44228_n2983_bF_buf74;
  wire u2__abc_44228_n2983_bF_buf75;
  wire u2__abc_44228_n2983_bF_buf76;
  wire u2__abc_44228_n2983_bF_buf77;
  wire u2__abc_44228_n2983_bF_buf78;
  wire u2__abc_44228_n2983_bF_buf79;
  wire u2__abc_44228_n2983_bF_buf8;
  wire u2__abc_44228_n2983_bF_buf80;
  wire u2__abc_44228_n2983_bF_buf81;
  wire u2__abc_44228_n2983_bF_buf82;
  wire u2__abc_44228_n2983_bF_buf83;
  wire u2__abc_44228_n2983_bF_buf84;
  wire u2__abc_44228_n2983_bF_buf85;
  wire u2__abc_44228_n2983_bF_buf86;
  wire u2__abc_44228_n2983_bF_buf87;
  wire u2__abc_44228_n2983_bF_buf88;
  wire u2__abc_44228_n2983_bF_buf89;
  wire u2__abc_44228_n2983_bF_buf9;
  wire u2__abc_44228_n2983_bF_buf90;
  wire u2__abc_44228_n2983_bF_buf91;
  wire u2__abc_44228_n2983_bF_buf92;
  wire u2__abc_44228_n2983_bF_buf93;
  wire u2__abc_44228_n2983_bF_buf94;
  wire u2__abc_44228_n2983_bF_buf95;
  wire u2__abc_44228_n2983_bF_buf96;
  wire u2__abc_44228_n2983_bF_buf97;
  wire u2__abc_44228_n2983_bF_buf98;
  wire u2__abc_44228_n2983_bF_buf99;
  wire u2__abc_44228_n2983_hier0_bF_buf0;
  wire u2__abc_44228_n2983_hier0_bF_buf1;
  wire u2__abc_44228_n2983_hier0_bF_buf10;
  wire u2__abc_44228_n2983_hier0_bF_buf2;
  wire u2__abc_44228_n2983_hier0_bF_buf3;
  wire u2__abc_44228_n2983_hier0_bF_buf4;
  wire u2__abc_44228_n2983_hier0_bF_buf5;
  wire u2__abc_44228_n2983_hier0_bF_buf6;
  wire u2__abc_44228_n2983_hier0_bF_buf7;
  wire u2__abc_44228_n2983_hier0_bF_buf8;
  wire u2__abc_44228_n2983_hier0_bF_buf9;
  wire u2__abc_44228_n2984;
  wire u2__abc_44228_n2984_bF_buf0;
  wire u2__abc_44228_n2984_bF_buf1;
  wire u2__abc_44228_n2984_bF_buf10;
  wire u2__abc_44228_n2984_bF_buf11;
  wire u2__abc_44228_n2984_bF_buf12;
  wire u2__abc_44228_n2984_bF_buf13;
  wire u2__abc_44228_n2984_bF_buf14;
  wire u2__abc_44228_n2984_bF_buf2;
  wire u2__abc_44228_n2984_bF_buf3;
  wire u2__abc_44228_n2984_bF_buf4;
  wire u2__abc_44228_n2984_bF_buf5;
  wire u2__abc_44228_n2984_bF_buf6;
  wire u2__abc_44228_n2984_bF_buf7;
  wire u2__abc_44228_n2984_bF_buf8;
  wire u2__abc_44228_n2984_bF_buf9;
  wire u2__abc_44228_n2985;
  wire u2__abc_44228_n2986;
  wire u2__abc_44228_n2987;
  wire u2__abc_44228_n2987_bF_buf0;
  wire u2__abc_44228_n2987_bF_buf1;
  wire u2__abc_44228_n2987_bF_buf10;
  wire u2__abc_44228_n2987_bF_buf11;
  wire u2__abc_44228_n2987_bF_buf12;
  wire u2__abc_44228_n2987_bF_buf13;
  wire u2__abc_44228_n2987_bF_buf14;
  wire u2__abc_44228_n2987_bF_buf2;
  wire u2__abc_44228_n2987_bF_buf3;
  wire u2__abc_44228_n2987_bF_buf4;
  wire u2__abc_44228_n2987_bF_buf5;
  wire u2__abc_44228_n2987_bF_buf6;
  wire u2__abc_44228_n2987_bF_buf7;
  wire u2__abc_44228_n2987_bF_buf8;
  wire u2__abc_44228_n2987_bF_buf9;
  wire u2__abc_44228_n2988;
  wire u2__abc_44228_n2988_bF_buf0;
  wire u2__abc_44228_n2988_bF_buf1;
  wire u2__abc_44228_n2988_bF_buf10;
  wire u2__abc_44228_n2988_bF_buf11;
  wire u2__abc_44228_n2988_bF_buf12;
  wire u2__abc_44228_n2988_bF_buf13;
  wire u2__abc_44228_n2988_bF_buf2;
  wire u2__abc_44228_n2988_bF_buf3;
  wire u2__abc_44228_n2988_bF_buf4;
  wire u2__abc_44228_n2988_bF_buf5;
  wire u2__abc_44228_n2988_bF_buf6;
  wire u2__abc_44228_n2988_bF_buf7;
  wire u2__abc_44228_n2988_bF_buf8;
  wire u2__abc_44228_n2988_bF_buf9;
  wire u2__abc_44228_n2989;
  wire u2__abc_44228_n2989_bF_buf0;
  wire u2__abc_44228_n2989_bF_buf1;
  wire u2__abc_44228_n2989_bF_buf2;
  wire u2__abc_44228_n2989_bF_buf3;
  wire u2__abc_44228_n2990;
  wire u2__abc_44228_n2992;
  wire u2__abc_44228_n2993;
  wire u2__abc_44228_n2995;
  wire u2__abc_44228_n2996;
  wire u2__abc_44228_n2997;
  wire u2__abc_44228_n2998;
  wire u2__abc_44228_n2999;
  wire u2__abc_44228_n3001;
  wire u2__abc_44228_n3002;
  wire u2__abc_44228_n3003;
  wire u2__abc_44228_n3004;
  wire u2__abc_44228_n3005;
  wire u2__abc_44228_n3006;
  wire u2__abc_44228_n3008;
  wire u2__abc_44228_n3009;
  wire u2__abc_44228_n3010;
  wire u2__abc_44228_n3011;
  wire u2__abc_44228_n3012;
  wire u2__abc_44228_n3013;
  wire u2__abc_44228_n3014;
  wire u2__abc_44228_n3015;
  wire u2__abc_44228_n3016;
  wire u2__abc_44228_n3018;
  wire u2__abc_44228_n3019;
  wire u2__abc_44228_n3020;
  wire u2__abc_44228_n3021;
  wire u2__abc_44228_n3022;
  wire u2__abc_44228_n3023;
  wire u2__abc_44228_n3025;
  wire u2__abc_44228_n3026;
  wire u2__abc_44228_n3027;
  wire u2__abc_44228_n3028;
  wire u2__abc_44228_n3029;
  wire u2__abc_44228_n3030;
  wire u2__abc_44228_n3032;
  wire u2__abc_44228_n3033;
  wire u2__abc_44228_n3034;
  wire u2__abc_44228_n3035;
  wire u2__abc_44228_n3036;
  wire u2__abc_44228_n3037;
  wire u2__abc_44228_n3039;
  wire u2__abc_44228_n3040;
  wire u2__abc_44228_n3041;
  wire u2__abc_44228_n3042;
  wire u2__abc_44228_n3043;
  wire u2__abc_44228_n3044;
  wire u2__abc_44228_n3045;
  wire u2__abc_44228_n3047;
  wire u2__abc_44228_n3048;
  wire u2__abc_44228_n3049;
  wire u2__abc_44228_n3050;
  wire u2__abc_44228_n3051;
  wire u2__abc_44228_n3052;
  wire u2__abc_44228_n3053;
  wire u2__abc_44228_n3054;
  wire u2__abc_44228_n3055;
  wire u2__abc_44228_n3056;
  wire u2__abc_44228_n3058;
  wire u2__abc_44228_n3059;
  wire u2__abc_44228_n3060;
  wire u2__abc_44228_n3061;
  wire u2__abc_44228_n3062;
  wire u2__abc_44228_n3062_bF_buf0;
  wire u2__abc_44228_n3062_bF_buf1;
  wire u2__abc_44228_n3062_bF_buf10;
  wire u2__abc_44228_n3062_bF_buf11;
  wire u2__abc_44228_n3062_bF_buf12;
  wire u2__abc_44228_n3062_bF_buf13;
  wire u2__abc_44228_n3062_bF_buf14;
  wire u2__abc_44228_n3062_bF_buf15;
  wire u2__abc_44228_n3062_bF_buf16;
  wire u2__abc_44228_n3062_bF_buf17;
  wire u2__abc_44228_n3062_bF_buf18;
  wire u2__abc_44228_n3062_bF_buf19;
  wire u2__abc_44228_n3062_bF_buf2;
  wire u2__abc_44228_n3062_bF_buf20;
  wire u2__abc_44228_n3062_bF_buf21;
  wire u2__abc_44228_n3062_bF_buf22;
  wire u2__abc_44228_n3062_bF_buf23;
  wire u2__abc_44228_n3062_bF_buf24;
  wire u2__abc_44228_n3062_bF_buf25;
  wire u2__abc_44228_n3062_bF_buf26;
  wire u2__abc_44228_n3062_bF_buf27;
  wire u2__abc_44228_n3062_bF_buf28;
  wire u2__abc_44228_n3062_bF_buf29;
  wire u2__abc_44228_n3062_bF_buf3;
  wire u2__abc_44228_n3062_bF_buf30;
  wire u2__abc_44228_n3062_bF_buf31;
  wire u2__abc_44228_n3062_bF_buf32;
  wire u2__abc_44228_n3062_bF_buf33;
  wire u2__abc_44228_n3062_bF_buf34;
  wire u2__abc_44228_n3062_bF_buf35;
  wire u2__abc_44228_n3062_bF_buf36;
  wire u2__abc_44228_n3062_bF_buf37;
  wire u2__abc_44228_n3062_bF_buf38;
  wire u2__abc_44228_n3062_bF_buf39;
  wire u2__abc_44228_n3062_bF_buf4;
  wire u2__abc_44228_n3062_bF_buf40;
  wire u2__abc_44228_n3062_bF_buf41;
  wire u2__abc_44228_n3062_bF_buf42;
  wire u2__abc_44228_n3062_bF_buf43;
  wire u2__abc_44228_n3062_bF_buf44;
  wire u2__abc_44228_n3062_bF_buf45;
  wire u2__abc_44228_n3062_bF_buf46;
  wire u2__abc_44228_n3062_bF_buf47;
  wire u2__abc_44228_n3062_bF_buf48;
  wire u2__abc_44228_n3062_bF_buf49;
  wire u2__abc_44228_n3062_bF_buf5;
  wire u2__abc_44228_n3062_bF_buf50;
  wire u2__abc_44228_n3062_bF_buf51;
  wire u2__abc_44228_n3062_bF_buf52;
  wire u2__abc_44228_n3062_bF_buf53;
  wire u2__abc_44228_n3062_bF_buf54;
  wire u2__abc_44228_n3062_bF_buf55;
  wire u2__abc_44228_n3062_bF_buf56;
  wire u2__abc_44228_n3062_bF_buf57;
  wire u2__abc_44228_n3062_bF_buf58;
  wire u2__abc_44228_n3062_bF_buf59;
  wire u2__abc_44228_n3062_bF_buf6;
  wire u2__abc_44228_n3062_bF_buf60;
  wire u2__abc_44228_n3062_bF_buf61;
  wire u2__abc_44228_n3062_bF_buf62;
  wire u2__abc_44228_n3062_bF_buf63;
  wire u2__abc_44228_n3062_bF_buf64;
  wire u2__abc_44228_n3062_bF_buf65;
  wire u2__abc_44228_n3062_bF_buf66;
  wire u2__abc_44228_n3062_bF_buf67;
  wire u2__abc_44228_n3062_bF_buf68;
  wire u2__abc_44228_n3062_bF_buf69;
  wire u2__abc_44228_n3062_bF_buf7;
  wire u2__abc_44228_n3062_bF_buf70;
  wire u2__abc_44228_n3062_bF_buf71;
  wire u2__abc_44228_n3062_bF_buf72;
  wire u2__abc_44228_n3062_bF_buf73;
  wire u2__abc_44228_n3062_bF_buf74;
  wire u2__abc_44228_n3062_bF_buf75;
  wire u2__abc_44228_n3062_bF_buf76;
  wire u2__abc_44228_n3062_bF_buf77;
  wire u2__abc_44228_n3062_bF_buf78;
  wire u2__abc_44228_n3062_bF_buf79;
  wire u2__abc_44228_n3062_bF_buf8;
  wire u2__abc_44228_n3062_bF_buf80;
  wire u2__abc_44228_n3062_bF_buf81;
  wire u2__abc_44228_n3062_bF_buf82;
  wire u2__abc_44228_n3062_bF_buf83;
  wire u2__abc_44228_n3062_bF_buf84;
  wire u2__abc_44228_n3062_bF_buf85;
  wire u2__abc_44228_n3062_bF_buf86;
  wire u2__abc_44228_n3062_bF_buf87;
  wire u2__abc_44228_n3062_bF_buf88;
  wire u2__abc_44228_n3062_bF_buf89;
  wire u2__abc_44228_n3062_bF_buf9;
  wire u2__abc_44228_n3062_bF_buf90;
  wire u2__abc_44228_n3062_bF_buf91;
  wire u2__abc_44228_n3062_bF_buf92;
  wire u2__abc_44228_n3062_hier0_bF_buf0;
  wire u2__abc_44228_n3062_hier0_bF_buf1;
  wire u2__abc_44228_n3062_hier0_bF_buf2;
  wire u2__abc_44228_n3062_hier0_bF_buf3;
  wire u2__abc_44228_n3062_hier0_bF_buf4;
  wire u2__abc_44228_n3062_hier0_bF_buf5;
  wire u2__abc_44228_n3062_hier0_bF_buf6;
  wire u2__abc_44228_n3062_hier0_bF_buf7;
  wire u2__abc_44228_n3062_hier0_bF_buf8;
  wire u2__abc_44228_n3063;
  wire u2__abc_44228_n3064;
  wire u2__abc_44228_n3065;
  wire u2__abc_44228_n3066;
  wire u2__abc_44228_n3067;
  wire u2__abc_44228_n3068;
  wire u2__abc_44228_n3069;
  wire u2__abc_44228_n3070;
  wire u2__abc_44228_n3071;
  wire u2__abc_44228_n3072;
  wire u2__abc_44228_n3073;
  wire u2__abc_44228_n3074;
  wire u2__abc_44228_n3075;
  wire u2__abc_44228_n3076;
  wire u2__abc_44228_n3077;
  wire u2__abc_44228_n3078;
  wire u2__abc_44228_n3079;
  wire u2__abc_44228_n3080;
  wire u2__abc_44228_n3081;
  wire u2__abc_44228_n3082;
  wire u2__abc_44228_n3083;
  wire u2__abc_44228_n3084;
  wire u2__abc_44228_n3085;
  wire u2__abc_44228_n3086;
  wire u2__abc_44228_n3087;
  wire u2__abc_44228_n3088;
  wire u2__abc_44228_n3089;
  wire u2__abc_44228_n3090;
  wire u2__abc_44228_n3091;
  wire u2__abc_44228_n3092;
  wire u2__abc_44228_n3093;
  wire u2__abc_44228_n3094;
  wire u2__abc_44228_n3095;
  wire u2__abc_44228_n3096;
  wire u2__abc_44228_n3097;
  wire u2__abc_44228_n3098;
  wire u2__abc_44228_n3099;
  wire u2__abc_44228_n3100;
  wire u2__abc_44228_n3101;
  wire u2__abc_44228_n3102;
  wire u2__abc_44228_n3103;
  wire u2__abc_44228_n3104;
  wire u2__abc_44228_n3105;
  wire u2__abc_44228_n3106;
  wire u2__abc_44228_n3107;
  wire u2__abc_44228_n3108;
  wire u2__abc_44228_n3109;
  wire u2__abc_44228_n3110;
  wire u2__abc_44228_n3111;
  wire u2__abc_44228_n3112;
  wire u2__abc_44228_n3113;
  wire u2__abc_44228_n3114;
  wire u2__abc_44228_n3115;
  wire u2__abc_44228_n3116;
  wire u2__abc_44228_n3117;
  wire u2__abc_44228_n3118;
  wire u2__abc_44228_n3119;
  wire u2__abc_44228_n3120;
  wire u2__abc_44228_n3121;
  wire u2__abc_44228_n3122;
  wire u2__abc_44228_n3123;
  wire u2__abc_44228_n3124;
  wire u2__abc_44228_n3125;
  wire u2__abc_44228_n3126;
  wire u2__abc_44228_n3127;
  wire u2__abc_44228_n3128;
  wire u2__abc_44228_n3129;
  wire u2__abc_44228_n3130;
  wire u2__abc_44228_n3131;
  wire u2__abc_44228_n3132;
  wire u2__abc_44228_n3133;
  wire u2__abc_44228_n3134;
  wire u2__abc_44228_n3135;
  wire u2__abc_44228_n3136;
  wire u2__abc_44228_n3137;
  wire u2__abc_44228_n3138;
  wire u2__abc_44228_n3139;
  wire u2__abc_44228_n3140;
  wire u2__abc_44228_n3141;
  wire u2__abc_44228_n3142;
  wire u2__abc_44228_n3143;
  wire u2__abc_44228_n3144;
  wire u2__abc_44228_n3145;
  wire u2__abc_44228_n3146;
  wire u2__abc_44228_n3147;
  wire u2__abc_44228_n3148;
  wire u2__abc_44228_n3149;
  wire u2__abc_44228_n3150;
  wire u2__abc_44228_n3151;
  wire u2__abc_44228_n3152;
  wire u2__abc_44228_n3153;
  wire u2__abc_44228_n3154;
  wire u2__abc_44228_n3155;
  wire u2__abc_44228_n3156;
  wire u2__abc_44228_n3157;
  wire u2__abc_44228_n3158;
  wire u2__abc_44228_n3159;
  wire u2__abc_44228_n3160;
  wire u2__abc_44228_n3161;
  wire u2__abc_44228_n3162;
  wire u2__abc_44228_n3163;
  wire u2__abc_44228_n3164;
  wire u2__abc_44228_n3165;
  wire u2__abc_44228_n3166;
  wire u2__abc_44228_n3167;
  wire u2__abc_44228_n3168;
  wire u2__abc_44228_n3169;
  wire u2__abc_44228_n3170;
  wire u2__abc_44228_n3171;
  wire u2__abc_44228_n3172;
  wire u2__abc_44228_n3173;
  wire u2__abc_44228_n3174;
  wire u2__abc_44228_n3175;
  wire u2__abc_44228_n3176;
  wire u2__abc_44228_n3177;
  wire u2__abc_44228_n3178;
  wire u2__abc_44228_n3179;
  wire u2__abc_44228_n3180;
  wire u2__abc_44228_n3181;
  wire u2__abc_44228_n3182;
  wire u2__abc_44228_n3183;
  wire u2__abc_44228_n3184;
  wire u2__abc_44228_n3185;
  wire u2__abc_44228_n3186;
  wire u2__abc_44228_n3187;
  wire u2__abc_44228_n3188;
  wire u2__abc_44228_n3189;
  wire u2__abc_44228_n3190;
  wire u2__abc_44228_n3191;
  wire u2__abc_44228_n3192;
  wire u2__abc_44228_n3193;
  wire u2__abc_44228_n3194;
  wire u2__abc_44228_n3195;
  wire u2__abc_44228_n3196;
  wire u2__abc_44228_n3197;
  wire u2__abc_44228_n3198;
  wire u2__abc_44228_n3199;
  wire u2__abc_44228_n3200;
  wire u2__abc_44228_n3201;
  wire u2__abc_44228_n3202;
  wire u2__abc_44228_n3203;
  wire u2__abc_44228_n3204;
  wire u2__abc_44228_n3205;
  wire u2__abc_44228_n3206;
  wire u2__abc_44228_n3207;
  wire u2__abc_44228_n3208;
  wire u2__abc_44228_n3209;
  wire u2__abc_44228_n3210;
  wire u2__abc_44228_n3211;
  wire u2__abc_44228_n3212;
  wire u2__abc_44228_n3213;
  wire u2__abc_44228_n3214;
  wire u2__abc_44228_n3215;
  wire u2__abc_44228_n3216;
  wire u2__abc_44228_n3217;
  wire u2__abc_44228_n3218;
  wire u2__abc_44228_n3219;
  wire u2__abc_44228_n3220;
  wire u2__abc_44228_n3221;
  wire u2__abc_44228_n3222;
  wire u2__abc_44228_n3223;
  wire u2__abc_44228_n3224;
  wire u2__abc_44228_n3225;
  wire u2__abc_44228_n3226;
  wire u2__abc_44228_n3227;
  wire u2__abc_44228_n3228;
  wire u2__abc_44228_n3229;
  wire u2__abc_44228_n3230;
  wire u2__abc_44228_n3231;
  wire u2__abc_44228_n3232;
  wire u2__abc_44228_n3233;
  wire u2__abc_44228_n3234;
  wire u2__abc_44228_n3235;
  wire u2__abc_44228_n3236;
  wire u2__abc_44228_n3237;
  wire u2__abc_44228_n3238;
  wire u2__abc_44228_n3239;
  wire u2__abc_44228_n3240;
  wire u2__abc_44228_n3241;
  wire u2__abc_44228_n3242;
  wire u2__abc_44228_n3243;
  wire u2__abc_44228_n3244;
  wire u2__abc_44228_n3245;
  wire u2__abc_44228_n3246;
  wire u2__abc_44228_n3247;
  wire u2__abc_44228_n3248;
  wire u2__abc_44228_n3249;
  wire u2__abc_44228_n3250;
  wire u2__abc_44228_n3251;
  wire u2__abc_44228_n3252;
  wire u2__abc_44228_n3253;
  wire u2__abc_44228_n3254;
  wire u2__abc_44228_n3255;
  wire u2__abc_44228_n3256;
  wire u2__abc_44228_n3257;
  wire u2__abc_44228_n3258;
  wire u2__abc_44228_n3259;
  wire u2__abc_44228_n3260;
  wire u2__abc_44228_n3261;
  wire u2__abc_44228_n3262;
  wire u2__abc_44228_n3263;
  wire u2__abc_44228_n3264;
  wire u2__abc_44228_n3265;
  wire u2__abc_44228_n3266;
  wire u2__abc_44228_n3267;
  wire u2__abc_44228_n3268;
  wire u2__abc_44228_n3269;
  wire u2__abc_44228_n3270;
  wire u2__abc_44228_n3271;
  wire u2__abc_44228_n3272;
  wire u2__abc_44228_n3273;
  wire u2__abc_44228_n3274;
  wire u2__abc_44228_n3275;
  wire u2__abc_44228_n3276;
  wire u2__abc_44228_n3277;
  wire u2__abc_44228_n3278;
  wire u2__abc_44228_n3279;
  wire u2__abc_44228_n3280;
  wire u2__abc_44228_n3281;
  wire u2__abc_44228_n3282;
  wire u2__abc_44228_n3283;
  wire u2__abc_44228_n3284;
  wire u2__abc_44228_n3285;
  wire u2__abc_44228_n3286;
  wire u2__abc_44228_n3287;
  wire u2__abc_44228_n3288;
  wire u2__abc_44228_n3289;
  wire u2__abc_44228_n3290;
  wire u2__abc_44228_n3291;
  wire u2__abc_44228_n3292;
  wire u2__abc_44228_n3293;
  wire u2__abc_44228_n3294;
  wire u2__abc_44228_n3295;
  wire u2__abc_44228_n3296;
  wire u2__abc_44228_n3297;
  wire u2__abc_44228_n3298;
  wire u2__abc_44228_n3299;
  wire u2__abc_44228_n3300;
  wire u2__abc_44228_n3301;
  wire u2__abc_44228_n3302;
  wire u2__abc_44228_n3303;
  wire u2__abc_44228_n3304;
  wire u2__abc_44228_n3305;
  wire u2__abc_44228_n3306;
  wire u2__abc_44228_n3307;
  wire u2__abc_44228_n3308;
  wire u2__abc_44228_n3309;
  wire u2__abc_44228_n3310;
  wire u2__abc_44228_n3311;
  wire u2__abc_44228_n3312;
  wire u2__abc_44228_n3313;
  wire u2__abc_44228_n3314;
  wire u2__abc_44228_n3315;
  wire u2__abc_44228_n3316;
  wire u2__abc_44228_n3317;
  wire u2__abc_44228_n3318;
  wire u2__abc_44228_n3319;
  wire u2__abc_44228_n3320;
  wire u2__abc_44228_n3321;
  wire u2__abc_44228_n3322;
  wire u2__abc_44228_n3323;
  wire u2__abc_44228_n3324;
  wire u2__abc_44228_n3325;
  wire u2__abc_44228_n3326;
  wire u2__abc_44228_n3327;
  wire u2__abc_44228_n3328;
  wire u2__abc_44228_n3329;
  wire u2__abc_44228_n3330;
  wire u2__abc_44228_n3331;
  wire u2__abc_44228_n3332;
  wire u2__abc_44228_n3333;
  wire u2__abc_44228_n3334;
  wire u2__abc_44228_n3335;
  wire u2__abc_44228_n3336;
  wire u2__abc_44228_n3337;
  wire u2__abc_44228_n3338;
  wire u2__abc_44228_n3339;
  wire u2__abc_44228_n3340;
  wire u2__abc_44228_n3341;
  wire u2__abc_44228_n3342;
  wire u2__abc_44228_n3343;
  wire u2__abc_44228_n3344;
  wire u2__abc_44228_n3345;
  wire u2__abc_44228_n3346;
  wire u2__abc_44228_n3347;
  wire u2__abc_44228_n3348;
  wire u2__abc_44228_n3349;
  wire u2__abc_44228_n3350;
  wire u2__abc_44228_n3351;
  wire u2__abc_44228_n3352;
  wire u2__abc_44228_n3353;
  wire u2__abc_44228_n3354;
  wire u2__abc_44228_n3355;
  wire u2__abc_44228_n3356;
  wire u2__abc_44228_n3357;
  wire u2__abc_44228_n3358;
  wire u2__abc_44228_n3359;
  wire u2__abc_44228_n3360;
  wire u2__abc_44228_n3361;
  wire u2__abc_44228_n3362;
  wire u2__abc_44228_n3363;
  wire u2__abc_44228_n3364;
  wire u2__abc_44228_n3365;
  wire u2__abc_44228_n3366;
  wire u2__abc_44228_n3367;
  wire u2__abc_44228_n3368;
  wire u2__abc_44228_n3369;
  wire u2__abc_44228_n3370;
  wire u2__abc_44228_n3371;
  wire u2__abc_44228_n3372;
  wire u2__abc_44228_n3373;
  wire u2__abc_44228_n3374;
  wire u2__abc_44228_n3375;
  wire u2__abc_44228_n3376;
  wire u2__abc_44228_n3377;
  wire u2__abc_44228_n3378;
  wire u2__abc_44228_n3379;
  wire u2__abc_44228_n3380;
  wire u2__abc_44228_n3381;
  wire u2__abc_44228_n3382;
  wire u2__abc_44228_n3383;
  wire u2__abc_44228_n3384;
  wire u2__abc_44228_n3385;
  wire u2__abc_44228_n3386;
  wire u2__abc_44228_n3387;
  wire u2__abc_44228_n3388;
  wire u2__abc_44228_n3389;
  wire u2__abc_44228_n3390;
  wire u2__abc_44228_n3391;
  wire u2__abc_44228_n3392;
  wire u2__abc_44228_n3393;
  wire u2__abc_44228_n3394;
  wire u2__abc_44228_n3395;
  wire u2__abc_44228_n3396;
  wire u2__abc_44228_n3397;
  wire u2__abc_44228_n3398;
  wire u2__abc_44228_n3399;
  wire u2__abc_44228_n3400;
  wire u2__abc_44228_n3401;
  wire u2__abc_44228_n3402;
  wire u2__abc_44228_n3403;
  wire u2__abc_44228_n3404;
  wire u2__abc_44228_n3405;
  wire u2__abc_44228_n3406;
  wire u2__abc_44228_n3407;
  wire u2__abc_44228_n3408;
  wire u2__abc_44228_n3409;
  wire u2__abc_44228_n3410;
  wire u2__abc_44228_n3411;
  wire u2__abc_44228_n3412;
  wire u2__abc_44228_n3413;
  wire u2__abc_44228_n3414;
  wire u2__abc_44228_n3415;
  wire u2__abc_44228_n3416;
  wire u2__abc_44228_n3417;
  wire u2__abc_44228_n3418;
  wire u2__abc_44228_n3419;
  wire u2__abc_44228_n3420;
  wire u2__abc_44228_n3421;
  wire u2__abc_44228_n3422;
  wire u2__abc_44228_n3423;
  wire u2__abc_44228_n3424;
  wire u2__abc_44228_n3425;
  wire u2__abc_44228_n3426;
  wire u2__abc_44228_n3427;
  wire u2__abc_44228_n3428;
  wire u2__abc_44228_n3429;
  wire u2__abc_44228_n3430;
  wire u2__abc_44228_n3431;
  wire u2__abc_44228_n3432;
  wire u2__abc_44228_n3433;
  wire u2__abc_44228_n3434;
  wire u2__abc_44228_n3435;
  wire u2__abc_44228_n3436;
  wire u2__abc_44228_n3437;
  wire u2__abc_44228_n3438;
  wire u2__abc_44228_n3439_1;
  wire u2__abc_44228_n3440;
  wire u2__abc_44228_n3441;
  wire u2__abc_44228_n3442;
  wire u2__abc_44228_n3443;
  wire u2__abc_44228_n3444;
  wire u2__abc_44228_n3445;
  wire u2__abc_44228_n3446;
  wire u2__abc_44228_n3447;
  wire u2__abc_44228_n3448;
  wire u2__abc_44228_n3449_1;
  wire u2__abc_44228_n3450;
  wire u2__abc_44228_n3451;
  wire u2__abc_44228_n3452;
  wire u2__abc_44228_n3453;
  wire u2__abc_44228_n3454;
  wire u2__abc_44228_n3455;
  wire u2__abc_44228_n3456;
  wire u2__abc_44228_n3457_1;
  wire u2__abc_44228_n3458;
  wire u2__abc_44228_n3459;
  wire u2__abc_44228_n3460;
  wire u2__abc_44228_n3461;
  wire u2__abc_44228_n3462;
  wire u2__abc_44228_n3463;
  wire u2__abc_44228_n3464;
  wire u2__abc_44228_n3465;
  wire u2__abc_44228_n3466;
  wire u2__abc_44228_n3467_1;
  wire u2__abc_44228_n3468;
  wire u2__abc_44228_n3469;
  wire u2__abc_44228_n3470;
  wire u2__abc_44228_n3471;
  wire u2__abc_44228_n3472;
  wire u2__abc_44228_n3473;
  wire u2__abc_44228_n3474;
  wire u2__abc_44228_n3475_1;
  wire u2__abc_44228_n3476;
  wire u2__abc_44228_n3477;
  wire u2__abc_44228_n3478;
  wire u2__abc_44228_n3479;
  wire u2__abc_44228_n3480;
  wire u2__abc_44228_n3481;
  wire u2__abc_44228_n3482;
  wire u2__abc_44228_n3483;
  wire u2__abc_44228_n3484_1;
  wire u2__abc_44228_n3485;
  wire u2__abc_44228_n3486;
  wire u2__abc_44228_n3487;
  wire u2__abc_44228_n3488;
  wire u2__abc_44228_n3489;
  wire u2__abc_44228_n3490;
  wire u2__abc_44228_n3491;
  wire u2__abc_44228_n3492;
  wire u2__abc_44228_n3493;
  wire u2__abc_44228_n3494;
  wire u2__abc_44228_n3495_1;
  wire u2__abc_44228_n3496;
  wire u2__abc_44228_n3497;
  wire u2__abc_44228_n3498;
  wire u2__abc_44228_n3499;
  wire u2__abc_44228_n3500;
  wire u2__abc_44228_n3501;
  wire u2__abc_44228_n3502;
  wire u2__abc_44228_n3503;
  wire u2__abc_44228_n3504;
  wire u2__abc_44228_n3505_1;
  wire u2__abc_44228_n3506;
  wire u2__abc_44228_n3507;
  wire u2__abc_44228_n3508;
  wire u2__abc_44228_n3509;
  wire u2__abc_44228_n3510;
  wire u2__abc_44228_n3511;
  wire u2__abc_44228_n3512;
  wire u2__abc_44228_n3513_1;
  wire u2__abc_44228_n3514;
  wire u2__abc_44228_n3515;
  wire u2__abc_44228_n3516;
  wire u2__abc_44228_n3517;
  wire u2__abc_44228_n3518;
  wire u2__abc_44228_n3519;
  wire u2__abc_44228_n3520;
  wire u2__abc_44228_n3521;
  wire u2__abc_44228_n3522;
  wire u2__abc_44228_n3523_1;
  wire u2__abc_44228_n3524;
  wire u2__abc_44228_n3525;
  wire u2__abc_44228_n3526;
  wire u2__abc_44228_n3527;
  wire u2__abc_44228_n3528;
  wire u2__abc_44228_n3529;
  wire u2__abc_44228_n3530;
  wire u2__abc_44228_n3531;
  wire u2__abc_44228_n3532_1;
  wire u2__abc_44228_n3533;
  wire u2__abc_44228_n3534;
  wire u2__abc_44228_n3535;
  wire u2__abc_44228_n3536;
  wire u2__abc_44228_n3537;
  wire u2__abc_44228_n3538;
  wire u2__abc_44228_n3539;
  wire u2__abc_44228_n3540;
  wire u2__abc_44228_n3541_1;
  wire u2__abc_44228_n3542;
  wire u2__abc_44228_n3543;
  wire u2__abc_44228_n3544;
  wire u2__abc_44228_n3545;
  wire u2__abc_44228_n3546;
  wire u2__abc_44228_n3547;
  wire u2__abc_44228_n3548;
  wire u2__abc_44228_n3549;
  wire u2__abc_44228_n3550;
  wire u2__abc_44228_n3551;
  wire u2__abc_44228_n3552_1;
  wire u2__abc_44228_n3553;
  wire u2__abc_44228_n3554;
  wire u2__abc_44228_n3555;
  wire u2__abc_44228_n3556;
  wire u2__abc_44228_n3557;
  wire u2__abc_44228_n3558;
  wire u2__abc_44228_n3559;
  wire u2__abc_44228_n3560;
  wire u2__abc_44228_n3561;
  wire u2__abc_44228_n3562_1;
  wire u2__abc_44228_n3563;
  wire u2__abc_44228_n3564;
  wire u2__abc_44228_n3565;
  wire u2__abc_44228_n3566;
  wire u2__abc_44228_n3567;
  wire u2__abc_44228_n3568;
  wire u2__abc_44228_n3569;
  wire u2__abc_44228_n3570;
  wire u2__abc_44228_n3571_1;
  wire u2__abc_44228_n3572;
  wire u2__abc_44228_n3573;
  wire u2__abc_44228_n3574;
  wire u2__abc_44228_n3575;
  wire u2__abc_44228_n3576;
  wire u2__abc_44228_n3577;
  wire u2__abc_44228_n3578;
  wire u2__abc_44228_n3579;
  wire u2__abc_44228_n3580_1;
  wire u2__abc_44228_n3581;
  wire u2__abc_44228_n3582;
  wire u2__abc_44228_n3583;
  wire u2__abc_44228_n3584;
  wire u2__abc_44228_n3585;
  wire u2__abc_44228_n3586;
  wire u2__abc_44228_n3587;
  wire u2__abc_44228_n3588_1;
  wire u2__abc_44228_n3589;
  wire u2__abc_44228_n3590;
  wire u2__abc_44228_n3591;
  wire u2__abc_44228_n3592;
  wire u2__abc_44228_n3593;
  wire u2__abc_44228_n3594;
  wire u2__abc_44228_n3595;
  wire u2__abc_44228_n3596;
  wire u2__abc_44228_n3597_1;
  wire u2__abc_44228_n3598;
  wire u2__abc_44228_n3599;
  wire u2__abc_44228_n3600;
  wire u2__abc_44228_n3601;
  wire u2__abc_44228_n3602;
  wire u2__abc_44228_n3603;
  wire u2__abc_44228_n3604;
  wire u2__abc_44228_n3605;
  wire u2__abc_44228_n3606;
  wire u2__abc_44228_n3607;
  wire u2__abc_44228_n3608_1;
  wire u2__abc_44228_n3609;
  wire u2__abc_44228_n3610;
  wire u2__abc_44228_n3611;
  wire u2__abc_44228_n3612;
  wire u2__abc_44228_n3613;
  wire u2__abc_44228_n3614;
  wire u2__abc_44228_n3615;
  wire u2__abc_44228_n3616;
  wire u2__abc_44228_n3617_1;
  wire u2__abc_44228_n3618;
  wire u2__abc_44228_n3619;
  wire u2__abc_44228_n3620;
  wire u2__abc_44228_n3621;
  wire u2__abc_44228_n3622;
  wire u2__abc_44228_n3623;
  wire u2__abc_44228_n3624;
  wire u2__abc_44228_n3625;
  wire u2__abc_44228_n3626;
  wire u2__abc_44228_n3627_1;
  wire u2__abc_44228_n3628;
  wire u2__abc_44228_n3629;
  wire u2__abc_44228_n3630;
  wire u2__abc_44228_n3631;
  wire u2__abc_44228_n3632;
  wire u2__abc_44228_n3633;
  wire u2__abc_44228_n3634;
  wire u2__abc_44228_n3635;
  wire u2__abc_44228_n3636;
  wire u2__abc_44228_n3637_1;
  wire u2__abc_44228_n3638;
  wire u2__abc_44228_n3639;
  wire u2__abc_44228_n3640;
  wire u2__abc_44228_n3641;
  wire u2__abc_44228_n3642;
  wire u2__abc_44228_n3643;
  wire u2__abc_44228_n3644;
  wire u2__abc_44228_n3645;
  wire u2__abc_44228_n3646;
  wire u2__abc_44228_n3647_1;
  wire u2__abc_44228_n3648;
  wire u2__abc_44228_n3649;
  wire u2__abc_44228_n3650;
  wire u2__abc_44228_n3651;
  wire u2__abc_44228_n3652;
  wire u2__abc_44228_n3653;
  wire u2__abc_44228_n3654;
  wire u2__abc_44228_n3655;
  wire u2__abc_44228_n3656_1;
  wire u2__abc_44228_n3657;
  wire u2__abc_44228_n3658;
  wire u2__abc_44228_n3659;
  wire u2__abc_44228_n3660;
  wire u2__abc_44228_n3661;
  wire u2__abc_44228_n3662;
  wire u2__abc_44228_n3663;
  wire u2__abc_44228_n3664;
  wire u2__abc_44228_n3665;
  wire u2__abc_44228_n3666_1;
  wire u2__abc_44228_n3667;
  wire u2__abc_44228_n3668;
  wire u2__abc_44228_n3669;
  wire u2__abc_44228_n3670;
  wire u2__abc_44228_n3671;
  wire u2__abc_44228_n3672;
  wire u2__abc_44228_n3673;
  wire u2__abc_44228_n3674;
  wire u2__abc_44228_n3675_1;
  wire u2__abc_44228_n3676;
  wire u2__abc_44228_n3677;
  wire u2__abc_44228_n3678;
  wire u2__abc_44228_n3679;
  wire u2__abc_44228_n3680;
  wire u2__abc_44228_n3681;
  wire u2__abc_44228_n3682;
  wire u2__abc_44228_n3683;
  wire u2__abc_44228_n3684;
  wire u2__abc_44228_n3685_1;
  wire u2__abc_44228_n3686;
  wire u2__abc_44228_n3687;
  wire u2__abc_44228_n3688;
  wire u2__abc_44228_n3689;
  wire u2__abc_44228_n3690;
  wire u2__abc_44228_n3691;
  wire u2__abc_44228_n3692;
  wire u2__abc_44228_n3693;
  wire u2__abc_44228_n3694_1;
  wire u2__abc_44228_n3695;
  wire u2__abc_44228_n3696;
  wire u2__abc_44228_n3697;
  wire u2__abc_44228_n3698;
  wire u2__abc_44228_n3699;
  wire u2__abc_44228_n3700;
  wire u2__abc_44228_n3701;
  wire u2__abc_44228_n3702;
  wire u2__abc_44228_n3703;
  wire u2__abc_44228_n3704_1;
  wire u2__abc_44228_n3705;
  wire u2__abc_44228_n3706;
  wire u2__abc_44228_n3707;
  wire u2__abc_44228_n3708;
  wire u2__abc_44228_n3709;
  wire u2__abc_44228_n3710;
  wire u2__abc_44228_n3711;
  wire u2__abc_44228_n3712;
  wire u2__abc_44228_n3713;
  wire u2__abc_44228_n3714_1;
  wire u2__abc_44228_n3715;
  wire u2__abc_44228_n3716;
  wire u2__abc_44228_n3717;
  wire u2__abc_44228_n3718;
  wire u2__abc_44228_n3719;
  wire u2__abc_44228_n3720;
  wire u2__abc_44228_n3721;
  wire u2__abc_44228_n3722;
  wire u2__abc_44228_n3723_1;
  wire u2__abc_44228_n3724;
  wire u2__abc_44228_n3725;
  wire u2__abc_44228_n3726;
  wire u2__abc_44228_n3727;
  wire u2__abc_44228_n3728;
  wire u2__abc_44228_n3729;
  wire u2__abc_44228_n3730;
  wire u2__abc_44228_n3731;
  wire u2__abc_44228_n3732_1;
  wire u2__abc_44228_n3733;
  wire u2__abc_44228_n3734;
  wire u2__abc_44228_n3735;
  wire u2__abc_44228_n3736;
  wire u2__abc_44228_n3737;
  wire u2__abc_44228_n3738;
  wire u2__abc_44228_n3739;
  wire u2__abc_44228_n3740_1;
  wire u2__abc_44228_n3741;
  wire u2__abc_44228_n3742;
  wire u2__abc_44228_n3743;
  wire u2__abc_44228_n3744;
  wire u2__abc_44228_n3745;
  wire u2__abc_44228_n3746;
  wire u2__abc_44228_n3747;
  wire u2__abc_44228_n3748;
  wire u2__abc_44228_n3749;
  wire u2__abc_44228_n3750_1;
  wire u2__abc_44228_n3751;
  wire u2__abc_44228_n3752;
  wire u2__abc_44228_n3753;
  wire u2__abc_44228_n3754;
  wire u2__abc_44228_n3755;
  wire u2__abc_44228_n3756;
  wire u2__abc_44228_n3757;
  wire u2__abc_44228_n3758;
  wire u2__abc_44228_n3759_1;
  wire u2__abc_44228_n3760;
  wire u2__abc_44228_n3761;
  wire u2__abc_44228_n3762;
  wire u2__abc_44228_n3763;
  wire u2__abc_44228_n3764;
  wire u2__abc_44228_n3765;
  wire u2__abc_44228_n3766;
  wire u2__abc_44228_n3767;
  wire u2__abc_44228_n3768_1;
  wire u2__abc_44228_n3769;
  wire u2__abc_44228_n3770;
  wire u2__abc_44228_n3771;
  wire u2__abc_44228_n3772;
  wire u2__abc_44228_n3773;
  wire u2__abc_44228_n3774;
  wire u2__abc_44228_n3775;
  wire u2__abc_44228_n3776;
  wire u2__abc_44228_n3777;
  wire u2__abc_44228_n3778;
  wire u2__abc_44228_n3779_1;
  wire u2__abc_44228_n3780;
  wire u2__abc_44228_n3781;
  wire u2__abc_44228_n3782;
  wire u2__abc_44228_n3783;
  wire u2__abc_44228_n3784;
  wire u2__abc_44228_n3785;
  wire u2__abc_44228_n3786;
  wire u2__abc_44228_n3787;
  wire u2__abc_44228_n3788;
  wire u2__abc_44228_n3789_1;
  wire u2__abc_44228_n3790;
  wire u2__abc_44228_n3791;
  wire u2__abc_44228_n3792;
  wire u2__abc_44228_n3793;
  wire u2__abc_44228_n3794;
  wire u2__abc_44228_n3795;
  wire u2__abc_44228_n3796;
  wire u2__abc_44228_n3797;
  wire u2__abc_44228_n3798_1;
  wire u2__abc_44228_n3799;
  wire u2__abc_44228_n3800;
  wire u2__abc_44228_n3801;
  wire u2__abc_44228_n3802;
  wire u2__abc_44228_n3803;
  wire u2__abc_44228_n3804;
  wire u2__abc_44228_n3805;
  wire u2__abc_44228_n3806;
  wire u2__abc_44228_n3807_1;
  wire u2__abc_44228_n3808;
  wire u2__abc_44228_n3809;
  wire u2__abc_44228_n3810;
  wire u2__abc_44228_n3811;
  wire u2__abc_44228_n3812;
  wire u2__abc_44228_n3813;
  wire u2__abc_44228_n3814;
  wire u2__abc_44228_n3815;
  wire u2__abc_44228_n3816_1;
  wire u2__abc_44228_n3817;
  wire u2__abc_44228_n3818;
  wire u2__abc_44228_n3819;
  wire u2__abc_44228_n3820;
  wire u2__abc_44228_n3821;
  wire u2__abc_44228_n3822;
  wire u2__abc_44228_n3823;
  wire u2__abc_44228_n3824;
  wire u2__abc_44228_n3825_1;
  wire u2__abc_44228_n3826;
  wire u2__abc_44228_n3827;
  wire u2__abc_44228_n3828;
  wire u2__abc_44228_n3829;
  wire u2__abc_44228_n3830;
  wire u2__abc_44228_n3831;
  wire u2__abc_44228_n3832;
  wire u2__abc_44228_n3833;
  wire u2__abc_44228_n3834;
  wire u2__abc_44228_n3835_1;
  wire u2__abc_44228_n3836;
  wire u2__abc_44228_n3837;
  wire u2__abc_44228_n3838;
  wire u2__abc_44228_n3839;
  wire u2__abc_44228_n3840;
  wire u2__abc_44228_n3841;
  wire u2__abc_44228_n3842;
  wire u2__abc_44228_n3843;
  wire u2__abc_44228_n3844_1;
  wire u2__abc_44228_n3845;
  wire u2__abc_44228_n3846;
  wire u2__abc_44228_n3847;
  wire u2__abc_44228_n3848;
  wire u2__abc_44228_n3849;
  wire u2__abc_44228_n3850;
  wire u2__abc_44228_n3851;
  wire u2__abc_44228_n3852;
  wire u2__abc_44228_n3853;
  wire u2__abc_44228_n3854_1;
  wire u2__abc_44228_n3855;
  wire u2__abc_44228_n3856;
  wire u2__abc_44228_n3857;
  wire u2__abc_44228_n3858;
  wire u2__abc_44228_n3859;
  wire u2__abc_44228_n3860;
  wire u2__abc_44228_n3861;
  wire u2__abc_44228_n3862;
  wire u2__abc_44228_n3863;
  wire u2__abc_44228_n3864_1;
  wire u2__abc_44228_n3865;
  wire u2__abc_44228_n3866;
  wire u2__abc_44228_n3867;
  wire u2__abc_44228_n3868;
  wire u2__abc_44228_n3869;
  wire u2__abc_44228_n3870;
  wire u2__abc_44228_n3871;
  wire u2__abc_44228_n3872;
  wire u2__abc_44228_n3873_1;
  wire u2__abc_44228_n3874;
  wire u2__abc_44228_n3875;
  wire u2__abc_44228_n3876;
  wire u2__abc_44228_n3877;
  wire u2__abc_44228_n3878;
  wire u2__abc_44228_n3879;
  wire u2__abc_44228_n3880;
  wire u2__abc_44228_n3881;
  wire u2__abc_44228_n3882_1;
  wire u2__abc_44228_n3883;
  wire u2__abc_44228_n3884;
  wire u2__abc_44228_n3885;
  wire u2__abc_44228_n3886;
  wire u2__abc_44228_n3887;
  wire u2__abc_44228_n3888;
  wire u2__abc_44228_n3889;
  wire u2__abc_44228_n3890;
  wire u2__abc_44228_n3891;
  wire u2__abc_44228_n3892;
  wire u2__abc_44228_n3893_1;
  wire u2__abc_44228_n3894;
  wire u2__abc_44228_n3895;
  wire u2__abc_44228_n3896;
  wire u2__abc_44228_n3897;
  wire u2__abc_44228_n3898;
  wire u2__abc_44228_n3899;
  wire u2__abc_44228_n3900;
  wire u2__abc_44228_n3901;
  wire u2__abc_44228_n3902;
  wire u2__abc_44228_n3903_1;
  wire u2__abc_44228_n3904;
  wire u2__abc_44228_n3905;
  wire u2__abc_44228_n3906;
  wire u2__abc_44228_n3907;
  wire u2__abc_44228_n3908;
  wire u2__abc_44228_n3909;
  wire u2__abc_44228_n3910;
  wire u2__abc_44228_n3911;
  wire u2__abc_44228_n3912_1;
  wire u2__abc_44228_n3913;
  wire u2__abc_44228_n3914;
  wire u2__abc_44228_n3915;
  wire u2__abc_44228_n3916;
  wire u2__abc_44228_n3917;
  wire u2__abc_44228_n3918;
  wire u2__abc_44228_n3919;
  wire u2__abc_44228_n3920;
  wire u2__abc_44228_n3921_1;
  wire u2__abc_44228_n3922;
  wire u2__abc_44228_n3923;
  wire u2__abc_44228_n3924;
  wire u2__abc_44228_n3925;
  wire u2__abc_44228_n3926;
  wire u2__abc_44228_n3927;
  wire u2__abc_44228_n3928;
  wire u2__abc_44228_n3929;
  wire u2__abc_44228_n3930_1;
  wire u2__abc_44228_n3931;
  wire u2__abc_44228_n3932;
  wire u2__abc_44228_n3933;
  wire u2__abc_44228_n3934;
  wire u2__abc_44228_n3935;
  wire u2__abc_44228_n3936;
  wire u2__abc_44228_n3937;
  wire u2__abc_44228_n3938;
  wire u2__abc_44228_n3939;
  wire u2__abc_44228_n3940_1;
  wire u2__abc_44228_n3941;
  wire u2__abc_44228_n3942;
  wire u2__abc_44228_n3943;
  wire u2__abc_44228_n3944;
  wire u2__abc_44228_n3945;
  wire u2__abc_44228_n3946;
  wire u2__abc_44228_n3947;
  wire u2__abc_44228_n3948;
  wire u2__abc_44228_n3949_1;
  wire u2__abc_44228_n3950;
  wire u2__abc_44228_n3951;
  wire u2__abc_44228_n3952;
  wire u2__abc_44228_n3953;
  wire u2__abc_44228_n3954;
  wire u2__abc_44228_n3955;
  wire u2__abc_44228_n3956;
  wire u2__abc_44228_n3957;
  wire u2__abc_44228_n3958_1;
  wire u2__abc_44228_n3959;
  wire u2__abc_44228_n3960;
  wire u2__abc_44228_n3961;
  wire u2__abc_44228_n3962;
  wire u2__abc_44228_n3963;
  wire u2__abc_44228_n3964;
  wire u2__abc_44228_n3965;
  wire u2__abc_44228_n3966;
  wire u2__abc_44228_n3967_1;
  wire u2__abc_44228_n3968;
  wire u2__abc_44228_n3969;
  wire u2__abc_44228_n3970;
  wire u2__abc_44228_n3971;
  wire u2__abc_44228_n3972;
  wire u2__abc_44228_n3973;
  wire u2__abc_44228_n3974;
  wire u2__abc_44228_n3975;
  wire u2__abc_44228_n3976_1;
  wire u2__abc_44228_n3977;
  wire u2__abc_44228_n3978;
  wire u2__abc_44228_n3979;
  wire u2__abc_44228_n3980;
  wire u2__abc_44228_n3981;
  wire u2__abc_44228_n3982;
  wire u2__abc_44228_n3983;
  wire u2__abc_44228_n3984;
  wire u2__abc_44228_n3985;
  wire u2__abc_44228_n3986_1;
  wire u2__abc_44228_n3987;
  wire u2__abc_44228_n3988;
  wire u2__abc_44228_n3989;
  wire u2__abc_44228_n3990;
  wire u2__abc_44228_n3991;
  wire u2__abc_44228_n3992;
  wire u2__abc_44228_n3993;
  wire u2__abc_44228_n3994;
  wire u2__abc_44228_n3995_1;
  wire u2__abc_44228_n3996;
  wire u2__abc_44228_n3997;
  wire u2__abc_44228_n3998;
  wire u2__abc_44228_n3999;
  wire u2__abc_44228_n4000;
  wire u2__abc_44228_n4001;
  wire u2__abc_44228_n4002;
  wire u2__abc_44228_n4003;
  wire u2__abc_44228_n4004;
  wire u2__abc_44228_n4005_1;
  wire u2__abc_44228_n4006;
  wire u2__abc_44228_n4007;
  wire u2__abc_44228_n4008;
  wire u2__abc_44228_n4009;
  wire u2__abc_44228_n4010;
  wire u2__abc_44228_n4011;
  wire u2__abc_44228_n4012;
  wire u2__abc_44228_n4013;
  wire u2__abc_44228_n4014;
  wire u2__abc_44228_n4015_1;
  wire u2__abc_44228_n4016;
  wire u2__abc_44228_n4017;
  wire u2__abc_44228_n4018;
  wire u2__abc_44228_n4019;
  wire u2__abc_44228_n4020;
  wire u2__abc_44228_n4021;
  wire u2__abc_44228_n4022;
  wire u2__abc_44228_n4023;
  wire u2__abc_44228_n4024_1;
  wire u2__abc_44228_n4025;
  wire u2__abc_44228_n4026;
  wire u2__abc_44228_n4027;
  wire u2__abc_44228_n4028;
  wire u2__abc_44228_n4029;
  wire u2__abc_44228_n4030;
  wire u2__abc_44228_n4031;
  wire u2__abc_44228_n4032;
  wire u2__abc_44228_n4033_1;
  wire u2__abc_44228_n4034;
  wire u2__abc_44228_n4035;
  wire u2__abc_44228_n4036;
  wire u2__abc_44228_n4037;
  wire u2__abc_44228_n4038;
  wire u2__abc_44228_n4039;
  wire u2__abc_44228_n4040;
  wire u2__abc_44228_n4041_1;
  wire u2__abc_44228_n4042;
  wire u2__abc_44228_n4043;
  wire u2__abc_44228_n4044;
  wire u2__abc_44228_n4045;
  wire u2__abc_44228_n4046;
  wire u2__abc_44228_n4047;
  wire u2__abc_44228_n4048;
  wire u2__abc_44228_n4049;
  wire u2__abc_44228_n4050_1;
  wire u2__abc_44228_n4051;
  wire u2__abc_44228_n4052;
  wire u2__abc_44228_n4053;
  wire u2__abc_44228_n4054;
  wire u2__abc_44228_n4055;
  wire u2__abc_44228_n4056;
  wire u2__abc_44228_n4057;
  wire u2__abc_44228_n4058;
  wire u2__abc_44228_n4059;
  wire u2__abc_44228_n4060;
  wire u2__abc_44228_n4061_1;
  wire u2__abc_44228_n4062;
  wire u2__abc_44228_n4063;
  wire u2__abc_44228_n4064;
  wire u2__abc_44228_n4065;
  wire u2__abc_44228_n4066;
  wire u2__abc_44228_n4067;
  wire u2__abc_44228_n4068;
  wire u2__abc_44228_n4069;
  wire u2__abc_44228_n4070_1;
  wire u2__abc_44228_n4071;
  wire u2__abc_44228_n4072;
  wire u2__abc_44228_n4073;
  wire u2__abc_44228_n4074;
  wire u2__abc_44228_n4075;
  wire u2__abc_44228_n4076;
  wire u2__abc_44228_n4077;
  wire u2__abc_44228_n4078;
  wire u2__abc_44228_n4079;
  wire u2__abc_44228_n4080_1;
  wire u2__abc_44228_n4081;
  wire u2__abc_44228_n4082;
  wire u2__abc_44228_n4083;
  wire u2__abc_44228_n4084;
  wire u2__abc_44228_n4085;
  wire u2__abc_44228_n4086;
  wire u2__abc_44228_n4087;
  wire u2__abc_44228_n4088;
  wire u2__abc_44228_n4089;
  wire u2__abc_44228_n4090_1;
  wire u2__abc_44228_n4091;
  wire u2__abc_44228_n4092;
  wire u2__abc_44228_n4093;
  wire u2__abc_44228_n4094;
  wire u2__abc_44228_n4095;
  wire u2__abc_44228_n4096;
  wire u2__abc_44228_n4097;
  wire u2__abc_44228_n4098;
  wire u2__abc_44228_n4099;
  wire u2__abc_44228_n4100_1;
  wire u2__abc_44228_n4101;
  wire u2__abc_44228_n4102;
  wire u2__abc_44228_n4103;
  wire u2__abc_44228_n4104;
  wire u2__abc_44228_n4105;
  wire u2__abc_44228_n4106;
  wire u2__abc_44228_n4107;
  wire u2__abc_44228_n4108;
  wire u2__abc_44228_n4109_1;
  wire u2__abc_44228_n4110;
  wire u2__abc_44228_n4111;
  wire u2__abc_44228_n4112;
  wire u2__abc_44228_n4113;
  wire u2__abc_44228_n4114;
  wire u2__abc_44228_n4115;
  wire u2__abc_44228_n4116;
  wire u2__abc_44228_n4117;
  wire u2__abc_44228_n4118;
  wire u2__abc_44228_n4119_1;
  wire u2__abc_44228_n4120;
  wire u2__abc_44228_n4121;
  wire u2__abc_44228_n4122;
  wire u2__abc_44228_n4123;
  wire u2__abc_44228_n4124;
  wire u2__abc_44228_n4125;
  wire u2__abc_44228_n4126;
  wire u2__abc_44228_n4127;
  wire u2__abc_44228_n4128_1;
  wire u2__abc_44228_n4129;
  wire u2__abc_44228_n4130;
  wire u2__abc_44228_n4131;
  wire u2__abc_44228_n4132;
  wire u2__abc_44228_n4133;
  wire u2__abc_44228_n4134;
  wire u2__abc_44228_n4135;
  wire u2__abc_44228_n4136;
  wire u2__abc_44228_n4137;
  wire u2__abc_44228_n4138_1;
  wire u2__abc_44228_n4139;
  wire u2__abc_44228_n4140;
  wire u2__abc_44228_n4141;
  wire u2__abc_44228_n4142;
  wire u2__abc_44228_n4143;
  wire u2__abc_44228_n4144;
  wire u2__abc_44228_n4145;
  wire u2__abc_44228_n4146;
  wire u2__abc_44228_n4147_1;
  wire u2__abc_44228_n4148;
  wire u2__abc_44228_n4149;
  wire u2__abc_44228_n4150;
  wire u2__abc_44228_n4151;
  wire u2__abc_44228_n4152;
  wire u2__abc_44228_n4153;
  wire u2__abc_44228_n4154;
  wire u2__abc_44228_n4155;
  wire u2__abc_44228_n4156;
  wire u2__abc_44228_n4157_1;
  wire u2__abc_44228_n4158;
  wire u2__abc_44228_n4159;
  wire u2__abc_44228_n4160;
  wire u2__abc_44228_n4161;
  wire u2__abc_44228_n4162;
  wire u2__abc_44228_n4163;
  wire u2__abc_44228_n4164;
  wire u2__abc_44228_n4165;
  wire u2__abc_44228_n4166;
  wire u2__abc_44228_n4167_1;
  wire u2__abc_44228_n4168;
  wire u2__abc_44228_n4169;
  wire u2__abc_44228_n4170;
  wire u2__abc_44228_n4171;
  wire u2__abc_44228_n4172;
  wire u2__abc_44228_n4173;
  wire u2__abc_44228_n4174;
  wire u2__abc_44228_n4175;
  wire u2__abc_44228_n4176_1;
  wire u2__abc_44228_n4177;
  wire u2__abc_44228_n4178;
  wire u2__abc_44228_n4179;
  wire u2__abc_44228_n4180;
  wire u2__abc_44228_n4181;
  wire u2__abc_44228_n4182;
  wire u2__abc_44228_n4183;
  wire u2__abc_44228_n4184;
  wire u2__abc_44228_n4185_1;
  wire u2__abc_44228_n4186;
  wire u2__abc_44228_n4187;
  wire u2__abc_44228_n4188;
  wire u2__abc_44228_n4189;
  wire u2__abc_44228_n4190;
  wire u2__abc_44228_n4191;
  wire u2__abc_44228_n4192;
  wire u2__abc_44228_n4193;
  wire u2__abc_44228_n4194;
  wire u2__abc_44228_n4195_1;
  wire u2__abc_44228_n4196;
  wire u2__abc_44228_n4197;
  wire u2__abc_44228_n4198;
  wire u2__abc_44228_n4199;
  wire u2__abc_44228_n4200;
  wire u2__abc_44228_n4201;
  wire u2__abc_44228_n4202;
  wire u2__abc_44228_n4203;
  wire u2__abc_44228_n4204;
  wire u2__abc_44228_n4205_1;
  wire u2__abc_44228_n4206;
  wire u2__abc_44228_n4207;
  wire u2__abc_44228_n4208;
  wire u2__abc_44228_n4209;
  wire u2__abc_44228_n4210;
  wire u2__abc_44228_n4211;
  wire u2__abc_44228_n4212;
  wire u2__abc_44228_n4213;
  wire u2__abc_44228_n4214;
  wire u2__abc_44228_n4215_1;
  wire u2__abc_44228_n4216;
  wire u2__abc_44228_n4217;
  wire u2__abc_44228_n4218;
  wire u2__abc_44228_n4219;
  wire u2__abc_44228_n4220;
  wire u2__abc_44228_n4221;
  wire u2__abc_44228_n4222;
  wire u2__abc_44228_n4223;
  wire u2__abc_44228_n4224_1;
  wire u2__abc_44228_n4225;
  wire u2__abc_44228_n4226;
  wire u2__abc_44228_n4227;
  wire u2__abc_44228_n4228;
  wire u2__abc_44228_n4229;
  wire u2__abc_44228_n4230;
  wire u2__abc_44228_n4231;
  wire u2__abc_44228_n4232;
  wire u2__abc_44228_n4233_1;
  wire u2__abc_44228_n4234;
  wire u2__abc_44228_n4235;
  wire u2__abc_44228_n4236;
  wire u2__abc_44228_n4237;
  wire u2__abc_44228_n4238;
  wire u2__abc_44228_n4239;
  wire u2__abc_44228_n4240;
  wire u2__abc_44228_n4241;
  wire u2__abc_44228_n4242;
  wire u2__abc_44228_n4243_1;
  wire u2__abc_44228_n4244;
  wire u2__abc_44228_n4245;
  wire u2__abc_44228_n4246;
  wire u2__abc_44228_n4247;
  wire u2__abc_44228_n4248;
  wire u2__abc_44228_n4249;
  wire u2__abc_44228_n4250;
  wire u2__abc_44228_n4251;
  wire u2__abc_44228_n4252;
  wire u2__abc_44228_n4253_1;
  wire u2__abc_44228_n4254;
  wire u2__abc_44228_n4255;
  wire u2__abc_44228_n4256;
  wire u2__abc_44228_n4257;
  wire u2__abc_44228_n4258;
  wire u2__abc_44228_n4259;
  wire u2__abc_44228_n4260;
  wire u2__abc_44228_n4261;
  wire u2__abc_44228_n4262_1;
  wire u2__abc_44228_n4263;
  wire u2__abc_44228_n4264;
  wire u2__abc_44228_n4265;
  wire u2__abc_44228_n4266;
  wire u2__abc_44228_n4267;
  wire u2__abc_44228_n4268;
  wire u2__abc_44228_n4269;
  wire u2__abc_44228_n4270;
  wire u2__abc_44228_n4271;
  wire u2__abc_44228_n4272_1;
  wire u2__abc_44228_n4273;
  wire u2__abc_44228_n4274;
  wire u2__abc_44228_n4275;
  wire u2__abc_44228_n4276;
  wire u2__abc_44228_n4277;
  wire u2__abc_44228_n4278;
  wire u2__abc_44228_n4279;
  wire u2__abc_44228_n4280;
  wire u2__abc_44228_n4281_1;
  wire u2__abc_44228_n4282;
  wire u2__abc_44228_n4283;
  wire u2__abc_44228_n4284;
  wire u2__abc_44228_n4285;
  wire u2__abc_44228_n4286;
  wire u2__abc_44228_n4287;
  wire u2__abc_44228_n4288;
  wire u2__abc_44228_n4289;
  wire u2__abc_44228_n4290;
  wire u2__abc_44228_n4291_1;
  wire u2__abc_44228_n4292;
  wire u2__abc_44228_n4293;
  wire u2__abc_44228_n4294;
  wire u2__abc_44228_n4295;
  wire u2__abc_44228_n4296;
  wire u2__abc_44228_n4297;
  wire u2__abc_44228_n4298;
  wire u2__abc_44228_n4299;
  wire u2__abc_44228_n4300_1;
  wire u2__abc_44228_n4301;
  wire u2__abc_44228_n4302;
  wire u2__abc_44228_n4303;
  wire u2__abc_44228_n4304;
  wire u2__abc_44228_n4305;
  wire u2__abc_44228_n4306;
  wire u2__abc_44228_n4307;
  wire u2__abc_44228_n4308;
  wire u2__abc_44228_n4309;
  wire u2__abc_44228_n4310_1;
  wire u2__abc_44228_n4311;
  wire u2__abc_44228_n4312;
  wire u2__abc_44228_n4313;
  wire u2__abc_44228_n4314;
  wire u2__abc_44228_n4315;
  wire u2__abc_44228_n4316;
  wire u2__abc_44228_n4317;
  wire u2__abc_44228_n4318;
  wire u2__abc_44228_n4319;
  wire u2__abc_44228_n4320_1;
  wire u2__abc_44228_n4321;
  wire u2__abc_44228_n4322;
  wire u2__abc_44228_n4323;
  wire u2__abc_44228_n4324;
  wire u2__abc_44228_n4325;
  wire u2__abc_44228_n4326;
  wire u2__abc_44228_n4327;
  wire u2__abc_44228_n4328;
  wire u2__abc_44228_n4329_1;
  wire u2__abc_44228_n4330;
  wire u2__abc_44228_n4331;
  wire u2__abc_44228_n4332;
  wire u2__abc_44228_n4333;
  wire u2__abc_44228_n4334;
  wire u2__abc_44228_n4335;
  wire u2__abc_44228_n4336;
  wire u2__abc_44228_n4337;
  wire u2__abc_44228_n4338_1;
  wire u2__abc_44228_n4339;
  wire u2__abc_44228_n4340;
  wire u2__abc_44228_n4341;
  wire u2__abc_44228_n4342;
  wire u2__abc_44228_n4343;
  wire u2__abc_44228_n4344;
  wire u2__abc_44228_n4345;
  wire u2__abc_44228_n4346;
  wire u2__abc_44228_n4347;
  wire u2__abc_44228_n4348;
  wire u2__abc_44228_n4349_1;
  wire u2__abc_44228_n4350;
  wire u2__abc_44228_n4351;
  wire u2__abc_44228_n4352;
  wire u2__abc_44228_n4353;
  wire u2__abc_44228_n4354;
  wire u2__abc_44228_n4355;
  wire u2__abc_44228_n4356;
  wire u2__abc_44228_n4357;
  wire u2__abc_44228_n4358;
  wire u2__abc_44228_n4359_1;
  wire u2__abc_44228_n4360;
  wire u2__abc_44228_n4361;
  wire u2__abc_44228_n4362;
  wire u2__abc_44228_n4363;
  wire u2__abc_44228_n4364;
  wire u2__abc_44228_n4365;
  wire u2__abc_44228_n4366;
  wire u2__abc_44228_n4367;
  wire u2__abc_44228_n4368_1;
  wire u2__abc_44228_n4369;
  wire u2__abc_44228_n4370;
  wire u2__abc_44228_n4371;
  wire u2__abc_44228_n4372;
  wire u2__abc_44228_n4373;
  wire u2__abc_44228_n4374;
  wire u2__abc_44228_n4375;
  wire u2__abc_44228_n4376;
  wire u2__abc_44228_n4377_1;
  wire u2__abc_44228_n4378;
  wire u2__abc_44228_n4379;
  wire u2__abc_44228_n4380;
  wire u2__abc_44228_n4381;
  wire u2__abc_44228_n4382;
  wire u2__abc_44228_n4383;
  wire u2__abc_44228_n4384;
  wire u2__abc_44228_n4385;
  wire u2__abc_44228_n4386_1;
  wire u2__abc_44228_n4387;
  wire u2__abc_44228_n4388;
  wire u2__abc_44228_n4389;
  wire u2__abc_44228_n4390;
  wire u2__abc_44228_n4391;
  wire u2__abc_44228_n4392;
  wire u2__abc_44228_n4393;
  wire u2__abc_44228_n4394;
  wire u2__abc_44228_n4395;
  wire u2__abc_44228_n4396_1;
  wire u2__abc_44228_n4397;
  wire u2__abc_44228_n4398;
  wire u2__abc_44228_n4399;
  wire u2__abc_44228_n4400;
  wire u2__abc_44228_n4401;
  wire u2__abc_44228_n4402;
  wire u2__abc_44228_n4403;
  wire u2__abc_44228_n4404;
  wire u2__abc_44228_n4405_1;
  wire u2__abc_44228_n4406;
  wire u2__abc_44228_n4407;
  wire u2__abc_44228_n4408;
  wire u2__abc_44228_n4409;
  wire u2__abc_44228_n4410;
  wire u2__abc_44228_n4411;
  wire u2__abc_44228_n4412;
  wire u2__abc_44228_n4413;
  wire u2__abc_44228_n4414_1;
  wire u2__abc_44228_n4415;
  wire u2__abc_44228_n4416;
  wire u2__abc_44228_n4417;
  wire u2__abc_44228_n4418;
  wire u2__abc_44228_n4419;
  wire u2__abc_44228_n4420;
  wire u2__abc_44228_n4421;
  wire u2__abc_44228_n4422;
  wire u2__abc_44228_n4423_1;
  wire u2__abc_44228_n4424;
  wire u2__abc_44228_n4425;
  wire u2__abc_44228_n4426;
  wire u2__abc_44228_n4427;
  wire u2__abc_44228_n4428;
  wire u2__abc_44228_n4429;
  wire u2__abc_44228_n4430;
  wire u2__abc_44228_n4431;
  wire u2__abc_44228_n4432_1;
  wire u2__abc_44228_n4433;
  wire u2__abc_44228_n4434;
  wire u2__abc_44228_n4435;
  wire u2__abc_44228_n4436;
  wire u2__abc_44228_n4437;
  wire u2__abc_44228_n4438;
  wire u2__abc_44228_n4439;
  wire u2__abc_44228_n4440;
  wire u2__abc_44228_n4441;
  wire u2__abc_44228_n4442_1;
  wire u2__abc_44228_n4443;
  wire u2__abc_44228_n4444;
  wire u2__abc_44228_n4445;
  wire u2__abc_44228_n4446;
  wire u2__abc_44228_n4447;
  wire u2__abc_44228_n4448;
  wire u2__abc_44228_n4449;
  wire u2__abc_44228_n4450;
  wire u2__abc_44228_n4451_1;
  wire u2__abc_44228_n4452;
  wire u2__abc_44228_n4453;
  wire u2__abc_44228_n4454;
  wire u2__abc_44228_n4455;
  wire u2__abc_44228_n4456;
  wire u2__abc_44228_n4457;
  wire u2__abc_44228_n4458;
  wire u2__abc_44228_n4459;
  wire u2__abc_44228_n4460;
  wire u2__abc_44228_n4461_1;
  wire u2__abc_44228_n4462;
  wire u2__abc_44228_n4463;
  wire u2__abc_44228_n4464;
  wire u2__abc_44228_n4465;
  wire u2__abc_44228_n4466;
  wire u2__abc_44228_n4467;
  wire u2__abc_44228_n4468;
  wire u2__abc_44228_n4469;
  wire u2__abc_44228_n4470;
  wire u2__abc_44228_n4471_1;
  wire u2__abc_44228_n4472;
  wire u2__abc_44228_n4473;
  wire u2__abc_44228_n4474;
  wire u2__abc_44228_n4475;
  wire u2__abc_44228_n4476;
  wire u2__abc_44228_n4477;
  wire u2__abc_44228_n4478;
  wire u2__abc_44228_n4479;
  wire u2__abc_44228_n4480_1;
  wire u2__abc_44228_n4481;
  wire u2__abc_44228_n4482;
  wire u2__abc_44228_n4483;
  wire u2__abc_44228_n4484;
  wire u2__abc_44228_n4485;
  wire u2__abc_44228_n4486;
  wire u2__abc_44228_n4487;
  wire u2__abc_44228_n4488;
  wire u2__abc_44228_n4489_1;
  wire u2__abc_44228_n4490;
  wire u2__abc_44228_n4491;
  wire u2__abc_44228_n4492;
  wire u2__abc_44228_n4493;
  wire u2__abc_44228_n4494;
  wire u2__abc_44228_n4495;
  wire u2__abc_44228_n4496;
  wire u2__abc_44228_n4497;
  wire u2__abc_44228_n4498_1;
  wire u2__abc_44228_n4499;
  wire u2__abc_44228_n4500;
  wire u2__abc_44228_n4501;
  wire u2__abc_44228_n4502;
  wire u2__abc_44228_n4503;
  wire u2__abc_44228_n4504;
  wire u2__abc_44228_n4505;
  wire u2__abc_44228_n4506;
  wire u2__abc_44228_n4507;
  wire u2__abc_44228_n4508_1;
  wire u2__abc_44228_n4509;
  wire u2__abc_44228_n4510;
  wire u2__abc_44228_n4511;
  wire u2__abc_44228_n4512;
  wire u2__abc_44228_n4513;
  wire u2__abc_44228_n4514;
  wire u2__abc_44228_n4515;
  wire u2__abc_44228_n4516;
  wire u2__abc_44228_n4517_1;
  wire u2__abc_44228_n4518;
  wire u2__abc_44228_n4519;
  wire u2__abc_44228_n4520;
  wire u2__abc_44228_n4521;
  wire u2__abc_44228_n4522;
  wire u2__abc_44228_n4523;
  wire u2__abc_44228_n4524;
  wire u2__abc_44228_n4525;
  wire u2__abc_44228_n4526_1;
  wire u2__abc_44228_n4527;
  wire u2__abc_44228_n4528;
  wire u2__abc_44228_n4529;
  wire u2__abc_44228_n4530;
  wire u2__abc_44228_n4531;
  wire u2__abc_44228_n4532;
  wire u2__abc_44228_n4533;
  wire u2__abc_44228_n4534;
  wire u2__abc_44228_n4535_1;
  wire u2__abc_44228_n4536;
  wire u2__abc_44228_n4537;
  wire u2__abc_44228_n4538;
  wire u2__abc_44228_n4539;
  wire u2__abc_44228_n4540;
  wire u2__abc_44228_n4541;
  wire u2__abc_44228_n4542;
  wire u2__abc_44228_n4543;
  wire u2__abc_44228_n4544;
  wire u2__abc_44228_n4545_1;
  wire u2__abc_44228_n4546;
  wire u2__abc_44228_n4547;
  wire u2__abc_44228_n4548;
  wire u2__abc_44228_n4549;
  wire u2__abc_44228_n4550;
  wire u2__abc_44228_n4551;
  wire u2__abc_44228_n4552;
  wire u2__abc_44228_n4553;
  wire u2__abc_44228_n4554_1;
  wire u2__abc_44228_n4555;
  wire u2__abc_44228_n4556;
  wire u2__abc_44228_n4557;
  wire u2__abc_44228_n4558;
  wire u2__abc_44228_n4559;
  wire u2__abc_44228_n4560;
  wire u2__abc_44228_n4561;
  wire u2__abc_44228_n4562;
  wire u2__abc_44228_n4563_1;
  wire u2__abc_44228_n4564;
  wire u2__abc_44228_n4565;
  wire u2__abc_44228_n4566;
  wire u2__abc_44228_n4567;
  wire u2__abc_44228_n4568;
  wire u2__abc_44228_n4569;
  wire u2__abc_44228_n4570;
  wire u2__abc_44228_n4571;
  wire u2__abc_44228_n4572_1;
  wire u2__abc_44228_n4573;
  wire u2__abc_44228_n4574;
  wire u2__abc_44228_n4575;
  wire u2__abc_44228_n4576;
  wire u2__abc_44228_n4577;
  wire u2__abc_44228_n4578;
  wire u2__abc_44228_n4579;
  wire u2__abc_44228_n4580;
  wire u2__abc_44228_n4581_1;
  wire u2__abc_44228_n4582;
  wire u2__abc_44228_n4583;
  wire u2__abc_44228_n4584;
  wire u2__abc_44228_n4585;
  wire u2__abc_44228_n4586;
  wire u2__abc_44228_n4587;
  wire u2__abc_44228_n4588;
  wire u2__abc_44228_n4589;
  wire u2__abc_44228_n4590;
  wire u2__abc_44228_n4591_1;
  wire u2__abc_44228_n4592;
  wire u2__abc_44228_n4593;
  wire u2__abc_44228_n4594;
  wire u2__abc_44228_n4595;
  wire u2__abc_44228_n4596;
  wire u2__abc_44228_n4597;
  wire u2__abc_44228_n4598;
  wire u2__abc_44228_n4599;
  wire u2__abc_44228_n4600_1;
  wire u2__abc_44228_n4601;
  wire u2__abc_44228_n4602;
  wire u2__abc_44228_n4603;
  wire u2__abc_44228_n4604;
  wire u2__abc_44228_n4605;
  wire u2__abc_44228_n4606;
  wire u2__abc_44228_n4607;
  wire u2__abc_44228_n4608;
  wire u2__abc_44228_n4609;
  wire u2__abc_44228_n4610_1;
  wire u2__abc_44228_n4611;
  wire u2__abc_44228_n4612;
  wire u2__abc_44228_n4613;
  wire u2__abc_44228_n4614;
  wire u2__abc_44228_n4615;
  wire u2__abc_44228_n4616;
  wire u2__abc_44228_n4617;
  wire u2__abc_44228_n4618;
  wire u2__abc_44228_n4619;
  wire u2__abc_44228_n4620_1;
  wire u2__abc_44228_n4621;
  wire u2__abc_44228_n4622;
  wire u2__abc_44228_n4623;
  wire u2__abc_44228_n4624;
  wire u2__abc_44228_n4625;
  wire u2__abc_44228_n4626;
  wire u2__abc_44228_n4627;
  wire u2__abc_44228_n4628;
  wire u2__abc_44228_n4629_1;
  wire u2__abc_44228_n4630;
  wire u2__abc_44228_n4631;
  wire u2__abc_44228_n4632;
  wire u2__abc_44228_n4633;
  wire u2__abc_44228_n4634;
  wire u2__abc_44228_n4635;
  wire u2__abc_44228_n4636;
  wire u2__abc_44228_n4637;
  wire u2__abc_44228_n4638_1;
  wire u2__abc_44228_n4639;
  wire u2__abc_44228_n4640;
  wire u2__abc_44228_n4641;
  wire u2__abc_44228_n4642;
  wire u2__abc_44228_n4643;
  wire u2__abc_44228_n4644;
  wire u2__abc_44228_n4645;
  wire u2__abc_44228_n4646_1;
  wire u2__abc_44228_n4647;
  wire u2__abc_44228_n4648;
  wire u2__abc_44228_n4649;
  wire u2__abc_44228_n4650;
  wire u2__abc_44228_n4651;
  wire u2__abc_44228_n4652;
  wire u2__abc_44228_n4653;
  wire u2__abc_44228_n4654;
  wire u2__abc_44228_n4655;
  wire u2__abc_44228_n4656_1;
  wire u2__abc_44228_n4657;
  wire u2__abc_44228_n4658;
  wire u2__abc_44228_n4659;
  wire u2__abc_44228_n4660;
  wire u2__abc_44228_n4661;
  wire u2__abc_44228_n4662;
  wire u2__abc_44228_n4663;
  wire u2__abc_44228_n4664;
  wire u2__abc_44228_n4665_1;
  wire u2__abc_44228_n4666;
  wire u2__abc_44228_n4667;
  wire u2__abc_44228_n4668;
  wire u2__abc_44228_n4669;
  wire u2__abc_44228_n4670;
  wire u2__abc_44228_n4671;
  wire u2__abc_44228_n4672;
  wire u2__abc_44228_n4673;
  wire u2__abc_44228_n4674_1;
  wire u2__abc_44228_n4675;
  wire u2__abc_44228_n4676;
  wire u2__abc_44228_n4677;
  wire u2__abc_44228_n4678;
  wire u2__abc_44228_n4679;
  wire u2__abc_44228_n4680;
  wire u2__abc_44228_n4681;
  wire u2__abc_44228_n4682;
  wire u2__abc_44228_n4683;
  wire u2__abc_44228_n4684;
  wire u2__abc_44228_n4685_1;
  wire u2__abc_44228_n4686;
  wire u2__abc_44228_n4687;
  wire u2__abc_44228_n4688;
  wire u2__abc_44228_n4689;
  wire u2__abc_44228_n4690;
  wire u2__abc_44228_n4691;
  wire u2__abc_44228_n4692;
  wire u2__abc_44228_n4693;
  wire u2__abc_44228_n4694;
  wire u2__abc_44228_n4695_1;
  wire u2__abc_44228_n4696;
  wire u2__abc_44228_n4697;
  wire u2__abc_44228_n4698;
  wire u2__abc_44228_n4699;
  wire u2__abc_44228_n4700;
  wire u2__abc_44228_n4701;
  wire u2__abc_44228_n4702;
  wire u2__abc_44228_n4703;
  wire u2__abc_44228_n4704_1;
  wire u2__abc_44228_n4705;
  wire u2__abc_44228_n4706;
  wire u2__abc_44228_n4707;
  wire u2__abc_44228_n4708;
  wire u2__abc_44228_n4709;
  wire u2__abc_44228_n4710;
  wire u2__abc_44228_n4711;
  wire u2__abc_44228_n4712;
  wire u2__abc_44228_n4713_1;
  wire u2__abc_44228_n4714;
  wire u2__abc_44228_n4715;
  wire u2__abc_44228_n4716;
  wire u2__abc_44228_n4717;
  wire u2__abc_44228_n4718;
  wire u2__abc_44228_n4719;
  wire u2__abc_44228_n4720;
  wire u2__abc_44228_n4721;
  wire u2__abc_44228_n4722_1;
  wire u2__abc_44228_n4723;
  wire u2__abc_44228_n4724;
  wire u2__abc_44228_n4725;
  wire u2__abc_44228_n4726;
  wire u2__abc_44228_n4727;
  wire u2__abc_44228_n4728;
  wire u2__abc_44228_n4729;
  wire u2__abc_44228_n4730;
  wire u2__abc_44228_n4731_1;
  wire u2__abc_44228_n4732;
  wire u2__abc_44228_n4733;
  wire u2__abc_44228_n4734;
  wire u2__abc_44228_n4735;
  wire u2__abc_44228_n4736;
  wire u2__abc_44228_n4737;
  wire u2__abc_44228_n4738;
  wire u2__abc_44228_n4739;
  wire u2__abc_44228_n4740;
  wire u2__abc_44228_n4741_1;
  wire u2__abc_44228_n4742;
  wire u2__abc_44228_n4743;
  wire u2__abc_44228_n4744;
  wire u2__abc_44228_n4745;
  wire u2__abc_44228_n4746;
  wire u2__abc_44228_n4747;
  wire u2__abc_44228_n4748;
  wire u2__abc_44228_n4749;
  wire u2__abc_44228_n4750_1;
  wire u2__abc_44228_n4751;
  wire u2__abc_44228_n4752;
  wire u2__abc_44228_n4753;
  wire u2__abc_44228_n4754;
  wire u2__abc_44228_n4755;
  wire u2__abc_44228_n4756;
  wire u2__abc_44228_n4757;
  wire u2__abc_44228_n4758;
  wire u2__abc_44228_n4759;
  wire u2__abc_44228_n4760_1;
  wire u2__abc_44228_n4761;
  wire u2__abc_44228_n4762;
  wire u2__abc_44228_n4763;
  wire u2__abc_44228_n4764;
  wire u2__abc_44228_n4765;
  wire u2__abc_44228_n4766;
  wire u2__abc_44228_n4767;
  wire u2__abc_44228_n4768;
  wire u2__abc_44228_n4769;
  wire u2__abc_44228_n4770_1;
  wire u2__abc_44228_n4771;
  wire u2__abc_44228_n4772;
  wire u2__abc_44228_n4773;
  wire u2__abc_44228_n4774;
  wire u2__abc_44228_n4775;
  wire u2__abc_44228_n4776;
  wire u2__abc_44228_n4777;
  wire u2__abc_44228_n4778;
  wire u2__abc_44228_n4779_1;
  wire u2__abc_44228_n4780;
  wire u2__abc_44228_n4781;
  wire u2__abc_44228_n4782;
  wire u2__abc_44228_n4783;
  wire u2__abc_44228_n4784;
  wire u2__abc_44228_n4785;
  wire u2__abc_44228_n4786;
  wire u2__abc_44228_n4787;
  wire u2__abc_44228_n4788_1;
  wire u2__abc_44228_n4789;
  wire u2__abc_44228_n4790;
  wire u2__abc_44228_n4791;
  wire u2__abc_44228_n4792;
  wire u2__abc_44228_n4793;
  wire u2__abc_44228_n4794;
  wire u2__abc_44228_n4795;
  wire u2__abc_44228_n4796;
  wire u2__abc_44228_n4797;
  wire u2__abc_44228_n4798;
  wire u2__abc_44228_n4799_1;
  wire u2__abc_44228_n4800;
  wire u2__abc_44228_n4801;
  wire u2__abc_44228_n4802;
  wire u2__abc_44228_n4803;
  wire u2__abc_44228_n4804;
  wire u2__abc_44228_n4805;
  wire u2__abc_44228_n4806;
  wire u2__abc_44228_n4807;
  wire u2__abc_44228_n4808;
  wire u2__abc_44228_n4809_1;
  wire u2__abc_44228_n4810;
  wire u2__abc_44228_n4811;
  wire u2__abc_44228_n4812;
  wire u2__abc_44228_n4813;
  wire u2__abc_44228_n4814;
  wire u2__abc_44228_n4815;
  wire u2__abc_44228_n4816;
  wire u2__abc_44228_n4817;
  wire u2__abc_44228_n4818_1;
  wire u2__abc_44228_n4819;
  wire u2__abc_44228_n4820;
  wire u2__abc_44228_n4821;
  wire u2__abc_44228_n4822;
  wire u2__abc_44228_n4823;
  wire u2__abc_44228_n4824;
  wire u2__abc_44228_n4825;
  wire u2__abc_44228_n4826;
  wire u2__abc_44228_n4827_1;
  wire u2__abc_44228_n4828;
  wire u2__abc_44228_n4829;
  wire u2__abc_44228_n4830;
  wire u2__abc_44228_n4831;
  wire u2__abc_44228_n4832;
  wire u2__abc_44228_n4833;
  wire u2__abc_44228_n4834;
  wire u2__abc_44228_n4835;
  wire u2__abc_44228_n4836_1;
  wire u2__abc_44228_n4837;
  wire u2__abc_44228_n4838;
  wire u2__abc_44228_n4839;
  wire u2__abc_44228_n4840;
  wire u2__abc_44228_n4841;
  wire u2__abc_44228_n4842;
  wire u2__abc_44228_n4843;
  wire u2__abc_44228_n4844;
  wire u2__abc_44228_n4845;
  wire u2__abc_44228_n4846_1;
  wire u2__abc_44228_n4847;
  wire u2__abc_44228_n4848;
  wire u2__abc_44228_n4849;
  wire u2__abc_44228_n4850;
  wire u2__abc_44228_n4851;
  wire u2__abc_44228_n4852;
  wire u2__abc_44228_n4853;
  wire u2__abc_44228_n4854;
  wire u2__abc_44228_n4855_1;
  wire u2__abc_44228_n4856;
  wire u2__abc_44228_n4857;
  wire u2__abc_44228_n4858;
  wire u2__abc_44228_n4859;
  wire u2__abc_44228_n4860;
  wire u2__abc_44228_n4861;
  wire u2__abc_44228_n4862;
  wire u2__abc_44228_n4863;
  wire u2__abc_44228_n4864_1;
  wire u2__abc_44228_n4865;
  wire u2__abc_44228_n4866;
  wire u2__abc_44228_n4867;
  wire u2__abc_44228_n4868;
  wire u2__abc_44228_n4869;
  wire u2__abc_44228_n4870;
  wire u2__abc_44228_n4871;
  wire u2__abc_44228_n4872;
  wire u2__abc_44228_n4873_1;
  wire u2__abc_44228_n4874;
  wire u2__abc_44228_n4875;
  wire u2__abc_44228_n4876;
  wire u2__abc_44228_n4877;
  wire u2__abc_44228_n4878;
  wire u2__abc_44228_n4879;
  wire u2__abc_44228_n4880;
  wire u2__abc_44228_n4881;
  wire u2__abc_44228_n4882_1;
  wire u2__abc_44228_n4883;
  wire u2__abc_44228_n4884;
  wire u2__abc_44228_n4885;
  wire u2__abc_44228_n4886;
  wire u2__abc_44228_n4887;
  wire u2__abc_44228_n4888;
  wire u2__abc_44228_n4889;
  wire u2__abc_44228_n4890;
  wire u2__abc_44228_n4891;
  wire u2__abc_44228_n4892_1;
  wire u2__abc_44228_n4893;
  wire u2__abc_44228_n4894;
  wire u2__abc_44228_n4895;
  wire u2__abc_44228_n4896;
  wire u2__abc_44228_n4897;
  wire u2__abc_44228_n4898;
  wire u2__abc_44228_n4899;
  wire u2__abc_44228_n4900;
  wire u2__abc_44228_n4901_1;
  wire u2__abc_44228_n4902;
  wire u2__abc_44228_n4903;
  wire u2__abc_44228_n4904;
  wire u2__abc_44228_n4905;
  wire u2__abc_44228_n4906;
  wire u2__abc_44228_n4907;
  wire u2__abc_44228_n4908;
  wire u2__abc_44228_n4909;
  wire u2__abc_44228_n4910;
  wire u2__abc_44228_n4911_1;
  wire u2__abc_44228_n4912;
  wire u2__abc_44228_n4913;
  wire u2__abc_44228_n4914;
  wire u2__abc_44228_n4915;
  wire u2__abc_44228_n4916;
  wire u2__abc_44228_n4917;
  wire u2__abc_44228_n4918;
  wire u2__abc_44228_n4919;
  wire u2__abc_44228_n4920;
  wire u2__abc_44228_n4921_1;
  wire u2__abc_44228_n4922;
  wire u2__abc_44228_n4923;
  wire u2__abc_44228_n4924;
  wire u2__abc_44228_n4925;
  wire u2__abc_44228_n4926;
  wire u2__abc_44228_n4927;
  wire u2__abc_44228_n4928;
  wire u2__abc_44228_n4929;
  wire u2__abc_44228_n4930_1;
  wire u2__abc_44228_n4931;
  wire u2__abc_44228_n4932;
  wire u2__abc_44228_n4933;
  wire u2__abc_44228_n4934;
  wire u2__abc_44228_n4935;
  wire u2__abc_44228_n4936;
  wire u2__abc_44228_n4937;
  wire u2__abc_44228_n4938;
  wire u2__abc_44228_n4939_1;
  wire u2__abc_44228_n4940;
  wire u2__abc_44228_n4941;
  wire u2__abc_44228_n4942;
  wire u2__abc_44228_n4943;
  wire u2__abc_44228_n4944;
  wire u2__abc_44228_n4945;
  wire u2__abc_44228_n4946;
  wire u2__abc_44228_n4947;
  wire u2__abc_44228_n4948_1;
  wire u2__abc_44228_n4949;
  wire u2__abc_44228_n4950;
  wire u2__abc_44228_n4951;
  wire u2__abc_44228_n4952;
  wire u2__abc_44228_n4953;
  wire u2__abc_44228_n4954;
  wire u2__abc_44228_n4955;
  wire u2__abc_44228_n4956;
  wire u2__abc_44228_n4957_1;
  wire u2__abc_44228_n4958;
  wire u2__abc_44228_n4959;
  wire u2__abc_44228_n4960;
  wire u2__abc_44228_n4961;
  wire u2__abc_44228_n4962;
  wire u2__abc_44228_n4963;
  wire u2__abc_44228_n4964;
  wire u2__abc_44228_n4965;
  wire u2__abc_44228_n4966;
  wire u2__abc_44228_n4967_1;
  wire u2__abc_44228_n4968;
  wire u2__abc_44228_n4969;
  wire u2__abc_44228_n4970;
  wire u2__abc_44228_n4971;
  wire u2__abc_44228_n4972;
  wire u2__abc_44228_n4973;
  wire u2__abc_44228_n4974;
  wire u2__abc_44228_n4975;
  wire u2__abc_44228_n4976_1;
  wire u2__abc_44228_n4977;
  wire u2__abc_44228_n4978;
  wire u2__abc_44228_n4979;
  wire u2__abc_44228_n4980;
  wire u2__abc_44228_n4981;
  wire u2__abc_44228_n4982;
  wire u2__abc_44228_n4983;
  wire u2__abc_44228_n4984;
  wire u2__abc_44228_n4985;
  wire u2__abc_44228_n4986_1;
  wire u2__abc_44228_n4987;
  wire u2__abc_44228_n4988;
  wire u2__abc_44228_n4989;
  wire u2__abc_44228_n4990;
  wire u2__abc_44228_n4991;
  wire u2__abc_44228_n4992;
  wire u2__abc_44228_n4993;
  wire u2__abc_44228_n4994;
  wire u2__abc_44228_n4995;
  wire u2__abc_44228_n4996_1;
  wire u2__abc_44228_n4997;
  wire u2__abc_44228_n4998;
  wire u2__abc_44228_n4999;
  wire u2__abc_44228_n5000;
  wire u2__abc_44228_n5001;
  wire u2__abc_44228_n5002;
  wire u2__abc_44228_n5003;
  wire u2__abc_44228_n5004;
  wire u2__abc_44228_n5005_1;
  wire u2__abc_44228_n5006;
  wire u2__abc_44228_n5007;
  wire u2__abc_44228_n5008;
  wire u2__abc_44228_n5009;
  wire u2__abc_44228_n5010;
  wire u2__abc_44228_n5011;
  wire u2__abc_44228_n5012;
  wire u2__abc_44228_n5013;
  wire u2__abc_44228_n5014_1;
  wire u2__abc_44228_n5015;
  wire u2__abc_44228_n5016;
  wire u2__abc_44228_n5017;
  wire u2__abc_44228_n5018;
  wire u2__abc_44228_n5019;
  wire u2__abc_44228_n5020;
  wire u2__abc_44228_n5021;
  wire u2__abc_44228_n5022;
  wire u2__abc_44228_n5023_1;
  wire u2__abc_44228_n5024;
  wire u2__abc_44228_n5025;
  wire u2__abc_44228_n5026;
  wire u2__abc_44228_n5027;
  wire u2__abc_44228_n5028;
  wire u2__abc_44228_n5029;
  wire u2__abc_44228_n5030;
  wire u2__abc_44228_n5031;
  wire u2__abc_44228_n5032_1;
  wire u2__abc_44228_n5033;
  wire u2__abc_44228_n5034;
  wire u2__abc_44228_n5035;
  wire u2__abc_44228_n5036;
  wire u2__abc_44228_n5037;
  wire u2__abc_44228_n5038;
  wire u2__abc_44228_n5039;
  wire u2__abc_44228_n5040;
  wire u2__abc_44228_n5041;
  wire u2__abc_44228_n5042_1;
  wire u2__abc_44228_n5043;
  wire u2__abc_44228_n5044;
  wire u2__abc_44228_n5045;
  wire u2__abc_44228_n5046;
  wire u2__abc_44228_n5047;
  wire u2__abc_44228_n5048;
  wire u2__abc_44228_n5049;
  wire u2__abc_44228_n5050;
  wire u2__abc_44228_n5051_1;
  wire u2__abc_44228_n5052;
  wire u2__abc_44228_n5053;
  wire u2__abc_44228_n5054;
  wire u2__abc_44228_n5055;
  wire u2__abc_44228_n5056;
  wire u2__abc_44228_n5057;
  wire u2__abc_44228_n5058;
  wire u2__abc_44228_n5059;
  wire u2__abc_44228_n5060;
  wire u2__abc_44228_n5061_1;
  wire u2__abc_44228_n5062;
  wire u2__abc_44228_n5063;
  wire u2__abc_44228_n5064;
  wire u2__abc_44228_n5065;
  wire u2__abc_44228_n5066;
  wire u2__abc_44228_n5067;
  wire u2__abc_44228_n5068;
  wire u2__abc_44228_n5069;
  wire u2__abc_44228_n5070;
  wire u2__abc_44228_n5071_1;
  wire u2__abc_44228_n5072;
  wire u2__abc_44228_n5073;
  wire u2__abc_44228_n5074;
  wire u2__abc_44228_n5075;
  wire u2__abc_44228_n5076;
  wire u2__abc_44228_n5077;
  wire u2__abc_44228_n5078;
  wire u2__abc_44228_n5079;
  wire u2__abc_44228_n5080_1;
  wire u2__abc_44228_n5081;
  wire u2__abc_44228_n5082;
  wire u2__abc_44228_n5083;
  wire u2__abc_44228_n5084;
  wire u2__abc_44228_n5085;
  wire u2__abc_44228_n5086;
  wire u2__abc_44228_n5087;
  wire u2__abc_44228_n5088;
  wire u2__abc_44228_n5089_1;
  wire u2__abc_44228_n5090;
  wire u2__abc_44228_n5091;
  wire u2__abc_44228_n5092;
  wire u2__abc_44228_n5093;
  wire u2__abc_44228_n5094;
  wire u2__abc_44228_n5095;
  wire u2__abc_44228_n5096;
  wire u2__abc_44228_n5097;
  wire u2__abc_44228_n5098;
  wire u2__abc_44228_n5099_1;
  wire u2__abc_44228_n5100;
  wire u2__abc_44228_n5101;
  wire u2__abc_44228_n5102;
  wire u2__abc_44228_n5103;
  wire u2__abc_44228_n5104;
  wire u2__abc_44228_n5105;
  wire u2__abc_44228_n5106;
  wire u2__abc_44228_n5107;
  wire u2__abc_44228_n5108;
  wire u2__abc_44228_n5109_1;
  wire u2__abc_44228_n5110;
  wire u2__abc_44228_n5111;
  wire u2__abc_44228_n5112;
  wire u2__abc_44228_n5113;
  wire u2__abc_44228_n5114;
  wire u2__abc_44228_n5115;
  wire u2__abc_44228_n5116;
  wire u2__abc_44228_n5117;
  wire u2__abc_44228_n5118_1;
  wire u2__abc_44228_n5119;
  wire u2__abc_44228_n5120;
  wire u2__abc_44228_n5121;
  wire u2__abc_44228_n5122;
  wire u2__abc_44228_n5123;
  wire u2__abc_44228_n5124;
  wire u2__abc_44228_n5125;
  wire u2__abc_44228_n5126;
  wire u2__abc_44228_n5127_1;
  wire u2__abc_44228_n5128;
  wire u2__abc_44228_n5129;
  wire u2__abc_44228_n5130;
  wire u2__abc_44228_n5131;
  wire u2__abc_44228_n5132;
  wire u2__abc_44228_n5133;
  wire u2__abc_44228_n5134;
  wire u2__abc_44228_n5135;
  wire u2__abc_44228_n5136_1;
  wire u2__abc_44228_n5137;
  wire u2__abc_44228_n5138;
  wire u2__abc_44228_n5139;
  wire u2__abc_44228_n5140;
  wire u2__abc_44228_n5141;
  wire u2__abc_44228_n5142;
  wire u2__abc_44228_n5143;
  wire u2__abc_44228_n5144;
  wire u2__abc_44228_n5145;
  wire u2__abc_44228_n5146_1;
  wire u2__abc_44228_n5147;
  wire u2__abc_44228_n5148;
  wire u2__abc_44228_n5149;
  wire u2__abc_44228_n5150;
  wire u2__abc_44228_n5151;
  wire u2__abc_44228_n5152;
  wire u2__abc_44228_n5153;
  wire u2__abc_44228_n5154;
  wire u2__abc_44228_n5155_1;
  wire u2__abc_44228_n5156;
  wire u2__abc_44228_n5157;
  wire u2__abc_44228_n5158;
  wire u2__abc_44228_n5159;
  wire u2__abc_44228_n5160;
  wire u2__abc_44228_n5161;
  wire u2__abc_44228_n5162;
  wire u2__abc_44228_n5163;
  wire u2__abc_44228_n5164_1;
  wire u2__abc_44228_n5165;
  wire u2__abc_44228_n5166;
  wire u2__abc_44228_n5167;
  wire u2__abc_44228_n5168;
  wire u2__abc_44228_n5169;
  wire u2__abc_44228_n5170;
  wire u2__abc_44228_n5171;
  wire u2__abc_44228_n5172;
  wire u2__abc_44228_n5173_1;
  wire u2__abc_44228_n5174;
  wire u2__abc_44228_n5175;
  wire u2__abc_44228_n5176;
  wire u2__abc_44228_n5177;
  wire u2__abc_44228_n5178;
  wire u2__abc_44228_n5179;
  wire u2__abc_44228_n5180;
  wire u2__abc_44228_n5181;
  wire u2__abc_44228_n5182_1;
  wire u2__abc_44228_n5183;
  wire u2__abc_44228_n5184;
  wire u2__abc_44228_n5185;
  wire u2__abc_44228_n5186;
  wire u2__abc_44228_n5187;
  wire u2__abc_44228_n5188;
  wire u2__abc_44228_n5189;
  wire u2__abc_44228_n5190;
  wire u2__abc_44228_n5191;
  wire u2__abc_44228_n5192_1;
  wire u2__abc_44228_n5193;
  wire u2__abc_44228_n5194;
  wire u2__abc_44228_n5195;
  wire u2__abc_44228_n5196;
  wire u2__abc_44228_n5197;
  wire u2__abc_44228_n5198;
  wire u2__abc_44228_n5199;
  wire u2__abc_44228_n5200;
  wire u2__abc_44228_n5201_1;
  wire u2__abc_44228_n5202;
  wire u2__abc_44228_n5203;
  wire u2__abc_44228_n5204;
  wire u2__abc_44228_n5205;
  wire u2__abc_44228_n5206;
  wire u2__abc_44228_n5207;
  wire u2__abc_44228_n5208;
  wire u2__abc_44228_n5209;
  wire u2__abc_44228_n5210;
  wire u2__abc_44228_n5211_1;
  wire u2__abc_44228_n5212;
  wire u2__abc_44228_n5213;
  wire u2__abc_44228_n5214;
  wire u2__abc_44228_n5215;
  wire u2__abc_44228_n5216;
  wire u2__abc_44228_n5217;
  wire u2__abc_44228_n5218;
  wire u2__abc_44228_n5219;
  wire u2__abc_44228_n5220;
  wire u2__abc_44228_n5221_1;
  wire u2__abc_44228_n5222;
  wire u2__abc_44228_n5223;
  wire u2__abc_44228_n5224;
  wire u2__abc_44228_n5225;
  wire u2__abc_44228_n5226;
  wire u2__abc_44228_n5227;
  wire u2__abc_44228_n5228;
  wire u2__abc_44228_n5229;
  wire u2__abc_44228_n5230_1;
  wire u2__abc_44228_n5231;
  wire u2__abc_44228_n5232;
  wire u2__abc_44228_n5233;
  wire u2__abc_44228_n5234;
  wire u2__abc_44228_n5235;
  wire u2__abc_44228_n5236;
  wire u2__abc_44228_n5237;
  wire u2__abc_44228_n5238;
  wire u2__abc_44228_n5239_1;
  wire u2__abc_44228_n5240;
  wire u2__abc_44228_n5241;
  wire u2__abc_44228_n5242;
  wire u2__abc_44228_n5243;
  wire u2__abc_44228_n5244;
  wire u2__abc_44228_n5245;
  wire u2__abc_44228_n5246;
  wire u2__abc_44228_n5247;
  wire u2__abc_44228_n5248;
  wire u2__abc_44228_n5249;
  wire u2__abc_44228_n5250_1;
  wire u2__abc_44228_n5251;
  wire u2__abc_44228_n5252;
  wire u2__abc_44228_n5253;
  wire u2__abc_44228_n5254;
  wire u2__abc_44228_n5255;
  wire u2__abc_44228_n5256;
  wire u2__abc_44228_n5257;
  wire u2__abc_44228_n5258;
  wire u2__abc_44228_n5259;
  wire u2__abc_44228_n5260_1;
  wire u2__abc_44228_n5261;
  wire u2__abc_44228_n5262;
  wire u2__abc_44228_n5263;
  wire u2__abc_44228_n5264;
  wire u2__abc_44228_n5265;
  wire u2__abc_44228_n5266;
  wire u2__abc_44228_n5267;
  wire u2__abc_44228_n5268;
  wire u2__abc_44228_n5269_1;
  wire u2__abc_44228_n5270;
  wire u2__abc_44228_n5271;
  wire u2__abc_44228_n5272;
  wire u2__abc_44228_n5273;
  wire u2__abc_44228_n5274;
  wire u2__abc_44228_n5275;
  wire u2__abc_44228_n5276;
  wire u2__abc_44228_n5277;
  wire u2__abc_44228_n5278_1;
  wire u2__abc_44228_n5279;
  wire u2__abc_44228_n5280;
  wire u2__abc_44228_n5281;
  wire u2__abc_44228_n5282;
  wire u2__abc_44228_n5283;
  wire u2__abc_44228_n5284;
  wire u2__abc_44228_n5285;
  wire u2__abc_44228_n5286;
  wire u2__abc_44228_n5287_1;
  wire u2__abc_44228_n5288;
  wire u2__abc_44228_n5289;
  wire u2__abc_44228_n5290;
  wire u2__abc_44228_n5291;
  wire u2__abc_44228_n5292;
  wire u2__abc_44228_n5293;
  wire u2__abc_44228_n5294;
  wire u2__abc_44228_n5295;
  wire u2__abc_44228_n5296;
  wire u2__abc_44228_n5297_1;
  wire u2__abc_44228_n5298;
  wire u2__abc_44228_n5299;
  wire u2__abc_44228_n5300;
  wire u2__abc_44228_n5301;
  wire u2__abc_44228_n5302;
  wire u2__abc_44228_n5303;
  wire u2__abc_44228_n5304;
  wire u2__abc_44228_n5305;
  wire u2__abc_44228_n5306_1;
  wire u2__abc_44228_n5307;
  wire u2__abc_44228_n5308;
  wire u2__abc_44228_n5309;
  wire u2__abc_44228_n5310;
  wire u2__abc_44228_n5311;
  wire u2__abc_44228_n5312;
  wire u2__abc_44228_n5313;
  wire u2__abc_44228_n5314;
  wire u2__abc_44228_n5315_1;
  wire u2__abc_44228_n5316;
  wire u2__abc_44228_n5317;
  wire u2__abc_44228_n5318;
  wire u2__abc_44228_n5319;
  wire u2__abc_44228_n5320;
  wire u2__abc_44228_n5321;
  wire u2__abc_44228_n5322;
  wire u2__abc_44228_n5323;
  wire u2__abc_44228_n5324_1;
  wire u2__abc_44228_n5325;
  wire u2__abc_44228_n5326;
  wire u2__abc_44228_n5327;
  wire u2__abc_44228_n5328;
  wire u2__abc_44228_n5329;
  wire u2__abc_44228_n5330;
  wire u2__abc_44228_n5331;
  wire u2__abc_44228_n5332;
  wire u2__abc_44228_n5333_1;
  wire u2__abc_44228_n5334;
  wire u2__abc_44228_n5335;
  wire u2__abc_44228_n5336;
  wire u2__abc_44228_n5337;
  wire u2__abc_44228_n5338;
  wire u2__abc_44228_n5339;
  wire u2__abc_44228_n5340;
  wire u2__abc_44228_n5341;
  wire u2__abc_44228_n5342;
  wire u2__abc_44228_n5343_1;
  wire u2__abc_44228_n5344;
  wire u2__abc_44228_n5345;
  wire u2__abc_44228_n5346;
  wire u2__abc_44228_n5347;
  wire u2__abc_44228_n5348;
  wire u2__abc_44228_n5349;
  wire u2__abc_44228_n5350;
  wire u2__abc_44228_n5351;
  wire u2__abc_44228_n5352_1;
  wire u2__abc_44228_n5353;
  wire u2__abc_44228_n5354;
  wire u2__abc_44228_n5355;
  wire u2__abc_44228_n5356;
  wire u2__abc_44228_n5357;
  wire u2__abc_44228_n5358;
  wire u2__abc_44228_n5359;
  wire u2__abc_44228_n5360;
  wire u2__abc_44228_n5361;
  wire u2__abc_44228_n5362_1;
  wire u2__abc_44228_n5363;
  wire u2__abc_44228_n5364;
  wire u2__abc_44228_n5365;
  wire u2__abc_44228_n5366;
  wire u2__abc_44228_n5367;
  wire u2__abc_44228_n5368;
  wire u2__abc_44228_n5369;
  wire u2__abc_44228_n5370;
  wire u2__abc_44228_n5371;
  wire u2__abc_44228_n5372_1;
  wire u2__abc_44228_n5373;
  wire u2__abc_44228_n5374;
  wire u2__abc_44228_n5375;
  wire u2__abc_44228_n5376;
  wire u2__abc_44228_n5377;
  wire u2__abc_44228_n5378;
  wire u2__abc_44228_n5379;
  wire u2__abc_44228_n5380;
  wire u2__abc_44228_n5381_1;
  wire u2__abc_44228_n5382;
  wire u2__abc_44228_n5383;
  wire u2__abc_44228_n5384;
  wire u2__abc_44228_n5385;
  wire u2__abc_44228_n5386;
  wire u2__abc_44228_n5387;
  wire u2__abc_44228_n5388;
  wire u2__abc_44228_n5389;
  wire u2__abc_44228_n5390_1;
  wire u2__abc_44228_n5391;
  wire u2__abc_44228_n5392;
  wire u2__abc_44228_n5393;
  wire u2__abc_44228_n5394;
  wire u2__abc_44228_n5395;
  wire u2__abc_44228_n5396;
  wire u2__abc_44228_n5397;
  wire u2__abc_44228_n5398;
  wire u2__abc_44228_n5399;
  wire u2__abc_44228_n5400_1;
  wire u2__abc_44228_n5401;
  wire u2__abc_44228_n5402;
  wire u2__abc_44228_n5403;
  wire u2__abc_44228_n5404;
  wire u2__abc_44228_n5405;
  wire u2__abc_44228_n5406;
  wire u2__abc_44228_n5407;
  wire u2__abc_44228_n5408;
  wire u2__abc_44228_n5409;
  wire u2__abc_44228_n5410_1;
  wire u2__abc_44228_n5411;
  wire u2__abc_44228_n5412;
  wire u2__abc_44228_n5413;
  wire u2__abc_44228_n5414;
  wire u2__abc_44228_n5415;
  wire u2__abc_44228_n5416;
  wire u2__abc_44228_n5417;
  wire u2__abc_44228_n5418;
  wire u2__abc_44228_n5419_1;
  wire u2__abc_44228_n5420;
  wire u2__abc_44228_n5421;
  wire u2__abc_44228_n5422;
  wire u2__abc_44228_n5423;
  wire u2__abc_44228_n5424;
  wire u2__abc_44228_n5425;
  wire u2__abc_44228_n5426;
  wire u2__abc_44228_n5427;
  wire u2__abc_44228_n5428_1;
  wire u2__abc_44228_n5429;
  wire u2__abc_44228_n5430;
  wire u2__abc_44228_n5431;
  wire u2__abc_44228_n5432;
  wire u2__abc_44228_n5433;
  wire u2__abc_44228_n5434;
  wire u2__abc_44228_n5435;
  wire u2__abc_44228_n5436;
  wire u2__abc_44228_n5437_1;
  wire u2__abc_44228_n5438;
  wire u2__abc_44228_n5439;
  wire u2__abc_44228_n5440;
  wire u2__abc_44228_n5441;
  wire u2__abc_44228_n5442;
  wire u2__abc_44228_n5443;
  wire u2__abc_44228_n5444;
  wire u2__abc_44228_n5445;
  wire u2__abc_44228_n5446;
  wire u2__abc_44228_n5447_1;
  wire u2__abc_44228_n5448;
  wire u2__abc_44228_n5449;
  wire u2__abc_44228_n5450;
  wire u2__abc_44228_n5451;
  wire u2__abc_44228_n5452;
  wire u2__abc_44228_n5453;
  wire u2__abc_44228_n5454;
  wire u2__abc_44228_n5455;
  wire u2__abc_44228_n5456_1;
  wire u2__abc_44228_n5457;
  wire u2__abc_44228_n5458;
  wire u2__abc_44228_n5459;
  wire u2__abc_44228_n5460;
  wire u2__abc_44228_n5461;
  wire u2__abc_44228_n5462;
  wire u2__abc_44228_n5463;
  wire u2__abc_44228_n5464;
  wire u2__abc_44228_n5465_1;
  wire u2__abc_44228_n5466;
  wire u2__abc_44228_n5467;
  wire u2__abc_44228_n5468;
  wire u2__abc_44228_n5469;
  wire u2__abc_44228_n5470;
  wire u2__abc_44228_n5471;
  wire u2__abc_44228_n5472;
  wire u2__abc_44228_n5473;
  wire u2__abc_44228_n5474_1;
  wire u2__abc_44228_n5475;
  wire u2__abc_44228_n5476;
  wire u2__abc_44228_n5477;
  wire u2__abc_44228_n5478;
  wire u2__abc_44228_n5479;
  wire u2__abc_44228_n5480;
  wire u2__abc_44228_n5481;
  wire u2__abc_44228_n5482;
  wire u2__abc_44228_n5483_1;
  wire u2__abc_44228_n5484;
  wire u2__abc_44228_n5485;
  wire u2__abc_44228_n5486;
  wire u2__abc_44228_n5487;
  wire u2__abc_44228_n5488;
  wire u2__abc_44228_n5489;
  wire u2__abc_44228_n5490;
  wire u2__abc_44228_n5491;
  wire u2__abc_44228_n5492;
  wire u2__abc_44228_n5493_1;
  wire u2__abc_44228_n5494;
  wire u2__abc_44228_n5495;
  wire u2__abc_44228_n5496;
  wire u2__abc_44228_n5497;
  wire u2__abc_44228_n5498;
  wire u2__abc_44228_n5499;
  wire u2__abc_44228_n5500;
  wire u2__abc_44228_n5501;
  wire u2__abc_44228_n5502_1;
  wire u2__abc_44228_n5503;
  wire u2__abc_44228_n5504;
  wire u2__abc_44228_n5505;
  wire u2__abc_44228_n5506;
  wire u2__abc_44228_n5507;
  wire u2__abc_44228_n5508;
  wire u2__abc_44228_n5509;
  wire u2__abc_44228_n5510;
  wire u2__abc_44228_n5511;
  wire u2__abc_44228_n5512_1;
  wire u2__abc_44228_n5513;
  wire u2__abc_44228_n5514;
  wire u2__abc_44228_n5515;
  wire u2__abc_44228_n5516;
  wire u2__abc_44228_n5517;
  wire u2__abc_44228_n5518;
  wire u2__abc_44228_n5519;
  wire u2__abc_44228_n5520;
  wire u2__abc_44228_n5521;
  wire u2__abc_44228_n5522_1;
  wire u2__abc_44228_n5523;
  wire u2__abc_44228_n5524;
  wire u2__abc_44228_n5525;
  wire u2__abc_44228_n5526;
  wire u2__abc_44228_n5527;
  wire u2__abc_44228_n5528;
  wire u2__abc_44228_n5529;
  wire u2__abc_44228_n5530;
  wire u2__abc_44228_n5531_1;
  wire u2__abc_44228_n5532;
  wire u2__abc_44228_n5533;
  wire u2__abc_44228_n5534;
  wire u2__abc_44228_n5535;
  wire u2__abc_44228_n5536;
  wire u2__abc_44228_n5537;
  wire u2__abc_44228_n5538;
  wire u2__abc_44228_n5539;
  wire u2__abc_44228_n5540_1;
  wire u2__abc_44228_n5541;
  wire u2__abc_44228_n5542;
  wire u2__abc_44228_n5543;
  wire u2__abc_44228_n5544;
  wire u2__abc_44228_n5545;
  wire u2__abc_44228_n5546;
  wire u2__abc_44228_n5547;
  wire u2__abc_44228_n5548;
  wire u2__abc_44228_n5549_1;
  wire u2__abc_44228_n5550;
  wire u2__abc_44228_n5551;
  wire u2__abc_44228_n5552;
  wire u2__abc_44228_n5553;
  wire u2__abc_44228_n5554;
  wire u2__abc_44228_n5555;
  wire u2__abc_44228_n5556;
  wire u2__abc_44228_n5557;
  wire u2__abc_44228_n5558_1;
  wire u2__abc_44228_n5559;
  wire u2__abc_44228_n5560;
  wire u2__abc_44228_n5561;
  wire u2__abc_44228_n5562;
  wire u2__abc_44228_n5563;
  wire u2__abc_44228_n5564;
  wire u2__abc_44228_n5565;
  wire u2__abc_44228_n5566;
  wire u2__abc_44228_n5567;
  wire u2__abc_44228_n5568_1;
  wire u2__abc_44228_n5569;
  wire u2__abc_44228_n5570;
  wire u2__abc_44228_n5571;
  wire u2__abc_44228_n5572;
  wire u2__abc_44228_n5573;
  wire u2__abc_44228_n5574;
  wire u2__abc_44228_n5575;
  wire u2__abc_44228_n5576;
  wire u2__abc_44228_n5577_1;
  wire u2__abc_44228_n5578;
  wire u2__abc_44228_n5579;
  wire u2__abc_44228_n5580;
  wire u2__abc_44228_n5581;
  wire u2__abc_44228_n5582;
  wire u2__abc_44228_n5583;
  wire u2__abc_44228_n5584;
  wire u2__abc_44228_n5585;
  wire u2__abc_44228_n5586;
  wire u2__abc_44228_n5587_1;
  wire u2__abc_44228_n5588;
  wire u2__abc_44228_n5589;
  wire u2__abc_44228_n5590;
  wire u2__abc_44228_n5591;
  wire u2__abc_44228_n5592;
  wire u2__abc_44228_n5593;
  wire u2__abc_44228_n5594;
  wire u2__abc_44228_n5595;
  wire u2__abc_44228_n5596;
  wire u2__abc_44228_n5597_1;
  wire u2__abc_44228_n5598;
  wire u2__abc_44228_n5599;
  wire u2__abc_44228_n5600;
  wire u2__abc_44228_n5601;
  wire u2__abc_44228_n5602;
  wire u2__abc_44228_n5603;
  wire u2__abc_44228_n5604;
  wire u2__abc_44228_n5605;
  wire u2__abc_44228_n5606_1;
  wire u2__abc_44228_n5607;
  wire u2__abc_44228_n5608;
  wire u2__abc_44228_n5609;
  wire u2__abc_44228_n5610;
  wire u2__abc_44228_n5611;
  wire u2__abc_44228_n5612;
  wire u2__abc_44228_n5613;
  wire u2__abc_44228_n5614;
  wire u2__abc_44228_n5615_1;
  wire u2__abc_44228_n5616;
  wire u2__abc_44228_n5617;
  wire u2__abc_44228_n5618;
  wire u2__abc_44228_n5619;
  wire u2__abc_44228_n5620;
  wire u2__abc_44228_n5621;
  wire u2__abc_44228_n5622;
  wire u2__abc_44228_n5623;
  wire u2__abc_44228_n5624_1;
  wire u2__abc_44228_n5625;
  wire u2__abc_44228_n5626;
  wire u2__abc_44228_n5627;
  wire u2__abc_44228_n5628;
  wire u2__abc_44228_n5629;
  wire u2__abc_44228_n5630;
  wire u2__abc_44228_n5631;
  wire u2__abc_44228_n5632;
  wire u2__abc_44228_n5633_1;
  wire u2__abc_44228_n5634;
  wire u2__abc_44228_n5635;
  wire u2__abc_44228_n5636;
  wire u2__abc_44228_n5637;
  wire u2__abc_44228_n5638;
  wire u2__abc_44228_n5639;
  wire u2__abc_44228_n5640;
  wire u2__abc_44228_n5641;
  wire u2__abc_44228_n5642;
  wire u2__abc_44228_n5643_1;
  wire u2__abc_44228_n5644;
  wire u2__abc_44228_n5645;
  wire u2__abc_44228_n5646;
  wire u2__abc_44228_n5647;
  wire u2__abc_44228_n5648;
  wire u2__abc_44228_n5649;
  wire u2__abc_44228_n5650;
  wire u2__abc_44228_n5651;
  wire u2__abc_44228_n5652_1;
  wire u2__abc_44228_n5653;
  wire u2__abc_44228_n5654;
  wire u2__abc_44228_n5655;
  wire u2__abc_44228_n5656;
  wire u2__abc_44228_n5657;
  wire u2__abc_44228_n5658;
  wire u2__abc_44228_n5659;
  wire u2__abc_44228_n5660;
  wire u2__abc_44228_n5661;
  wire u2__abc_44228_n5662_1;
  wire u2__abc_44228_n5663;
  wire u2__abc_44228_n5664;
  wire u2__abc_44228_n5665;
  wire u2__abc_44228_n5666;
  wire u2__abc_44228_n5667;
  wire u2__abc_44228_n5668;
  wire u2__abc_44228_n5669;
  wire u2__abc_44228_n5670;
  wire u2__abc_44228_n5671;
  wire u2__abc_44228_n5672_1;
  wire u2__abc_44228_n5673;
  wire u2__abc_44228_n5674;
  wire u2__abc_44228_n5675;
  wire u2__abc_44228_n5676;
  wire u2__abc_44228_n5677;
  wire u2__abc_44228_n5678;
  wire u2__abc_44228_n5679;
  wire u2__abc_44228_n5680;
  wire u2__abc_44228_n5681_1;
  wire u2__abc_44228_n5682;
  wire u2__abc_44228_n5683;
  wire u2__abc_44228_n5684;
  wire u2__abc_44228_n5685;
  wire u2__abc_44228_n5686;
  wire u2__abc_44228_n5687;
  wire u2__abc_44228_n5688;
  wire u2__abc_44228_n5689;
  wire u2__abc_44228_n5690_1;
  wire u2__abc_44228_n5691;
  wire u2__abc_44228_n5692;
  wire u2__abc_44228_n5693;
  wire u2__abc_44228_n5694;
  wire u2__abc_44228_n5695;
  wire u2__abc_44228_n5696;
  wire u2__abc_44228_n5697;
  wire u2__abc_44228_n5698;
  wire u2__abc_44228_n5699;
  wire u2__abc_44228_n5700_1;
  wire u2__abc_44228_n5701;
  wire u2__abc_44228_n5702;
  wire u2__abc_44228_n5703;
  wire u2__abc_44228_n5704;
  wire u2__abc_44228_n5705;
  wire u2__abc_44228_n5706;
  wire u2__abc_44228_n5707;
  wire u2__abc_44228_n5708;
  wire u2__abc_44228_n5709;
  wire u2__abc_44228_n5710_1;
  wire u2__abc_44228_n5711;
  wire u2__abc_44228_n5712;
  wire u2__abc_44228_n5713;
  wire u2__abc_44228_n5714;
  wire u2__abc_44228_n5715;
  wire u2__abc_44228_n5716;
  wire u2__abc_44228_n5717;
  wire u2__abc_44228_n5718;
  wire u2__abc_44228_n5719_1;
  wire u2__abc_44228_n5720;
  wire u2__abc_44228_n5721;
  wire u2__abc_44228_n5722;
  wire u2__abc_44228_n5723;
  wire u2__abc_44228_n5724;
  wire u2__abc_44228_n5725;
  wire u2__abc_44228_n5726;
  wire u2__abc_44228_n5727;
  wire u2__abc_44228_n5728_1;
  wire u2__abc_44228_n5729;
  wire u2__abc_44228_n5730;
  wire u2__abc_44228_n5731;
  wire u2__abc_44228_n5732;
  wire u2__abc_44228_n5733;
  wire u2__abc_44228_n5734;
  wire u2__abc_44228_n5735;
  wire u2__abc_44228_n5736;
  wire u2__abc_44228_n5737_1;
  wire u2__abc_44228_n5738;
  wire u2__abc_44228_n5739;
  wire u2__abc_44228_n5740;
  wire u2__abc_44228_n5741;
  wire u2__abc_44228_n5742;
  wire u2__abc_44228_n5743;
  wire u2__abc_44228_n5744;
  wire u2__abc_44228_n5745;
  wire u2__abc_44228_n5746;
  wire u2__abc_44228_n5747_1;
  wire u2__abc_44228_n5748;
  wire u2__abc_44228_n5749;
  wire u2__abc_44228_n5750;
  wire u2__abc_44228_n5751;
  wire u2__abc_44228_n5752;
  wire u2__abc_44228_n5753;
  wire u2__abc_44228_n5754;
  wire u2__abc_44228_n5755;
  wire u2__abc_44228_n5756_1;
  wire u2__abc_44228_n5757;
  wire u2__abc_44228_n5758;
  wire u2__abc_44228_n5759;
  wire u2__abc_44228_n5760;
  wire u2__abc_44228_n5761;
  wire u2__abc_44228_n5762;
  wire u2__abc_44228_n5763;
  wire u2__abc_44228_n5764;
  wire u2__abc_44228_n5765_1;
  wire u2__abc_44228_n5766;
  wire u2__abc_44228_n5767;
  wire u2__abc_44228_n5768;
  wire u2__abc_44228_n5769;
  wire u2__abc_44228_n5770;
  wire u2__abc_44228_n5771;
  wire u2__abc_44228_n5772;
  wire u2__abc_44228_n5773;
  wire u2__abc_44228_n5774_1;
  wire u2__abc_44228_n5775;
  wire u2__abc_44228_n5776;
  wire u2__abc_44228_n5777;
  wire u2__abc_44228_n5778;
  wire u2__abc_44228_n5779;
  wire u2__abc_44228_n5780;
  wire u2__abc_44228_n5781;
  wire u2__abc_44228_n5782;
  wire u2__abc_44228_n5783_1;
  wire u2__abc_44228_n5784;
  wire u2__abc_44228_n5785;
  wire u2__abc_44228_n5786;
  wire u2__abc_44228_n5787;
  wire u2__abc_44228_n5788;
  wire u2__abc_44228_n5789;
  wire u2__abc_44228_n5790;
  wire u2__abc_44228_n5791;
  wire u2__abc_44228_n5792;
  wire u2__abc_44228_n5793_1;
  wire u2__abc_44228_n5794;
  wire u2__abc_44228_n5795;
  wire u2__abc_44228_n5796;
  wire u2__abc_44228_n5797;
  wire u2__abc_44228_n5798;
  wire u2__abc_44228_n5799;
  wire u2__abc_44228_n5800;
  wire u2__abc_44228_n5801;
  wire u2__abc_44228_n5802_1;
  wire u2__abc_44228_n5803;
  wire u2__abc_44228_n5804;
  wire u2__abc_44228_n5805;
  wire u2__abc_44228_n5806;
  wire u2__abc_44228_n5807;
  wire u2__abc_44228_n5808;
  wire u2__abc_44228_n5809;
  wire u2__abc_44228_n5810;
  wire u2__abc_44228_n5811;
  wire u2__abc_44228_n5812_1;
  wire u2__abc_44228_n5813;
  wire u2__abc_44228_n5814;
  wire u2__abc_44228_n5815;
  wire u2__abc_44228_n5816;
  wire u2__abc_44228_n5817;
  wire u2__abc_44228_n5818;
  wire u2__abc_44228_n5819;
  wire u2__abc_44228_n5820;
  wire u2__abc_44228_n5821;
  wire u2__abc_44228_n5822_1;
  wire u2__abc_44228_n5823;
  wire u2__abc_44228_n5824;
  wire u2__abc_44228_n5825;
  wire u2__abc_44228_n5826;
  wire u2__abc_44228_n5827;
  wire u2__abc_44228_n5828;
  wire u2__abc_44228_n5829;
  wire u2__abc_44228_n5830_1;
  wire u2__abc_44228_n5831;
  wire u2__abc_44228_n5832;
  wire u2__abc_44228_n5833;
  wire u2__abc_44228_n5834;
  wire u2__abc_44228_n5835;
  wire u2__abc_44228_n5836;
  wire u2__abc_44228_n5837;
  wire u2__abc_44228_n5838_1;
  wire u2__abc_44228_n5839;
  wire u2__abc_44228_n5840;
  wire u2__abc_44228_n5841;
  wire u2__abc_44228_n5842;
  wire u2__abc_44228_n5843;
  wire u2__abc_44228_n5844;
  wire u2__abc_44228_n5845_1;
  wire u2__abc_44228_n5846;
  wire u2__abc_44228_n5847;
  wire u2__abc_44228_n5848;
  wire u2__abc_44228_n5849;
  wire u2__abc_44228_n5850;
  wire u2__abc_44228_n5851;
  wire u2__abc_44228_n5852;
  wire u2__abc_44228_n5853;
  wire u2__abc_44228_n5854_1;
  wire u2__abc_44228_n5855;
  wire u2__abc_44228_n5856;
  wire u2__abc_44228_n5857;
  wire u2__abc_44228_n5858;
  wire u2__abc_44228_n5859;
  wire u2__abc_44228_n5860;
  wire u2__abc_44228_n5861;
  wire u2__abc_44228_n5862;
  wire u2__abc_44228_n5863_1;
  wire u2__abc_44228_n5864;
  wire u2__abc_44228_n5865;
  wire u2__abc_44228_n5866;
  wire u2__abc_44228_n5867;
  wire u2__abc_44228_n5868;
  wire u2__abc_44228_n5869;
  wire u2__abc_44228_n5870;
  wire u2__abc_44228_n5871;
  wire u2__abc_44228_n5872;
  wire u2__abc_44228_n5873_1;
  wire u2__abc_44228_n5874;
  wire u2__abc_44228_n5875;
  wire u2__abc_44228_n5876;
  wire u2__abc_44228_n5877;
  wire u2__abc_44228_n5878;
  wire u2__abc_44228_n5879;
  wire u2__abc_44228_n5880;
  wire u2__abc_44228_n5881;
  wire u2__abc_44228_n5882;
  wire u2__abc_44228_n5883_1;
  wire u2__abc_44228_n5884;
  wire u2__abc_44228_n5885;
  wire u2__abc_44228_n5886;
  wire u2__abc_44228_n5887;
  wire u2__abc_44228_n5888;
  wire u2__abc_44228_n5889;
  wire u2__abc_44228_n5890;
  wire u2__abc_44228_n5891;
  wire u2__abc_44228_n5892_1;
  wire u2__abc_44228_n5893;
  wire u2__abc_44228_n5894;
  wire u2__abc_44228_n5895;
  wire u2__abc_44228_n5896;
  wire u2__abc_44228_n5897;
  wire u2__abc_44228_n5898;
  wire u2__abc_44228_n5899;
  wire u2__abc_44228_n5900;
  wire u2__abc_44228_n5901_1;
  wire u2__abc_44228_n5902;
  wire u2__abc_44228_n5903;
  wire u2__abc_44228_n5904;
  wire u2__abc_44228_n5905;
  wire u2__abc_44228_n5906;
  wire u2__abc_44228_n5907;
  wire u2__abc_44228_n5908;
  wire u2__abc_44228_n5909;
  wire u2__abc_44228_n5910;
  wire u2__abc_44228_n5911_1;
  wire u2__abc_44228_n5912;
  wire u2__abc_44228_n5913;
  wire u2__abc_44228_n5914;
  wire u2__abc_44228_n5915;
  wire u2__abc_44228_n5916;
  wire u2__abc_44228_n5917;
  wire u2__abc_44228_n5918;
  wire u2__abc_44228_n5919;
  wire u2__abc_44228_n5920_1;
  wire u2__abc_44228_n5921;
  wire u2__abc_44228_n5922;
  wire u2__abc_44228_n5923;
  wire u2__abc_44228_n5924;
  wire u2__abc_44228_n5925;
  wire u2__abc_44228_n5926;
  wire u2__abc_44228_n5927;
  wire u2__abc_44228_n5928;
  wire u2__abc_44228_n5929;
  wire u2__abc_44228_n5930_1;
  wire u2__abc_44228_n5931;
  wire u2__abc_44228_n5932;
  wire u2__abc_44228_n5933;
  wire u2__abc_44228_n5934;
  wire u2__abc_44228_n5935;
  wire u2__abc_44228_n5936;
  wire u2__abc_44228_n5937;
  wire u2__abc_44228_n5938_1;
  wire u2__abc_44228_n5939;
  wire u2__abc_44228_n5940;
  wire u2__abc_44228_n5941;
  wire u2__abc_44228_n5942;
  wire u2__abc_44228_n5943;
  wire u2__abc_44228_n5944;
  wire u2__abc_44228_n5945;
  wire u2__abc_44228_n5946;
  wire u2__abc_44228_n5947;
  wire u2__abc_44228_n5948_1;
  wire u2__abc_44228_n5949;
  wire u2__abc_44228_n5950;
  wire u2__abc_44228_n5951;
  wire u2__abc_44228_n5952;
  wire u2__abc_44228_n5953;
  wire u2__abc_44228_n5954;
  wire u2__abc_44228_n5955;
  wire u2__abc_44228_n5956;
  wire u2__abc_44228_n5957_1;
  wire u2__abc_44228_n5958;
  wire u2__abc_44228_n5959;
  wire u2__abc_44228_n5960;
  wire u2__abc_44228_n5961;
  wire u2__abc_44228_n5962;
  wire u2__abc_44228_n5963;
  wire u2__abc_44228_n5964;
  wire u2__abc_44228_n5965;
  wire u2__abc_44228_n5966_1;
  wire u2__abc_44228_n5967;
  wire u2__abc_44228_n5968;
  wire u2__abc_44228_n5969;
  wire u2__abc_44228_n5970;
  wire u2__abc_44228_n5971;
  wire u2__abc_44228_n5972;
  wire u2__abc_44228_n5973;
  wire u2__abc_44228_n5974;
  wire u2__abc_44228_n5975_1;
  wire u2__abc_44228_n5976;
  wire u2__abc_44228_n5977;
  wire u2__abc_44228_n5978;
  wire u2__abc_44228_n5979;
  wire u2__abc_44228_n5980;
  wire u2__abc_44228_n5981;
  wire u2__abc_44228_n5982;
  wire u2__abc_44228_n5983;
  wire u2__abc_44228_n5984;
  wire u2__abc_44228_n5985_1;
  wire u2__abc_44228_n5986;
  wire u2__abc_44228_n5987;
  wire u2__abc_44228_n5988;
  wire u2__abc_44228_n5989;
  wire u2__abc_44228_n5990;
  wire u2__abc_44228_n5991;
  wire u2__abc_44228_n5992;
  wire u2__abc_44228_n5993;
  wire u2__abc_44228_n5994_1;
  wire u2__abc_44228_n5995;
  wire u2__abc_44228_n5996;
  wire u2__abc_44228_n5997;
  wire u2__abc_44228_n5998;
  wire u2__abc_44228_n5999;
  wire u2__abc_44228_n6000;
  wire u2__abc_44228_n6001;
  wire u2__abc_44228_n6002;
  wire u2__abc_44228_n6003_1;
  wire u2__abc_44228_n6004;
  wire u2__abc_44228_n6005;
  wire u2__abc_44228_n6006;
  wire u2__abc_44228_n6007;
  wire u2__abc_44228_n6008;
  wire u2__abc_44228_n6009;
  wire u2__abc_44228_n6010;
  wire u2__abc_44228_n6011;
  wire u2__abc_44228_n6012_1;
  wire u2__abc_44228_n6013;
  wire u2__abc_44228_n6014;
  wire u2__abc_44228_n6015;
  wire u2__abc_44228_n6016;
  wire u2__abc_44228_n6017;
  wire u2__abc_44228_n6018;
  wire u2__abc_44228_n6019;
  wire u2__abc_44228_n6020;
  wire u2__abc_44228_n6021;
  wire u2__abc_44228_n6022_1;
  wire u2__abc_44228_n6023;
  wire u2__abc_44228_n6024;
  wire u2__abc_44228_n6025;
  wire u2__abc_44228_n6026;
  wire u2__abc_44228_n6027;
  wire u2__abc_44228_n6028;
  wire u2__abc_44228_n6029;
  wire u2__abc_44228_n6030;
  wire u2__abc_44228_n6031_1;
  wire u2__abc_44228_n6032;
  wire u2__abc_44228_n6033;
  wire u2__abc_44228_n6034;
  wire u2__abc_44228_n6035;
  wire u2__abc_44228_n6036;
  wire u2__abc_44228_n6037;
  wire u2__abc_44228_n6038;
  wire u2__abc_44228_n6039;
  wire u2__abc_44228_n6040_1;
  wire u2__abc_44228_n6041;
  wire u2__abc_44228_n6042;
  wire u2__abc_44228_n6043;
  wire u2__abc_44228_n6044;
  wire u2__abc_44228_n6045;
  wire u2__abc_44228_n6046;
  wire u2__abc_44228_n6047;
  wire u2__abc_44228_n6048;
  wire u2__abc_44228_n6049_1;
  wire u2__abc_44228_n6050;
  wire u2__abc_44228_n6051;
  wire u2__abc_44228_n6052;
  wire u2__abc_44228_n6053;
  wire u2__abc_44228_n6054;
  wire u2__abc_44228_n6055;
  wire u2__abc_44228_n6056;
  wire u2__abc_44228_n6057;
  wire u2__abc_44228_n6058;
  wire u2__abc_44228_n6059_1;
  wire u2__abc_44228_n6060;
  wire u2__abc_44228_n6061;
  wire u2__abc_44228_n6062;
  wire u2__abc_44228_n6063;
  wire u2__abc_44228_n6064;
  wire u2__abc_44228_n6065;
  wire u2__abc_44228_n6066;
  wire u2__abc_44228_n6067;
  wire u2__abc_44228_n6068_1;
  wire u2__abc_44228_n6069;
  wire u2__abc_44228_n6070;
  wire u2__abc_44228_n6071;
  wire u2__abc_44228_n6072;
  wire u2__abc_44228_n6073;
  wire u2__abc_44228_n6074;
  wire u2__abc_44228_n6075;
  wire u2__abc_44228_n6076;
  wire u2__abc_44228_n6077;
  wire u2__abc_44228_n6078_1;
  wire u2__abc_44228_n6079;
  wire u2__abc_44228_n6080;
  wire u2__abc_44228_n6081;
  wire u2__abc_44228_n6082;
  wire u2__abc_44228_n6083;
  wire u2__abc_44228_n6084;
  wire u2__abc_44228_n6085;
  wire u2__abc_44228_n6086_1;
  wire u2__abc_44228_n6087;
  wire u2__abc_44228_n6088;
  wire u2__abc_44228_n6089;
  wire u2__abc_44228_n6090;
  wire u2__abc_44228_n6091;
  wire u2__abc_44228_n6092;
  wire u2__abc_44228_n6093;
  wire u2__abc_44228_n6094;
  wire u2__abc_44228_n6095;
  wire u2__abc_44228_n6096_1;
  wire u2__abc_44228_n6097;
  wire u2__abc_44228_n6098;
  wire u2__abc_44228_n6099;
  wire u2__abc_44228_n6100;
  wire u2__abc_44228_n6101;
  wire u2__abc_44228_n6102;
  wire u2__abc_44228_n6103;
  wire u2__abc_44228_n6104_1;
  wire u2__abc_44228_n6105;
  wire u2__abc_44228_n6106;
  wire u2__abc_44228_n6107;
  wire u2__abc_44228_n6108;
  wire u2__abc_44228_n6109;
  wire u2__abc_44228_n6110;
  wire u2__abc_44228_n6111;
  wire u2__abc_44228_n6112;
  wire u2__abc_44228_n6113_1;
  wire u2__abc_44228_n6114;
  wire u2__abc_44228_n6115;
  wire u2__abc_44228_n6116;
  wire u2__abc_44228_n6117;
  wire u2__abc_44228_n6118;
  wire u2__abc_44228_n6119;
  wire u2__abc_44228_n6120;
  wire u2__abc_44228_n6121;
  wire u2__abc_44228_n6122_1;
  wire u2__abc_44228_n6123;
  wire u2__abc_44228_n6124;
  wire u2__abc_44228_n6125;
  wire u2__abc_44228_n6126;
  wire u2__abc_44228_n6127;
  wire u2__abc_44228_n6128;
  wire u2__abc_44228_n6129;
  wire u2__abc_44228_n6130;
  wire u2__abc_44228_n6131;
  wire u2__abc_44228_n6132_1;
  wire u2__abc_44228_n6133;
  wire u2__abc_44228_n6134;
  wire u2__abc_44228_n6135;
  wire u2__abc_44228_n6136;
  wire u2__abc_44228_n6137;
  wire u2__abc_44228_n6138;
  wire u2__abc_44228_n6139;
  wire u2__abc_44228_n6140;
  wire u2__abc_44228_n6141_1;
  wire u2__abc_44228_n6142;
  wire u2__abc_44228_n6143;
  wire u2__abc_44228_n6144;
  wire u2__abc_44228_n6145;
  wire u2__abc_44228_n6146;
  wire u2__abc_44228_n6147;
  wire u2__abc_44228_n6148;
  wire u2__abc_44228_n6149;
  wire u2__abc_44228_n6150;
  wire u2__abc_44228_n6151_1;
  wire u2__abc_44228_n6152;
  wire u2__abc_44228_n6153;
  wire u2__abc_44228_n6154;
  wire u2__abc_44228_n6155;
  wire u2__abc_44228_n6156;
  wire u2__abc_44228_n6157;
  wire u2__abc_44228_n6158;
  wire u2__abc_44228_n6159_1;
  wire u2__abc_44228_n6160;
  wire u2__abc_44228_n6161;
  wire u2__abc_44228_n6162;
  wire u2__abc_44228_n6163;
  wire u2__abc_44228_n6164;
  wire u2__abc_44228_n6165;
  wire u2__abc_44228_n6166;
  wire u2__abc_44228_n6167;
  wire u2__abc_44228_n6168;
  wire u2__abc_44228_n6169_1;
  wire u2__abc_44228_n6170;
  wire u2__abc_44228_n6171;
  wire u2__abc_44228_n6172;
  wire u2__abc_44228_n6173;
  wire u2__abc_44228_n6174;
  wire u2__abc_44228_n6175;
  wire u2__abc_44228_n6176;
  wire u2__abc_44228_n6177;
  wire u2__abc_44228_n6178_1;
  wire u2__abc_44228_n6179;
  wire u2__abc_44228_n6180;
  wire u2__abc_44228_n6181;
  wire u2__abc_44228_n6182;
  wire u2__abc_44228_n6183;
  wire u2__abc_44228_n6184;
  wire u2__abc_44228_n6185;
  wire u2__abc_44228_n6186;
  wire u2__abc_44228_n6187_1;
  wire u2__abc_44228_n6188;
  wire u2__abc_44228_n6189;
  wire u2__abc_44228_n6190;
  wire u2__abc_44228_n6191;
  wire u2__abc_44228_n6192;
  wire u2__abc_44228_n6193;
  wire u2__abc_44228_n6194;
  wire u2__abc_44228_n6195;
  wire u2__abc_44228_n6196_1;
  wire u2__abc_44228_n6197;
  wire u2__abc_44228_n6198;
  wire u2__abc_44228_n6199;
  wire u2__abc_44228_n6200;
  wire u2__abc_44228_n6201;
  wire u2__abc_44228_n6202;
  wire u2__abc_44228_n6203;
  wire u2__abc_44228_n6204;
  wire u2__abc_44228_n6205;
  wire u2__abc_44228_n6206_1;
  wire u2__abc_44228_n6207;
  wire u2__abc_44228_n6208;
  wire u2__abc_44228_n6209;
  wire u2__abc_44228_n6210;
  wire u2__abc_44228_n6211;
  wire u2__abc_44228_n6212;
  wire u2__abc_44228_n6213;
  wire u2__abc_44228_n6214_1;
  wire u2__abc_44228_n6215;
  wire u2__abc_44228_n6216;
  wire u2__abc_44228_n6217;
  wire u2__abc_44228_n6218;
  wire u2__abc_44228_n6219;
  wire u2__abc_44228_n6220;
  wire u2__abc_44228_n6221;
  wire u2__abc_44228_n6222;
  wire u2__abc_44228_n6223;
  wire u2__abc_44228_n6224_1;
  wire u2__abc_44228_n6225;
  wire u2__abc_44228_n6226;
  wire u2__abc_44228_n6227;
  wire u2__abc_44228_n6228;
  wire u2__abc_44228_n6229;
  wire u2__abc_44228_n6230;
  wire u2__abc_44228_n6231;
  wire u2__abc_44228_n6232_1;
  wire u2__abc_44228_n6233;
  wire u2__abc_44228_n6234;
  wire u2__abc_44228_n6235;
  wire u2__abc_44228_n6236;
  wire u2__abc_44228_n6237;
  wire u2__abc_44228_n6238;
  wire u2__abc_44228_n6239;
  wire u2__abc_44228_n6240;
  wire u2__abc_44228_n6241;
  wire u2__abc_44228_n6242_1;
  wire u2__abc_44228_n6243;
  wire u2__abc_44228_n6244;
  wire u2__abc_44228_n6245;
  wire u2__abc_44228_n6246;
  wire u2__abc_44228_n6247;
  wire u2__abc_44228_n6248;
  wire u2__abc_44228_n6249;
  wire u2__abc_44228_n6250;
  wire u2__abc_44228_n6251_1;
  wire u2__abc_44228_n6252;
  wire u2__abc_44228_n6253;
  wire u2__abc_44228_n6254;
  wire u2__abc_44228_n6255;
  wire u2__abc_44228_n6256;
  wire u2__abc_44228_n6257;
  wire u2__abc_44228_n6258;
  wire u2__abc_44228_n6259;
  wire u2__abc_44228_n6260_1;
  wire u2__abc_44228_n6261;
  wire u2__abc_44228_n6262;
  wire u2__abc_44228_n6263;
  wire u2__abc_44228_n6264;
  wire u2__abc_44228_n6265;
  wire u2__abc_44228_n6266;
  wire u2__abc_44228_n6267;
  wire u2__abc_44228_n6268;
  wire u2__abc_44228_n6269_1;
  wire u2__abc_44228_n6270;
  wire u2__abc_44228_n6271;
  wire u2__abc_44228_n6272;
  wire u2__abc_44228_n6273;
  wire u2__abc_44228_n6274;
  wire u2__abc_44228_n6275;
  wire u2__abc_44228_n6276;
  wire u2__abc_44228_n6277;
  wire u2__abc_44228_n6278;
  wire u2__abc_44228_n6279_1;
  wire u2__abc_44228_n6280;
  wire u2__abc_44228_n6281;
  wire u2__abc_44228_n6282;
  wire u2__abc_44228_n6283;
  wire u2__abc_44228_n6284;
  wire u2__abc_44228_n6285;
  wire u2__abc_44228_n6286;
  wire u2__abc_44228_n6287_1;
  wire u2__abc_44228_n6288;
  wire u2__abc_44228_n6289;
  wire u2__abc_44228_n6290;
  wire u2__abc_44228_n6291;
  wire u2__abc_44228_n6292;
  wire u2__abc_44228_n6293;
  wire u2__abc_44228_n6294;
  wire u2__abc_44228_n6295;
  wire u2__abc_44228_n6296_1;
  wire u2__abc_44228_n6297;
  wire u2__abc_44228_n6298;
  wire u2__abc_44228_n6299;
  wire u2__abc_44228_n6300;
  wire u2__abc_44228_n6301;
  wire u2__abc_44228_n6302;
  wire u2__abc_44228_n6303;
  wire u2__abc_44228_n6304;
  wire u2__abc_44228_n6305_1;
  wire u2__abc_44228_n6306;
  wire u2__abc_44228_n6307;
  wire u2__abc_44228_n6308;
  wire u2__abc_44228_n6309;
  wire u2__abc_44228_n6310;
  wire u2__abc_44228_n6311;
  wire u2__abc_44228_n6312;
  wire u2__abc_44228_n6313;
  wire u2__abc_44228_n6314;
  wire u2__abc_44228_n6315_1;
  wire u2__abc_44228_n6316;
  wire u2__abc_44228_n6317;
  wire u2__abc_44228_n6318;
  wire u2__abc_44228_n6319;
  wire u2__abc_44228_n6320;
  wire u2__abc_44228_n6321;
  wire u2__abc_44228_n6322;
  wire u2__abc_44228_n6323;
  wire u2__abc_44228_n6324_1;
  wire u2__abc_44228_n6325;
  wire u2__abc_44228_n6326;
  wire u2__abc_44228_n6327;
  wire u2__abc_44228_n6328;
  wire u2__abc_44228_n6329;
  wire u2__abc_44228_n6330;
  wire u2__abc_44228_n6331;
  wire u2__abc_44228_n6332;
  wire u2__abc_44228_n6333_1;
  wire u2__abc_44228_n6334;
  wire u2__abc_44228_n6335;
  wire u2__abc_44228_n6336;
  wire u2__abc_44228_n6337;
  wire u2__abc_44228_n6338;
  wire u2__abc_44228_n6339;
  wire u2__abc_44228_n6340;
  wire u2__abc_44228_n6341;
  wire u2__abc_44228_n6342_1;
  wire u2__abc_44228_n6343;
  wire u2__abc_44228_n6344;
  wire u2__abc_44228_n6345;
  wire u2__abc_44228_n6346;
  wire u2__abc_44228_n6347;
  wire u2__abc_44228_n6348;
  wire u2__abc_44228_n6349;
  wire u2__abc_44228_n6350;
  wire u2__abc_44228_n6351;
  wire u2__abc_44228_n6352_1;
  wire u2__abc_44228_n6353;
  wire u2__abc_44228_n6354;
  wire u2__abc_44228_n6355;
  wire u2__abc_44228_n6356;
  wire u2__abc_44228_n6357;
  wire u2__abc_44228_n6358;
  wire u2__abc_44228_n6359;
  wire u2__abc_44228_n6360;
  wire u2__abc_44228_n6361_1;
  wire u2__abc_44228_n6362;
  wire u2__abc_44228_n6363;
  wire u2__abc_44228_n6364;
  wire u2__abc_44228_n6365;
  wire u2__abc_44228_n6366;
  wire u2__abc_44228_n6367;
  wire u2__abc_44228_n6368;
  wire u2__abc_44228_n6369;
  wire u2__abc_44228_n6370;
  wire u2__abc_44228_n6371_1;
  wire u2__abc_44228_n6372;
  wire u2__abc_44228_n6373;
  wire u2__abc_44228_n6374;
  wire u2__abc_44228_n6375;
  wire u2__abc_44228_n6376;
  wire u2__abc_44228_n6377;
  wire u2__abc_44228_n6378;
  wire u2__abc_44228_n6379_1;
  wire u2__abc_44228_n6380;
  wire u2__abc_44228_n6381;
  wire u2__abc_44228_n6382;
  wire u2__abc_44228_n6383;
  wire u2__abc_44228_n6384;
  wire u2__abc_44228_n6385;
  wire u2__abc_44228_n6386;
  wire u2__abc_44228_n6387;
  wire u2__abc_44228_n6388;
  wire u2__abc_44228_n6389_1;
  wire u2__abc_44228_n6390;
  wire u2__abc_44228_n6391;
  wire u2__abc_44228_n6392;
  wire u2__abc_44228_n6393;
  wire u2__abc_44228_n6394;
  wire u2__abc_44228_n6395;
  wire u2__abc_44228_n6396;
  wire u2__abc_44228_n6397_1;
  wire u2__abc_44228_n6398;
  wire u2__abc_44228_n6399;
  wire u2__abc_44228_n6400;
  wire u2__abc_44228_n6401;
  wire u2__abc_44228_n6402;
  wire u2__abc_44228_n6403;
  wire u2__abc_44228_n6404;
  wire u2__abc_44228_n6405;
  wire u2__abc_44228_n6406_1;
  wire u2__abc_44228_n6407;
  wire u2__abc_44228_n6408;
  wire u2__abc_44228_n6409;
  wire u2__abc_44228_n6410;
  wire u2__abc_44228_n6411;
  wire u2__abc_44228_n6412;
  wire u2__abc_44228_n6413;
  wire u2__abc_44228_n6414;
  wire u2__abc_44228_n6415_1;
  wire u2__abc_44228_n6416;
  wire u2__abc_44228_n6417;
  wire u2__abc_44228_n6418;
  wire u2__abc_44228_n6419;
  wire u2__abc_44228_n6420;
  wire u2__abc_44228_n6421;
  wire u2__abc_44228_n6422;
  wire u2__abc_44228_n6423;
  wire u2__abc_44228_n6424;
  wire u2__abc_44228_n6425_1;
  wire u2__abc_44228_n6426;
  wire u2__abc_44228_n6427;
  wire u2__abc_44228_n6428;
  wire u2__abc_44228_n6429;
  wire u2__abc_44228_n6430;
  wire u2__abc_44228_n6431;
  wire u2__abc_44228_n6432;
  wire u2__abc_44228_n6433;
  wire u2__abc_44228_n6434;
  wire u2__abc_44228_n6435_1;
  wire u2__abc_44228_n6436;
  wire u2__abc_44228_n6437;
  wire u2__abc_44228_n6438;
  wire u2__abc_44228_n6439;
  wire u2__abc_44228_n6440;
  wire u2__abc_44228_n6441;
  wire u2__abc_44228_n6442;
  wire u2__abc_44228_n6443;
  wire u2__abc_44228_n6444;
  wire u2__abc_44228_n6445_1;
  wire u2__abc_44228_n6446;
  wire u2__abc_44228_n6447;
  wire u2__abc_44228_n6448;
  wire u2__abc_44228_n6449;
  wire u2__abc_44228_n6450;
  wire u2__abc_44228_n6451;
  wire u2__abc_44228_n6452;
  wire u2__abc_44228_n6453_1;
  wire u2__abc_44228_n6454;
  wire u2__abc_44228_n6455;
  wire u2__abc_44228_n6456;
  wire u2__abc_44228_n6457;
  wire u2__abc_44228_n6458;
  wire u2__abc_44228_n6459;
  wire u2__abc_44228_n6460;
  wire u2__abc_44228_n6461;
  wire u2__abc_44228_n6462;
  wire u2__abc_44228_n6463_1;
  wire u2__abc_44228_n6464;
  wire u2__abc_44228_n6465;
  wire u2__abc_44228_n6466;
  wire u2__abc_44228_n6467;
  wire u2__abc_44228_n6468;
  wire u2__abc_44228_n6469;
  wire u2__abc_44228_n6470;
  wire u2__abc_44228_n6471_1;
  wire u2__abc_44228_n6472;
  wire u2__abc_44228_n6473;
  wire u2__abc_44228_n6474;
  wire u2__abc_44228_n6475;
  wire u2__abc_44228_n6476;
  wire u2__abc_44228_n6477;
  wire u2__abc_44228_n6478;
  wire u2__abc_44228_n6479;
  wire u2__abc_44228_n6480_1;
  wire u2__abc_44228_n6481;
  wire u2__abc_44228_n6482;
  wire u2__abc_44228_n6483;
  wire u2__abc_44228_n6484;
  wire u2__abc_44228_n6485;
  wire u2__abc_44228_n6486;
  wire u2__abc_44228_n6487;
  wire u2__abc_44228_n6488;
  wire u2__abc_44228_n6489_1;
  wire u2__abc_44228_n6490;
  wire u2__abc_44228_n6491;
  wire u2__abc_44228_n6492;
  wire u2__abc_44228_n6493;
  wire u2__abc_44228_n6494;
  wire u2__abc_44228_n6495;
  wire u2__abc_44228_n6496;
  wire u2__abc_44228_n6497;
  wire u2__abc_44228_n6498;
  wire u2__abc_44228_n6499_1;
  wire u2__abc_44228_n6500;
  wire u2__abc_44228_n6501;
  wire u2__abc_44228_n6502;
  wire u2__abc_44228_n6503;
  wire u2__abc_44228_n6504;
  wire u2__abc_44228_n6505;
  wire u2__abc_44228_n6506;
  wire u2__abc_44228_n6507_1;
  wire u2__abc_44228_n6508;
  wire u2__abc_44228_n6509;
  wire u2__abc_44228_n6510;
  wire u2__abc_44228_n6511;
  wire u2__abc_44228_n6512;
  wire u2__abc_44228_n6513;
  wire u2__abc_44228_n6514;
  wire u2__abc_44228_n6515;
  wire u2__abc_44228_n6516;
  wire u2__abc_44228_n6517_1;
  wire u2__abc_44228_n6518;
  wire u2__abc_44228_n6519;
  wire u2__abc_44228_n6520;
  wire u2__abc_44228_n6521;
  wire u2__abc_44228_n6522;
  wire u2__abc_44228_n6523;
  wire u2__abc_44228_n6524;
  wire u2__abc_44228_n6525_1;
  wire u2__abc_44228_n6526;
  wire u2__abc_44228_n6527;
  wire u2__abc_44228_n6528;
  wire u2__abc_44228_n6529;
  wire u2__abc_44228_n6530;
  wire u2__abc_44228_n6531;
  wire u2__abc_44228_n6532;
  wire u2__abc_44228_n6533;
  wire u2__abc_44228_n6534;
  wire u2__abc_44228_n6535_1;
  wire u2__abc_44228_n6536;
  wire u2__abc_44228_n6537;
  wire u2__abc_44228_n6538;
  wire u2__abc_44228_n6539;
  wire u2__abc_44228_n6540;
  wire u2__abc_44228_n6541;
  wire u2__abc_44228_n6542;
  wire u2__abc_44228_n6543_1;
  wire u2__abc_44228_n6544;
  wire u2__abc_44228_n6545;
  wire u2__abc_44228_n6546;
  wire u2__abc_44228_n6547;
  wire u2__abc_44228_n6548;
  wire u2__abc_44228_n6549;
  wire u2__abc_44228_n6550;
  wire u2__abc_44228_n6551;
  wire u2__abc_44228_n6552_1;
  wire u2__abc_44228_n6553;
  wire u2__abc_44228_n6554;
  wire u2__abc_44228_n6555;
  wire u2__abc_44228_n6556;
  wire u2__abc_44228_n6557;
  wire u2__abc_44228_n6558;
  wire u2__abc_44228_n6559;
  wire u2__abc_44228_n6560;
  wire u2__abc_44228_n6561_1;
  wire u2__abc_44228_n6562;
  wire u2__abc_44228_n6563;
  wire u2__abc_44228_n6564;
  wire u2__abc_44228_n6565;
  wire u2__abc_44228_n6566;
  wire u2__abc_44228_n6567;
  wire u2__abc_44228_n6568;
  wire u2__abc_44228_n6569;
  wire u2__abc_44228_n6570;
  wire u2__abc_44228_n6571_1;
  wire u2__abc_44228_n6572;
  wire u2__abc_44228_n6573;
  wire u2__abc_44228_n6574;
  wire u2__abc_44228_n6575;
  wire u2__abc_44228_n6576;
  wire u2__abc_44228_n6577;
  wire u2__abc_44228_n6578;
  wire u2__abc_44228_n6579_1;
  wire u2__abc_44228_n6580;
  wire u2__abc_44228_n6581;
  wire u2__abc_44228_n6582;
  wire u2__abc_44228_n6583;
  wire u2__abc_44228_n6584;
  wire u2__abc_44228_n6585;
  wire u2__abc_44228_n6586;
  wire u2__abc_44228_n6587;
  wire u2__abc_44228_n6588_1;
  wire u2__abc_44228_n6589;
  wire u2__abc_44228_n6590;
  wire u2__abc_44228_n6591;
  wire u2__abc_44228_n6592;
  wire u2__abc_44228_n6593;
  wire u2__abc_44228_n6594;
  wire u2__abc_44228_n6595;
  wire u2__abc_44228_n6596;
  wire u2__abc_44228_n6597_1;
  wire u2__abc_44228_n6598;
  wire u2__abc_44228_n6599;
  wire u2__abc_44228_n6600;
  wire u2__abc_44228_n6601;
  wire u2__abc_44228_n6602;
  wire u2__abc_44228_n6603;
  wire u2__abc_44228_n6604;
  wire u2__abc_44228_n6605;
  wire u2__abc_44228_n6606;
  wire u2__abc_44228_n6607_1;
  wire u2__abc_44228_n6608;
  wire u2__abc_44228_n6609;
  wire u2__abc_44228_n6610;
  wire u2__abc_44228_n6611;
  wire u2__abc_44228_n6612;
  wire u2__abc_44228_n6613;
  wire u2__abc_44228_n6614;
  wire u2__abc_44228_n6615;
  wire u2__abc_44228_n6616_1;
  wire u2__abc_44228_n6617;
  wire u2__abc_44228_n6618;
  wire u2__abc_44228_n6619;
  wire u2__abc_44228_n6620;
  wire u2__abc_44228_n6621;
  wire u2__abc_44228_n6622;
  wire u2__abc_44228_n6623;
  wire u2__abc_44228_n6624;
  wire u2__abc_44228_n6625_1;
  wire u2__abc_44228_n6626;
  wire u2__abc_44228_n6627;
  wire u2__abc_44228_n6628;
  wire u2__abc_44228_n6629;
  wire u2__abc_44228_n6630;
  wire u2__abc_44228_n6631;
  wire u2__abc_44228_n6632;
  wire u2__abc_44228_n6633;
  wire u2__abc_44228_n6634_1;
  wire u2__abc_44228_n6635;
  wire u2__abc_44228_n6636;
  wire u2__abc_44228_n6637;
  wire u2__abc_44228_n6638;
  wire u2__abc_44228_n6639;
  wire u2__abc_44228_n6640;
  wire u2__abc_44228_n6641;
  wire u2__abc_44228_n6642;
  wire u2__abc_44228_n6643;
  wire u2__abc_44228_n6644_1;
  wire u2__abc_44228_n6645;
  wire u2__abc_44228_n6646;
  wire u2__abc_44228_n6647;
  wire u2__abc_44228_n6648;
  wire u2__abc_44228_n6649;
  wire u2__abc_44228_n6650;
  wire u2__abc_44228_n6651;
  wire u2__abc_44228_n6652;
  wire u2__abc_44228_n6653_1;
  wire u2__abc_44228_n6654;
  wire u2__abc_44228_n6655;
  wire u2__abc_44228_n6656;
  wire u2__abc_44228_n6657;
  wire u2__abc_44228_n6658;
  wire u2__abc_44228_n6659;
  wire u2__abc_44228_n6660;
  wire u2__abc_44228_n6661;
  wire u2__abc_44228_n6662;
  wire u2__abc_44228_n6663_1;
  wire u2__abc_44228_n6664;
  wire u2__abc_44228_n6665;
  wire u2__abc_44228_n6666;
  wire u2__abc_44228_n6667;
  wire u2__abc_44228_n6668;
  wire u2__abc_44228_n6669;
  wire u2__abc_44228_n6670;
  wire u2__abc_44228_n6671_1;
  wire u2__abc_44228_n6672;
  wire u2__abc_44228_n6673;
  wire u2__abc_44228_n6674;
  wire u2__abc_44228_n6675;
  wire u2__abc_44228_n6676;
  wire u2__abc_44228_n6677;
  wire u2__abc_44228_n6678;
  wire u2__abc_44228_n6679;
  wire u2__abc_44228_n6680;
  wire u2__abc_44228_n6681_1;
  wire u2__abc_44228_n6682;
  wire u2__abc_44228_n6683;
  wire u2__abc_44228_n6684;
  wire u2__abc_44228_n6685;
  wire u2__abc_44228_n6686;
  wire u2__abc_44228_n6687;
  wire u2__abc_44228_n6688;
  wire u2__abc_44228_n6689_1;
  wire u2__abc_44228_n6690;
  wire u2__abc_44228_n6691;
  wire u2__abc_44228_n6692;
  wire u2__abc_44228_n6693;
  wire u2__abc_44228_n6694;
  wire u2__abc_44228_n6695;
  wire u2__abc_44228_n6696;
  wire u2__abc_44228_n6697;
  wire u2__abc_44228_n6698_1;
  wire u2__abc_44228_n6699;
  wire u2__abc_44228_n6700;
  wire u2__abc_44228_n6701;
  wire u2__abc_44228_n6702;
  wire u2__abc_44228_n6703;
  wire u2__abc_44228_n6704;
  wire u2__abc_44228_n6705;
  wire u2__abc_44228_n6706;
  wire u2__abc_44228_n6707_1;
  wire u2__abc_44228_n6708;
  wire u2__abc_44228_n6709;
  wire u2__abc_44228_n6710;
  wire u2__abc_44228_n6711;
  wire u2__abc_44228_n6712;
  wire u2__abc_44228_n6713;
  wire u2__abc_44228_n6714;
  wire u2__abc_44228_n6715;
  wire u2__abc_44228_n6716;
  wire u2__abc_44228_n6717_1;
  wire u2__abc_44228_n6718;
  wire u2__abc_44228_n6719;
  wire u2__abc_44228_n6720;
  wire u2__abc_44228_n6721;
  wire u2__abc_44228_n6722;
  wire u2__abc_44228_n6723;
  wire u2__abc_44228_n6724;
  wire u2__abc_44228_n6725_1;
  wire u2__abc_44228_n6726;
  wire u2__abc_44228_n6727;
  wire u2__abc_44228_n6728;
  wire u2__abc_44228_n6729;
  wire u2__abc_44228_n6730;
  wire u2__abc_44228_n6731;
  wire u2__abc_44228_n6732;
  wire u2__abc_44228_n6733;
  wire u2__abc_44228_n6734;
  wire u2__abc_44228_n6735_1;
  wire u2__abc_44228_n6736;
  wire u2__abc_44228_n6737;
  wire u2__abc_44228_n6738;
  wire u2__abc_44228_n6739;
  wire u2__abc_44228_n6740;
  wire u2__abc_44228_n6741;
  wire u2__abc_44228_n6742;
  wire u2__abc_44228_n6743_1;
  wire u2__abc_44228_n6744;
  wire u2__abc_44228_n6745;
  wire u2__abc_44228_n6746;
  wire u2__abc_44228_n6747;
  wire u2__abc_44228_n6748;
  wire u2__abc_44228_n6749;
  wire u2__abc_44228_n6750;
  wire u2__abc_44228_n6751;
  wire u2__abc_44228_n6752;
  wire u2__abc_44228_n6753_1;
  wire u2__abc_44228_n6754;
  wire u2__abc_44228_n6755;
  wire u2__abc_44228_n6756;
  wire u2__abc_44228_n6757;
  wire u2__abc_44228_n6758;
  wire u2__abc_44228_n6759;
  wire u2__abc_44228_n6760;
  wire u2__abc_44228_n6761_1;
  wire u2__abc_44228_n6762;
  wire u2__abc_44228_n6763;
  wire u2__abc_44228_n6764;
  wire u2__abc_44228_n6765;
  wire u2__abc_44228_n6766;
  wire u2__abc_44228_n6767;
  wire u2__abc_44228_n6768;
  wire u2__abc_44228_n6769;
  wire u2__abc_44228_n6770_1;
  wire u2__abc_44228_n6771;
  wire u2__abc_44228_n6772;
  wire u2__abc_44228_n6773;
  wire u2__abc_44228_n6774;
  wire u2__abc_44228_n6775;
  wire u2__abc_44228_n6776;
  wire u2__abc_44228_n6777;
  wire u2__abc_44228_n6778;
  wire u2__abc_44228_n6779_1;
  wire u2__abc_44228_n6780;
  wire u2__abc_44228_n6781;
  wire u2__abc_44228_n6782;
  wire u2__abc_44228_n6783;
  wire u2__abc_44228_n6784;
  wire u2__abc_44228_n6785;
  wire u2__abc_44228_n6786;
  wire u2__abc_44228_n6787;
  wire u2__abc_44228_n6788;
  wire u2__abc_44228_n6789_1;
  wire u2__abc_44228_n6790;
  wire u2__abc_44228_n6791;
  wire u2__abc_44228_n6792;
  wire u2__abc_44228_n6793;
  wire u2__abc_44228_n6794;
  wire u2__abc_44228_n6795;
  wire u2__abc_44228_n6796;
  wire u2__abc_44228_n6797_1;
  wire u2__abc_44228_n6798;
  wire u2__abc_44228_n6799;
  wire u2__abc_44228_n6800;
  wire u2__abc_44228_n6801;
  wire u2__abc_44228_n6802;
  wire u2__abc_44228_n6803;
  wire u2__abc_44228_n6804;
  wire u2__abc_44228_n6805;
  wire u2__abc_44228_n6806;
  wire u2__abc_44228_n6807_1;
  wire u2__abc_44228_n6808;
  wire u2__abc_44228_n6809;
  wire u2__abc_44228_n6810;
  wire u2__abc_44228_n6811;
  wire u2__abc_44228_n6812;
  wire u2__abc_44228_n6813;
  wire u2__abc_44228_n6814;
  wire u2__abc_44228_n6815_1;
  wire u2__abc_44228_n6816;
  wire u2__abc_44228_n6817;
  wire u2__abc_44228_n6818;
  wire u2__abc_44228_n6819;
  wire u2__abc_44228_n6820;
  wire u2__abc_44228_n6821;
  wire u2__abc_44228_n6822;
  wire u2__abc_44228_n6823;
  wire u2__abc_44228_n6824;
  wire u2__abc_44228_n6825_1;
  wire u2__abc_44228_n6826;
  wire u2__abc_44228_n6827;
  wire u2__abc_44228_n6828;
  wire u2__abc_44228_n6829;
  wire u2__abc_44228_n6830;
  wire u2__abc_44228_n6831;
  wire u2__abc_44228_n6832;
  wire u2__abc_44228_n6833_1;
  wire u2__abc_44228_n6834;
  wire u2__abc_44228_n6835;
  wire u2__abc_44228_n6836;
  wire u2__abc_44228_n6837;
  wire u2__abc_44228_n6838;
  wire u2__abc_44228_n6839;
  wire u2__abc_44228_n6840;
  wire u2__abc_44228_n6841;
  wire u2__abc_44228_n6842_1;
  wire u2__abc_44228_n6843;
  wire u2__abc_44228_n6844;
  wire u2__abc_44228_n6845;
  wire u2__abc_44228_n6846;
  wire u2__abc_44228_n6847;
  wire u2__abc_44228_n6848;
  wire u2__abc_44228_n6849;
  wire u2__abc_44228_n6850;
  wire u2__abc_44228_n6851_1;
  wire u2__abc_44228_n6852;
  wire u2__abc_44228_n6853;
  wire u2__abc_44228_n6854;
  wire u2__abc_44228_n6855;
  wire u2__abc_44228_n6856;
  wire u2__abc_44228_n6857;
  wire u2__abc_44228_n6858;
  wire u2__abc_44228_n6859;
  wire u2__abc_44228_n6860;
  wire u2__abc_44228_n6861_1;
  wire u2__abc_44228_n6862;
  wire u2__abc_44228_n6863;
  wire u2__abc_44228_n6864;
  wire u2__abc_44228_n6865;
  wire u2__abc_44228_n6866;
  wire u2__abc_44228_n6867;
  wire u2__abc_44228_n6868;
  wire u2__abc_44228_n6869_1;
  wire u2__abc_44228_n6870;
  wire u2__abc_44228_n6871;
  wire u2__abc_44228_n6872;
  wire u2__abc_44228_n6873;
  wire u2__abc_44228_n6874;
  wire u2__abc_44228_n6875;
  wire u2__abc_44228_n6876;
  wire u2__abc_44228_n6877;
  wire u2__abc_44228_n6878_1;
  wire u2__abc_44228_n6879;
  wire u2__abc_44228_n6880;
  wire u2__abc_44228_n6881;
  wire u2__abc_44228_n6882;
  wire u2__abc_44228_n6883;
  wire u2__abc_44228_n6884;
  wire u2__abc_44228_n6885;
  wire u2__abc_44228_n6886;
  wire u2__abc_44228_n6887_1;
  wire u2__abc_44228_n6888;
  wire u2__abc_44228_n6889;
  wire u2__abc_44228_n6890;
  wire u2__abc_44228_n6891;
  wire u2__abc_44228_n6892;
  wire u2__abc_44228_n6893;
  wire u2__abc_44228_n6894;
  wire u2__abc_44228_n6895;
  wire u2__abc_44228_n6896;
  wire u2__abc_44228_n6897_1;
  wire u2__abc_44228_n6898;
  wire u2__abc_44228_n6899;
  wire u2__abc_44228_n6900;
  wire u2__abc_44228_n6901;
  wire u2__abc_44228_n6902;
  wire u2__abc_44228_n6903;
  wire u2__abc_44228_n6904;
  wire u2__abc_44228_n6905;
  wire u2__abc_44228_n6906_1;
  wire u2__abc_44228_n6907;
  wire u2__abc_44228_n6908;
  wire u2__abc_44228_n6909;
  wire u2__abc_44228_n6910;
  wire u2__abc_44228_n6911;
  wire u2__abc_44228_n6912;
  wire u2__abc_44228_n6913;
  wire u2__abc_44228_n6914;
  wire u2__abc_44228_n6915_1;
  wire u2__abc_44228_n6916;
  wire u2__abc_44228_n6917;
  wire u2__abc_44228_n6918;
  wire u2__abc_44228_n6919;
  wire u2__abc_44228_n6920;
  wire u2__abc_44228_n6921;
  wire u2__abc_44228_n6922;
  wire u2__abc_44228_n6923;
  wire u2__abc_44228_n6924_1;
  wire u2__abc_44228_n6925;
  wire u2__abc_44228_n6926;
  wire u2__abc_44228_n6927;
  wire u2__abc_44228_n6928;
  wire u2__abc_44228_n6929;
  wire u2__abc_44228_n6930;
  wire u2__abc_44228_n6931;
  wire u2__abc_44228_n6932;
  wire u2__abc_44228_n6933;
  wire u2__abc_44228_n6934_1;
  wire u2__abc_44228_n6935;
  wire u2__abc_44228_n6936;
  wire u2__abc_44228_n6937;
  wire u2__abc_44228_n6938;
  wire u2__abc_44228_n6939;
  wire u2__abc_44228_n6940;
  wire u2__abc_44228_n6941;
  wire u2__abc_44228_n6942;
  wire u2__abc_44228_n6943_1;
  wire u2__abc_44228_n6944;
  wire u2__abc_44228_n6945;
  wire u2__abc_44228_n6946;
  wire u2__abc_44228_n6947;
  wire u2__abc_44228_n6948;
  wire u2__abc_44228_n6949;
  wire u2__abc_44228_n6950;
  wire u2__abc_44228_n6951;
  wire u2__abc_44228_n6952;
  wire u2__abc_44228_n6953_1;
  wire u2__abc_44228_n6954;
  wire u2__abc_44228_n6955;
  wire u2__abc_44228_n6956;
  wire u2__abc_44228_n6957;
  wire u2__abc_44228_n6958;
  wire u2__abc_44228_n6959;
  wire u2__abc_44228_n6960;
  wire u2__abc_44228_n6961_1;
  wire u2__abc_44228_n6962;
  wire u2__abc_44228_n6963;
  wire u2__abc_44228_n6964;
  wire u2__abc_44228_n6965;
  wire u2__abc_44228_n6966;
  wire u2__abc_44228_n6967;
  wire u2__abc_44228_n6968;
  wire u2__abc_44228_n6969;
  wire u2__abc_44228_n6970;
  wire u2__abc_44228_n6971_1;
  wire u2__abc_44228_n6972;
  wire u2__abc_44228_n6973;
  wire u2__abc_44228_n6974;
  wire u2__abc_44228_n6975;
  wire u2__abc_44228_n6976;
  wire u2__abc_44228_n6977;
  wire u2__abc_44228_n6978;
  wire u2__abc_44228_n6979_1;
  wire u2__abc_44228_n6980;
  wire u2__abc_44228_n6981;
  wire u2__abc_44228_n6982;
  wire u2__abc_44228_n6983;
  wire u2__abc_44228_n6984;
  wire u2__abc_44228_n6985;
  wire u2__abc_44228_n6986;
  wire u2__abc_44228_n6987;
  wire u2__abc_44228_n6988_1;
  wire u2__abc_44228_n6989;
  wire u2__abc_44228_n6990;
  wire u2__abc_44228_n6991;
  wire u2__abc_44228_n6992;
  wire u2__abc_44228_n6993;
  wire u2__abc_44228_n6994;
  wire u2__abc_44228_n6995;
  wire u2__abc_44228_n6996;
  wire u2__abc_44228_n6997_1;
  wire u2__abc_44228_n6998;
  wire u2__abc_44228_n6999;
  wire u2__abc_44228_n7000;
  wire u2__abc_44228_n7001;
  wire u2__abc_44228_n7002;
  wire u2__abc_44228_n7003;
  wire u2__abc_44228_n7004;
  wire u2__abc_44228_n7005;
  wire u2__abc_44228_n7006;
  wire u2__abc_44228_n7007_1;
  wire u2__abc_44228_n7008;
  wire u2__abc_44228_n7009;
  wire u2__abc_44228_n7010;
  wire u2__abc_44228_n7011;
  wire u2__abc_44228_n7012;
  wire u2__abc_44228_n7013;
  wire u2__abc_44228_n7014_1;
  wire u2__abc_44228_n7015;
  wire u2__abc_44228_n7016;
  wire u2__abc_44228_n7017;
  wire u2__abc_44228_n7018;
  wire u2__abc_44228_n7019;
  wire u2__abc_44228_n7020;
  wire u2__abc_44228_n7021;
  wire u2__abc_44228_n7022_1;
  wire u2__abc_44228_n7023;
  wire u2__abc_44228_n7024;
  wire u2__abc_44228_n7025;
  wire u2__abc_44228_n7026;
  wire u2__abc_44228_n7027;
  wire u2__abc_44228_n7028;
  wire u2__abc_44228_n7029;
  wire u2__abc_44228_n7030;
  wire u2__abc_44228_n7031;
  wire u2__abc_44228_n7032_1;
  wire u2__abc_44228_n7033;
  wire u2__abc_44228_n7034;
  wire u2__abc_44228_n7035;
  wire u2__abc_44228_n7036;
  wire u2__abc_44228_n7037;
  wire u2__abc_44228_n7038;
  wire u2__abc_44228_n7039;
  wire u2__abc_44228_n7040;
  wire u2__abc_44228_n7041;
  wire u2__abc_44228_n7042_1;
  wire u2__abc_44228_n7043;
  wire u2__abc_44228_n7044;
  wire u2__abc_44228_n7045;
  wire u2__abc_44228_n7046;
  wire u2__abc_44228_n7047;
  wire u2__abc_44228_n7048;
  wire u2__abc_44228_n7049;
  wire u2__abc_44228_n7050_1;
  wire u2__abc_44228_n7051;
  wire u2__abc_44228_n7052;
  wire u2__abc_44228_n7053;
  wire u2__abc_44228_n7054;
  wire u2__abc_44228_n7055;
  wire u2__abc_44228_n7056;
  wire u2__abc_44228_n7057;
  wire u2__abc_44228_n7058;
  wire u2__abc_44228_n7059_1;
  wire u2__abc_44228_n7060;
  wire u2__abc_44228_n7061;
  wire u2__abc_44228_n7062;
  wire u2__abc_44228_n7063;
  wire u2__abc_44228_n7064;
  wire u2__abc_44228_n7065;
  wire u2__abc_44228_n7066;
  wire u2__abc_44228_n7067;
  wire u2__abc_44228_n7068_1;
  wire u2__abc_44228_n7069;
  wire u2__abc_44228_n7070;
  wire u2__abc_44228_n7071;
  wire u2__abc_44228_n7072;
  wire u2__abc_44228_n7073;
  wire u2__abc_44228_n7074;
  wire u2__abc_44228_n7075;
  wire u2__abc_44228_n7076;
  wire u2__abc_44228_n7077;
  wire u2__abc_44228_n7078_1;
  wire u2__abc_44228_n7079;
  wire u2__abc_44228_n7080;
  wire u2__abc_44228_n7081;
  wire u2__abc_44228_n7082;
  wire u2__abc_44228_n7083;
  wire u2__abc_44228_n7084;
  wire u2__abc_44228_n7085;
  wire u2__abc_44228_n7086;
  wire u2__abc_44228_n7087;
  wire u2__abc_44228_n7088_1;
  wire u2__abc_44228_n7089;
  wire u2__abc_44228_n7090;
  wire u2__abc_44228_n7091;
  wire u2__abc_44228_n7092;
  wire u2__abc_44228_n7093;
  wire u2__abc_44228_n7094;
  wire u2__abc_44228_n7095;
  wire u2__abc_44228_n7096;
  wire u2__abc_44228_n7097;
  wire u2__abc_44228_n7098_1;
  wire u2__abc_44228_n7099;
  wire u2__abc_44228_n7100;
  wire u2__abc_44228_n7101;
  wire u2__abc_44228_n7102;
  wire u2__abc_44228_n7103;
  wire u2__abc_44228_n7104;
  wire u2__abc_44228_n7105;
  wire u2__abc_44228_n7106_1;
  wire u2__abc_44228_n7107;
  wire u2__abc_44228_n7108;
  wire u2__abc_44228_n7109;
  wire u2__abc_44228_n7110;
  wire u2__abc_44228_n7111;
  wire u2__abc_44228_n7112;
  wire u2__abc_44228_n7113;
  wire u2__abc_44228_n7114;
  wire u2__abc_44228_n7115;
  wire u2__abc_44228_n7116_1;
  wire u2__abc_44228_n7117;
  wire u2__abc_44228_n7118;
  wire u2__abc_44228_n7119;
  wire u2__abc_44228_n7120;
  wire u2__abc_44228_n7121;
  wire u2__abc_44228_n7122;
  wire u2__abc_44228_n7123;
  wire u2__abc_44228_n7124;
  wire u2__abc_44228_n7125_1;
  wire u2__abc_44228_n7126;
  wire u2__abc_44228_n7127;
  wire u2__abc_44228_n7128;
  wire u2__abc_44228_n7129;
  wire u2__abc_44228_n7130;
  wire u2__abc_44228_n7131;
  wire u2__abc_44228_n7132;
  wire u2__abc_44228_n7133;
  wire u2__abc_44228_n7134_1;
  wire u2__abc_44228_n7135;
  wire u2__abc_44228_n7136;
  wire u2__abc_44228_n7137;
  wire u2__abc_44228_n7138;
  wire u2__abc_44228_n7139;
  wire u2__abc_44228_n7140;
  wire u2__abc_44228_n7141;
  wire u2__abc_44228_n7142;
  wire u2__abc_44228_n7143_1;
  wire u2__abc_44228_n7144;
  wire u2__abc_44228_n7145;
  wire u2__abc_44228_n7146;
  wire u2__abc_44228_n7147;
  wire u2__abc_44228_n7148;
  wire u2__abc_44228_n7149;
  wire u2__abc_44228_n7150;
  wire u2__abc_44228_n7151;
  wire u2__abc_44228_n7152;
  wire u2__abc_44228_n7153_1;
  wire u2__abc_44228_n7154;
  wire u2__abc_44228_n7155;
  wire u2__abc_44228_n7156;
  wire u2__abc_44228_n7157;
  wire u2__abc_44228_n7158;
  wire u2__abc_44228_n7159;
  wire u2__abc_44228_n7160;
  wire u2__abc_44228_n7161_1;
  wire u2__abc_44228_n7162;
  wire u2__abc_44228_n7163;
  wire u2__abc_44228_n7164;
  wire u2__abc_44228_n7165;
  wire u2__abc_44228_n7166;
  wire u2__abc_44228_n7167;
  wire u2__abc_44228_n7168;
  wire u2__abc_44228_n7169;
  wire u2__abc_44228_n7170_1;
  wire u2__abc_44228_n7171;
  wire u2__abc_44228_n7172;
  wire u2__abc_44228_n7173;
  wire u2__abc_44228_n7174;
  wire u2__abc_44228_n7175;
  wire u2__abc_44228_n7176;
  wire u2__abc_44228_n7177;
  wire u2__abc_44228_n7178;
  wire u2__abc_44228_n7179_1;
  wire u2__abc_44228_n7180;
  wire u2__abc_44228_n7181;
  wire u2__abc_44228_n7182;
  wire u2__abc_44228_n7183;
  wire u2__abc_44228_n7184;
  wire u2__abc_44228_n7185;
  wire u2__abc_44228_n7186;
  wire u2__abc_44228_n7187;
  wire u2__abc_44228_n7188;
  wire u2__abc_44228_n7189_1;
  wire u2__abc_44228_n7190;
  wire u2__abc_44228_n7191;
  wire u2__abc_44228_n7192;
  wire u2__abc_44228_n7193;
  wire u2__abc_44228_n7194;
  wire u2__abc_44228_n7195;
  wire u2__abc_44228_n7196;
  wire u2__abc_44228_n7197_1;
  wire u2__abc_44228_n7198;
  wire u2__abc_44228_n7199;
  wire u2__abc_44228_n7200;
  wire u2__abc_44228_n7201;
  wire u2__abc_44228_n7202;
  wire u2__abc_44228_n7203;
  wire u2__abc_44228_n7204;
  wire u2__abc_44228_n7205;
  wire u2__abc_44228_n7206_1;
  wire u2__abc_44228_n7207;
  wire u2__abc_44228_n7208;
  wire u2__abc_44228_n7209;
  wire u2__abc_44228_n7210;
  wire u2__abc_44228_n7211;
  wire u2__abc_44228_n7212;
  wire u2__abc_44228_n7213;
  wire u2__abc_44228_n7214;
  wire u2__abc_44228_n7215_1;
  wire u2__abc_44228_n7216;
  wire u2__abc_44228_n7217;
  wire u2__abc_44228_n7218;
  wire u2__abc_44228_n7219;
  wire u2__abc_44228_n7220;
  wire u2__abc_44228_n7221;
  wire u2__abc_44228_n7222;
  wire u2__abc_44228_n7223;
  wire u2__abc_44228_n7224;
  wire u2__abc_44228_n7225_1;
  wire u2__abc_44228_n7226;
  wire u2__abc_44228_n7227;
  wire u2__abc_44228_n7228;
  wire u2__abc_44228_n7229;
  wire u2__abc_44228_n7230;
  wire u2__abc_44228_n7231;
  wire u2__abc_44228_n7232;
  wire u2__abc_44228_n7233;
  wire u2__abc_44228_n7234_1;
  wire u2__abc_44228_n7235;
  wire u2__abc_44228_n7236;
  wire u2__abc_44228_n7237;
  wire u2__abc_44228_n7238;
  wire u2__abc_44228_n7239;
  wire u2__abc_44228_n7240;
  wire u2__abc_44228_n7241;
  wire u2__abc_44228_n7242;
  wire u2__abc_44228_n7243;
  wire u2__abc_44228_n7244_1;
  wire u2__abc_44228_n7245;
  wire u2__abc_44228_n7246;
  wire u2__abc_44228_n7247;
  wire u2__abc_44228_n7248;
  wire u2__abc_44228_n7249;
  wire u2__abc_44228_n7250;
  wire u2__abc_44228_n7251;
  wire u2__abc_44228_n7252_1;
  wire u2__abc_44228_n7253;
  wire u2__abc_44228_n7254;
  wire u2__abc_44228_n7255;
  wire u2__abc_44228_n7256;
  wire u2__abc_44228_n7257;
  wire u2__abc_44228_n7258;
  wire u2__abc_44228_n7259;
  wire u2__abc_44228_n7260;
  wire u2__abc_44228_n7261;
  wire u2__abc_44228_n7262_1;
  wire u2__abc_44228_n7263;
  wire u2__abc_44228_n7264;
  wire u2__abc_44228_n7265;
  wire u2__abc_44228_n7266;
  wire u2__abc_44228_n7267;
  wire u2__abc_44228_n7268;
  wire u2__abc_44228_n7269;
  wire u2__abc_44228_n7270;
  wire u2__abc_44228_n7271_1;
  wire u2__abc_44228_n7272;
  wire u2__abc_44228_n7273;
  wire u2__abc_44228_n7274;
  wire u2__abc_44228_n7275;
  wire u2__abc_44228_n7276;
  wire u2__abc_44228_n7277;
  wire u2__abc_44228_n7278;
  wire u2__abc_44228_n7279;
  wire u2__abc_44228_n7280_1;
  wire u2__abc_44228_n7281;
  wire u2__abc_44228_n7282;
  wire u2__abc_44228_n7283;
  wire u2__abc_44228_n7284;
  wire u2__abc_44228_n7285;
  wire u2__abc_44228_n7286;
  wire u2__abc_44228_n7287;
  wire u2__abc_44228_n7288;
  wire u2__abc_44228_n7289_1;
  wire u2__abc_44228_n7290;
  wire u2__abc_44228_n7291;
  wire u2__abc_44228_n7292;
  wire u2__abc_44228_n7293;
  wire u2__abc_44228_n7294;
  wire u2__abc_44228_n7295;
  wire u2__abc_44228_n7296;
  wire u2__abc_44228_n7297;
  wire u2__abc_44228_n7298;
  wire u2__abc_44228_n7299_1;
  wire u2__abc_44228_n7300;
  wire u2__abc_44228_n7301;
  wire u2__abc_44228_n7302;
  wire u2__abc_44228_n7303;
  wire u2__abc_44228_n7304;
  wire u2__abc_44228_n7305;
  wire u2__abc_44228_n7306;
  wire u2__abc_44228_n7307;
  wire u2__abc_44228_n7308;
  wire u2__abc_44228_n7309_1;
  wire u2__abc_44228_n7310;
  wire u2__abc_44228_n7311;
  wire u2__abc_44228_n7312;
  wire u2__abc_44228_n7313;
  wire u2__abc_44228_n7314;
  wire u2__abc_44228_n7315;
  wire u2__abc_44228_n7316;
  wire u2__abc_44228_n7317;
  wire u2__abc_44228_n7318;
  wire u2__abc_44228_n7319_1;
  wire u2__abc_44228_n7320;
  wire u2__abc_44228_n7321;
  wire u2__abc_44228_n7322;
  wire u2__abc_44228_n7323;
  wire u2__abc_44228_n7324;
  wire u2__abc_44228_n7325;
  wire u2__abc_44228_n7326;
  wire u2__abc_44228_n7327_1;
  wire u2__abc_44228_n7328;
  wire u2__abc_44228_n7329;
  wire u2__abc_44228_n7330;
  wire u2__abc_44228_n7331;
  wire u2__abc_44228_n7332;
  wire u2__abc_44228_n7333;
  wire u2__abc_44228_n7334;
  wire u2__abc_44228_n7335;
  wire u2__abc_44228_n7336;
  wire u2__abc_44228_n7337_1;
  wire u2__abc_44228_n7338;
  wire u2__abc_44228_n7339;
  wire u2__abc_44228_n7340;
  wire u2__abc_44228_n7341;
  wire u2__abc_44228_n7342;
  wire u2__abc_44228_n7343;
  wire u2__abc_44228_n7344;
  wire u2__abc_44228_n7345;
  wire u2__abc_44228_n7346_1;
  wire u2__abc_44228_n7347;
  wire u2__abc_44228_n7348;
  wire u2__abc_44228_n7349;
  wire u2__abc_44228_n7350;
  wire u2__abc_44228_n7351;
  wire u2__abc_44228_n7352;
  wire u2__abc_44228_n7353;
  wire u2__abc_44228_n7354;
  wire u2__abc_44228_n7355_1;
  wire u2__abc_44228_n7356;
  wire u2__abc_44228_n7357;
  wire u2__abc_44228_n7358;
  wire u2__abc_44228_n7359;
  wire u2__abc_44228_n7360;
  wire u2__abc_44228_n7361;
  wire u2__abc_44228_n7362;
  wire u2__abc_44228_n7363;
  wire u2__abc_44228_n7364_1;
  wire u2__abc_44228_n7365;
  wire u2__abc_44228_n7366;
  wire u2__abc_44228_n7367;
  wire u2__abc_44228_n7368;
  wire u2__abc_44228_n7369;
  wire u2__abc_44228_n7370;
  wire u2__abc_44228_n7371;
  wire u2__abc_44228_n7372;
  wire u2__abc_44228_n7373;
  wire u2__abc_44228_n7374_1;
  wire u2__abc_44228_n7375;
  wire u2__abc_44228_n7376;
  wire u2__abc_44228_n7377;
  wire u2__abc_44228_n7378;
  wire u2__abc_44228_n7379;
  wire u2__abc_44228_n7380;
  wire u2__abc_44228_n7381;
  wire u2__abc_44228_n7382_1;
  wire u2__abc_44228_n7383;
  wire u2__abc_44228_n7384;
  wire u2__abc_44228_n7385;
  wire u2__abc_44228_n7386;
  wire u2__abc_44228_n7387;
  wire u2__abc_44228_n7388;
  wire u2__abc_44228_n7389;
  wire u2__abc_44228_n7390;
  wire u2__abc_44228_n7391;
  wire u2__abc_44228_n7392_1;
  wire u2__abc_44228_n7393;
  wire u2__abc_44228_n7394;
  wire u2__abc_44228_n7395;
  wire u2__abc_44228_n7396;
  wire u2__abc_44228_n7397;
  wire u2__abc_44228_n7398;
  wire u2__abc_44228_n7399;
  wire u2__abc_44228_n7400_1;
  wire u2__abc_44228_n7401;
  wire u2__abc_44228_n7402;
  wire u2__abc_44228_n7403;
  wire u2__abc_44228_n7404;
  wire u2__abc_44228_n7405;
  wire u2__abc_44228_n7406;
  wire u2__abc_44228_n7407;
  wire u2__abc_44228_n7408;
  wire u2__abc_44228_n7409;
  wire u2__abc_44228_n7410_1;
  wire u2__abc_44228_n7411;
  wire u2__abc_44228_n7412;
  wire u2__abc_44228_n7413;
  wire u2__abc_44228_n7414;
  wire u2__abc_44228_n7415;
  wire u2__abc_44228_n7416;
  wire u2__abc_44228_n7417;
  wire u2__abc_44228_n7418;
  wire u2__abc_44228_n7419_1;
  wire u2__abc_44228_n7420;
  wire u2__abc_44228_n7421;
  wire u2__abc_44228_n7422;
  wire u2__abc_44228_n7423;
  wire u2__abc_44228_n7424;
  wire u2__abc_44228_n7425;
  wire u2__abc_44228_n7426;
  wire u2__abc_44228_n7427;
  wire u2__abc_44228_n7428_1;
  wire u2__abc_44228_n7429;
  wire u2__abc_44228_n7430;
  wire u2__abc_44228_n7431;
  wire u2__abc_44228_n7432;
  wire u2__abc_44228_n7433;
  wire u2__abc_44228_n7434;
  wire u2__abc_44228_n7435;
  wire u2__abc_44228_n7436;
  wire u2__abc_44228_n7437_1;
  wire u2__abc_44228_n7438;
  wire u2__abc_44228_n7439;
  wire u2__abc_44228_n7440;
  wire u2__abc_44228_n7441;
  wire u2__abc_44228_n7442;
  wire u2__abc_44228_n7443;
  wire u2__abc_44228_n7444;
  wire u2__abc_44228_n7445;
  wire u2__abc_44228_n7446;
  wire u2__abc_44228_n7447_1;
  wire u2__abc_44228_n7448;
  wire u2__abc_44228_n7449;
  wire u2__abc_44228_n7450;
  wire u2__abc_44228_n7451;
  wire u2__abc_44228_n7452;
  wire u2__abc_44228_n7453;
  wire u2__abc_44228_n7454;
  wire u2__abc_44228_n7455_1;
  wire u2__abc_44228_n7456;
  wire u2__abc_44228_n7457;
  wire u2__abc_44228_n7458;
  wire u2__abc_44228_n7459;
  wire u2__abc_44228_n7460;
  wire u2__abc_44228_n7461;
  wire u2__abc_44228_n7462;
  wire u2__abc_44228_n7463;
  wire u2__abc_44228_n7464_1;
  wire u2__abc_44228_n7465;
  wire u2__abc_44228_n7466;
  wire u2__abc_44228_n7467;
  wire u2__abc_44228_n7468;
  wire u2__abc_44228_n7469;
  wire u2__abc_44228_n7470;
  wire u2__abc_44228_n7471;
  wire u2__abc_44228_n7472;
  wire u2__abc_44228_n7473_1;
  wire u2__abc_44228_n7474;
  wire u2__abc_44228_n7475;
  wire u2__abc_44228_n7476;
  wire u2__abc_44228_n7477;
  wire u2__abc_44228_n7478;
  wire u2__abc_44228_n7479;
  wire u2__abc_44228_n7480;
  wire u2__abc_44228_n7481;
  wire u2__abc_44228_n7482;
  wire u2__abc_44228_n7483_1;
  wire u2__abc_44228_n7484;
  wire u2__abc_44228_n7485;
  wire u2__abc_44228_n7486;
  wire u2__abc_44228_n7487;
  wire u2__abc_44228_n7488;
  wire u2__abc_44228_n7489;
  wire u2__abc_44228_n7490;
  wire u2__abc_44228_n7491;
  wire u2__abc_44228_n7492;
  wire u2__abc_44228_n7493_1;
  wire u2__abc_44228_n7494;
  wire u2__abc_44228_n7495;
  wire u2__abc_44228_n7496;
  wire u2__abc_44228_n7497;
  wire u2__abc_44228_n7498;
  wire u2__abc_44228_n7499;
  wire u2__abc_44228_n7500;
  wire u2__abc_44228_n7501;
  wire u2__abc_44228_n7502_1;
  wire u2__abc_44228_n7503;
  wire u2__abc_44228_n7504;
  wire u2__abc_44228_n7505;
  wire u2__abc_44228_n7506;
  wire u2__abc_44228_n7507;
  wire u2__abc_44228_n7508;
  wire u2__abc_44228_n7509;
  wire u2__abc_44228_n7510;
  wire u2__abc_44228_n7511_1;
  wire u2__abc_44228_n7512;
  wire u2__abc_44228_n7513;
  wire u2__abc_44228_n7514;
  wire u2__abc_44228_n7515;
  wire u2__abc_44228_n7516;
  wire u2__abc_44228_n7517;
  wire u2__abc_44228_n7518;
  wire u2__abc_44228_n7519;
  wire u2__abc_44228_n7520;
  wire u2__abc_44228_n7521_1;
  wire u2__abc_44228_n7522;
  wire u2__abc_44228_n7523;
  wire u2__abc_44228_n7524;
  wire u2__abc_44228_n7525;
  wire u2__abc_44228_n7526;
  wire u2__abc_44228_n7527;
  wire u2__abc_44228_n7528;
  wire u2__abc_44228_n7529;
  wire u2__abc_44228_n7530_1;
  wire u2__abc_44228_n7531;
  wire u2__abc_44228_n7532;
  wire u2__abc_44228_n7533;
  wire u2__abc_44228_n7534;
  wire u2__abc_44228_n7535;
  wire u2__abc_44228_n7536;
  wire u2__abc_44228_n7537;
  wire u2__abc_44228_n7538;
  wire u2__abc_44228_n7539;
  wire u2__abc_44228_n7540_1;
  wire u2__abc_44228_n7541;
  wire u2__abc_44228_n7542;
  wire u2__abc_44228_n7543;
  wire u2__abc_44228_n7544;
  wire u2__abc_44228_n7545;
  wire u2__abc_44228_n7546;
  wire u2__abc_44228_n7547;
  wire u2__abc_44228_n7547_bF_buf0;
  wire u2__abc_44228_n7547_bF_buf1;
  wire u2__abc_44228_n7547_bF_buf10;
  wire u2__abc_44228_n7547_bF_buf11;
  wire u2__abc_44228_n7547_bF_buf12;
  wire u2__abc_44228_n7547_bF_buf13;
  wire u2__abc_44228_n7547_bF_buf14;
  wire u2__abc_44228_n7547_bF_buf15;
  wire u2__abc_44228_n7547_bF_buf16;
  wire u2__abc_44228_n7547_bF_buf17;
  wire u2__abc_44228_n7547_bF_buf18;
  wire u2__abc_44228_n7547_bF_buf19;
  wire u2__abc_44228_n7547_bF_buf2;
  wire u2__abc_44228_n7547_bF_buf20;
  wire u2__abc_44228_n7547_bF_buf21;
  wire u2__abc_44228_n7547_bF_buf22;
  wire u2__abc_44228_n7547_bF_buf23;
  wire u2__abc_44228_n7547_bF_buf24;
  wire u2__abc_44228_n7547_bF_buf25;
  wire u2__abc_44228_n7547_bF_buf26;
  wire u2__abc_44228_n7547_bF_buf27;
  wire u2__abc_44228_n7547_bF_buf28;
  wire u2__abc_44228_n7547_bF_buf29;
  wire u2__abc_44228_n7547_bF_buf3;
  wire u2__abc_44228_n7547_bF_buf30;
  wire u2__abc_44228_n7547_bF_buf31;
  wire u2__abc_44228_n7547_bF_buf32;
  wire u2__abc_44228_n7547_bF_buf33;
  wire u2__abc_44228_n7547_bF_buf34;
  wire u2__abc_44228_n7547_bF_buf35;
  wire u2__abc_44228_n7547_bF_buf36;
  wire u2__abc_44228_n7547_bF_buf37;
  wire u2__abc_44228_n7547_bF_buf38;
  wire u2__abc_44228_n7547_bF_buf39;
  wire u2__abc_44228_n7547_bF_buf4;
  wire u2__abc_44228_n7547_bF_buf40;
  wire u2__abc_44228_n7547_bF_buf41;
  wire u2__abc_44228_n7547_bF_buf42;
  wire u2__abc_44228_n7547_bF_buf43;
  wire u2__abc_44228_n7547_bF_buf44;
  wire u2__abc_44228_n7547_bF_buf45;
  wire u2__abc_44228_n7547_bF_buf46;
  wire u2__abc_44228_n7547_bF_buf47;
  wire u2__abc_44228_n7547_bF_buf48;
  wire u2__abc_44228_n7547_bF_buf49;
  wire u2__abc_44228_n7547_bF_buf5;
  wire u2__abc_44228_n7547_bF_buf50;
  wire u2__abc_44228_n7547_bF_buf51;
  wire u2__abc_44228_n7547_bF_buf52;
  wire u2__abc_44228_n7547_bF_buf53;
  wire u2__abc_44228_n7547_bF_buf54;
  wire u2__abc_44228_n7547_bF_buf55;
  wire u2__abc_44228_n7547_bF_buf56;
  wire u2__abc_44228_n7547_bF_buf57;
  wire u2__abc_44228_n7547_bF_buf6;
  wire u2__abc_44228_n7547_bF_buf7;
  wire u2__abc_44228_n7547_bF_buf8;
  wire u2__abc_44228_n7547_bF_buf9;
  wire u2__abc_44228_n7547_hier0_bF_buf0;
  wire u2__abc_44228_n7547_hier0_bF_buf1;
  wire u2__abc_44228_n7547_hier0_bF_buf2;
  wire u2__abc_44228_n7547_hier0_bF_buf3;
  wire u2__abc_44228_n7547_hier0_bF_buf4;
  wire u2__abc_44228_n7547_hier0_bF_buf5;
  wire u2__abc_44228_n7547_hier0_bF_buf6;
  wire u2__abc_44228_n7548_1;
  wire u2__abc_44228_n7548_1_bF_buf0;
  wire u2__abc_44228_n7548_1_bF_buf1;
  wire u2__abc_44228_n7548_1_bF_buf10;
  wire u2__abc_44228_n7548_1_bF_buf11;
  wire u2__abc_44228_n7548_1_bF_buf12;
  wire u2__abc_44228_n7548_1_bF_buf13;
  wire u2__abc_44228_n7548_1_bF_buf14;
  wire u2__abc_44228_n7548_1_bF_buf15;
  wire u2__abc_44228_n7548_1_bF_buf16;
  wire u2__abc_44228_n7548_1_bF_buf17;
  wire u2__abc_44228_n7548_1_bF_buf18;
  wire u2__abc_44228_n7548_1_bF_buf19;
  wire u2__abc_44228_n7548_1_bF_buf2;
  wire u2__abc_44228_n7548_1_bF_buf20;
  wire u2__abc_44228_n7548_1_bF_buf21;
  wire u2__abc_44228_n7548_1_bF_buf22;
  wire u2__abc_44228_n7548_1_bF_buf23;
  wire u2__abc_44228_n7548_1_bF_buf24;
  wire u2__abc_44228_n7548_1_bF_buf25;
  wire u2__abc_44228_n7548_1_bF_buf26;
  wire u2__abc_44228_n7548_1_bF_buf27;
  wire u2__abc_44228_n7548_1_bF_buf28;
  wire u2__abc_44228_n7548_1_bF_buf29;
  wire u2__abc_44228_n7548_1_bF_buf3;
  wire u2__abc_44228_n7548_1_bF_buf30;
  wire u2__abc_44228_n7548_1_bF_buf31;
  wire u2__abc_44228_n7548_1_bF_buf32;
  wire u2__abc_44228_n7548_1_bF_buf33;
  wire u2__abc_44228_n7548_1_bF_buf34;
  wire u2__abc_44228_n7548_1_bF_buf35;
  wire u2__abc_44228_n7548_1_bF_buf36;
  wire u2__abc_44228_n7548_1_bF_buf37;
  wire u2__abc_44228_n7548_1_bF_buf38;
  wire u2__abc_44228_n7548_1_bF_buf39;
  wire u2__abc_44228_n7548_1_bF_buf4;
  wire u2__abc_44228_n7548_1_bF_buf40;
  wire u2__abc_44228_n7548_1_bF_buf41;
  wire u2__abc_44228_n7548_1_bF_buf42;
  wire u2__abc_44228_n7548_1_bF_buf43;
  wire u2__abc_44228_n7548_1_bF_buf44;
  wire u2__abc_44228_n7548_1_bF_buf45;
  wire u2__abc_44228_n7548_1_bF_buf46;
  wire u2__abc_44228_n7548_1_bF_buf47;
  wire u2__abc_44228_n7548_1_bF_buf48;
  wire u2__abc_44228_n7548_1_bF_buf49;
  wire u2__abc_44228_n7548_1_bF_buf5;
  wire u2__abc_44228_n7548_1_bF_buf50;
  wire u2__abc_44228_n7548_1_bF_buf51;
  wire u2__abc_44228_n7548_1_bF_buf52;
  wire u2__abc_44228_n7548_1_bF_buf53;
  wire u2__abc_44228_n7548_1_bF_buf54;
  wire u2__abc_44228_n7548_1_bF_buf55;
  wire u2__abc_44228_n7548_1_bF_buf56;
  wire u2__abc_44228_n7548_1_bF_buf57;
  wire u2__abc_44228_n7548_1_bF_buf6;
  wire u2__abc_44228_n7548_1_bF_buf7;
  wire u2__abc_44228_n7548_1_bF_buf8;
  wire u2__abc_44228_n7548_1_bF_buf9;
  wire u2__abc_44228_n7548_1_hier0_bF_buf0;
  wire u2__abc_44228_n7548_1_hier0_bF_buf1;
  wire u2__abc_44228_n7548_1_hier0_bF_buf2;
  wire u2__abc_44228_n7548_1_hier0_bF_buf3;
  wire u2__abc_44228_n7548_1_hier0_bF_buf4;
  wire u2__abc_44228_n7548_1_hier0_bF_buf5;
  wire u2__abc_44228_n7548_1_hier0_bF_buf6;
  wire u2__abc_44228_n7549;
  wire u2__abc_44228_n7550;
  wire u2__abc_44228_n7551;
  wire u2__abc_44228_n7552;
  wire u2__abc_44228_n7553;
  wire u2__abc_44228_n7554;
  wire u2__abc_44228_n7555;
  wire u2__abc_44228_n7556;
  wire u2__abc_44228_n7557;
  wire u2__abc_44228_n7558_1;
  wire u2__abc_44228_n7559;
  wire u2__abc_44228_n7561;
  wire u2__abc_44228_n7562;
  wire u2__abc_44228_n7563;
  wire u2__abc_44228_n7564;
  wire u2__abc_44228_n7565;
  wire u2__abc_44228_n7566;
  wire u2__abc_44228_n7567_1;
  wire u2__abc_44228_n7568;
  wire u2__abc_44228_n7569;
  wire u2__abc_44228_n7570;
  wire u2__abc_44228_n7571;
  wire u2__abc_44228_n7572;
  wire u2__abc_44228_n7573;
  wire u2__abc_44228_n7575;
  wire u2__abc_44228_n7576_1;
  wire u2__abc_44228_n7577;
  wire u2__abc_44228_n7578;
  wire u2__abc_44228_n7579;
  wire u2__abc_44228_n7580;
  wire u2__abc_44228_n7581;
  wire u2__abc_44228_n7582;
  wire u2__abc_44228_n7583;
  wire u2__abc_44228_n7584;
  wire u2__abc_44228_n7585;
  wire u2__abc_44228_n7586_1;
  wire u2__abc_44228_n7587;
  wire u2__abc_44228_n7588;
  wire u2__abc_44228_n7589;
  wire u2__abc_44228_n7591;
  wire u2__abc_44228_n7592;
  wire u2__abc_44228_n7593;
  wire u2__abc_44228_n7594;
  wire u2__abc_44228_n7595;
  wire u2__abc_44228_n7596;
  wire u2__abc_44228_n7597_1;
  wire u2__abc_44228_n7598;
  wire u2__abc_44228_n7599;
  wire u2__abc_44228_n7600;
  wire u2__abc_44228_n7601;
  wire u2__abc_44228_n7602;
  wire u2__abc_44228_n7603;
  wire u2__abc_44228_n7604;
  wire u2__abc_44228_n7605_1;
  wire u2__abc_44228_n7606;
  wire u2__abc_44228_n7607;
  wire u2__abc_44228_n7609;
  wire u2__abc_44228_n7610;
  wire u2__abc_44228_n7611;
  wire u2__abc_44228_n7612;
  wire u2__abc_44228_n7613;
  wire u2__abc_44228_n7614;
  wire u2__abc_44228_n7615_1;
  wire u2__abc_44228_n7616_1;
  wire u2__abc_44228_n7617;
  wire u2__abc_44228_n7618;
  wire u2__abc_44228_n7619;
  wire u2__abc_44228_n7620;
  wire u2__abc_44228_n7621;
  wire u2__abc_44228_n7622_1;
  wire u2__abc_44228_n7624;
  wire u2__abc_44228_n7625;
  wire u2__abc_44228_n7626;
  wire u2__abc_44228_n7627;
  wire u2__abc_44228_n7628;
  wire u2__abc_44228_n7629_1;
  wire u2__abc_44228_n7630_1;
  wire u2__abc_44228_n7631;
  wire u2__abc_44228_n7632;
  wire u2__abc_44228_n7633;
  wire u2__abc_44228_n7634;
  wire u2__abc_44228_n7635;
  wire u2__abc_44228_n7636_1;
  wire u2__abc_44228_n7637_1;
  wire u2__abc_44228_n7638;
  wire u2__abc_44228_n7639;
  wire u2__abc_44228_n7641;
  wire u2__abc_44228_n7642;
  wire u2__abc_44228_n7643_1;
  wire u2__abc_44228_n7644_1;
  wire u2__abc_44228_n7645;
  wire u2__abc_44228_n7646;
  wire u2__abc_44228_n7647;
  wire u2__abc_44228_n7648;
  wire u2__abc_44228_n7649;
  wire u2__abc_44228_n7650_1;
  wire u2__abc_44228_n7651_1;
  wire u2__abc_44228_n7652;
  wire u2__abc_44228_n7653;
  wire u2__abc_44228_n7654;
  wire u2__abc_44228_n7655;
  wire u2__abc_44228_n7656;
  wire u2__abc_44228_n7658_1;
  wire u2__abc_44228_n7659;
  wire u2__abc_44228_n7660;
  wire u2__abc_44228_n7661;
  wire u2__abc_44228_n7662;
  wire u2__abc_44228_n7663;
  wire u2__abc_44228_n7664_1;
  wire u2__abc_44228_n7665_1;
  wire u2__abc_44228_n7666;
  wire u2__abc_44228_n7667;
  wire u2__abc_44228_n7668;
  wire u2__abc_44228_n7669;
  wire u2__abc_44228_n7670;
  wire u2__abc_44228_n7671_1;
  wire u2__abc_44228_n7672_1;
  wire u2__abc_44228_n7673;
  wire u2__abc_44228_n7675;
  wire u2__abc_44228_n7676;
  wire u2__abc_44228_n7677;
  wire u2__abc_44228_n7678_1;
  wire u2__abc_44228_n7679_1;
  wire u2__abc_44228_n7680;
  wire u2__abc_44228_n7681;
  wire u2__abc_44228_n7682;
  wire u2__abc_44228_n7683;
  wire u2__abc_44228_n7684;
  wire u2__abc_44228_n7685_1;
  wire u2__abc_44228_n7686_1;
  wire u2__abc_44228_n7687;
  wire u2__abc_44228_n7688;
  wire u2__abc_44228_n7690;
  wire u2__abc_44228_n7691;
  wire u2__abc_44228_n7692_1;
  wire u2__abc_44228_n7693_1;
  wire u2__abc_44228_n7694;
  wire u2__abc_44228_n7695;
  wire u2__abc_44228_n7696;
  wire u2__abc_44228_n7697;
  wire u2__abc_44228_n7698;
  wire u2__abc_44228_n7699_1;
  wire u2__abc_44228_n7700_1;
  wire u2__abc_44228_n7701;
  wire u2__abc_44228_n7702;
  wire u2__abc_44228_n7703;
  wire u2__abc_44228_n7704;
  wire u2__abc_44228_n7705;
  wire u2__abc_44228_n7707_1;
  wire u2__abc_44228_n7708;
  wire u2__abc_44228_n7709;
  wire u2__abc_44228_n7710;
  wire u2__abc_44228_n7711;
  wire u2__abc_44228_n7712;
  wire u2__abc_44228_n7713_1;
  wire u2__abc_44228_n7714_1;
  wire u2__abc_44228_n7715;
  wire u2__abc_44228_n7716;
  wire u2__abc_44228_n7717;
  wire u2__abc_44228_n7718;
  wire u2__abc_44228_n7719;
  wire u2__abc_44228_n7720_1;
  wire u2__abc_44228_n7721_1;
  wire u2__abc_44228_n7722;
  wire u2__abc_44228_n7724;
  wire u2__abc_44228_n7725;
  wire u2__abc_44228_n7726;
  wire u2__abc_44228_n7727_1;
  wire u2__abc_44228_n7728_1;
  wire u2__abc_44228_n7729;
  wire u2__abc_44228_n7730;
  wire u2__abc_44228_n7731;
  wire u2__abc_44228_n7732;
  wire u2__abc_44228_n7733;
  wire u2__abc_44228_n7734_1;
  wire u2__abc_44228_n7735_1;
  wire u2__abc_44228_n7736;
  wire u2__abc_44228_n7737;
  wire u2__abc_44228_n7738;
  wire u2__abc_44228_n7739;
  wire u2__abc_44228_n7741_1;
  wire u2__abc_44228_n7742_1;
  wire u2__abc_44228_n7743;
  wire u2__abc_44228_n7744;
  wire u2__abc_44228_n7745;
  wire u2__abc_44228_n7746;
  wire u2__abc_44228_n7747;
  wire u2__abc_44228_n7748_1;
  wire u2__abc_44228_n7749_1;
  wire u2__abc_44228_n7750;
  wire u2__abc_44228_n7751;
  wire u2__abc_44228_n7752;
  wire u2__abc_44228_n7753;
  wire u2__abc_44228_n7754;
  wire u2__abc_44228_n7755_1;
  wire u2__abc_44228_n7756_1;
  wire u2__abc_44228_n7758;
  wire u2__abc_44228_n7759;
  wire u2__abc_44228_n7760;
  wire u2__abc_44228_n7761;
  wire u2__abc_44228_n7762_1;
  wire u2__abc_44228_n7763_1;
  wire u2__abc_44228_n7764;
  wire u2__abc_44228_n7765;
  wire u2__abc_44228_n7766;
  wire u2__abc_44228_n7767;
  wire u2__abc_44228_n7768;
  wire u2__abc_44228_n7769_1;
  wire u2__abc_44228_n7770_1;
  wire u2__abc_44228_n7771;
  wire u2__abc_44228_n7772;
  wire u2__abc_44228_n7773;
  wire u2__abc_44228_n7775;
  wire u2__abc_44228_n7776_1;
  wire u2__abc_44228_n7777_1;
  wire u2__abc_44228_n7778;
  wire u2__abc_44228_n7779;
  wire u2__abc_44228_n7780;
  wire u2__abc_44228_n7781;
  wire u2__abc_44228_n7782;
  wire u2__abc_44228_n7783_1;
  wire u2__abc_44228_n7784_1;
  wire u2__abc_44228_n7785;
  wire u2__abc_44228_n7786;
  wire u2__abc_44228_n7787;
  wire u2__abc_44228_n7788;
  wire u2__abc_44228_n7789;
  wire u2__abc_44228_n7790_1;
  wire u2__abc_44228_n7792;
  wire u2__abc_44228_n7793;
  wire u2__abc_44228_n7794;
  wire u2__abc_44228_n7795;
  wire u2__abc_44228_n7796;
  wire u2__abc_44228_n7797_1;
  wire u2__abc_44228_n7798_1;
  wire u2__abc_44228_n7799;
  wire u2__abc_44228_n7800;
  wire u2__abc_44228_n7801;
  wire u2__abc_44228_n7802;
  wire u2__abc_44228_n7803;
  wire u2__abc_44228_n7804_1;
  wire u2__abc_44228_n7805_1;
  wire u2__abc_44228_n7806;
  wire u2__abc_44228_n7807;
  wire u2__abc_44228_n7809;
  wire u2__abc_44228_n7810;
  wire u2__abc_44228_n7811_1;
  wire u2__abc_44228_n7812_1;
  wire u2__abc_44228_n7813;
  wire u2__abc_44228_n7814;
  wire u2__abc_44228_n7815;
  wire u2__abc_44228_n7816;
  wire u2__abc_44228_n7817;
  wire u2__abc_44228_n7818_1;
  wire u2__abc_44228_n7819_1;
  wire u2__abc_44228_n7820;
  wire u2__abc_44228_n7821;
  wire u2__abc_44228_n7822;
  wire u2__abc_44228_n7824;
  wire u2__abc_44228_n7825_1;
  wire u2__abc_44228_n7826_1;
  wire u2__abc_44228_n7827;
  wire u2__abc_44228_n7828;
  wire u2__abc_44228_n7829;
  wire u2__abc_44228_n7830;
  wire u2__abc_44228_n7831;
  wire u2__abc_44228_n7832_1;
  wire u2__abc_44228_n7833_1;
  wire u2__abc_44228_n7834;
  wire u2__abc_44228_n7835;
  wire u2__abc_44228_n7836;
  wire u2__abc_44228_n7837;
  wire u2__abc_44228_n7838;
  wire u2__abc_44228_n7839_1;
  wire u2__abc_44228_n7841;
  wire u2__abc_44228_n7842;
  wire u2__abc_44228_n7843;
  wire u2__abc_44228_n7844;
  wire u2__abc_44228_n7845_1;
  wire u2__abc_44228_n7846;
  wire u2__abc_44228_n7847;
  wire u2__abc_44228_n7848;
  wire u2__abc_44228_n7849;
  wire u2__abc_44228_n7850_1;
  wire u2__abc_44228_n7851_1;
  wire u2__abc_44228_n7852;
  wire u2__abc_44228_n7853;
  wire u2__abc_44228_n7854;
  wire u2__abc_44228_n7855;
  wire u2__abc_44228_n7856_1;
  wire u2__abc_44228_n7858;
  wire u2__abc_44228_n7859;
  wire u2__abc_44228_n7860;
  wire u2__abc_44228_n7861_1;
  wire u2__abc_44228_n7862_1;
  wire u2__abc_44228_n7863;
  wire u2__abc_44228_n7864;
  wire u2__abc_44228_n7865;
  wire u2__abc_44228_n7866;
  wire u2__abc_44228_n7867_1;
  wire u2__abc_44228_n7868;
  wire u2__abc_44228_n7869;
  wire u2__abc_44228_n7870;
  wire u2__abc_44228_n7871;
  wire u2__abc_44228_n7872_1;
  wire u2__abc_44228_n7873_1;
  wire u2__abc_44228_n7875;
  wire u2__abc_44228_n7876;
  wire u2__abc_44228_n7877;
  wire u2__abc_44228_n7878_1;
  wire u2__abc_44228_n7879;
  wire u2__abc_44228_n7880;
  wire u2__abc_44228_n7881;
  wire u2__abc_44228_n7882;
  wire u2__abc_44228_n7883_1;
  wire u2__abc_44228_n7884_1;
  wire u2__abc_44228_n7885;
  wire u2__abc_44228_n7886;
  wire u2__abc_44228_n7887;
  wire u2__abc_44228_n7888;
  wire u2__abc_44228_n7889_1;
  wire u2__abc_44228_n7890;
  wire u2__abc_44228_n7892;
  wire u2__abc_44228_n7893;
  wire u2__abc_44228_n7894_1;
  wire u2__abc_44228_n7895_1;
  wire u2__abc_44228_n7896;
  wire u2__abc_44228_n7897;
  wire u2__abc_44228_n7898;
  wire u2__abc_44228_n7899;
  wire u2__abc_44228_n7900_1;
  wire u2__abc_44228_n7901;
  wire u2__abc_44228_n7902;
  wire u2__abc_44228_n7903;
  wire u2__abc_44228_n7904;
  wire u2__abc_44228_n7905_1;
  wire u2__abc_44228_n7906_1;
  wire u2__abc_44228_n7907;
  wire u2__abc_44228_n7909;
  wire u2__abc_44228_n7910;
  wire u2__abc_44228_n7911_1;
  wire u2__abc_44228_n7912;
  wire u2__abc_44228_n7913;
  wire u2__abc_44228_n7914;
  wire u2__abc_44228_n7915;
  wire u2__abc_44228_n7916_1;
  wire u2__abc_44228_n7917_1;
  wire u2__abc_44228_n7918;
  wire u2__abc_44228_n7919;
  wire u2__abc_44228_n7920;
  wire u2__abc_44228_n7921;
  wire u2__abc_44228_n7922_1;
  wire u2__abc_44228_n7923;
  wire u2__abc_44228_n7924;
  wire u2__abc_44228_n7926;
  wire u2__abc_44228_n7927_1;
  wire u2__abc_44228_n7928_1;
  wire u2__abc_44228_n7929;
  wire u2__abc_44228_n7930;
  wire u2__abc_44228_n7931;
  wire u2__abc_44228_n7932;
  wire u2__abc_44228_n7933_1;
  wire u2__abc_44228_n7934;
  wire u2__abc_44228_n7935;
  wire u2__abc_44228_n7936;
  wire u2__abc_44228_n7937;
  wire u2__abc_44228_n7938_1;
  wire u2__abc_44228_n7939_1;
  wire u2__abc_44228_n7940;
  wire u2__abc_44228_n7941;
  wire u2__abc_44228_n7943;
  wire u2__abc_44228_n7944_1;
  wire u2__abc_44228_n7945;
  wire u2__abc_44228_n7946;
  wire u2__abc_44228_n7947;
  wire u2__abc_44228_n7948;
  wire u2__abc_44228_n7949_1;
  wire u2__abc_44228_n7950_1;
  wire u2__abc_44228_n7951;
  wire u2__abc_44228_n7952;
  wire u2__abc_44228_n7953;
  wire u2__abc_44228_n7954;
  wire u2__abc_44228_n7955_1;
  wire u2__abc_44228_n7956;
  wire u2__abc_44228_n7957;
  wire u2__abc_44228_n7958;
  wire u2__abc_44228_n7960_1;
  wire u2__abc_44228_n7961_1;
  wire u2__abc_44228_n7962;
  wire u2__abc_44228_n7963;
  wire u2__abc_44228_n7964;
  wire u2__abc_44228_n7965;
  wire u2__abc_44228_n7966_1;
  wire u2__abc_44228_n7967;
  wire u2__abc_44228_n7968;
  wire u2__abc_44228_n7969;
  wire u2__abc_44228_n7970;
  wire u2__abc_44228_n7971_1;
  wire u2__abc_44228_n7972_1;
  wire u2__abc_44228_n7973;
  wire u2__abc_44228_n7974;
  wire u2__abc_44228_n7975;
  wire u2__abc_44228_n7977_1;
  wire u2__abc_44228_n7978;
  wire u2__abc_44228_n7979;
  wire u2__abc_44228_n7980;
  wire u2__abc_44228_n7981;
  wire u2__abc_44228_n7982_1;
  wire u2__abc_44228_n7983_1;
  wire u2__abc_44228_n7984;
  wire u2__abc_44228_n7985;
  wire u2__abc_44228_n7986;
  wire u2__abc_44228_n7987;
  wire u2__abc_44228_n7988_1;
  wire u2__abc_44228_n7989;
  wire u2__abc_44228_n7990;
  wire u2__abc_44228_n7991;
  wire u2__abc_44228_n7992;
  wire u2__abc_44228_n7994_1;
  wire u2__abc_44228_n7995;
  wire u2__abc_44228_n7996;
  wire u2__abc_44228_n7997;
  wire u2__abc_44228_n7998;
  wire u2__abc_44228_n7999_1;
  wire u2__abc_44228_n8000;
  wire u2__abc_44228_n8001;
  wire u2__abc_44228_n8002;
  wire u2__abc_44228_n8003;
  wire u2__abc_44228_n8004_1;
  wire u2__abc_44228_n8005_1;
  wire u2__abc_44228_n8006;
  wire u2__abc_44228_n8007;
  wire u2__abc_44228_n8008;
  wire u2__abc_44228_n8009;
  wire u2__abc_44228_n8011;
  wire u2__abc_44228_n8012;
  wire u2__abc_44228_n8013;
  wire u2__abc_44228_n8014;
  wire u2__abc_44228_n8015_1;
  wire u2__abc_44228_n8016_1;
  wire u2__abc_44228_n8017;
  wire u2__abc_44228_n8018;
  wire u2__abc_44228_n8019;
  wire u2__abc_44228_n8020;
  wire u2__abc_44228_n8021_1;
  wire u2__abc_44228_n8022;
  wire u2__abc_44228_n8023;
  wire u2__abc_44228_n8024;
  wire u2__abc_44228_n8025;
  wire u2__abc_44228_n8026_1;
  wire u2__abc_44228_n8027_1;
  wire u2__abc_44228_n8029;
  wire u2__abc_44228_n8030;
  wire u2__abc_44228_n8031;
  wire u2__abc_44228_n8032_1;
  wire u2__abc_44228_n8033;
  wire u2__abc_44228_n8034;
  wire u2__abc_44228_n8035;
  wire u2__abc_44228_n8036;
  wire u2__abc_44228_n8037_1;
  wire u2__abc_44228_n8038_1;
  wire u2__abc_44228_n8039;
  wire u2__abc_44228_n8040;
  wire u2__abc_44228_n8041;
  wire u2__abc_44228_n8042;
  wire u2__abc_44228_n8043_1;
  wire u2__abc_44228_n8044;
  wire u2__abc_44228_n8046;
  wire u2__abc_44228_n8047;
  wire u2__abc_44228_n8048_1;
  wire u2__abc_44228_n8049_1;
  wire u2__abc_44228_n8050;
  wire u2__abc_44228_n8051;
  wire u2__abc_44228_n8052;
  wire u2__abc_44228_n8053;
  wire u2__abc_44228_n8054_1;
  wire u2__abc_44228_n8055;
  wire u2__abc_44228_n8056;
  wire u2__abc_44228_n8057;
  wire u2__abc_44228_n8058;
  wire u2__abc_44228_n8059_1;
  wire u2__abc_44228_n8060_1;
  wire u2__abc_44228_n8061;
  wire u2__abc_44228_n8062;
  wire u2__abc_44228_n8064;
  wire u2__abc_44228_n8065_1;
  wire u2__abc_44228_n8066;
  wire u2__abc_44228_n8067;
  wire u2__abc_44228_n8068;
  wire u2__abc_44228_n8069;
  wire u2__abc_44228_n8070_1;
  wire u2__abc_44228_n8071_1;
  wire u2__abc_44228_n8072;
  wire u2__abc_44228_n8073;
  wire u2__abc_44228_n8074;
  wire u2__abc_44228_n8075;
  wire u2__abc_44228_n8076_1;
  wire u2__abc_44228_n8077;
  wire u2__abc_44228_n8078;
  wire u2__abc_44228_n8079;
  wire u2__abc_44228_n8081_1;
  wire u2__abc_44228_n8082_1;
  wire u2__abc_44228_n8083;
  wire u2__abc_44228_n8084;
  wire u2__abc_44228_n8085;
  wire u2__abc_44228_n8086;
  wire u2__abc_44228_n8087_1;
  wire u2__abc_44228_n8088;
  wire u2__abc_44228_n8089;
  wire u2__abc_44228_n8090;
  wire u2__abc_44228_n8091;
  wire u2__abc_44228_n8092_1;
  wire u2__abc_44228_n8093_1;
  wire u2__abc_44228_n8094;
  wire u2__abc_44228_n8096;
  wire u2__abc_44228_n8097;
  wire u2__abc_44228_n8098_1;
  wire u2__abc_44228_n8099;
  wire u2__abc_44228_n8100;
  wire u2__abc_44228_n8101;
  wire u2__abc_44228_n8102;
  wire u2__abc_44228_n8103_1;
  wire u2__abc_44228_n8104_1;
  wire u2__abc_44228_n8105;
  wire u2__abc_44228_n8106;
  wire u2__abc_44228_n8107;
  wire u2__abc_44228_n8108;
  wire u2__abc_44228_n8109_1;
  wire u2__abc_44228_n8110;
  wire u2__abc_44228_n8111;
  wire u2__abc_44228_n8113;
  wire u2__abc_44228_n8114_1;
  wire u2__abc_44228_n8115_1;
  wire u2__abc_44228_n8116;
  wire u2__abc_44228_n8117;
  wire u2__abc_44228_n8118;
  wire u2__abc_44228_n8119;
  wire u2__abc_44228_n8120_1;
  wire u2__abc_44228_n8121;
  wire u2__abc_44228_n8122;
  wire u2__abc_44228_n8123;
  wire u2__abc_44228_n8124;
  wire u2__abc_44228_n8125_1;
  wire u2__abc_44228_n8126_1;
  wire u2__abc_44228_n8127;
  wire u2__abc_44228_n8128;
  wire u2__abc_44228_n8130;
  wire u2__abc_44228_n8131_1;
  wire u2__abc_44228_n8132;
  wire u2__abc_44228_n8133;
  wire u2__abc_44228_n8134;
  wire u2__abc_44228_n8135;
  wire u2__abc_44228_n8136_1;
  wire u2__abc_44228_n8137_1;
  wire u2__abc_44228_n8138;
  wire u2__abc_44228_n8139;
  wire u2__abc_44228_n8140;
  wire u2__abc_44228_n8141;
  wire u2__abc_44228_n8142_1;
  wire u2__abc_44228_n8143;
  wire u2__abc_44228_n8144;
  wire u2__abc_44228_n8145;
  wire u2__abc_44228_n8147_1;
  wire u2__abc_44228_n8148_1;
  wire u2__abc_44228_n8149;
  wire u2__abc_44228_n8150;
  wire u2__abc_44228_n8151;
  wire u2__abc_44228_n8152;
  wire u2__abc_44228_n8153_1;
  wire u2__abc_44228_n8154;
  wire u2__abc_44228_n8155;
  wire u2__abc_44228_n8156;
  wire u2__abc_44228_n8157;
  wire u2__abc_44228_n8158_1;
  wire u2__abc_44228_n8159_1;
  wire u2__abc_44228_n8160;
  wire u2__abc_44228_n8161;
  wire u2__abc_44228_n8162;
  wire u2__abc_44228_n8164_1;
  wire u2__abc_44228_n8165;
  wire u2__abc_44228_n8166;
  wire u2__abc_44228_n8167;
  wire u2__abc_44228_n8168;
  wire u2__abc_44228_n8169_1;
  wire u2__abc_44228_n8170_1;
  wire u2__abc_44228_n8171;
  wire u2__abc_44228_n8172;
  wire u2__abc_44228_n8173;
  wire u2__abc_44228_n8174;
  wire u2__abc_44228_n8175_1;
  wire u2__abc_44228_n8176;
  wire u2__abc_44228_n8177;
  wire u2__abc_44228_n8178;
  wire u2__abc_44228_n8179;
  wire u2__abc_44228_n8181_1;
  wire u2__abc_44228_n8182;
  wire u2__abc_44228_n8183;
  wire u2__abc_44228_n8184;
  wire u2__abc_44228_n8185;
  wire u2__abc_44228_n8186_1;
  wire u2__abc_44228_n8187;
  wire u2__abc_44228_n8188;
  wire u2__abc_44228_n8189;
  wire u2__abc_44228_n8190;
  wire u2__abc_44228_n8191_1;
  wire u2__abc_44228_n8192_1;
  wire u2__abc_44228_n8193;
  wire u2__abc_44228_n8194;
  wire u2__abc_44228_n8195;
  wire u2__abc_44228_n8196;
  wire u2__abc_44228_n8197_1;
  wire u2__abc_44228_n8199;
  wire u2__abc_44228_n8200;
  wire u2__abc_44228_n8201;
  wire u2__abc_44228_n8202_1;
  wire u2__abc_44228_n8203_1;
  wire u2__abc_44228_n8204;
  wire u2__abc_44228_n8205;
  wire u2__abc_44228_n8206;
  wire u2__abc_44228_n8207;
  wire u2__abc_44228_n8208_1;
  wire u2__abc_44228_n8209;
  wire u2__abc_44228_n8209_bF_buf0;
  wire u2__abc_44228_n8209_bF_buf1;
  wire u2__abc_44228_n8209_bF_buf2;
  wire u2__abc_44228_n8209_bF_buf3;
  wire u2__abc_44228_n8209_bF_buf4;
  wire u2__abc_44228_n8209_bF_buf5;
  wire u2__abc_44228_n8209_bF_buf6;
  wire u2__abc_44228_n8209_bF_buf7;
  wire u2__abc_44228_n8209_bF_buf8;
  wire u2__abc_44228_n8209_bF_buf9;
  wire u2__abc_44228_n8210;
  wire u2__abc_44228_n8211;
  wire u2__abc_44228_n8212;
  wire u2__abc_44228_n8213_1;
  wire u2__abc_44228_n8214_1;
  wire u2__abc_44228_n8215;
  wire u2__abc_44228_n8216;
  wire u2__abc_44228_n8217;
  wire u2__abc_44228_n8219_1;
  wire u2__abc_44228_n8220;
  wire u2__abc_44228_n8221;
  wire u2__abc_44228_n8222;
  wire u2__abc_44228_n8223;
  wire u2__abc_44228_n8224_1;
  wire u2__abc_44228_n8225_1;
  wire u2__abc_44228_n8226;
  wire u2__abc_44228_n8227;
  wire u2__abc_44228_n8228;
  wire u2__abc_44228_n8229;
  wire u2__abc_44228_n8230_1;
  wire u2__abc_44228_n8231;
  wire u2__abc_44228_n8232;
  wire u2__abc_44228_n8233;
  wire u2__abc_44228_n8234;
  wire u2__abc_44228_n8236_1;
  wire u2__abc_44228_n8237;
  wire u2__abc_44228_n8238;
  wire u2__abc_44228_n8239;
  wire u2__abc_44228_n8240;
  wire u2__abc_44228_n8241_1;
  wire u2__abc_44228_n8242;
  wire u2__abc_44228_n8243;
  wire u2__abc_44228_n8244;
  wire u2__abc_44228_n8245;
  wire u2__abc_44228_n8246_1;
  wire u2__abc_44228_n8247_1;
  wire u2__abc_44228_n8248;
  wire u2__abc_44228_n8249;
  wire u2__abc_44228_n8250;
  wire u2__abc_44228_n8251;
  wire u2__abc_44228_n8253;
  wire u2__abc_44228_n8254;
  wire u2__abc_44228_n8255;
  wire u2__abc_44228_n8256;
  wire u2__abc_44228_n8257_1;
  wire u2__abc_44228_n8258_1;
  wire u2__abc_44228_n8259;
  wire u2__abc_44228_n8260;
  wire u2__abc_44228_n8261;
  wire u2__abc_44228_n8262;
  wire u2__abc_44228_n8263_1;
  wire u2__abc_44228_n8264;
  wire u2__abc_44228_n8265;
  wire u2__abc_44228_n8266;
  wire u2__abc_44228_n8267;
  wire u2__abc_44228_n8268_1;
  wire u2__abc_44228_n8270;
  wire u2__abc_44228_n8271;
  wire u2__abc_44228_n8272;
  wire u2__abc_44228_n8273;
  wire u2__abc_44228_n8274_1;
  wire u2__abc_44228_n8275;
  wire u2__abc_44228_n8276;
  wire u2__abc_44228_n8277;
  wire u2__abc_44228_n8278;
  wire u2__abc_44228_n8279_1;
  wire u2__abc_44228_n8280_1;
  wire u2__abc_44228_n8281;
  wire u2__abc_44228_n8282;
  wire u2__abc_44228_n8283;
  wire u2__abc_44228_n8284;
  wire u2__abc_44228_n8285_1;
  wire u2__abc_44228_n8287;
  wire u2__abc_44228_n8288;
  wire u2__abc_44228_n8289;
  wire u2__abc_44228_n8290_1;
  wire u2__abc_44228_n8291_1;
  wire u2__abc_44228_n8292;
  wire u2__abc_44228_n8293;
  wire u2__abc_44228_n8294;
  wire u2__abc_44228_n8295;
  wire u2__abc_44228_n8296_1;
  wire u2__abc_44228_n8297;
  wire u2__abc_44228_n8298;
  wire u2__abc_44228_n8299;
  wire u2__abc_44228_n8300;
  wire u2__abc_44228_n8301_1;
  wire u2__abc_44228_n8302_1;
  wire u2__abc_44228_n8303;
  wire u2__abc_44228_n8305;
  wire u2__abc_44228_n8306;
  wire u2__abc_44228_n8307_1;
  wire u2__abc_44228_n8308;
  wire u2__abc_44228_n8309;
  wire u2__abc_44228_n8310;
  wire u2__abc_44228_n8311;
  wire u2__abc_44228_n8312_1;
  wire u2__abc_44228_n8313_1;
  wire u2__abc_44228_n8314;
  wire u2__abc_44228_n8315;
  wire u2__abc_44228_n8316;
  wire u2__abc_44228_n8317;
  wire u2__abc_44228_n8318_1;
  wire u2__abc_44228_n8319;
  wire u2__abc_44228_n8320;
  wire u2__abc_44228_n8322;
  wire u2__abc_44228_n8323_1;
  wire u2__abc_44228_n8324_1;
  wire u2__abc_44228_n8325;
  wire u2__abc_44228_n8326;
  wire u2__abc_44228_n8327;
  wire u2__abc_44228_n8328;
  wire u2__abc_44228_n8329_1;
  wire u2__abc_44228_n8330;
  wire u2__abc_44228_n8331;
  wire u2__abc_44228_n8332;
  wire u2__abc_44228_n8333;
  wire u2__abc_44228_n8334_1;
  wire u2__abc_44228_n8335_1;
  wire u2__abc_44228_n8336;
  wire u2__abc_44228_n8337;
  wire u2__abc_44228_n8338;
  wire u2__abc_44228_n8340_1;
  wire u2__abc_44228_n8341;
  wire u2__abc_44228_n8342;
  wire u2__abc_44228_n8343;
  wire u2__abc_44228_n8344;
  wire u2__abc_44228_n8345_1;
  wire u2__abc_44228_n8346_1;
  wire u2__abc_44228_n8347;
  wire u2__abc_44228_n8348;
  wire u2__abc_44228_n8349;
  wire u2__abc_44228_n8350;
  wire u2__abc_44228_n8351_1;
  wire u2__abc_44228_n8352;
  wire u2__abc_44228_n8353;
  wire u2__abc_44228_n8354;
  wire u2__abc_44228_n8355;
  wire u2__abc_44228_n8357_1;
  wire u2__abc_44228_n8358;
  wire u2__abc_44228_n8359;
  wire u2__abc_44228_n8360;
  wire u2__abc_44228_n8361;
  wire u2__abc_44228_n8362_1;
  wire u2__abc_44228_n8363;
  wire u2__abc_44228_n8364;
  wire u2__abc_44228_n8365;
  wire u2__abc_44228_n8366;
  wire u2__abc_44228_n8367_1;
  wire u2__abc_44228_n8368_1;
  wire u2__abc_44228_n8369;
  wire u2__abc_44228_n8370;
  wire u2__abc_44228_n8371;
  wire u2__abc_44228_n8372;
  wire u2__abc_44228_n8374;
  wire u2__abc_44228_n8375;
  wire u2__abc_44228_n8376;
  wire u2__abc_44228_n8377;
  wire u2__abc_44228_n8378_1;
  wire u2__abc_44228_n8379_1;
  wire u2__abc_44228_n8380;
  wire u2__abc_44228_n8381;
  wire u2__abc_44228_n8382;
  wire u2__abc_44228_n8383;
  wire u2__abc_44228_n8384_1;
  wire u2__abc_44228_n8385;
  wire u2__abc_44228_n8386;
  wire u2__abc_44228_n8387;
  wire u2__abc_44228_n8388;
  wire u2__abc_44228_n8389_1;
  wire u2__abc_44228_n8391;
  wire u2__abc_44228_n8392;
  wire u2__abc_44228_n8393;
  wire u2__abc_44228_n8394;
  wire u2__abc_44228_n8395_1;
  wire u2__abc_44228_n8396;
  wire u2__abc_44228_n8397;
  wire u2__abc_44228_n8398;
  wire u2__abc_44228_n8399;
  wire u2__abc_44228_n8400_1;
  wire u2__abc_44228_n8401_1;
  wire u2__abc_44228_n8402;
  wire u2__abc_44228_n8403;
  wire u2__abc_44228_n8404;
  wire u2__abc_44228_n8405;
  wire u2__abc_44228_n8406_1;
  wire u2__abc_44228_n8408;
  wire u2__abc_44228_n8409;
  wire u2__abc_44228_n8410;
  wire u2__abc_44228_n8411_1;
  wire u2__abc_44228_n8412_1;
  wire u2__abc_44228_n8413;
  wire u2__abc_44228_n8414;
  wire u2__abc_44228_n8415;
  wire u2__abc_44228_n8416;
  wire u2__abc_44228_n8417_1;
  wire u2__abc_44228_n8418;
  wire u2__abc_44228_n8419;
  wire u2__abc_44228_n8420;
  wire u2__abc_44228_n8421;
  wire u2__abc_44228_n8422_1;
  wire u2__abc_44228_n8423_1;
  wire u2__abc_44228_n8425;
  wire u2__abc_44228_n8426;
  wire u2__abc_44228_n8427;
  wire u2__abc_44228_n8428_1;
  wire u2__abc_44228_n8429;
  wire u2__abc_44228_n8430;
  wire u2__abc_44228_n8431;
  wire u2__abc_44228_n8432;
  wire u2__abc_44228_n8433_1;
  wire u2__abc_44228_n8434_1;
  wire u2__abc_44228_n8435;
  wire u2__abc_44228_n8436;
  wire u2__abc_44228_n8437;
  wire u2__abc_44228_n8438;
  wire u2__abc_44228_n8439_1;
  wire u2__abc_44228_n8440;
  wire u2__abc_44228_n8442;
  wire u2__abc_44228_n8443;
  wire u2__abc_44228_n8444_1;
  wire u2__abc_44228_n8445_1;
  wire u2__abc_44228_n8446;
  wire u2__abc_44228_n8447;
  wire u2__abc_44228_n8448;
  wire u2__abc_44228_n8449;
  wire u2__abc_44228_n8450_1;
  wire u2__abc_44228_n8451;
  wire u2__abc_44228_n8452;
  wire u2__abc_44228_n8453;
  wire u2__abc_44228_n8454;
  wire u2__abc_44228_n8455_1;
  wire u2__abc_44228_n8456_1;
  wire u2__abc_44228_n8457;
  wire u2__abc_44228_n8459;
  wire u2__abc_44228_n8460;
  wire u2__abc_44228_n8461_1;
  wire u2__abc_44228_n8462;
  wire u2__abc_44228_n8463;
  wire u2__abc_44228_n8464;
  wire u2__abc_44228_n8465;
  wire u2__abc_44228_n8466_1;
  wire u2__abc_44228_n8467_1;
  wire u2__abc_44228_n8468;
  wire u2__abc_44228_n8469;
  wire u2__abc_44228_n8470;
  wire u2__abc_44228_n8471;
  wire u2__abc_44228_n8472_1;
  wire u2__abc_44228_n8473;
  wire u2__abc_44228_n8474;
  wire u2__abc_44228_n8475;
  wire u2__abc_44228_n8477_1;
  wire u2__abc_44228_n8478_1;
  wire u2__abc_44228_n8479;
  wire u2__abc_44228_n8480;
  wire u2__abc_44228_n8481;
  wire u2__abc_44228_n8482;
  wire u2__abc_44228_n8483_1;
  wire u2__abc_44228_n8484;
  wire u2__abc_44228_n8485;
  wire u2__abc_44228_n8486;
  wire u2__abc_44228_n8487;
  wire u2__abc_44228_n8488_1;
  wire u2__abc_44228_n8489_1;
  wire u2__abc_44228_n8490;
  wire u2__abc_44228_n8491;
  wire u2__abc_44228_n8492;
  wire u2__abc_44228_n8494_1;
  wire u2__abc_44228_n8495;
  wire u2__abc_44228_n8496;
  wire u2__abc_44228_n8497;
  wire u2__abc_44228_n8498;
  wire u2__abc_44228_n8499_1;
  wire u2__abc_44228_n8500_1;
  wire u2__abc_44228_n8501;
  wire u2__abc_44228_n8502;
  wire u2__abc_44228_n8503;
  wire u2__abc_44228_n8504;
  wire u2__abc_44228_n8505_1;
  wire u2__abc_44228_n8506;
  wire u2__abc_44228_n8507;
  wire u2__abc_44228_n8508;
  wire u2__abc_44228_n8509;
  wire u2__abc_44228_n8511_1;
  wire u2__abc_44228_n8512;
  wire u2__abc_44228_n8513;
  wire u2__abc_44228_n8514;
  wire u2__abc_44228_n8515;
  wire u2__abc_44228_n8516_1;
  wire u2__abc_44228_n8517;
  wire u2__abc_44228_n8518;
  wire u2__abc_44228_n8519;
  wire u2__abc_44228_n8520;
  wire u2__abc_44228_n8521_1;
  wire u2__abc_44228_n8522_1;
  wire u2__abc_44228_n8523;
  wire u2__abc_44228_n8524;
  wire u2__abc_44228_n8525;
  wire u2__abc_44228_n8526;
  wire u2__abc_44228_n8528;
  wire u2__abc_44228_n8529;
  wire u2__abc_44228_n8530;
  wire u2__abc_44228_n8531;
  wire u2__abc_44228_n8532_1;
  wire u2__abc_44228_n8533_1;
  wire u2__abc_44228_n8534;
  wire u2__abc_44228_n8535;
  wire u2__abc_44228_n8536;
  wire u2__abc_44228_n8537;
  wire u2__abc_44228_n8538_1;
  wire u2__abc_44228_n8539;
  wire u2__abc_44228_n8540;
  wire u2__abc_44228_n8541;
  wire u2__abc_44228_n8542;
  wire u2__abc_44228_n8543_1;
  wire u2__abc_44228_n8545;
  wire u2__abc_44228_n8546;
  wire u2__abc_44228_n8547;
  wire u2__abc_44228_n8548;
  wire u2__abc_44228_n8549_1;
  wire u2__abc_44228_n8550;
  wire u2__abc_44228_n8551;
  wire u2__abc_44228_n8552;
  wire u2__abc_44228_n8553;
  wire u2__abc_44228_n8554_1;
  wire u2__abc_44228_n8555_1;
  wire u2__abc_44228_n8556;
  wire u2__abc_44228_n8557;
  wire u2__abc_44228_n8558;
  wire u2__abc_44228_n8559;
  wire u2__abc_44228_n8560_1;
  wire u2__abc_44228_n8562;
  wire u2__abc_44228_n8563;
  wire u2__abc_44228_n8564;
  wire u2__abc_44228_n8565_1;
  wire u2__abc_44228_n8566_1;
  wire u2__abc_44228_n8567;
  wire u2__abc_44228_n8568;
  wire u2__abc_44228_n8569;
  wire u2__abc_44228_n8570;
  wire u2__abc_44228_n8571_1;
  wire u2__abc_44228_n8572;
  wire u2__abc_44228_n8573;
  wire u2__abc_44228_n8574;
  wire u2__abc_44228_n8575;
  wire u2__abc_44228_n8576_1;
  wire u2__abc_44228_n8577_1;
  wire u2__abc_44228_n8578;
  wire u2__abc_44228_n8580;
  wire u2__abc_44228_n8581;
  wire u2__abc_44228_n8582_1;
  wire u2__abc_44228_n8583;
  wire u2__abc_44228_n8584;
  wire u2__abc_44228_n8585;
  wire u2__abc_44228_n8586;
  wire u2__abc_44228_n8587_1;
  wire u2__abc_44228_n8588_1;
  wire u2__abc_44228_n8589;
  wire u2__abc_44228_n8590;
  wire u2__abc_44228_n8591;
  wire u2__abc_44228_n8592;
  wire u2__abc_44228_n8593_1;
  wire u2__abc_44228_n8594;
  wire u2__abc_44228_n8595;
  wire u2__abc_44228_n8597;
  wire u2__abc_44228_n8598_1;
  wire u2__abc_44228_n8599_1;
  wire u2__abc_44228_n8600;
  wire u2__abc_44228_n8601;
  wire u2__abc_44228_n8602;
  wire u2__abc_44228_n8603;
  wire u2__abc_44228_n8604_1;
  wire u2__abc_44228_n8605;
  wire u2__abc_44228_n8606;
  wire u2__abc_44228_n8607;
  wire u2__abc_44228_n8608;
  wire u2__abc_44228_n8609_1;
  wire u2__abc_44228_n8610_1;
  wire u2__abc_44228_n8611;
  wire u2__abc_44228_n8612;
  wire u2__abc_44228_n8613;
  wire u2__abc_44228_n8615_1;
  wire u2__abc_44228_n8616;
  wire u2__abc_44228_n8617;
  wire u2__abc_44228_n8618;
  wire u2__abc_44228_n8619;
  wire u2__abc_44228_n8620_1;
  wire u2__abc_44228_n8621_1;
  wire u2__abc_44228_n8622;
  wire u2__abc_44228_n8623;
  wire u2__abc_44228_n8624;
  wire u2__abc_44228_n8625;
  wire u2__abc_44228_n8626_1;
  wire u2__abc_44228_n8627;
  wire u2__abc_44228_n8628;
  wire u2__abc_44228_n8629;
  wire u2__abc_44228_n8630;
  wire u2__abc_44228_n8632_1;
  wire u2__abc_44228_n8633;
  wire u2__abc_44228_n8634;
  wire u2__abc_44228_n8635;
  wire u2__abc_44228_n8636;
  wire u2__abc_44228_n8637_1;
  wire u2__abc_44228_n8638;
  wire u2__abc_44228_n8639;
  wire u2__abc_44228_n8640;
  wire u2__abc_44228_n8641;
  wire u2__abc_44228_n8642_1;
  wire u2__abc_44228_n8643_1;
  wire u2__abc_44228_n8644;
  wire u2__abc_44228_n8645;
  wire u2__abc_44228_n8647;
  wire u2__abc_44228_n8648_1;
  wire u2__abc_44228_n8649;
  wire u2__abc_44228_n8650;
  wire u2__abc_44228_n8651;
  wire u2__abc_44228_n8652;
  wire u2__abc_44228_n8653_1;
  wire u2__abc_44228_n8654_1;
  wire u2__abc_44228_n8655;
  wire u2__abc_44228_n8656;
  wire u2__abc_44228_n8657;
  wire u2__abc_44228_n8658;
  wire u2__abc_44228_n8659_1;
  wire u2__abc_44228_n8660;
  wire u2__abc_44228_n8661;
  wire u2__abc_44228_n8662;
  wire u2__abc_44228_n8664_1;
  wire u2__abc_44228_n8665_1;
  wire u2__abc_44228_n8666;
  wire u2__abc_44228_n8667;
  wire u2__abc_44228_n8668;
  wire u2__abc_44228_n8669;
  wire u2__abc_44228_n8670_1;
  wire u2__abc_44228_n8671;
  wire u2__abc_44228_n8672;
  wire u2__abc_44228_n8673;
  wire u2__abc_44228_n8674;
  wire u2__abc_44228_n8675_1;
  wire u2__abc_44228_n8676_1;
  wire u2__abc_44228_n8677;
  wire u2__abc_44228_n8678;
  wire u2__abc_44228_n8679;
  wire u2__abc_44228_n8681_1;
  wire u2__abc_44228_n8682;
  wire u2__abc_44228_n8683;
  wire u2__abc_44228_n8684;
  wire u2__abc_44228_n8685;
  wire u2__abc_44228_n8686_1;
  wire u2__abc_44228_n8687_1;
  wire u2__abc_44228_n8688;
  wire u2__abc_44228_n8689;
  wire u2__abc_44228_n8690;
  wire u2__abc_44228_n8691;
  wire u2__abc_44228_n8692_1;
  wire u2__abc_44228_n8693;
  wire u2__abc_44228_n8694;
  wire u2__abc_44228_n8695;
  wire u2__abc_44228_n8696;
  wire u2__abc_44228_n8698_1;
  wire u2__abc_44228_n8699;
  wire u2__abc_44228_n8700;
  wire u2__abc_44228_n8701;
  wire u2__abc_44228_n8702;
  wire u2__abc_44228_n8703_1;
  wire u2__abc_44228_n8704;
  wire u2__abc_44228_n8705;
  wire u2__abc_44228_n8706;
  wire u2__abc_44228_n8707;
  wire u2__abc_44228_n8708_1;
  wire u2__abc_44228_n8709_1;
  wire u2__abc_44228_n8710;
  wire u2__abc_44228_n8711;
  wire u2__abc_44228_n8712;
  wire u2__abc_44228_n8713;
  wire u2__abc_44228_n8715;
  wire u2__abc_44228_n8716;
  wire u2__abc_44228_n8717;
  wire u2__abc_44228_n8718;
  wire u2__abc_44228_n8719_1;
  wire u2__abc_44228_n8720_1;
  wire u2__abc_44228_n8721;
  wire u2__abc_44228_n8722;
  wire u2__abc_44228_n8723;
  wire u2__abc_44228_n8724;
  wire u2__abc_44228_n8725_1;
  wire u2__abc_44228_n8726;
  wire u2__abc_44228_n8727;
  wire u2__abc_44228_n8728;
  wire u2__abc_44228_n8729;
  wire u2__abc_44228_n8730_1;
  wire u2__abc_44228_n8732;
  wire u2__abc_44228_n8733;
  wire u2__abc_44228_n8734;
  wire u2__abc_44228_n8735;
  wire u2__abc_44228_n8736_1;
  wire u2__abc_44228_n8737;
  wire u2__abc_44228_n8738;
  wire u2__abc_44228_n8739;
  wire u2__abc_44228_n8740;
  wire u2__abc_44228_n8741_1;
  wire u2__abc_44228_n8742_1;
  wire u2__abc_44228_n8743;
  wire u2__abc_44228_n8744;
  wire u2__abc_44228_n8745;
  wire u2__abc_44228_n8746;
  wire u2__abc_44228_n8747_1;
  wire u2__abc_44228_n8749;
  wire u2__abc_44228_n8750;
  wire u2__abc_44228_n8751;
  wire u2__abc_44228_n8752_1;
  wire u2__abc_44228_n8753_1;
  wire u2__abc_44228_n8754;
  wire u2__abc_44228_n8755;
  wire u2__abc_44228_n8756;
  wire u2__abc_44228_n8757;
  wire u2__abc_44228_n8758_1;
  wire u2__abc_44228_n8759;
  wire u2__abc_44228_n8760;
  wire u2__abc_44228_n8761;
  wire u2__abc_44228_n8762;
  wire u2__abc_44228_n8763_1;
  wire u2__abc_44228_n8764_1;
  wire u2__abc_44228_n8766;
  wire u2__abc_44228_n8767;
  wire u2__abc_44228_n8768;
  wire u2__abc_44228_n8769_1;
  wire u2__abc_44228_n8770;
  wire u2__abc_44228_n8771;
  wire u2__abc_44228_n8772;
  wire u2__abc_44228_n8773;
  wire u2__abc_44228_n8774_1;
  wire u2__abc_44228_n8775_1;
  wire u2__abc_44228_n8776;
  wire u2__abc_44228_n8777;
  wire u2__abc_44228_n8778;
  wire u2__abc_44228_n8779;
  wire u2__abc_44228_n8780_1;
  wire u2__abc_44228_n8781;
  wire u2__abc_44228_n8783;
  wire u2__abc_44228_n8784;
  wire u2__abc_44228_n8785_1;
  wire u2__abc_44228_n8786_1;
  wire u2__abc_44228_n8787;
  wire u2__abc_44228_n8788;
  wire u2__abc_44228_n8789;
  wire u2__abc_44228_n8790;
  wire u2__abc_44228_n8791_1;
  wire u2__abc_44228_n8792;
  wire u2__abc_44228_n8793;
  wire u2__abc_44228_n8794;
  wire u2__abc_44228_n8795;
  wire u2__abc_44228_n8796_1;
  wire u2__abc_44228_n8797_1;
  wire u2__abc_44228_n8798;
  wire u2__abc_44228_n8800;
  wire u2__abc_44228_n8801;
  wire u2__abc_44228_n8802_1;
  wire u2__abc_44228_n8803;
  wire u2__abc_44228_n8804;
  wire u2__abc_44228_n8805;
  wire u2__abc_44228_n8806;
  wire u2__abc_44228_n8807_1;
  wire u2__abc_44228_n8808_1;
  wire u2__abc_44228_n8809;
  wire u2__abc_44228_n8810;
  wire u2__abc_44228_n8811;
  wire u2__abc_44228_n8812;
  wire u2__abc_44228_n8813_1;
  wire u2__abc_44228_n8814;
  wire u2__abc_44228_n8815;
  wire u2__abc_44228_n8817;
  wire u2__abc_44228_n8818_1;
  wire u2__abc_44228_n8819_1;
  wire u2__abc_44228_n8820;
  wire u2__abc_44228_n8821;
  wire u2__abc_44228_n8822;
  wire u2__abc_44228_n8823;
  wire u2__abc_44228_n8824_1;
  wire u2__abc_44228_n8825;
  wire u2__abc_44228_n8826;
  wire u2__abc_44228_n8827;
  wire u2__abc_44228_n8828;
  wire u2__abc_44228_n8829_1;
  wire u2__abc_44228_n8830_1;
  wire u2__abc_44228_n8831;
  wire u2__abc_44228_n8832;
  wire u2__abc_44228_n8834;
  wire u2__abc_44228_n8835_1;
  wire u2__abc_44228_n8836;
  wire u2__abc_44228_n8837;
  wire u2__abc_44228_n8838;
  wire u2__abc_44228_n8839;
  wire u2__abc_44228_n8840_1;
  wire u2__abc_44228_n8841_1;
  wire u2__abc_44228_n8842;
  wire u2__abc_44228_n8843;
  wire u2__abc_44228_n8844;
  wire u2__abc_44228_n8845;
  wire u2__abc_44228_n8846_1;
  wire u2__abc_44228_n8847;
  wire u2__abc_44228_n8848;
  wire u2__abc_44228_n8849;
  wire u2__abc_44228_n8850;
  wire u2__abc_44228_n8852_1;
  wire u2__abc_44228_n8853;
  wire u2__abc_44228_n8854;
  wire u2__abc_44228_n8855;
  wire u2__abc_44228_n8856;
  wire u2__abc_44228_n8857_1;
  wire u2__abc_44228_n8858;
  wire u2__abc_44228_n8859;
  wire u2__abc_44228_n8860;
  wire u2__abc_44228_n8861;
  wire u2__abc_44228_n8862_1;
  wire u2__abc_44228_n8863_1;
  wire u2__abc_44228_n8864;
  wire u2__abc_44228_n8865;
  wire u2__abc_44228_n8866;
  wire u2__abc_44228_n8867;
  wire u2__abc_44228_n8869;
  wire u2__abc_44228_n8870;
  wire u2__abc_44228_n8871;
  wire u2__abc_44228_n8872;
  wire u2__abc_44228_n8873_1;
  wire u2__abc_44228_n8874_1;
  wire u2__abc_44228_n8875;
  wire u2__abc_44228_n8876;
  wire u2__abc_44228_n8877;
  wire u2__abc_44228_n8878;
  wire u2__abc_44228_n8879_1;
  wire u2__abc_44228_n8880;
  wire u2__abc_44228_n8881;
  wire u2__abc_44228_n8882;
  wire u2__abc_44228_n8883;
  wire u2__abc_44228_n8884_1;
  wire u2__abc_44228_n8885_1;
  wire u2__abc_44228_n8887;
  wire u2__abc_44228_n8888;
  wire u2__abc_44228_n8889;
  wire u2__abc_44228_n8890_1;
  wire u2__abc_44228_n8891;
  wire u2__abc_44228_n8892;
  wire u2__abc_44228_n8893;
  wire u2__abc_44228_n8894;
  wire u2__abc_44228_n8895_1;
  wire u2__abc_44228_n8896_1;
  wire u2__abc_44228_n8897;
  wire u2__abc_44228_n8898;
  wire u2__abc_44228_n8899;
  wire u2__abc_44228_n8900;
  wire u2__abc_44228_n8901_1;
  wire u2__abc_44228_n8902;
  wire u2__abc_44228_n8903;
  wire u2__abc_44228_n8905;
  wire u2__abc_44228_n8906_1;
  wire u2__abc_44228_n8907_1;
  wire u2__abc_44228_n8908;
  wire u2__abc_44228_n8909;
  wire u2__abc_44228_n8910;
  wire u2__abc_44228_n8911;
  wire u2__abc_44228_n8912_1;
  wire u2__abc_44228_n8913;
  wire u2__abc_44228_n8914;
  wire u2__abc_44228_n8915;
  wire u2__abc_44228_n8916;
  wire u2__abc_44228_n8917_1;
  wire u2__abc_44228_n8918_1;
  wire u2__abc_44228_n8919;
  wire u2__abc_44228_n8920;
  wire u2__abc_44228_n8922;
  wire u2__abc_44228_n8923_1;
  wire u2__abc_44228_n8924;
  wire u2__abc_44228_n8925;
  wire u2__abc_44228_n8926;
  wire u2__abc_44228_n8927;
  wire u2__abc_44228_n8928_1;
  wire u2__abc_44228_n8929_1;
  wire u2__abc_44228_n8930;
  wire u2__abc_44228_n8931;
  wire u2__abc_44228_n8932;
  wire u2__abc_44228_n8933;
  wire u2__abc_44228_n8934_1;
  wire u2__abc_44228_n8935;
  wire u2__abc_44228_n8936;
  wire u2__abc_44228_n8937;
  wire u2__abc_44228_n8939_1;
  wire u2__abc_44228_n8940_1;
  wire u2__abc_44228_n8941;
  wire u2__abc_44228_n8942;
  wire u2__abc_44228_n8943;
  wire u2__abc_44228_n8944;
  wire u2__abc_44228_n8945_1;
  wire u2__abc_44228_n8946;
  wire u2__abc_44228_n8947;
  wire u2__abc_44228_n8948;
  wire u2__abc_44228_n8949;
  wire u2__abc_44228_n8950_1;
  wire u2__abc_44228_n8951_1;
  wire u2__abc_44228_n8952;
  wire u2__abc_44228_n8953;
  wire u2__abc_44228_n8954;
  wire u2__abc_44228_n8955;
  wire u2__abc_44228_n8957;
  wire u2__abc_44228_n8958;
  wire u2__abc_44228_n8959;
  wire u2__abc_44228_n8960;
  wire u2__abc_44228_n8961_1;
  wire u2__abc_44228_n8962_1;
  wire u2__abc_44228_n8963;
  wire u2__abc_44228_n8964;
  wire u2__abc_44228_n8965;
  wire u2__abc_44228_n8966;
  wire u2__abc_44228_n8967_1;
  wire u2__abc_44228_n8968;
  wire u2__abc_44228_n8969;
  wire u2__abc_44228_n8970;
  wire u2__abc_44228_n8971;
  wire u2__abc_44228_n8972_1;
  wire u2__abc_44228_n8974;
  wire u2__abc_44228_n8975;
  wire u2__abc_44228_n8976;
  wire u2__abc_44228_n8977;
  wire u2__abc_44228_n8978_1;
  wire u2__abc_44228_n8979;
  wire u2__abc_44228_n8980;
  wire u2__abc_44228_n8981;
  wire u2__abc_44228_n8982;
  wire u2__abc_44228_n8983_1;
  wire u2__abc_44228_n8984_1;
  wire u2__abc_44228_n8985;
  wire u2__abc_44228_n8986;
  wire u2__abc_44228_n8987;
  wire u2__abc_44228_n8988;
  wire u2__abc_44228_n8989_1;
  wire u2__abc_44228_n8991;
  wire u2__abc_44228_n8992;
  wire u2__abc_44228_n8993;
  wire u2__abc_44228_n8994_1;
  wire u2__abc_44228_n8995_1;
  wire u2__abc_44228_n8996;
  wire u2__abc_44228_n8997;
  wire u2__abc_44228_n8998;
  wire u2__abc_44228_n8999;
  wire u2__abc_44228_n9000_1;
  wire u2__abc_44228_n9001;
  wire u2__abc_44228_n9002;
  wire u2__abc_44228_n9003;
  wire u2__abc_44228_n9004;
  wire u2__abc_44228_n9005_1;
  wire u2__abc_44228_n9006_1;
  wire u2__abc_44228_n9008;
  wire u2__abc_44228_n9009;
  wire u2__abc_44228_n9010;
  wire u2__abc_44228_n9011_1;
  wire u2__abc_44228_n9012;
  wire u2__abc_44228_n9013;
  wire u2__abc_44228_n9014;
  wire u2__abc_44228_n9015;
  wire u2__abc_44228_n9016_1;
  wire u2__abc_44228_n9017_1;
  wire u2__abc_44228_n9018;
  wire u2__abc_44228_n9019;
  wire u2__abc_44228_n9020;
  wire u2__abc_44228_n9021;
  wire u2__abc_44228_n9022_1;
  wire u2__abc_44228_n9023;
  wire u2__abc_44228_n9025;
  wire u2__abc_44228_n9026;
  wire u2__abc_44228_n9027_1;
  wire u2__abc_44228_n9028_1;
  wire u2__abc_44228_n9029;
  wire u2__abc_44228_n9030;
  wire u2__abc_44228_n9031;
  wire u2__abc_44228_n9032;
  wire u2__abc_44228_n9033_1;
  wire u2__abc_44228_n9034;
  wire u2__abc_44228_n9035;
  wire u2__abc_44228_n9036;
  wire u2__abc_44228_n9037;
  wire u2__abc_44228_n9038_1;
  wire u2__abc_44228_n9039_1;
  wire u2__abc_44228_n9040;
  wire u2__abc_44228_n9042;
  wire u2__abc_44228_n9043;
  wire u2__abc_44228_n9044_1;
  wire u2__abc_44228_n9045;
  wire u2__abc_44228_n9046;
  wire u2__abc_44228_n9047;
  wire u2__abc_44228_n9048;
  wire u2__abc_44228_n9049_1;
  wire u2__abc_44228_n9050_1;
  wire u2__abc_44228_n9051;
  wire u2__abc_44228_n9052;
  wire u2__abc_44228_n9053;
  wire u2__abc_44228_n9054;
  wire u2__abc_44228_n9055_1;
  wire u2__abc_44228_n9056;
  wire u2__abc_44228_n9057;
  wire u2__abc_44228_n9059;
  wire u2__abc_44228_n9060_1;
  wire u2__abc_44228_n9061_1;
  wire u2__abc_44228_n9062;
  wire u2__abc_44228_n9063;
  wire u2__abc_44228_n9064;
  wire u2__abc_44228_n9065;
  wire u2__abc_44228_n9066_1;
  wire u2__abc_44228_n9067;
  wire u2__abc_44228_n9068;
  wire u2__abc_44228_n9069;
  wire u2__abc_44228_n9070;
  wire u2__abc_44228_n9071_1;
  wire u2__abc_44228_n9072_1;
  wire u2__abc_44228_n9073;
  wire u2__abc_44228_n9074;
  wire u2__abc_44228_n9076;
  wire u2__abc_44228_n9077_1;
  wire u2__abc_44228_n9078;
  wire u2__abc_44228_n9079;
  wire u2__abc_44228_n9080;
  wire u2__abc_44228_n9081;
  wire u2__abc_44228_n9082_1;
  wire u2__abc_44228_n9083_1;
  wire u2__abc_44228_n9084;
  wire u2__abc_44228_n9085;
  wire u2__abc_44228_n9086;
  wire u2__abc_44228_n9087;
  wire u2__abc_44228_n9088_1;
  wire u2__abc_44228_n9089;
  wire u2__abc_44228_n9090;
  wire u2__abc_44228_n9091;
  wire u2__abc_44228_n9092;
  wire u2__abc_44228_n9094_1;
  wire u2__abc_44228_n9095;
  wire u2__abc_44228_n9096;
  wire u2__abc_44228_n9097;
  wire u2__abc_44228_n9098;
  wire u2__abc_44228_n9099_1;
  wire u2__abc_44228_n9100;
  wire u2__abc_44228_n9101;
  wire u2__abc_44228_n9102;
  wire u2__abc_44228_n9103;
  wire u2__abc_44228_n9104_1;
  wire u2__abc_44228_n9105_1;
  wire u2__abc_44228_n9106;
  wire u2__abc_44228_n9107;
  wire u2__abc_44228_n9108;
  wire u2__abc_44228_n9109;
  wire u2__abc_44228_n9111;
  wire u2__abc_44228_n9112;
  wire u2__abc_44228_n9113;
  wire u2__abc_44228_n9114;
  wire u2__abc_44228_n9115_1;
  wire u2__abc_44228_n9116_1;
  wire u2__abc_44228_n9117;
  wire u2__abc_44228_n9118;
  wire u2__abc_44228_n9119;
  wire u2__abc_44228_n9120;
  wire u2__abc_44228_n9121_1;
  wire u2__abc_44228_n9122;
  wire u2__abc_44228_n9123;
  wire u2__abc_44228_n9124;
  wire u2__abc_44228_n9125;
  wire u2__abc_44228_n9126_1;
  wire u2__abc_44228_n9128;
  wire u2__abc_44228_n9129;
  wire u2__abc_44228_n9130;
  wire u2__abc_44228_n9131;
  wire u2__abc_44228_n9132_1;
  wire u2__abc_44228_n9133;
  wire u2__abc_44228_n9134;
  wire u2__abc_44228_n9135;
  wire u2__abc_44228_n9136;
  wire u2__abc_44228_n9137_1;
  wire u2__abc_44228_n9138_1;
  wire u2__abc_44228_n9139;
  wire u2__abc_44228_n9140;
  wire u2__abc_44228_n9141;
  wire u2__abc_44228_n9142;
  wire u2__abc_44228_n9143_1;
  wire u2__abc_44228_n9145;
  wire u2__abc_44228_n9146;
  wire u2__abc_44228_n9147;
  wire u2__abc_44228_n9148_1;
  wire u2__abc_44228_n9149_1;
  wire u2__abc_44228_n9150;
  wire u2__abc_44228_n9151;
  wire u2__abc_44228_n9152;
  wire u2__abc_44228_n9153;
  wire u2__abc_44228_n9154_1;
  wire u2__abc_44228_n9155;
  wire u2__abc_44228_n9156;
  wire u2__abc_44228_n9157;
  wire u2__abc_44228_n9158;
  wire u2__abc_44228_n9159_1;
  wire u2__abc_44228_n9160_1;
  wire u2__abc_44228_n9161;
  wire u2__abc_44228_n9163;
  wire u2__abc_44228_n9164;
  wire u2__abc_44228_n9165_1;
  wire u2__abc_44228_n9166;
  wire u2__abc_44228_n9167;
  wire u2__abc_44228_n9168;
  wire u2__abc_44228_n9169;
  wire u2__abc_44228_n9170_1;
  wire u2__abc_44228_n9171_1;
  wire u2__abc_44228_n9172;
  wire u2__abc_44228_n9173;
  wire u2__abc_44228_n9174;
  wire u2__abc_44228_n9175;
  wire u2__abc_44228_n9176_1;
  wire u2__abc_44228_n9177;
  wire u2__abc_44228_n9178;
  wire u2__abc_44228_n9180;
  wire u2__abc_44228_n9181_1;
  wire u2__abc_44228_n9182_1;
  wire u2__abc_44228_n9183;
  wire u2__abc_44228_n9184;
  wire u2__abc_44228_n9185;
  wire u2__abc_44228_n9186;
  wire u2__abc_44228_n9187_1;
  wire u2__abc_44228_n9188;
  wire u2__abc_44228_n9189;
  wire u2__abc_44228_n9190;
  wire u2__abc_44228_n9191;
  wire u2__abc_44228_n9192_1;
  wire u2__abc_44228_n9193_1;
  wire u2__abc_44228_n9194;
  wire u2__abc_44228_n9195;
  wire u2__abc_44228_n9197;
  wire u2__abc_44228_n9198_1;
  wire u2__abc_44228_n9199;
  wire u2__abc_44228_n9200;
  wire u2__abc_44228_n9201;
  wire u2__abc_44228_n9202;
  wire u2__abc_44228_n9203_1;
  wire u2__abc_44228_n9204_1;
  wire u2__abc_44228_n9205;
  wire u2__abc_44228_n9206;
  wire u2__abc_44228_n9207;
  wire u2__abc_44228_n9208;
  wire u2__abc_44228_n9209_1;
  wire u2__abc_44228_n9210;
  wire u2__abc_44228_n9211;
  wire u2__abc_44228_n9212;
  wire u2__abc_44228_n9214_1;
  wire u2__abc_44228_n9215_1;
  wire u2__abc_44228_n9216;
  wire u2__abc_44228_n9217;
  wire u2__abc_44228_n9218;
  wire u2__abc_44228_n9219;
  wire u2__abc_44228_n9220_1;
  wire u2__abc_44228_n9221;
  wire u2__abc_44228_n9222;
  wire u2__abc_44228_n9223;
  wire u2__abc_44228_n9224;
  wire u2__abc_44228_n9225_1;
  wire u2__abc_44228_n9226_1;
  wire u2__abc_44228_n9227;
  wire u2__abc_44228_n9228;
  wire u2__abc_44228_n9229;
  wire u2__abc_44228_n9230;
  wire u2__abc_44228_n9232;
  wire u2__abc_44228_n9233;
  wire u2__abc_44228_n9234;
  wire u2__abc_44228_n9235;
  wire u2__abc_44228_n9236_1;
  wire u2__abc_44228_n9237_1;
  wire u2__abc_44228_n9238;
  wire u2__abc_44228_n9239;
  wire u2__abc_44228_n9240;
  wire u2__abc_44228_n9241;
  wire u2__abc_44228_n9242_1;
  wire u2__abc_44228_n9243;
  wire u2__abc_44228_n9244;
  wire u2__abc_44228_n9245;
  wire u2__abc_44228_n9246;
  wire u2__abc_44228_n9247_1;
  wire u2__abc_44228_n9249;
  wire u2__abc_44228_n9250;
  wire u2__abc_44228_n9251;
  wire u2__abc_44228_n9252;
  wire u2__abc_44228_n9253_1;
  wire u2__abc_44228_n9254;
  wire u2__abc_44228_n9255;
  wire u2__abc_44228_n9256;
  wire u2__abc_44228_n9257;
  wire u2__abc_44228_n9258_1;
  wire u2__abc_44228_n9259_1;
  wire u2__abc_44228_n9260;
  wire u2__abc_44228_n9261;
  wire u2__abc_44228_n9262;
  wire u2__abc_44228_n9263;
  wire u2__abc_44228_n9264_1;
  wire u2__abc_44228_n9266;
  wire u2__abc_44228_n9267;
  wire u2__abc_44228_n9268;
  wire u2__abc_44228_n9269_1;
  wire u2__abc_44228_n9270_1;
  wire u2__abc_44228_n9271;
  wire u2__abc_44228_n9272;
  wire u2__abc_44228_n9273;
  wire u2__abc_44228_n9274;
  wire u2__abc_44228_n9275_1;
  wire u2__abc_44228_n9276;
  wire u2__abc_44228_n9277;
  wire u2__abc_44228_n9278;
  wire u2__abc_44228_n9279;
  wire u2__abc_44228_n9280_1;
  wire u2__abc_44228_n9281_1;
  wire u2__abc_44228_n9283;
  wire u2__abc_44228_n9284;
  wire u2__abc_44228_n9285;
  wire u2__abc_44228_n9286_1;
  wire u2__abc_44228_n9287;
  wire u2__abc_44228_n9288;
  wire u2__abc_44228_n9289;
  wire u2__abc_44228_n9290;
  wire u2__abc_44228_n9291_1;
  wire u2__abc_44228_n9292_1;
  wire u2__abc_44228_n9293;
  wire u2__abc_44228_n9294;
  wire u2__abc_44228_n9295;
  wire u2__abc_44228_n9296;
  wire u2__abc_44228_n9297_1;
  wire u2__abc_44228_n9298;
  wire u2__abc_44228_n9300;
  wire u2__abc_44228_n9301;
  wire u2__abc_44228_n9302_1;
  wire u2__abc_44228_n9303_1;
  wire u2__abc_44228_n9304;
  wire u2__abc_44228_n9305;
  wire u2__abc_44228_n9306;
  wire u2__abc_44228_n9307;
  wire u2__abc_44228_n9308_1;
  wire u2__abc_44228_n9309;
  wire u2__abc_44228_n9310;
  wire u2__abc_44228_n9311;
  wire u2__abc_44228_n9312;
  wire u2__abc_44228_n9313_1;
  wire u2__abc_44228_n9314_1;
  wire u2__abc_44228_n9315;
  wire u2__abc_44228_n9317;
  wire u2__abc_44228_n9318;
  wire u2__abc_44228_n9319_1;
  wire u2__abc_44228_n9320;
  wire u2__abc_44228_n9321;
  wire u2__abc_44228_n9322;
  wire u2__abc_44228_n9323;
  wire u2__abc_44228_n9324_1;
  wire u2__abc_44228_n9325_1;
  wire u2__abc_44228_n9326;
  wire u2__abc_44228_n9327;
  wire u2__abc_44228_n9328;
  wire u2__abc_44228_n9329;
  wire u2__abc_44228_n9330_1;
  wire u2__abc_44228_n9331;
  wire u2__abc_44228_n9332;
  wire u2__abc_44228_n9334;
  wire u2__abc_44228_n9335_1;
  wire u2__abc_44228_n9336_1;
  wire u2__abc_44228_n9337;
  wire u2__abc_44228_n9338;
  wire u2__abc_44228_n9339;
  wire u2__abc_44228_n9340;
  wire u2__abc_44228_n9341_1;
  wire u2__abc_44228_n9342;
  wire u2__abc_44228_n9343;
  wire u2__abc_44228_n9344;
  wire u2__abc_44228_n9345;
  wire u2__abc_44228_n9346_1;
  wire u2__abc_44228_n9347_1;
  wire u2__abc_44228_n9348;
  wire u2__abc_44228_n9349;
  wire u2__abc_44228_n9351;
  wire u2__abc_44228_n9352_1;
  wire u2__abc_44228_n9353;
  wire u2__abc_44228_n9354;
  wire u2__abc_44228_n9355;
  wire u2__abc_44228_n9356;
  wire u2__abc_44228_n9357_1;
  wire u2__abc_44228_n9358_1;
  wire u2__abc_44228_n9359;
  wire u2__abc_44228_n9360;
  wire u2__abc_44228_n9361;
  wire u2__abc_44228_n9362;
  wire u2__abc_44228_n9363_1;
  wire u2__abc_44228_n9364;
  wire u2__abc_44228_n9365;
  wire u2__abc_44228_n9366;
  wire u2__abc_44228_n9368_1;
  wire u2__abc_44228_n9369_1;
  wire u2__abc_44228_n9370;
  wire u2__abc_44228_n9371;
  wire u2__abc_44228_n9372;
  wire u2__abc_44228_n9373;
  wire u2__abc_44228_n9374_1;
  wire u2__abc_44228_n9375;
  wire u2__abc_44228_n9376;
  wire u2__abc_44228_n9377;
  wire u2__abc_44228_n9378;
  wire u2__abc_44228_n9379_1;
  wire u2__abc_44228_n9380_1;
  wire u2__abc_44228_n9381;
  wire u2__abc_44228_n9382;
  wire u2__abc_44228_n9383;
  wire u2__abc_44228_n9385_1;
  wire u2__abc_44228_n9386;
  wire u2__abc_44228_n9387;
  wire u2__abc_44228_n9388;
  wire u2__abc_44228_n9389;
  wire u2__abc_44228_n9390_1;
  wire u2__abc_44228_n9391_1;
  wire u2__abc_44228_n9392;
  wire u2__abc_44228_n9393;
  wire u2__abc_44228_n9394;
  wire u2__abc_44228_n9395;
  wire u2__abc_44228_n9396_1;
  wire u2__abc_44228_n9397;
  wire u2__abc_44228_n9398;
  wire u2__abc_44228_n9399;
  wire u2__abc_44228_n9400;
  wire u2__abc_44228_n9401_1;
  wire u2__abc_44228_n9403;
  wire u2__abc_44228_n9404;
  wire u2__abc_44228_n9405;
  wire u2__abc_44228_n9406;
  wire u2__abc_44228_n9407_1;
  wire u2__abc_44228_n9408;
  wire u2__abc_44228_n9409;
  wire u2__abc_44228_n9410;
  wire u2__abc_44228_n9411;
  wire u2__abc_44228_n9412_1;
  wire u2__abc_44228_n9413_1;
  wire u2__abc_44228_n9414;
  wire u2__abc_44228_n9415;
  wire u2__abc_44228_n9416;
  wire u2__abc_44228_n9417;
  wire u2__abc_44228_n9418_1;
  wire u2__abc_44228_n9420;
  wire u2__abc_44228_n9421;
  wire u2__abc_44228_n9422;
  wire u2__abc_44228_n9423_1;
  wire u2__abc_44228_n9424_1;
  wire u2__abc_44228_n9425;
  wire u2__abc_44228_n9426;
  wire u2__abc_44228_n9427;
  wire u2__abc_44228_n9428;
  wire u2__abc_44228_n9429_1;
  wire u2__abc_44228_n9430;
  wire u2__abc_44228_n9431;
  wire u2__abc_44228_n9432;
  wire u2__abc_44228_n9433;
  wire u2__abc_44228_n9434_1;
  wire u2__abc_44228_n9435_1;
  wire u2__abc_44228_n9436;
  wire u2__abc_44228_n9438;
  wire u2__abc_44228_n9439;
  wire u2__abc_44228_n9440_1;
  wire u2__abc_44228_n9441;
  wire u2__abc_44228_n9442;
  wire u2__abc_44228_n9443;
  wire u2__abc_44228_n9444;
  wire u2__abc_44228_n9445_1;
  wire u2__abc_44228_n9446_1;
  wire u2__abc_44228_n9447;
  wire u2__abc_44228_n9448;
  wire u2__abc_44228_n9449;
  wire u2__abc_44228_n9450;
  wire u2__abc_44228_n9451_1;
  wire u2__abc_44228_n9452;
  wire u2__abc_44228_n9453;
  wire u2__abc_44228_n9455;
  wire u2__abc_44228_n9456_1;
  wire u2__abc_44228_n9457_1;
  wire u2__abc_44228_n9458;
  wire u2__abc_44228_n9459;
  wire u2__abc_44228_n9460;
  wire u2__abc_44228_n9461;
  wire u2__abc_44228_n9462_1;
  wire u2__abc_44228_n9463;
  wire u2__abc_44228_n9464;
  wire u2__abc_44228_n9465;
  wire u2__abc_44228_n9466;
  wire u2__abc_44228_n9467_1;
  wire u2__abc_44228_n9468_1;
  wire u2__abc_44228_n9469;
  wire u2__abc_44228_n9470;
  wire u2__abc_44228_n9472;
  wire u2__abc_44228_n9473_1;
  wire u2__abc_44228_n9474;
  wire u2__abc_44228_n9475;
  wire u2__abc_44228_n9476;
  wire u2__abc_44228_n9477;
  wire u2__abc_44228_n9478_1;
  wire u2__abc_44228_n9479_1;
  wire u2__abc_44228_n9480;
  wire u2__abc_44228_n9481;
  wire u2__abc_44228_n9482;
  wire u2__abc_44228_n9483;
  wire u2__abc_44228_n9484_1;
  wire u2__abc_44228_n9485;
  wire u2__abc_44228_n9486;
  wire u2__abc_44228_n9487;
  wire u2__abc_44228_n9489_1;
  wire u2__abc_44228_n9490_1;
  wire u2__abc_44228_n9491;
  wire u2__abc_44228_n9492;
  wire u2__abc_44228_n9493;
  wire u2__abc_44228_n9494;
  wire u2__abc_44228_n9495_1;
  wire u2__abc_44228_n9496;
  wire u2__abc_44228_n9497;
  wire u2__abc_44228_n9498;
  wire u2__abc_44228_n9499;
  wire u2__abc_44228_n9500_1;
  wire u2__abc_44228_n9501_1;
  wire u2__abc_44228_n9502;
  wire u2__abc_44228_n9503;
  wire u2__abc_44228_n9504;
  wire u2__abc_44228_n9505;
  wire u2__abc_44228_n9507;
  wire u2__abc_44228_n9508;
  wire u2__abc_44228_n9509;
  wire u2__abc_44228_n9510;
  wire u2__abc_44228_n9511_1;
  wire u2__abc_44228_n9512_1;
  wire u2__abc_44228_n9513;
  wire u2__abc_44228_n9514;
  wire u2__abc_44228_n9515;
  wire u2__abc_44228_n9516;
  wire u2__abc_44228_n9517_1;
  wire u2__abc_44228_n9518;
  wire u2__abc_44228_n9519;
  wire u2__abc_44228_n9520;
  wire u2__abc_44228_n9521;
  wire u2__abc_44228_n9522_1;
  wire u2__abc_44228_n9524;
  wire u2__abc_44228_n9525;
  wire u2__abc_44228_n9526;
  wire u2__abc_44228_n9527;
  wire u2__abc_44228_n9528_1;
  wire u2__abc_44228_n9529;
  wire u2__abc_44228_n9530;
  wire u2__abc_44228_n9531;
  wire u2__abc_44228_n9532;
  wire u2__abc_44228_n9533_1;
  wire u2__abc_44228_n9534_1;
  wire u2__abc_44228_n9535;
  wire u2__abc_44228_n9536;
  wire u2__abc_44228_n9537;
  wire u2__abc_44228_n9538;
  wire u2__abc_44228_n9539_1;
  wire u2__abc_44228_n9541;
  wire u2__abc_44228_n9542;
  wire u2__abc_44228_n9543;
  wire u2__abc_44228_n9544_1;
  wire u2__abc_44228_n9545_1;
  wire u2__abc_44228_n9546;
  wire u2__abc_44228_n9547;
  wire u2__abc_44228_n9548;
  wire u2__abc_44228_n9549;
  wire u2__abc_44228_n9550_1;
  wire u2__abc_44228_n9551;
  wire u2__abc_44228_n9552;
  wire u2__abc_44228_n9553;
  wire u2__abc_44228_n9554;
  wire u2__abc_44228_n9555_1;
  wire u2__abc_44228_n9556_1;
  wire u2__abc_44228_n9558;
  wire u2__abc_44228_n9559;
  wire u2__abc_44228_n9560;
  wire u2__abc_44228_n9561_1;
  wire u2__abc_44228_n9562;
  wire u2__abc_44228_n9563;
  wire u2__abc_44228_n9564;
  wire u2__abc_44228_n9565;
  wire u2__abc_44228_n9566_1;
  wire u2__abc_44228_n9567_1;
  wire u2__abc_44228_n9568;
  wire u2__abc_44228_n9569;
  wire u2__abc_44228_n9570;
  wire u2__abc_44228_n9571;
  wire u2__abc_44228_n9572_1;
  wire u2__abc_44228_n9573;
  wire u2__abc_44228_n9575;
  wire u2__abc_44228_n9576;
  wire u2__abc_44228_n9577_1;
  wire u2__abc_44228_n9578_1;
  wire u2__abc_44228_n9579;
  wire u2__abc_44228_n9580;
  wire u2__abc_44228_n9581;
  wire u2__abc_44228_n9582;
  wire u2__abc_44228_n9583_1;
  wire u2__abc_44228_n9584;
  wire u2__abc_44228_n9585;
  wire u2__abc_44228_n9586;
  wire u2__abc_44228_n9587;
  wire u2__abc_44228_n9588_1;
  wire u2__abc_44228_n9589_1;
  wire u2__abc_44228_n9590;
  wire u2__abc_44228_n9592;
  wire u2__abc_44228_n9593;
  wire u2__abc_44228_n9594_1;
  wire u2__abc_44228_n9595;
  wire u2__abc_44228_n9596;
  wire u2__abc_44228_n9597;
  wire u2__abc_44228_n9598;
  wire u2__abc_44228_n9599_1;
  wire u2__abc_44228_n9600_1;
  wire u2__abc_44228_n9601;
  wire u2__abc_44228_n9602;
  wire u2__abc_44228_n9603;
  wire u2__abc_44228_n9604;
  wire u2__abc_44228_n9605_1;
  wire u2__abc_44228_n9606;
  wire u2__abc_44228_n9607;
  wire u2__abc_44228_n9609;
  wire u2__abc_44228_n9610_1;
  wire u2__abc_44228_n9611_1;
  wire u2__abc_44228_n9612;
  wire u2__abc_44228_n9613;
  wire u2__abc_44228_n9614;
  wire u2__abc_44228_n9615;
  wire u2__abc_44228_n9616_1;
  wire u2__abc_44228_n9617;
  wire u2__abc_44228_n9618;
  wire u2__abc_44228_n9619;
  wire u2__abc_44228_n9620;
  wire u2__abc_44228_n9621_1;
  wire u2__abc_44228_n9622_1;
  wire u2__abc_44228_n9623;
  wire u2__abc_44228_n9624;
  wire u2__abc_44228_n9626;
  wire u2__abc_44228_n9627_1;
  wire u2__abc_44228_n9628;
  wire u2__abc_44228_n9629;
  wire u2__abc_44228_n9630;
  wire u2__abc_44228_n9631;
  wire u2__abc_44228_n9632_1;
  wire u2__abc_44228_n9633_1;
  wire u2__abc_44228_n9634;
  wire u2__abc_44228_n9635;
  wire u2__abc_44228_n9636;
  wire u2__abc_44228_n9637;
  wire u2__abc_44228_n9638_1;
  wire u2__abc_44228_n9639;
  wire u2__abc_44228_n9640;
  wire u2__abc_44228_n9641;
  wire u2__abc_44228_n9643_1;
  wire u2__abc_44228_n9644_1;
  wire u2__abc_44228_n9645;
  wire u2__abc_44228_n9646;
  wire u2__abc_44228_n9647;
  wire u2__abc_44228_n9648;
  wire u2__abc_44228_n9649_1;
  wire u2__abc_44228_n9650;
  wire u2__abc_44228_n9651;
  wire u2__abc_44228_n9652;
  wire u2__abc_44228_n9653;
  wire u2__abc_44228_n9654_1;
  wire u2__abc_44228_n9655_1;
  wire u2__abc_44228_n9656;
  wire u2__abc_44228_n9657;
  wire u2__abc_44228_n9658;
  wire u2__abc_44228_n9660_1;
  wire u2__abc_44228_n9661;
  wire u2__abc_44228_n9662;
  wire u2__abc_44228_n9663;
  wire u2__abc_44228_n9664;
  wire u2__abc_44228_n9665_1;
  wire u2__abc_44228_n9666_1;
  wire u2__abc_44228_n9667;
  wire u2__abc_44228_n9668;
  wire u2__abc_44228_n9669;
  wire u2__abc_44228_n9670;
  wire u2__abc_44228_n9671_1;
  wire u2__abc_44228_n9672;
  wire u2__abc_44228_n9673;
  wire u2__abc_44228_n9674;
  wire u2__abc_44228_n9675;
  wire u2__abc_44228_n9677_1;
  wire u2__abc_44228_n9678;
  wire u2__abc_44228_n9679;
  wire u2__abc_44228_n9680;
  wire u2__abc_44228_n9681;
  wire u2__abc_44228_n9682_1;
  wire u2__abc_44228_n9683;
  wire u2__abc_44228_n9684;
  wire u2__abc_44228_n9685;
  wire u2__abc_44228_n9686;
  wire u2__abc_44228_n9687_1;
  wire u2__abc_44228_n9688_1;
  wire u2__abc_44228_n9689;
  wire u2__abc_44228_n9690;
  wire u2__abc_44228_n9691;
  wire u2__abc_44228_n9692;
  wire u2__abc_44228_n9694;
  wire u2__abc_44228_n9695;
  wire u2__abc_44228_n9696;
  wire u2__abc_44228_n9697;
  wire u2__abc_44228_n9698_1;
  wire u2__abc_44228_n9699_1;
  wire u2__abc_44228_n9700;
  wire u2__abc_44228_n9701;
  wire u2__abc_44228_n9702;
  wire u2__abc_44228_n9703;
  wire u2__abc_44228_n9704_1;
  wire u2__abc_44228_n9705;
  wire u2__abc_44228_n9706;
  wire u2__abc_44228_n9707;
  wire u2__abc_44228_n9708;
  wire u2__abc_44228_n9709_1;
  wire u2__abc_44228_n9710_1;
  wire u2__abc_44228_n9712;
  wire u2__abc_44228_n9713;
  wire u2__abc_44228_n9714;
  wire u2__abc_44228_n9715_1;
  wire u2__abc_44228_n9716;
  wire u2__abc_44228_n9717;
  wire u2__abc_44228_n9718;
  wire u2__abc_44228_n9719;
  wire u2__abc_44228_n9720_1;
  wire u2__abc_44228_n9721_1;
  wire u2__abc_44228_n9722;
  wire u2__abc_44228_n9723;
  wire u2__abc_44228_n9724;
  wire u2__abc_44228_n9725;
  wire u2__abc_44228_n9726_1;
  wire u2__abc_44228_n9727;
  wire u2__abc_44228_n9729;
  wire u2__abc_44228_n9730;
  wire u2__abc_44228_n9731_1;
  wire u2__abc_44228_n9732_1;
  wire u2__abc_44228_n9733;
  wire u2__abc_44228_n9734;
  wire u2__abc_44228_n9735;
  wire u2__abc_44228_n9736;
  wire u2__abc_44228_n9737_1;
  wire u2__abc_44228_n9738;
  wire u2__abc_44228_n9739;
  wire u2__abc_44228_n9740;
  wire u2__abc_44228_n9741;
  wire u2__abc_44228_n9742_1;
  wire u2__abc_44228_n9744;
  wire u2__abc_44228_n9745;
  wire u2__abc_44228_n9746;
  wire u2__abc_44228_n9747;
  wire u2__abc_44228_n9748_1;
  wire u2__abc_44228_n9749;
  wire u2__abc_44228_n9750;
  wire u2__abc_44228_n9751;
  wire u2__abc_44228_n9752;
  wire u2__abc_44228_n9753_1;
  wire u2__abc_44228_n9754_1;
  wire u2__abc_44228_n9755;
  wire u2__abc_44228_n9756;
  wire u2__abc_44228_n9757;
  wire u2__abc_44228_n9758;
  wire u2__abc_44228_n9759_1;
  wire u2__abc_44228_n9761;
  wire u2__abc_44228_n9762;
  wire u2__abc_44228_n9763;
  wire u2__abc_44228_n9764_1;
  wire u2__abc_44228_n9765_1;
  wire u2__abc_44228_n9766;
  wire u2__abc_44228_n9767;
  wire u2__abc_44228_n9768;
  wire u2__abc_44228_n9769;
  wire u2__abc_44228_n9770_1;
  wire u2__abc_44228_n9771;
  wire u2__abc_44228_n9772;
  wire u2__abc_44228_n9773;
  wire u2__abc_44228_n9774;
  wire u2__abc_44228_n9775_1;
  wire u2__abc_44228_n9776_1;
  wire u2__abc_44228_n9778;
  wire u2__abc_44228_n9779;
  wire u2__abc_44228_n9780;
  wire u2__abc_44228_n9781_1;
  wire u2__abc_44228_n9782;
  wire u2__abc_44228_n9783;
  wire u2__abc_44228_n9784;
  wire u2__abc_44228_n9785;
  wire u2__abc_44228_n9786_1;
  wire u2__abc_44228_n9787_1;
  wire u2__abc_44228_n9788;
  wire u2__abc_44228_n9789;
  wire u2__abc_44228_n9790;
  wire u2__abc_44228_n9791;
  wire u2__abc_44228_n9792_1;
  wire u2__abc_44228_n9793;
  wire u2__abc_44228_n9795;
  wire u2__abc_44228_n9796;
  wire u2__abc_44228_n9797_1;
  wire u2__abc_44228_n9798_1;
  wire u2__abc_44228_n9799;
  wire u2__abc_44228_n9800;
  wire u2__abc_44228_n9801;
  wire u2__abc_44228_n9802;
  wire u2__abc_44228_n9803_1;
  wire u2__abc_44228_n9804;
  wire u2__abc_44228_n9805;
  wire u2__abc_44228_n9806;
  wire u2__abc_44228_n9807;
  wire u2__abc_44228_n9808_1;
  wire u2__abc_44228_n9809_1;
  wire u2__abc_44228_n9810;
  wire u2__abc_44228_n9812;
  wire u2__abc_44228_n9813;
  wire u2__abc_44228_n9814_1;
  wire u2__abc_44228_n9815;
  wire u2__abc_44228_n9816;
  wire u2__abc_44228_n9817;
  wire u2__abc_44228_n9818;
  wire u2__abc_44228_n9819_1;
  wire u2__abc_44228_n9820_1;
  wire u2__abc_44228_n9821;
  wire u2__abc_44228_n9822;
  wire u2__abc_44228_n9823;
  wire u2__abc_44228_n9824;
  wire u2__abc_44228_n9825_1;
  wire u2__abc_44228_n9826;
  wire u2__abc_44228_n9827;
  wire u2__abc_44228_n9829;
  wire u2__abc_44228_n9830_1;
  wire u2__abc_44228_n9831_1;
  wire u2__abc_44228_n9832;
  wire u2__abc_44228_n9833;
  wire u2__abc_44228_n9834;
  wire u2__abc_44228_n9835;
  wire u2__abc_44228_n9836_1;
  wire u2__abc_44228_n9837;
  wire u2__abc_44228_n9838;
  wire u2__abc_44228_n9839;
  wire u2__abc_44228_n9840;
  wire u2__abc_44228_n9841_1;
  wire u2__abc_44228_n9842_1;
  wire u2__abc_44228_n9843;
  wire u2__abc_44228_n9844;
  wire u2__abc_44228_n9846;
  wire u2__abc_44228_n9847_1;
  wire u2__abc_44228_n9848;
  wire u2__abc_44228_n9849;
  wire u2__abc_44228_n9850;
  wire u2__abc_44228_n9851;
  wire u2__abc_44228_n9852_1;
  wire u2__abc_44228_n9853_1;
  wire u2__abc_44228_n9854;
  wire u2__abc_44228_n9855;
  wire u2__abc_44228_n9856;
  wire u2__abc_44228_n9857;
  wire u2__abc_44228_n9858_1;
  wire u2__abc_44228_n9859;
  wire u2__abc_44228_n9860;
  wire u2__abc_44228_n9861;
  wire u2__abc_44228_n9863_1;
  wire u2__abc_44228_n9864_1;
  wire u2__abc_44228_n9865;
  wire u2__abc_44228_n9866;
  wire u2__abc_44228_n9867;
  wire u2__abc_44228_n9868;
  wire u2__abc_44228_n9869_1;
  wire u2__abc_44228_n9870;
  wire u2__abc_44228_n9871;
  wire u2__abc_44228_n9872;
  wire u2__abc_44228_n9873;
  wire u2__abc_44228_n9874_1;
  wire u2__abc_44228_n9875_1;
  wire u2__abc_44228_n9876;
  wire u2__abc_44228_n9877;
  wire u2__abc_44228_n9878;
  wire u2__abc_44228_n9880_1;
  wire u2__abc_44228_n9881;
  wire u2__abc_44228_n9882;
  wire u2__abc_44228_n9883;
  wire u2__abc_44228_n9884;
  wire u2__abc_44228_n9885_1;
  wire u2__abc_44228_n9886_1;
  wire u2__abc_44228_n9887;
  wire u2__abc_44228_n9888;
  wire u2__abc_44228_n9889;
  wire u2__abc_44228_n9890;
  wire u2__abc_44228_n9891_1;
  wire u2__abc_44228_n9892;
  wire u2__abc_44228_n9893;
  wire u2__abc_44228_n9894;
  wire u2__abc_44228_n9895;
  wire u2__abc_44228_n9897_1;
  wire u2__abc_44228_n9898;
  wire u2__abc_44228_n9899;
  wire u2__abc_44228_n9900;
  wire u2__abc_44228_n9901;
  wire u2__abc_44228_n9902_1;
  wire u2__abc_44228_n9903;
  wire u2__abc_44228_n9904;
  wire u2__abc_44228_n9905;
  wire u2__abc_44228_n9906;
  wire u2__abc_44228_n9907_1;
  wire u2__abc_44228_n9908_1;
  wire u2__abc_44228_n9909;
  wire u2__abc_44228_n9910;
  wire u2__abc_44228_n9911;
  wire u2__abc_44228_n9912;
  wire u2__abc_44228_n9914;
  wire u2__abc_44228_n9915;
  wire u2__abc_44228_n9916;
  wire u2__abc_44228_n9917;
  wire u2__abc_44228_n9918_1;
  wire u2__abc_44228_n9919_1;
  wire u2__abc_44228_n9920;
  wire u2__abc_44228_n9921;
  wire u2__abc_44228_n9922;
  wire u2__abc_44228_n9923;
  wire u2__abc_44228_n9924_1;
  wire u2__abc_44228_n9925;
  wire u2__abc_44228_n9926;
  wire u2__abc_44228_n9927;
  wire u2__abc_44228_n9928;
  wire u2__abc_44228_n9929_1;
  wire u2__abc_44228_n9931;
  wire u2__abc_44228_n9932;
  wire u2__abc_44228_n9933;
  wire u2__abc_44228_n9934;
  wire u2__abc_44228_n9935_1;
  wire u2__abc_44228_n9936;
  wire u2__abc_44228_n9937;
  wire u2__abc_44228_n9938;
  wire u2__abc_44228_n9939;
  wire u2__abc_44228_n9940_1;
  wire u2__abc_44228_n9941_1;
  wire u2__abc_44228_n9942;
  wire u2__abc_44228_n9943;
  wire u2__abc_44228_n9944;
  wire u2__abc_44228_n9945;
  wire u2__abc_44228_n9946_1;
  wire u2__abc_44228_n9948;
  wire u2__abc_44228_n9949;
  wire u2__abc_44228_n9950;
  wire u2__abc_44228_n9951_1;
  wire u2__abc_44228_n9952_1;
  wire u2__abc_44228_n9953;
  wire u2__abc_44228_n9954;
  wire u2__abc_44228_n9955;
  wire u2__abc_44228_n9956;
  wire u2__abc_44228_n9957_1;
  wire u2__abc_44228_n9958;
  wire u2__abc_44228_n9959;
  wire u2__abc_44228_n9960;
  wire u2__abc_44228_n9961;
  wire u2__abc_44228_n9962_1;
  wire u2__abc_44228_n9963_1;
  wire u2__abc_44228_n9965;
  wire u2__abc_44228_n9966;
  wire u2__abc_44228_n9967;
  wire u2__abc_44228_n9968_1;
  wire u2__abc_44228_n9969;
  wire u2__abc_44228_n9970;
  wire u2__abc_44228_n9971;
  wire u2__abc_44228_n9972;
  wire u2__abc_44228_n9973_1;
  wire u2__abc_44228_n9974_1;
  wire u2__abc_44228_n9975;
  wire u2__abc_44228_n9976;
  wire u2__abc_44228_n9977;
  wire u2__abc_44228_n9978;
  wire u2__abc_44228_n9979_1;
  wire u2__abc_44228_n9980;
  wire u2__abc_44228_n9981;
  wire u2__abc_44228_n9983;
  wire u2__abc_44228_n9984_1;
  wire u2__abc_44228_n9985_1;
  wire u2__abc_44228_n9986;
  wire u2__abc_44228_n9987;
  wire u2__abc_44228_n9988;
  wire u2__abc_44228_n9989;
  wire u2__abc_44228_n9990_1;
  wire u2__abc_44228_n9991;
  wire u2__abc_44228_n9992;
  wire u2__abc_44228_n9993;
  wire u2__abc_44228_n9994;
  wire u2__abc_44228_n9995_1;
  wire u2__abc_44228_n9996_1;
  wire u2__abc_44228_n9997;
  wire u2__abc_44228_n9998;
  wire u2_cnt_0_;
  wire u2_cnt_0__FF_INPUT;
  wire u2_cnt_1_;
  wire u2_cnt_1__FF_INPUT;
  wire u2_cnt_2_;
  wire u2_cnt_2__FF_INPUT;
  wire u2_cnt_3_;
  wire u2_cnt_3__FF_INPUT;
  wire u2_cnt_4_;
  wire u2_cnt_4__FF_INPUT;
  wire u2_cnt_5_;
  wire u2_cnt_5__FF_INPUT;
  wire u2_cnt_6_;
  wire u2_cnt_6__FF_INPUT;
  wire u2_cnt_7_;
  wire u2_cnt_7__FF_INPUT;
  wire u2_o_226_;
  wire u2_o_227_;
  wire u2_o_228_;
  wire u2_o_229_;
  wire u2_o_230_;
  wire u2_o_231_;
  wire u2_o_232_;
  wire u2_o_233_;
  wire u2_o_234_;
  wire u2_o_235_;
  wire u2_o_236_;
  wire u2_o_237_;
  wire u2_o_238_;
  wire u2_o_239_;
  wire u2_o_240_;
  wire u2_o_241_;
  wire u2_o_242_;
  wire u2_o_243_;
  wire u2_o_244_;
  wire u2_o_245_;
  wire u2_o_246_;
  wire u2_o_247_;
  wire u2_o_248_;
  wire u2_o_249_;
  wire u2_o_250_;
  wire u2_o_251_;
  wire u2_o_252_;
  wire u2_o_253_;
  wire u2_o_254_;
  wire u2_o_255_;
  wire u2_o_256_;
  wire u2_o_257_;
  wire u2_o_258_;
  wire u2_o_259_;
  wire u2_o_260_;
  wire u2_o_261_;
  wire u2_o_262_;
  wire u2_o_263_;
  wire u2_o_264_;
  wire u2_o_265_;
  wire u2_o_266_;
  wire u2_o_267_;
  wire u2_o_268_;
  wire u2_o_269_;
  wire u2_o_270_;
  wire u2_o_271_;
  wire u2_o_272_;
  wire u2_o_273_;
  wire u2_o_274_;
  wire u2_o_275_;
  wire u2_o_276_;
  wire u2_o_277_;
  wire u2_o_278_;
  wire u2_o_279_;
  wire u2_o_280_;
  wire u2_o_281_;
  wire u2_o_282_;
  wire u2_o_283_;
  wire u2_o_284_;
  wire u2_o_285_;
  wire u2_o_286_;
  wire u2_o_287_;
  wire u2_o_288_;
  wire u2_o_289_;
  wire u2_o_290_;
  wire u2_o_291_;
  wire u2_o_292_;
  wire u2_o_293_;
  wire u2_o_294_;
  wire u2_o_295_;
  wire u2_o_296_;
  wire u2_o_297_;
  wire u2_o_298_;
  wire u2_o_299_;
  wire u2_o_300_;
  wire u2_o_301_;
  wire u2_o_302_;
  wire u2_o_303_;
  wire u2_o_304_;
  wire u2_o_305_;
  wire u2_o_306_;
  wire u2_o_307_;
  wire u2_o_308_;
  wire u2_o_309_;
  wire u2_o_310_;
  wire u2_o_311_;
  wire u2_o_312_;
  wire u2_o_313_;
  wire u2_o_314_;
  wire u2_o_315_;
  wire u2_o_316_;
  wire u2_o_317_;
  wire u2_o_318_;
  wire u2_o_319_;
  wire u2_o_320_;
  wire u2_o_321_;
  wire u2_o_322_;
  wire u2_o_323_;
  wire u2_o_324_;
  wire u2_o_325_;
  wire u2_o_326_;
  wire u2_o_327_;
  wire u2_o_328_;
  wire u2_o_329_;
  wire u2_o_330_;
  wire u2_o_331_;
  wire u2_o_332_;
  wire u2_o_333_;
  wire u2_o_334_;
  wire u2_o_335_;
  wire u2_o_336_;
  wire u2_o_337_;
  wire u2_o_338_;
  wire u2_o_339_;
  wire u2_o_340_;
  wire u2_o_341_;
  wire u2_o_342_;
  wire u2_o_343_;
  wire u2_o_344_;
  wire u2_o_345_;
  wire u2_o_346_;
  wire u2_o_347_;
  wire u2_o_348_;
  wire u2_o_349_;
  wire u2_o_350_;
  wire u2_o_351_;
  wire u2_o_352_;
  wire u2_o_353_;
  wire u2_o_354_;
  wire u2_o_355_;
  wire u2_o_356_;
  wire u2_o_357_;
  wire u2_o_358_;
  wire u2_o_359_;
  wire u2_o_360_;
  wire u2_o_361_;
  wire u2_o_362_;
  wire u2_o_363_;
  wire u2_o_364_;
  wire u2_o_365_;
  wire u2_o_366_;
  wire u2_o_367_;
  wire u2_o_368_;
  wire u2_o_369_;
  wire u2_o_370_;
  wire u2_o_371_;
  wire u2_o_372_;
  wire u2_o_373_;
  wire u2_o_374_;
  wire u2_o_375_;
  wire u2_o_376_;
  wire u2_o_377_;
  wire u2_o_378_;
  wire u2_o_379_;
  wire u2_o_380_;
  wire u2_o_381_;
  wire u2_o_382_;
  wire u2_o_383_;
  wire u2_o_384_;
  wire u2_o_385_;
  wire u2_o_386_;
  wire u2_o_387_;
  wire u2_o_388_;
  wire u2_o_389_;
  wire u2_o_390_;
  wire u2_o_391_;
  wire u2_o_392_;
  wire u2_o_393_;
  wire u2_o_394_;
  wire u2_o_395_;
  wire u2_o_396_;
  wire u2_o_397_;
  wire u2_o_398_;
  wire u2_o_399_;
  wire u2_o_400_;
  wire u2_o_401_;
  wire u2_o_402_;
  wire u2_o_403_;
  wire u2_o_404_;
  wire u2_o_405_;
  wire u2_o_406_;
  wire u2_o_407_;
  wire u2_o_408_;
  wire u2_o_409_;
  wire u2_o_410_;
  wire u2_o_411_;
  wire u2_o_412_;
  wire u2_o_413_;
  wire u2_o_414_;
  wire u2_o_415_;
  wire u2_o_416_;
  wire u2_o_417_;
  wire u2_o_418_;
  wire u2_o_419_;
  wire u2_o_420_;
  wire u2_o_421_;
  wire u2_o_422_;
  wire u2_o_423_;
  wire u2_o_424_;
  wire u2_o_425_;
  wire u2_o_426_;
  wire u2_o_427_;
  wire u2_o_428_;
  wire u2_o_429_;
  wire u2_o_430_;
  wire u2_o_431_;
  wire u2_o_432_;
  wire u2_o_433_;
  wire u2_o_434_;
  wire u2_o_435_;
  wire u2_o_436_;
  wire u2_o_437_;
  wire u2_o_438_;
  wire u2_o_439_;
  wire u2_o_440_;
  wire u2_o_441_;
  wire u2_o_442_;
  wire u2_o_443_;
  wire u2_o_444_;
  wire u2_o_445_;
  wire u2_o_446_;
  wire u2_o_447_;
  wire u2_o_448_;
  wire u2_o_449_;
  wire u2_remHiShift_0_;
  wire u2_remHiShift_1_;
  wire u2_remHi_0_;
  wire u2_remHi_0__FF_INPUT;
  wire u2_remHi_100_;
  wire u2_remHi_100__FF_INPUT;
  wire u2_remHi_101_;
  wire u2_remHi_101__FF_INPUT;
  wire u2_remHi_102_;
  wire u2_remHi_102__FF_INPUT;
  wire u2_remHi_103_;
  wire u2_remHi_103__FF_INPUT;
  wire u2_remHi_104_;
  wire u2_remHi_104__FF_INPUT;
  wire u2_remHi_105_;
  wire u2_remHi_105__FF_INPUT;
  wire u2_remHi_106_;
  wire u2_remHi_106__FF_INPUT;
  wire u2_remHi_107_;
  wire u2_remHi_107__FF_INPUT;
  wire u2_remHi_108_;
  wire u2_remHi_108__FF_INPUT;
  wire u2_remHi_109_;
  wire u2_remHi_109__FF_INPUT;
  wire u2_remHi_10_;
  wire u2_remHi_10__FF_INPUT;
  wire u2_remHi_110_;
  wire u2_remHi_110__FF_INPUT;
  wire u2_remHi_111_;
  wire u2_remHi_111__FF_INPUT;
  wire u2_remHi_112_;
  wire u2_remHi_112__FF_INPUT;
  wire u2_remHi_113_;
  wire u2_remHi_113__FF_INPUT;
  wire u2_remHi_114_;
  wire u2_remHi_114__FF_INPUT;
  wire u2_remHi_115_;
  wire u2_remHi_115__FF_INPUT;
  wire u2_remHi_116_;
  wire u2_remHi_116__FF_INPUT;
  wire u2_remHi_117_;
  wire u2_remHi_117__FF_INPUT;
  wire u2_remHi_118_;
  wire u2_remHi_118__FF_INPUT;
  wire u2_remHi_119_;
  wire u2_remHi_119__FF_INPUT;
  wire u2_remHi_11_;
  wire u2_remHi_11__FF_INPUT;
  wire u2_remHi_120_;
  wire u2_remHi_120__FF_INPUT;
  wire u2_remHi_121_;
  wire u2_remHi_121__FF_INPUT;
  wire u2_remHi_122_;
  wire u2_remHi_122__FF_INPUT;
  wire u2_remHi_123_;
  wire u2_remHi_123__FF_INPUT;
  wire u2_remHi_124_;
  wire u2_remHi_124__FF_INPUT;
  wire u2_remHi_125_;
  wire u2_remHi_125__FF_INPUT;
  wire u2_remHi_126_;
  wire u2_remHi_126__FF_INPUT;
  wire u2_remHi_127_;
  wire u2_remHi_127__FF_INPUT;
  wire u2_remHi_128_;
  wire u2_remHi_128__FF_INPUT;
  wire u2_remHi_129_;
  wire u2_remHi_129__FF_INPUT;
  wire u2_remHi_12_;
  wire u2_remHi_12__FF_INPUT;
  wire u2_remHi_130_;
  wire u2_remHi_130__FF_INPUT;
  wire u2_remHi_131_;
  wire u2_remHi_131__FF_INPUT;
  wire u2_remHi_132_;
  wire u2_remHi_132__FF_INPUT;
  wire u2_remHi_133_;
  wire u2_remHi_133__FF_INPUT;
  wire u2_remHi_134_;
  wire u2_remHi_134__FF_INPUT;
  wire u2_remHi_135_;
  wire u2_remHi_135__FF_INPUT;
  wire u2_remHi_136_;
  wire u2_remHi_136__FF_INPUT;
  wire u2_remHi_137_;
  wire u2_remHi_137__FF_INPUT;
  wire u2_remHi_138_;
  wire u2_remHi_138__FF_INPUT;
  wire u2_remHi_139_;
  wire u2_remHi_139__FF_INPUT;
  wire u2_remHi_13_;
  wire u2_remHi_13__FF_INPUT;
  wire u2_remHi_140_;
  wire u2_remHi_140__FF_INPUT;
  wire u2_remHi_141_;
  wire u2_remHi_141__FF_INPUT;
  wire u2_remHi_142_;
  wire u2_remHi_142__FF_INPUT;
  wire u2_remHi_143_;
  wire u2_remHi_143__FF_INPUT;
  wire u2_remHi_144_;
  wire u2_remHi_144__FF_INPUT;
  wire u2_remHi_145_;
  wire u2_remHi_145__FF_INPUT;
  wire u2_remHi_146_;
  wire u2_remHi_146__FF_INPUT;
  wire u2_remHi_147_;
  wire u2_remHi_147__FF_INPUT;
  wire u2_remHi_148_;
  wire u2_remHi_148__FF_INPUT;
  wire u2_remHi_149_;
  wire u2_remHi_149__FF_INPUT;
  wire u2_remHi_14_;
  wire u2_remHi_14__FF_INPUT;
  wire u2_remHi_150_;
  wire u2_remHi_150__FF_INPUT;
  wire u2_remHi_151_;
  wire u2_remHi_151__FF_INPUT;
  wire u2_remHi_152_;
  wire u2_remHi_152__FF_INPUT;
  wire u2_remHi_153_;
  wire u2_remHi_153__FF_INPUT;
  wire u2_remHi_154_;
  wire u2_remHi_154__FF_INPUT;
  wire u2_remHi_155_;
  wire u2_remHi_155__FF_INPUT;
  wire u2_remHi_156_;
  wire u2_remHi_156__FF_INPUT;
  wire u2_remHi_157_;
  wire u2_remHi_157__FF_INPUT;
  wire u2_remHi_158_;
  wire u2_remHi_158__FF_INPUT;
  wire u2_remHi_159_;
  wire u2_remHi_159__FF_INPUT;
  wire u2_remHi_15_;
  wire u2_remHi_15__FF_INPUT;
  wire u2_remHi_160_;
  wire u2_remHi_160__FF_INPUT;
  wire u2_remHi_161_;
  wire u2_remHi_161__FF_INPUT;
  wire u2_remHi_162_;
  wire u2_remHi_162__FF_INPUT;
  wire u2_remHi_163_;
  wire u2_remHi_163__FF_INPUT;
  wire u2_remHi_164_;
  wire u2_remHi_164__FF_INPUT;
  wire u2_remHi_165_;
  wire u2_remHi_165__FF_INPUT;
  wire u2_remHi_166_;
  wire u2_remHi_166__FF_INPUT;
  wire u2_remHi_167_;
  wire u2_remHi_167__FF_INPUT;
  wire u2_remHi_168_;
  wire u2_remHi_168__FF_INPUT;
  wire u2_remHi_169_;
  wire u2_remHi_169__FF_INPUT;
  wire u2_remHi_16_;
  wire u2_remHi_16__FF_INPUT;
  wire u2_remHi_170_;
  wire u2_remHi_170__FF_INPUT;
  wire u2_remHi_171_;
  wire u2_remHi_171__FF_INPUT;
  wire u2_remHi_172_;
  wire u2_remHi_172__FF_INPUT;
  wire u2_remHi_173_;
  wire u2_remHi_173__FF_INPUT;
  wire u2_remHi_174_;
  wire u2_remHi_174__FF_INPUT;
  wire u2_remHi_175_;
  wire u2_remHi_175__FF_INPUT;
  wire u2_remHi_176_;
  wire u2_remHi_176__FF_INPUT;
  wire u2_remHi_177_;
  wire u2_remHi_177__FF_INPUT;
  wire u2_remHi_178_;
  wire u2_remHi_178__FF_INPUT;
  wire u2_remHi_179_;
  wire u2_remHi_179__FF_INPUT;
  wire u2_remHi_17_;
  wire u2_remHi_17__FF_INPUT;
  wire u2_remHi_180_;
  wire u2_remHi_180__FF_INPUT;
  wire u2_remHi_181_;
  wire u2_remHi_181__FF_INPUT;
  wire u2_remHi_182_;
  wire u2_remHi_182__FF_INPUT;
  wire u2_remHi_183_;
  wire u2_remHi_183__FF_INPUT;
  wire u2_remHi_184_;
  wire u2_remHi_184__FF_INPUT;
  wire u2_remHi_185_;
  wire u2_remHi_185__FF_INPUT;
  wire u2_remHi_186_;
  wire u2_remHi_186__FF_INPUT;
  wire u2_remHi_187_;
  wire u2_remHi_187__FF_INPUT;
  wire u2_remHi_188_;
  wire u2_remHi_188__FF_INPUT;
  wire u2_remHi_189_;
  wire u2_remHi_189__FF_INPUT;
  wire u2_remHi_18_;
  wire u2_remHi_18__FF_INPUT;
  wire u2_remHi_190_;
  wire u2_remHi_190__FF_INPUT;
  wire u2_remHi_191_;
  wire u2_remHi_191__FF_INPUT;
  wire u2_remHi_192_;
  wire u2_remHi_192__FF_INPUT;
  wire u2_remHi_193_;
  wire u2_remHi_193__FF_INPUT;
  wire u2_remHi_194_;
  wire u2_remHi_194__FF_INPUT;
  wire u2_remHi_195_;
  wire u2_remHi_195__FF_INPUT;
  wire u2_remHi_196_;
  wire u2_remHi_196__FF_INPUT;
  wire u2_remHi_197_;
  wire u2_remHi_197__FF_INPUT;
  wire u2_remHi_198_;
  wire u2_remHi_198__FF_INPUT;
  wire u2_remHi_199_;
  wire u2_remHi_199__FF_INPUT;
  wire u2_remHi_19_;
  wire u2_remHi_19__FF_INPUT;
  wire u2_remHi_1_;
  wire u2_remHi_1__FF_INPUT;
  wire u2_remHi_200_;
  wire u2_remHi_200__FF_INPUT;
  wire u2_remHi_201_;
  wire u2_remHi_201__FF_INPUT;
  wire u2_remHi_202_;
  wire u2_remHi_202__FF_INPUT;
  wire u2_remHi_203_;
  wire u2_remHi_203__FF_INPUT;
  wire u2_remHi_204_;
  wire u2_remHi_204__FF_INPUT;
  wire u2_remHi_205_;
  wire u2_remHi_205__FF_INPUT;
  wire u2_remHi_206_;
  wire u2_remHi_206__FF_INPUT;
  wire u2_remHi_207_;
  wire u2_remHi_207__FF_INPUT;
  wire u2_remHi_208_;
  wire u2_remHi_208__FF_INPUT;
  wire u2_remHi_209_;
  wire u2_remHi_209__FF_INPUT;
  wire u2_remHi_20_;
  wire u2_remHi_20__FF_INPUT;
  wire u2_remHi_210_;
  wire u2_remHi_210__FF_INPUT;
  wire u2_remHi_211_;
  wire u2_remHi_211__FF_INPUT;
  wire u2_remHi_212_;
  wire u2_remHi_212__FF_INPUT;
  wire u2_remHi_213_;
  wire u2_remHi_213__FF_INPUT;
  wire u2_remHi_214_;
  wire u2_remHi_214__FF_INPUT;
  wire u2_remHi_215_;
  wire u2_remHi_215__FF_INPUT;
  wire u2_remHi_216_;
  wire u2_remHi_216__FF_INPUT;
  wire u2_remHi_217_;
  wire u2_remHi_217__FF_INPUT;
  wire u2_remHi_218_;
  wire u2_remHi_218__FF_INPUT;
  wire u2_remHi_219_;
  wire u2_remHi_219__FF_INPUT;
  wire u2_remHi_21_;
  wire u2_remHi_21__FF_INPUT;
  wire u2_remHi_220_;
  wire u2_remHi_220__FF_INPUT;
  wire u2_remHi_221_;
  wire u2_remHi_221__FF_INPUT;
  wire u2_remHi_222_;
  wire u2_remHi_222__FF_INPUT;
  wire u2_remHi_223_;
  wire u2_remHi_223__FF_INPUT;
  wire u2_remHi_224_;
  wire u2_remHi_224__FF_INPUT;
  wire u2_remHi_225_;
  wire u2_remHi_225__FF_INPUT;
  wire u2_remHi_226_;
  wire u2_remHi_226__FF_INPUT;
  wire u2_remHi_227_;
  wire u2_remHi_227__FF_INPUT;
  wire u2_remHi_228_;
  wire u2_remHi_228__FF_INPUT;
  wire u2_remHi_229_;
  wire u2_remHi_229__FF_INPUT;
  wire u2_remHi_22_;
  wire u2_remHi_22__FF_INPUT;
  wire u2_remHi_230_;
  wire u2_remHi_230__FF_INPUT;
  wire u2_remHi_231_;
  wire u2_remHi_231__FF_INPUT;
  wire u2_remHi_232_;
  wire u2_remHi_232__FF_INPUT;
  wire u2_remHi_233_;
  wire u2_remHi_233__FF_INPUT;
  wire u2_remHi_234_;
  wire u2_remHi_234__FF_INPUT;
  wire u2_remHi_235_;
  wire u2_remHi_235__FF_INPUT;
  wire u2_remHi_236_;
  wire u2_remHi_236__FF_INPUT;
  wire u2_remHi_237_;
  wire u2_remHi_237__FF_INPUT;
  wire u2_remHi_238_;
  wire u2_remHi_238__FF_INPUT;
  wire u2_remHi_239_;
  wire u2_remHi_239__FF_INPUT;
  wire u2_remHi_23_;
  wire u2_remHi_23__FF_INPUT;
  wire u2_remHi_240_;
  wire u2_remHi_240__FF_INPUT;
  wire u2_remHi_241_;
  wire u2_remHi_241__FF_INPUT;
  wire u2_remHi_242_;
  wire u2_remHi_242__FF_INPUT;
  wire u2_remHi_243_;
  wire u2_remHi_243__FF_INPUT;
  wire u2_remHi_244_;
  wire u2_remHi_244__FF_INPUT;
  wire u2_remHi_245_;
  wire u2_remHi_245__FF_INPUT;
  wire u2_remHi_246_;
  wire u2_remHi_246__FF_INPUT;
  wire u2_remHi_247_;
  wire u2_remHi_247__FF_INPUT;
  wire u2_remHi_248_;
  wire u2_remHi_248__FF_INPUT;
  wire u2_remHi_249_;
  wire u2_remHi_249__FF_INPUT;
  wire u2_remHi_24_;
  wire u2_remHi_24__FF_INPUT;
  wire u2_remHi_250_;
  wire u2_remHi_250__FF_INPUT;
  wire u2_remHi_251_;
  wire u2_remHi_251__FF_INPUT;
  wire u2_remHi_252_;
  wire u2_remHi_252__FF_INPUT;
  wire u2_remHi_253_;
  wire u2_remHi_253__FF_INPUT;
  wire u2_remHi_254_;
  wire u2_remHi_254__FF_INPUT;
  wire u2_remHi_255_;
  wire u2_remHi_255__FF_INPUT;
  wire u2_remHi_256_;
  wire u2_remHi_256__FF_INPUT;
  wire u2_remHi_257_;
  wire u2_remHi_257__FF_INPUT;
  wire u2_remHi_258_;
  wire u2_remHi_258__FF_INPUT;
  wire u2_remHi_259_;
  wire u2_remHi_259__FF_INPUT;
  wire u2_remHi_25_;
  wire u2_remHi_25__FF_INPUT;
  wire u2_remHi_260_;
  wire u2_remHi_260__FF_INPUT;
  wire u2_remHi_261_;
  wire u2_remHi_261__FF_INPUT;
  wire u2_remHi_262_;
  wire u2_remHi_262__FF_INPUT;
  wire u2_remHi_263_;
  wire u2_remHi_263__FF_INPUT;
  wire u2_remHi_264_;
  wire u2_remHi_264__FF_INPUT;
  wire u2_remHi_265_;
  wire u2_remHi_265__FF_INPUT;
  wire u2_remHi_266_;
  wire u2_remHi_266__FF_INPUT;
  wire u2_remHi_267_;
  wire u2_remHi_267__FF_INPUT;
  wire u2_remHi_268_;
  wire u2_remHi_268__FF_INPUT;
  wire u2_remHi_269_;
  wire u2_remHi_269__FF_INPUT;
  wire u2_remHi_26_;
  wire u2_remHi_26__FF_INPUT;
  wire u2_remHi_270_;
  wire u2_remHi_270__FF_INPUT;
  wire u2_remHi_271_;
  wire u2_remHi_271__FF_INPUT;
  wire u2_remHi_272_;
  wire u2_remHi_272__FF_INPUT;
  wire u2_remHi_273_;
  wire u2_remHi_273__FF_INPUT;
  wire u2_remHi_274_;
  wire u2_remHi_274__FF_INPUT;
  wire u2_remHi_275_;
  wire u2_remHi_275__FF_INPUT;
  wire u2_remHi_276_;
  wire u2_remHi_276__FF_INPUT;
  wire u2_remHi_277_;
  wire u2_remHi_277__FF_INPUT;
  wire u2_remHi_278_;
  wire u2_remHi_278__FF_INPUT;
  wire u2_remHi_279_;
  wire u2_remHi_279__FF_INPUT;
  wire u2_remHi_27_;
  wire u2_remHi_27__FF_INPUT;
  wire u2_remHi_280_;
  wire u2_remHi_280__FF_INPUT;
  wire u2_remHi_281_;
  wire u2_remHi_281__FF_INPUT;
  wire u2_remHi_282_;
  wire u2_remHi_282__FF_INPUT;
  wire u2_remHi_283_;
  wire u2_remHi_283__FF_INPUT;
  wire u2_remHi_284_;
  wire u2_remHi_284__FF_INPUT;
  wire u2_remHi_285_;
  wire u2_remHi_285__FF_INPUT;
  wire u2_remHi_286_;
  wire u2_remHi_286__FF_INPUT;
  wire u2_remHi_287_;
  wire u2_remHi_287__FF_INPUT;
  wire u2_remHi_288_;
  wire u2_remHi_288__FF_INPUT;
  wire u2_remHi_289_;
  wire u2_remHi_289__FF_INPUT;
  wire u2_remHi_28_;
  wire u2_remHi_28__FF_INPUT;
  wire u2_remHi_290_;
  wire u2_remHi_290__FF_INPUT;
  wire u2_remHi_291_;
  wire u2_remHi_291__FF_INPUT;
  wire u2_remHi_292_;
  wire u2_remHi_292__FF_INPUT;
  wire u2_remHi_293_;
  wire u2_remHi_293__FF_INPUT;
  wire u2_remHi_294_;
  wire u2_remHi_294__FF_INPUT;
  wire u2_remHi_295_;
  wire u2_remHi_295__FF_INPUT;
  wire u2_remHi_296_;
  wire u2_remHi_296__FF_INPUT;
  wire u2_remHi_297_;
  wire u2_remHi_297__FF_INPUT;
  wire u2_remHi_298_;
  wire u2_remHi_298__FF_INPUT;
  wire u2_remHi_299_;
  wire u2_remHi_299__FF_INPUT;
  wire u2_remHi_29_;
  wire u2_remHi_29__FF_INPUT;
  wire u2_remHi_2_;
  wire u2_remHi_2__FF_INPUT;
  wire u2_remHi_300_;
  wire u2_remHi_300__FF_INPUT;
  wire u2_remHi_301_;
  wire u2_remHi_301__FF_INPUT;
  wire u2_remHi_302_;
  wire u2_remHi_302__FF_INPUT;
  wire u2_remHi_303_;
  wire u2_remHi_303__FF_INPUT;
  wire u2_remHi_304_;
  wire u2_remHi_304__FF_INPUT;
  wire u2_remHi_305_;
  wire u2_remHi_305__FF_INPUT;
  wire u2_remHi_306_;
  wire u2_remHi_306__FF_INPUT;
  wire u2_remHi_307_;
  wire u2_remHi_307__FF_INPUT;
  wire u2_remHi_308_;
  wire u2_remHi_308__FF_INPUT;
  wire u2_remHi_309_;
  wire u2_remHi_309__FF_INPUT;
  wire u2_remHi_30_;
  wire u2_remHi_30__FF_INPUT;
  wire u2_remHi_310_;
  wire u2_remHi_310__FF_INPUT;
  wire u2_remHi_311_;
  wire u2_remHi_311__FF_INPUT;
  wire u2_remHi_312_;
  wire u2_remHi_312__FF_INPUT;
  wire u2_remHi_313_;
  wire u2_remHi_313__FF_INPUT;
  wire u2_remHi_314_;
  wire u2_remHi_314__FF_INPUT;
  wire u2_remHi_315_;
  wire u2_remHi_315__FF_INPUT;
  wire u2_remHi_316_;
  wire u2_remHi_316__FF_INPUT;
  wire u2_remHi_317_;
  wire u2_remHi_317__FF_INPUT;
  wire u2_remHi_318_;
  wire u2_remHi_318__FF_INPUT;
  wire u2_remHi_319_;
  wire u2_remHi_319__FF_INPUT;
  wire u2_remHi_31_;
  wire u2_remHi_31__FF_INPUT;
  wire u2_remHi_320_;
  wire u2_remHi_320__FF_INPUT;
  wire u2_remHi_321_;
  wire u2_remHi_321__FF_INPUT;
  wire u2_remHi_322_;
  wire u2_remHi_322__FF_INPUT;
  wire u2_remHi_323_;
  wire u2_remHi_323__FF_INPUT;
  wire u2_remHi_324_;
  wire u2_remHi_324__FF_INPUT;
  wire u2_remHi_325_;
  wire u2_remHi_325__FF_INPUT;
  wire u2_remHi_326_;
  wire u2_remHi_326__FF_INPUT;
  wire u2_remHi_327_;
  wire u2_remHi_327__FF_INPUT;
  wire u2_remHi_328_;
  wire u2_remHi_328__FF_INPUT;
  wire u2_remHi_329_;
  wire u2_remHi_329__FF_INPUT;
  wire u2_remHi_32_;
  wire u2_remHi_32__FF_INPUT;
  wire u2_remHi_330_;
  wire u2_remHi_330__FF_INPUT;
  wire u2_remHi_331_;
  wire u2_remHi_331__FF_INPUT;
  wire u2_remHi_332_;
  wire u2_remHi_332__FF_INPUT;
  wire u2_remHi_333_;
  wire u2_remHi_333__FF_INPUT;
  wire u2_remHi_334_;
  wire u2_remHi_334__FF_INPUT;
  wire u2_remHi_335_;
  wire u2_remHi_335__FF_INPUT;
  wire u2_remHi_336_;
  wire u2_remHi_336__FF_INPUT;
  wire u2_remHi_337_;
  wire u2_remHi_337__FF_INPUT;
  wire u2_remHi_338_;
  wire u2_remHi_338__FF_INPUT;
  wire u2_remHi_339_;
  wire u2_remHi_339__FF_INPUT;
  wire u2_remHi_33_;
  wire u2_remHi_33__FF_INPUT;
  wire u2_remHi_340_;
  wire u2_remHi_340__FF_INPUT;
  wire u2_remHi_341_;
  wire u2_remHi_341__FF_INPUT;
  wire u2_remHi_342_;
  wire u2_remHi_342__FF_INPUT;
  wire u2_remHi_343_;
  wire u2_remHi_343__FF_INPUT;
  wire u2_remHi_344_;
  wire u2_remHi_344__FF_INPUT;
  wire u2_remHi_345_;
  wire u2_remHi_345__FF_INPUT;
  wire u2_remHi_346_;
  wire u2_remHi_346__FF_INPUT;
  wire u2_remHi_347_;
  wire u2_remHi_347__FF_INPUT;
  wire u2_remHi_348_;
  wire u2_remHi_348__FF_INPUT;
  wire u2_remHi_349_;
  wire u2_remHi_349__FF_INPUT;
  wire u2_remHi_34_;
  wire u2_remHi_34__FF_INPUT;
  wire u2_remHi_350_;
  wire u2_remHi_350__FF_INPUT;
  wire u2_remHi_351_;
  wire u2_remHi_351__FF_INPUT;
  wire u2_remHi_352_;
  wire u2_remHi_352__FF_INPUT;
  wire u2_remHi_353_;
  wire u2_remHi_353__FF_INPUT;
  wire u2_remHi_354_;
  wire u2_remHi_354__FF_INPUT;
  wire u2_remHi_355_;
  wire u2_remHi_355__FF_INPUT;
  wire u2_remHi_356_;
  wire u2_remHi_356__FF_INPUT;
  wire u2_remHi_357_;
  wire u2_remHi_357__FF_INPUT;
  wire u2_remHi_358_;
  wire u2_remHi_358__FF_INPUT;
  wire u2_remHi_359_;
  wire u2_remHi_359__FF_INPUT;
  wire u2_remHi_35_;
  wire u2_remHi_35__FF_INPUT;
  wire u2_remHi_360_;
  wire u2_remHi_360__FF_INPUT;
  wire u2_remHi_361_;
  wire u2_remHi_361__FF_INPUT;
  wire u2_remHi_362_;
  wire u2_remHi_362__FF_INPUT;
  wire u2_remHi_363_;
  wire u2_remHi_363__FF_INPUT;
  wire u2_remHi_364_;
  wire u2_remHi_364__FF_INPUT;
  wire u2_remHi_365_;
  wire u2_remHi_365__FF_INPUT;
  wire u2_remHi_366_;
  wire u2_remHi_366__FF_INPUT;
  wire u2_remHi_367_;
  wire u2_remHi_367__FF_INPUT;
  wire u2_remHi_368_;
  wire u2_remHi_368__FF_INPUT;
  wire u2_remHi_369_;
  wire u2_remHi_369__FF_INPUT;
  wire u2_remHi_36_;
  wire u2_remHi_36__FF_INPUT;
  wire u2_remHi_370_;
  wire u2_remHi_370__FF_INPUT;
  wire u2_remHi_371_;
  wire u2_remHi_371__FF_INPUT;
  wire u2_remHi_372_;
  wire u2_remHi_372__FF_INPUT;
  wire u2_remHi_373_;
  wire u2_remHi_373__FF_INPUT;
  wire u2_remHi_374_;
  wire u2_remHi_374__FF_INPUT;
  wire u2_remHi_375_;
  wire u2_remHi_375__FF_INPUT;
  wire u2_remHi_376_;
  wire u2_remHi_376__FF_INPUT;
  wire u2_remHi_377_;
  wire u2_remHi_377__FF_INPUT;
  wire u2_remHi_378_;
  wire u2_remHi_378__FF_INPUT;
  wire u2_remHi_379_;
  wire u2_remHi_379__FF_INPUT;
  wire u2_remHi_37_;
  wire u2_remHi_37__FF_INPUT;
  wire u2_remHi_380_;
  wire u2_remHi_380__FF_INPUT;
  wire u2_remHi_381_;
  wire u2_remHi_381__FF_INPUT;
  wire u2_remHi_382_;
  wire u2_remHi_382__FF_INPUT;
  wire u2_remHi_383_;
  wire u2_remHi_383__FF_INPUT;
  wire u2_remHi_384_;
  wire u2_remHi_384__FF_INPUT;
  wire u2_remHi_385_;
  wire u2_remHi_385__FF_INPUT;
  wire u2_remHi_386_;
  wire u2_remHi_386__FF_INPUT;
  wire u2_remHi_387_;
  wire u2_remHi_387__FF_INPUT;
  wire u2_remHi_388_;
  wire u2_remHi_388__FF_INPUT;
  wire u2_remHi_389_;
  wire u2_remHi_389__FF_INPUT;
  wire u2_remHi_38_;
  wire u2_remHi_38__FF_INPUT;
  wire u2_remHi_390_;
  wire u2_remHi_390__FF_INPUT;
  wire u2_remHi_391_;
  wire u2_remHi_391__FF_INPUT;
  wire u2_remHi_392_;
  wire u2_remHi_392__FF_INPUT;
  wire u2_remHi_393_;
  wire u2_remHi_393__FF_INPUT;
  wire u2_remHi_394_;
  wire u2_remHi_394__FF_INPUT;
  wire u2_remHi_395_;
  wire u2_remHi_395__FF_INPUT;
  wire u2_remHi_396_;
  wire u2_remHi_396__FF_INPUT;
  wire u2_remHi_397_;
  wire u2_remHi_397__FF_INPUT;
  wire u2_remHi_398_;
  wire u2_remHi_398__FF_INPUT;
  wire u2_remHi_399_;
  wire u2_remHi_399__FF_INPUT;
  wire u2_remHi_39_;
  wire u2_remHi_39__FF_INPUT;
  wire u2_remHi_3_;
  wire u2_remHi_3__FF_INPUT;
  wire u2_remHi_400_;
  wire u2_remHi_400__FF_INPUT;
  wire u2_remHi_401_;
  wire u2_remHi_401__FF_INPUT;
  wire u2_remHi_402_;
  wire u2_remHi_402__FF_INPUT;
  wire u2_remHi_403_;
  wire u2_remHi_403__FF_INPUT;
  wire u2_remHi_404_;
  wire u2_remHi_404__FF_INPUT;
  wire u2_remHi_405_;
  wire u2_remHi_405__FF_INPUT;
  wire u2_remHi_406_;
  wire u2_remHi_406__FF_INPUT;
  wire u2_remHi_407_;
  wire u2_remHi_407__FF_INPUT;
  wire u2_remHi_408_;
  wire u2_remHi_408__FF_INPUT;
  wire u2_remHi_409_;
  wire u2_remHi_409__FF_INPUT;
  wire u2_remHi_40_;
  wire u2_remHi_40__FF_INPUT;
  wire u2_remHi_410_;
  wire u2_remHi_410__FF_INPUT;
  wire u2_remHi_411_;
  wire u2_remHi_411__FF_INPUT;
  wire u2_remHi_412_;
  wire u2_remHi_412__FF_INPUT;
  wire u2_remHi_413_;
  wire u2_remHi_413__FF_INPUT;
  wire u2_remHi_414_;
  wire u2_remHi_414__FF_INPUT;
  wire u2_remHi_415_;
  wire u2_remHi_415__FF_INPUT;
  wire u2_remHi_416_;
  wire u2_remHi_416__FF_INPUT;
  wire u2_remHi_417_;
  wire u2_remHi_417__FF_INPUT;
  wire u2_remHi_418_;
  wire u2_remHi_418__FF_INPUT;
  wire u2_remHi_419_;
  wire u2_remHi_419__FF_INPUT;
  wire u2_remHi_41_;
  wire u2_remHi_41__FF_INPUT;
  wire u2_remHi_420_;
  wire u2_remHi_420__FF_INPUT;
  wire u2_remHi_421_;
  wire u2_remHi_421__FF_INPUT;
  wire u2_remHi_422_;
  wire u2_remHi_422__FF_INPUT;
  wire u2_remHi_423_;
  wire u2_remHi_423__FF_INPUT;
  wire u2_remHi_424_;
  wire u2_remHi_424__FF_INPUT;
  wire u2_remHi_425_;
  wire u2_remHi_425__FF_INPUT;
  wire u2_remHi_426_;
  wire u2_remHi_426__FF_INPUT;
  wire u2_remHi_427_;
  wire u2_remHi_427__FF_INPUT;
  wire u2_remHi_428_;
  wire u2_remHi_428__FF_INPUT;
  wire u2_remHi_429_;
  wire u2_remHi_429__FF_INPUT;
  wire u2_remHi_42_;
  wire u2_remHi_42__FF_INPUT;
  wire u2_remHi_430_;
  wire u2_remHi_430__FF_INPUT;
  wire u2_remHi_431_;
  wire u2_remHi_431__FF_INPUT;
  wire u2_remHi_432_;
  wire u2_remHi_432__FF_INPUT;
  wire u2_remHi_433_;
  wire u2_remHi_433__FF_INPUT;
  wire u2_remHi_434_;
  wire u2_remHi_434__FF_INPUT;
  wire u2_remHi_435_;
  wire u2_remHi_435__FF_INPUT;
  wire u2_remHi_436_;
  wire u2_remHi_436__FF_INPUT;
  wire u2_remHi_437_;
  wire u2_remHi_437__FF_INPUT;
  wire u2_remHi_438_;
  wire u2_remHi_438__FF_INPUT;
  wire u2_remHi_439_;
  wire u2_remHi_439__FF_INPUT;
  wire u2_remHi_43_;
  wire u2_remHi_43__FF_INPUT;
  wire u2_remHi_440_;
  wire u2_remHi_440__FF_INPUT;
  wire u2_remHi_441_;
  wire u2_remHi_441__FF_INPUT;
  wire u2_remHi_442_;
  wire u2_remHi_442__FF_INPUT;
  wire u2_remHi_443_;
  wire u2_remHi_443__FF_INPUT;
  wire u2_remHi_444_;
  wire u2_remHi_444__FF_INPUT;
  wire u2_remHi_445_;
  wire u2_remHi_445__FF_INPUT;
  wire u2_remHi_446_;
  wire u2_remHi_446__FF_INPUT;
  wire u2_remHi_447_;
  wire u2_remHi_447__FF_INPUT;
  wire u2_remHi_448_;
  wire u2_remHi_448__FF_INPUT;
  wire u2_remHi_449_;
  wire u2_remHi_449__FF_INPUT;
  wire u2_remHi_44_;
  wire u2_remHi_44__FF_INPUT;
  wire u2_remHi_45_;
  wire u2_remHi_45__FF_INPUT;
  wire u2_remHi_46_;
  wire u2_remHi_46__FF_INPUT;
  wire u2_remHi_47_;
  wire u2_remHi_47__FF_INPUT;
  wire u2_remHi_48_;
  wire u2_remHi_48__FF_INPUT;
  wire u2_remHi_49_;
  wire u2_remHi_49__FF_INPUT;
  wire u2_remHi_4_;
  wire u2_remHi_4__FF_INPUT;
  wire u2_remHi_50_;
  wire u2_remHi_50__FF_INPUT;
  wire u2_remHi_51_;
  wire u2_remHi_51__FF_INPUT;
  wire u2_remHi_52_;
  wire u2_remHi_52__FF_INPUT;
  wire u2_remHi_53_;
  wire u2_remHi_53__FF_INPUT;
  wire u2_remHi_54_;
  wire u2_remHi_54__FF_INPUT;
  wire u2_remHi_55_;
  wire u2_remHi_55__FF_INPUT;
  wire u2_remHi_56_;
  wire u2_remHi_56__FF_INPUT;
  wire u2_remHi_57_;
  wire u2_remHi_57__FF_INPUT;
  wire u2_remHi_58_;
  wire u2_remHi_58__FF_INPUT;
  wire u2_remHi_59_;
  wire u2_remHi_59__FF_INPUT;
  wire u2_remHi_5_;
  wire u2_remHi_5__FF_INPUT;
  wire u2_remHi_60_;
  wire u2_remHi_60__FF_INPUT;
  wire u2_remHi_61_;
  wire u2_remHi_61__FF_INPUT;
  wire u2_remHi_62_;
  wire u2_remHi_62__FF_INPUT;
  wire u2_remHi_63_;
  wire u2_remHi_63__FF_INPUT;
  wire u2_remHi_64_;
  wire u2_remHi_64__FF_INPUT;
  wire u2_remHi_65_;
  wire u2_remHi_65__FF_INPUT;
  wire u2_remHi_66_;
  wire u2_remHi_66__FF_INPUT;
  wire u2_remHi_67_;
  wire u2_remHi_67__FF_INPUT;
  wire u2_remHi_68_;
  wire u2_remHi_68__FF_INPUT;
  wire u2_remHi_69_;
  wire u2_remHi_69__FF_INPUT;
  wire u2_remHi_6_;
  wire u2_remHi_6__FF_INPUT;
  wire u2_remHi_70_;
  wire u2_remHi_70__FF_INPUT;
  wire u2_remHi_71_;
  wire u2_remHi_71__FF_INPUT;
  wire u2_remHi_72_;
  wire u2_remHi_72__FF_INPUT;
  wire u2_remHi_73_;
  wire u2_remHi_73__FF_INPUT;
  wire u2_remHi_74_;
  wire u2_remHi_74__FF_INPUT;
  wire u2_remHi_75_;
  wire u2_remHi_75__FF_INPUT;
  wire u2_remHi_76_;
  wire u2_remHi_76__FF_INPUT;
  wire u2_remHi_77_;
  wire u2_remHi_77__FF_INPUT;
  wire u2_remHi_78_;
  wire u2_remHi_78__FF_INPUT;
  wire u2_remHi_79_;
  wire u2_remHi_79__FF_INPUT;
  wire u2_remHi_7_;
  wire u2_remHi_7__FF_INPUT;
  wire u2_remHi_80_;
  wire u2_remHi_80__FF_INPUT;
  wire u2_remHi_81_;
  wire u2_remHi_81__FF_INPUT;
  wire u2_remHi_82_;
  wire u2_remHi_82__FF_INPUT;
  wire u2_remHi_83_;
  wire u2_remHi_83__FF_INPUT;
  wire u2_remHi_84_;
  wire u2_remHi_84__FF_INPUT;
  wire u2_remHi_85_;
  wire u2_remHi_85__FF_INPUT;
  wire u2_remHi_86_;
  wire u2_remHi_86__FF_INPUT;
  wire u2_remHi_87_;
  wire u2_remHi_87__FF_INPUT;
  wire u2_remHi_88_;
  wire u2_remHi_88__FF_INPUT;
  wire u2_remHi_89_;
  wire u2_remHi_89__FF_INPUT;
  wire u2_remHi_8_;
  wire u2_remHi_8__FF_INPUT;
  wire u2_remHi_90_;
  wire u2_remHi_90__FF_INPUT;
  wire u2_remHi_91_;
  wire u2_remHi_91__FF_INPUT;
  wire u2_remHi_92_;
  wire u2_remHi_92__FF_INPUT;
  wire u2_remHi_93_;
  wire u2_remHi_93__FF_INPUT;
  wire u2_remHi_94_;
  wire u2_remHi_94__FF_INPUT;
  wire u2_remHi_95_;
  wire u2_remHi_95__FF_INPUT;
  wire u2_remHi_96_;
  wire u2_remHi_96__FF_INPUT;
  wire u2_remHi_97_;
  wire u2_remHi_97__FF_INPUT;
  wire u2_remHi_98_;
  wire u2_remHi_98__FF_INPUT;
  wire u2_remHi_99_;
  wire u2_remHi_99__FF_INPUT;
  wire u2_remHi_9_;
  wire u2_remHi_9__FF_INPUT;
  wire u2_remLo_0_;
  wire u2_remLo_0__FF_INPUT;
  wire u2_remLo_100_;
  wire u2_remLo_100__FF_INPUT;
  wire u2_remLo_101_;
  wire u2_remLo_101__FF_INPUT;
  wire u2_remLo_102_;
  wire u2_remLo_102__FF_INPUT;
  wire u2_remLo_103_;
  wire u2_remLo_103__FF_INPUT;
  wire u2_remLo_104_;
  wire u2_remLo_104__FF_INPUT;
  wire u2_remLo_105_;
  wire u2_remLo_105__FF_INPUT;
  wire u2_remLo_106_;
  wire u2_remLo_106__FF_INPUT;
  wire u2_remLo_107_;
  wire u2_remLo_107__FF_INPUT;
  wire u2_remLo_108_;
  wire u2_remLo_108__FF_INPUT;
  wire u2_remLo_109_;
  wire u2_remLo_109__FF_INPUT;
  wire u2_remLo_10_;
  wire u2_remLo_10__FF_INPUT;
  wire u2_remLo_110_;
  wire u2_remLo_110__FF_INPUT;
  wire u2_remLo_111_;
  wire u2_remLo_111__FF_INPUT;
  wire u2_remLo_112_;
  wire u2_remLo_112__FF_INPUT;
  wire u2_remLo_113_;
  wire u2_remLo_113__FF_INPUT;
  wire u2_remLo_114_;
  wire u2_remLo_114__FF_INPUT;
  wire u2_remLo_115_;
  wire u2_remLo_115__FF_INPUT;
  wire u2_remLo_116_;
  wire u2_remLo_116__FF_INPUT;
  wire u2_remLo_117_;
  wire u2_remLo_117__FF_INPUT;
  wire u2_remLo_118_;
  wire u2_remLo_118__FF_INPUT;
  wire u2_remLo_119_;
  wire u2_remLo_119__FF_INPUT;
  wire u2_remLo_11_;
  wire u2_remLo_11__FF_INPUT;
  wire u2_remLo_120_;
  wire u2_remLo_120__FF_INPUT;
  wire u2_remLo_121_;
  wire u2_remLo_121__FF_INPUT;
  wire u2_remLo_122_;
  wire u2_remLo_122__FF_INPUT;
  wire u2_remLo_123_;
  wire u2_remLo_123__FF_INPUT;
  wire u2_remLo_124_;
  wire u2_remLo_124__FF_INPUT;
  wire u2_remLo_125_;
  wire u2_remLo_125__FF_INPUT;
  wire u2_remLo_126_;
  wire u2_remLo_126__FF_INPUT;
  wire u2_remLo_127_;
  wire u2_remLo_127__FF_INPUT;
  wire u2_remLo_128_;
  wire u2_remLo_128__FF_INPUT;
  wire u2_remLo_129_;
  wire u2_remLo_129__FF_INPUT;
  wire u2_remLo_12_;
  wire u2_remLo_12__FF_INPUT;
  wire u2_remLo_130_;
  wire u2_remLo_130__FF_INPUT;
  wire u2_remLo_131_;
  wire u2_remLo_131__FF_INPUT;
  wire u2_remLo_132_;
  wire u2_remLo_132__FF_INPUT;
  wire u2_remLo_133_;
  wire u2_remLo_133__FF_INPUT;
  wire u2_remLo_134_;
  wire u2_remLo_134__FF_INPUT;
  wire u2_remLo_135_;
  wire u2_remLo_135__FF_INPUT;
  wire u2_remLo_136_;
  wire u2_remLo_136__FF_INPUT;
  wire u2_remLo_137_;
  wire u2_remLo_137__FF_INPUT;
  wire u2_remLo_138_;
  wire u2_remLo_138__FF_INPUT;
  wire u2_remLo_139_;
  wire u2_remLo_139__FF_INPUT;
  wire u2_remLo_13_;
  wire u2_remLo_13__FF_INPUT;
  wire u2_remLo_140_;
  wire u2_remLo_140__FF_INPUT;
  wire u2_remLo_141_;
  wire u2_remLo_141__FF_INPUT;
  wire u2_remLo_142_;
  wire u2_remLo_142__FF_INPUT;
  wire u2_remLo_143_;
  wire u2_remLo_143__FF_INPUT;
  wire u2_remLo_144_;
  wire u2_remLo_144__FF_INPUT;
  wire u2_remLo_145_;
  wire u2_remLo_145__FF_INPUT;
  wire u2_remLo_146_;
  wire u2_remLo_146__FF_INPUT;
  wire u2_remLo_147_;
  wire u2_remLo_147__FF_INPUT;
  wire u2_remLo_148_;
  wire u2_remLo_148__FF_INPUT;
  wire u2_remLo_149_;
  wire u2_remLo_149__FF_INPUT;
  wire u2_remLo_14_;
  wire u2_remLo_14__FF_INPUT;
  wire u2_remLo_150_;
  wire u2_remLo_150__FF_INPUT;
  wire u2_remLo_151_;
  wire u2_remLo_151__FF_INPUT;
  wire u2_remLo_152_;
  wire u2_remLo_152__FF_INPUT;
  wire u2_remLo_153_;
  wire u2_remLo_153__FF_INPUT;
  wire u2_remLo_154_;
  wire u2_remLo_154__FF_INPUT;
  wire u2_remLo_155_;
  wire u2_remLo_155__FF_INPUT;
  wire u2_remLo_156_;
  wire u2_remLo_156__FF_INPUT;
  wire u2_remLo_157_;
  wire u2_remLo_157__FF_INPUT;
  wire u2_remLo_158_;
  wire u2_remLo_158__FF_INPUT;
  wire u2_remLo_159_;
  wire u2_remLo_159__FF_INPUT;
  wire u2_remLo_15_;
  wire u2_remLo_15__FF_INPUT;
  wire u2_remLo_160_;
  wire u2_remLo_160__FF_INPUT;
  wire u2_remLo_161_;
  wire u2_remLo_161__FF_INPUT;
  wire u2_remLo_162_;
  wire u2_remLo_162__FF_INPUT;
  wire u2_remLo_163_;
  wire u2_remLo_163__FF_INPUT;
  wire u2_remLo_164_;
  wire u2_remLo_164__FF_INPUT;
  wire u2_remLo_165_;
  wire u2_remLo_165__FF_INPUT;
  wire u2_remLo_166_;
  wire u2_remLo_166__FF_INPUT;
  wire u2_remLo_167_;
  wire u2_remLo_167__FF_INPUT;
  wire u2_remLo_168_;
  wire u2_remLo_168__FF_INPUT;
  wire u2_remLo_169_;
  wire u2_remLo_169__FF_INPUT;
  wire u2_remLo_16_;
  wire u2_remLo_16__FF_INPUT;
  wire u2_remLo_170_;
  wire u2_remLo_170__FF_INPUT;
  wire u2_remLo_171_;
  wire u2_remLo_171__FF_INPUT;
  wire u2_remLo_172_;
  wire u2_remLo_172__FF_INPUT;
  wire u2_remLo_173_;
  wire u2_remLo_173__FF_INPUT;
  wire u2_remLo_174_;
  wire u2_remLo_174__FF_INPUT;
  wire u2_remLo_175_;
  wire u2_remLo_175__FF_INPUT;
  wire u2_remLo_176_;
  wire u2_remLo_176__FF_INPUT;
  wire u2_remLo_177_;
  wire u2_remLo_177__FF_INPUT;
  wire u2_remLo_178_;
  wire u2_remLo_178__FF_INPUT;
  wire u2_remLo_179_;
  wire u2_remLo_179__FF_INPUT;
  wire u2_remLo_17_;
  wire u2_remLo_17__FF_INPUT;
  wire u2_remLo_180_;
  wire u2_remLo_180__FF_INPUT;
  wire u2_remLo_181_;
  wire u2_remLo_181__FF_INPUT;
  wire u2_remLo_182_;
  wire u2_remLo_182__FF_INPUT;
  wire u2_remLo_183_;
  wire u2_remLo_183__FF_INPUT;
  wire u2_remLo_184_;
  wire u2_remLo_184__FF_INPUT;
  wire u2_remLo_185_;
  wire u2_remLo_185__FF_INPUT;
  wire u2_remLo_186_;
  wire u2_remLo_186__FF_INPUT;
  wire u2_remLo_187_;
  wire u2_remLo_187__FF_INPUT;
  wire u2_remLo_188_;
  wire u2_remLo_188__FF_INPUT;
  wire u2_remLo_189_;
  wire u2_remLo_189__FF_INPUT;
  wire u2_remLo_18_;
  wire u2_remLo_18__FF_INPUT;
  wire u2_remLo_190_;
  wire u2_remLo_190__FF_INPUT;
  wire u2_remLo_191_;
  wire u2_remLo_191__FF_INPUT;
  wire u2_remLo_192_;
  wire u2_remLo_192__FF_INPUT;
  wire u2_remLo_193_;
  wire u2_remLo_193__FF_INPUT;
  wire u2_remLo_194_;
  wire u2_remLo_194__FF_INPUT;
  wire u2_remLo_195_;
  wire u2_remLo_195__FF_INPUT;
  wire u2_remLo_196_;
  wire u2_remLo_196__FF_INPUT;
  wire u2_remLo_197_;
  wire u2_remLo_197__FF_INPUT;
  wire u2_remLo_198_;
  wire u2_remLo_198__FF_INPUT;
  wire u2_remLo_199_;
  wire u2_remLo_199__FF_INPUT;
  wire u2_remLo_19_;
  wire u2_remLo_19__FF_INPUT;
  wire u2_remLo_1_;
  wire u2_remLo_1__FF_INPUT;
  wire u2_remLo_200_;
  wire u2_remLo_200__FF_INPUT;
  wire u2_remLo_201_;
  wire u2_remLo_201__FF_INPUT;
  wire u2_remLo_202_;
  wire u2_remLo_202__FF_INPUT;
  wire u2_remLo_203_;
  wire u2_remLo_203__FF_INPUT;
  wire u2_remLo_204_;
  wire u2_remLo_204__FF_INPUT;
  wire u2_remLo_205_;
  wire u2_remLo_205__FF_INPUT;
  wire u2_remLo_206_;
  wire u2_remLo_206__FF_INPUT;
  wire u2_remLo_207_;
  wire u2_remLo_207__FF_INPUT;
  wire u2_remLo_208_;
  wire u2_remLo_208__FF_INPUT;
  wire u2_remLo_209_;
  wire u2_remLo_209__FF_INPUT;
  wire u2_remLo_20_;
  wire u2_remLo_20__FF_INPUT;
  wire u2_remLo_210_;
  wire u2_remLo_210__FF_INPUT;
  wire u2_remLo_211_;
  wire u2_remLo_211__FF_INPUT;
  wire u2_remLo_212_;
  wire u2_remLo_212__FF_INPUT;
  wire u2_remLo_213_;
  wire u2_remLo_213__FF_INPUT;
  wire u2_remLo_214_;
  wire u2_remLo_214__FF_INPUT;
  wire u2_remLo_215_;
  wire u2_remLo_215__FF_INPUT;
  wire u2_remLo_216_;
  wire u2_remLo_216__FF_INPUT;
  wire u2_remLo_217_;
  wire u2_remLo_217__FF_INPUT;
  wire u2_remLo_218_;
  wire u2_remLo_218__FF_INPUT;
  wire u2_remLo_219_;
  wire u2_remLo_219__FF_INPUT;
  wire u2_remLo_21_;
  wire u2_remLo_21__FF_INPUT;
  wire u2_remLo_220_;
  wire u2_remLo_220__FF_INPUT;
  wire u2_remLo_221_;
  wire u2_remLo_221__FF_INPUT;
  wire u2_remLo_222_;
  wire u2_remLo_222__FF_INPUT;
  wire u2_remLo_223_;
  wire u2_remLo_223__FF_INPUT;
  wire u2_remLo_224_;
  wire u2_remLo_224__FF_INPUT;
  wire u2_remLo_225_;
  wire u2_remLo_225__FF_INPUT;
  wire u2_remLo_226_;
  wire u2_remLo_226__FF_INPUT;
  wire u2_remLo_227_;
  wire u2_remLo_227__FF_INPUT;
  wire u2_remLo_228_;
  wire u2_remLo_228__FF_INPUT;
  wire u2_remLo_229_;
  wire u2_remLo_229__FF_INPUT;
  wire u2_remLo_22_;
  wire u2_remLo_22__FF_INPUT;
  wire u2_remLo_230_;
  wire u2_remLo_230__FF_INPUT;
  wire u2_remLo_231_;
  wire u2_remLo_231__FF_INPUT;
  wire u2_remLo_232_;
  wire u2_remLo_232__FF_INPUT;
  wire u2_remLo_233_;
  wire u2_remLo_233__FF_INPUT;
  wire u2_remLo_234_;
  wire u2_remLo_234__FF_INPUT;
  wire u2_remLo_235_;
  wire u2_remLo_235__FF_INPUT;
  wire u2_remLo_236_;
  wire u2_remLo_236__FF_INPUT;
  wire u2_remLo_237_;
  wire u2_remLo_237__FF_INPUT;
  wire u2_remLo_238_;
  wire u2_remLo_238__FF_INPUT;
  wire u2_remLo_239_;
  wire u2_remLo_239__FF_INPUT;
  wire u2_remLo_23_;
  wire u2_remLo_23__FF_INPUT;
  wire u2_remLo_240_;
  wire u2_remLo_240__FF_INPUT;
  wire u2_remLo_241_;
  wire u2_remLo_241__FF_INPUT;
  wire u2_remLo_242_;
  wire u2_remLo_242__FF_INPUT;
  wire u2_remLo_243_;
  wire u2_remLo_243__FF_INPUT;
  wire u2_remLo_244_;
  wire u2_remLo_244__FF_INPUT;
  wire u2_remLo_245_;
  wire u2_remLo_245__FF_INPUT;
  wire u2_remLo_246_;
  wire u2_remLo_246__FF_INPUT;
  wire u2_remLo_247_;
  wire u2_remLo_247__FF_INPUT;
  wire u2_remLo_248_;
  wire u2_remLo_248__FF_INPUT;
  wire u2_remLo_249_;
  wire u2_remLo_249__FF_INPUT;
  wire u2_remLo_24_;
  wire u2_remLo_24__FF_INPUT;
  wire u2_remLo_250_;
  wire u2_remLo_250__FF_INPUT;
  wire u2_remLo_251_;
  wire u2_remLo_251__FF_INPUT;
  wire u2_remLo_252_;
  wire u2_remLo_252__FF_INPUT;
  wire u2_remLo_253_;
  wire u2_remLo_253__FF_INPUT;
  wire u2_remLo_254_;
  wire u2_remLo_254__FF_INPUT;
  wire u2_remLo_255_;
  wire u2_remLo_255__FF_INPUT;
  wire u2_remLo_256_;
  wire u2_remLo_256__FF_INPUT;
  wire u2_remLo_257_;
  wire u2_remLo_257__FF_INPUT;
  wire u2_remLo_258_;
  wire u2_remLo_258__FF_INPUT;
  wire u2_remLo_259_;
  wire u2_remLo_259__FF_INPUT;
  wire u2_remLo_25_;
  wire u2_remLo_25__FF_INPUT;
  wire u2_remLo_260_;
  wire u2_remLo_260__FF_INPUT;
  wire u2_remLo_261_;
  wire u2_remLo_261__FF_INPUT;
  wire u2_remLo_262_;
  wire u2_remLo_262__FF_INPUT;
  wire u2_remLo_263_;
  wire u2_remLo_263__FF_INPUT;
  wire u2_remLo_264_;
  wire u2_remLo_264__FF_INPUT;
  wire u2_remLo_265_;
  wire u2_remLo_265__FF_INPUT;
  wire u2_remLo_266_;
  wire u2_remLo_266__FF_INPUT;
  wire u2_remLo_267_;
  wire u2_remLo_267__FF_INPUT;
  wire u2_remLo_268_;
  wire u2_remLo_268__FF_INPUT;
  wire u2_remLo_269_;
  wire u2_remLo_269__FF_INPUT;
  wire u2_remLo_26_;
  wire u2_remLo_26__FF_INPUT;
  wire u2_remLo_270_;
  wire u2_remLo_270__FF_INPUT;
  wire u2_remLo_271_;
  wire u2_remLo_271__FF_INPUT;
  wire u2_remLo_272_;
  wire u2_remLo_272__FF_INPUT;
  wire u2_remLo_273_;
  wire u2_remLo_273__FF_INPUT;
  wire u2_remLo_274_;
  wire u2_remLo_274__FF_INPUT;
  wire u2_remLo_275_;
  wire u2_remLo_275__FF_INPUT;
  wire u2_remLo_276_;
  wire u2_remLo_276__FF_INPUT;
  wire u2_remLo_277_;
  wire u2_remLo_277__FF_INPUT;
  wire u2_remLo_278_;
  wire u2_remLo_278__FF_INPUT;
  wire u2_remLo_279_;
  wire u2_remLo_279__FF_INPUT;
  wire u2_remLo_27_;
  wire u2_remLo_27__FF_INPUT;
  wire u2_remLo_280_;
  wire u2_remLo_280__FF_INPUT;
  wire u2_remLo_281_;
  wire u2_remLo_281__FF_INPUT;
  wire u2_remLo_282_;
  wire u2_remLo_282__FF_INPUT;
  wire u2_remLo_283_;
  wire u2_remLo_283__FF_INPUT;
  wire u2_remLo_284_;
  wire u2_remLo_284__FF_INPUT;
  wire u2_remLo_285_;
  wire u2_remLo_285__FF_INPUT;
  wire u2_remLo_286_;
  wire u2_remLo_286__FF_INPUT;
  wire u2_remLo_287_;
  wire u2_remLo_287__FF_INPUT;
  wire u2_remLo_288_;
  wire u2_remLo_288__FF_INPUT;
  wire u2_remLo_289_;
  wire u2_remLo_289__FF_INPUT;
  wire u2_remLo_28_;
  wire u2_remLo_28__FF_INPUT;
  wire u2_remLo_290_;
  wire u2_remLo_290__FF_INPUT;
  wire u2_remLo_291_;
  wire u2_remLo_291__FF_INPUT;
  wire u2_remLo_292_;
  wire u2_remLo_292__FF_INPUT;
  wire u2_remLo_293_;
  wire u2_remLo_293__FF_INPUT;
  wire u2_remLo_294_;
  wire u2_remLo_294__FF_INPUT;
  wire u2_remLo_295_;
  wire u2_remLo_295__FF_INPUT;
  wire u2_remLo_296_;
  wire u2_remLo_296__FF_INPUT;
  wire u2_remLo_297_;
  wire u2_remLo_297__FF_INPUT;
  wire u2_remLo_298_;
  wire u2_remLo_298__FF_INPUT;
  wire u2_remLo_299_;
  wire u2_remLo_299__FF_INPUT;
  wire u2_remLo_29_;
  wire u2_remLo_29__FF_INPUT;
  wire u2_remLo_2_;
  wire u2_remLo_2__FF_INPUT;
  wire u2_remLo_300_;
  wire u2_remLo_300__FF_INPUT;
  wire u2_remLo_301_;
  wire u2_remLo_301__FF_INPUT;
  wire u2_remLo_302_;
  wire u2_remLo_302__FF_INPUT;
  wire u2_remLo_303_;
  wire u2_remLo_303__FF_INPUT;
  wire u2_remLo_304_;
  wire u2_remLo_304__FF_INPUT;
  wire u2_remLo_305_;
  wire u2_remLo_305__FF_INPUT;
  wire u2_remLo_306_;
  wire u2_remLo_306__FF_INPUT;
  wire u2_remLo_307_;
  wire u2_remLo_307__FF_INPUT;
  wire u2_remLo_308_;
  wire u2_remLo_308__FF_INPUT;
  wire u2_remLo_309_;
  wire u2_remLo_309__FF_INPUT;
  wire u2_remLo_30_;
  wire u2_remLo_30__FF_INPUT;
  wire u2_remLo_310_;
  wire u2_remLo_310__FF_INPUT;
  wire u2_remLo_311_;
  wire u2_remLo_311__FF_INPUT;
  wire u2_remLo_312_;
  wire u2_remLo_312__FF_INPUT;
  wire u2_remLo_313_;
  wire u2_remLo_313__FF_INPUT;
  wire u2_remLo_314_;
  wire u2_remLo_314__FF_INPUT;
  wire u2_remLo_315_;
  wire u2_remLo_315__FF_INPUT;
  wire u2_remLo_316_;
  wire u2_remLo_316__FF_INPUT;
  wire u2_remLo_317_;
  wire u2_remLo_317__FF_INPUT;
  wire u2_remLo_318_;
  wire u2_remLo_318__FF_INPUT;
  wire u2_remLo_319_;
  wire u2_remLo_319__FF_INPUT;
  wire u2_remLo_31_;
  wire u2_remLo_31__FF_INPUT;
  wire u2_remLo_320_;
  wire u2_remLo_320__FF_INPUT;
  wire u2_remLo_321_;
  wire u2_remLo_321__FF_INPUT;
  wire u2_remLo_322_;
  wire u2_remLo_322__FF_INPUT;
  wire u2_remLo_323_;
  wire u2_remLo_323__FF_INPUT;
  wire u2_remLo_324_;
  wire u2_remLo_324__FF_INPUT;
  wire u2_remLo_325_;
  wire u2_remLo_325__FF_INPUT;
  wire u2_remLo_326_;
  wire u2_remLo_326__FF_INPUT;
  wire u2_remLo_327_;
  wire u2_remLo_327__FF_INPUT;
  wire u2_remLo_328_;
  wire u2_remLo_328__FF_INPUT;
  wire u2_remLo_329_;
  wire u2_remLo_329__FF_INPUT;
  wire u2_remLo_32_;
  wire u2_remLo_32__FF_INPUT;
  wire u2_remLo_330_;
  wire u2_remLo_330__FF_INPUT;
  wire u2_remLo_331_;
  wire u2_remLo_331__FF_INPUT;
  wire u2_remLo_332_;
  wire u2_remLo_332__FF_INPUT;
  wire u2_remLo_333_;
  wire u2_remLo_333__FF_INPUT;
  wire u2_remLo_334_;
  wire u2_remLo_334__FF_INPUT;
  wire u2_remLo_335_;
  wire u2_remLo_335__FF_INPUT;
  wire u2_remLo_336_;
  wire u2_remLo_336__FF_INPUT;
  wire u2_remLo_337_;
  wire u2_remLo_337__FF_INPUT;
  wire u2_remLo_338_;
  wire u2_remLo_338__FF_INPUT;
  wire u2_remLo_339_;
  wire u2_remLo_339__FF_INPUT;
  wire u2_remLo_33_;
  wire u2_remLo_33__FF_INPUT;
  wire u2_remLo_340_;
  wire u2_remLo_340__FF_INPUT;
  wire u2_remLo_341_;
  wire u2_remLo_341__FF_INPUT;
  wire u2_remLo_342_;
  wire u2_remLo_342__FF_INPUT;
  wire u2_remLo_343_;
  wire u2_remLo_343__FF_INPUT;
  wire u2_remLo_344_;
  wire u2_remLo_344__FF_INPUT;
  wire u2_remLo_345_;
  wire u2_remLo_345__FF_INPUT;
  wire u2_remLo_346_;
  wire u2_remLo_346__FF_INPUT;
  wire u2_remLo_347_;
  wire u2_remLo_347__FF_INPUT;
  wire u2_remLo_348_;
  wire u2_remLo_348__FF_INPUT;
  wire u2_remLo_349_;
  wire u2_remLo_349__FF_INPUT;
  wire u2_remLo_34_;
  wire u2_remLo_34__FF_INPUT;
  wire u2_remLo_350_;
  wire u2_remLo_350__FF_INPUT;
  wire u2_remLo_351_;
  wire u2_remLo_351__FF_INPUT;
  wire u2_remLo_352_;
  wire u2_remLo_352__FF_INPUT;
  wire u2_remLo_353_;
  wire u2_remLo_353__FF_INPUT;
  wire u2_remLo_354_;
  wire u2_remLo_354__FF_INPUT;
  wire u2_remLo_355_;
  wire u2_remLo_355__FF_INPUT;
  wire u2_remLo_356_;
  wire u2_remLo_356__FF_INPUT;
  wire u2_remLo_357_;
  wire u2_remLo_357__FF_INPUT;
  wire u2_remLo_358_;
  wire u2_remLo_358__FF_INPUT;
  wire u2_remLo_359_;
  wire u2_remLo_359__FF_INPUT;
  wire u2_remLo_35_;
  wire u2_remLo_35__FF_INPUT;
  wire u2_remLo_360_;
  wire u2_remLo_360__FF_INPUT;
  wire u2_remLo_361_;
  wire u2_remLo_361__FF_INPUT;
  wire u2_remLo_362_;
  wire u2_remLo_362__FF_INPUT;
  wire u2_remLo_363_;
  wire u2_remLo_363__FF_INPUT;
  wire u2_remLo_364_;
  wire u2_remLo_364__FF_INPUT;
  wire u2_remLo_365_;
  wire u2_remLo_365__FF_INPUT;
  wire u2_remLo_366_;
  wire u2_remLo_366__FF_INPUT;
  wire u2_remLo_367_;
  wire u2_remLo_367__FF_INPUT;
  wire u2_remLo_368_;
  wire u2_remLo_368__FF_INPUT;
  wire u2_remLo_369_;
  wire u2_remLo_369__FF_INPUT;
  wire u2_remLo_36_;
  wire u2_remLo_36__FF_INPUT;
  wire u2_remLo_370_;
  wire u2_remLo_370__FF_INPUT;
  wire u2_remLo_371_;
  wire u2_remLo_371__FF_INPUT;
  wire u2_remLo_372_;
  wire u2_remLo_372__FF_INPUT;
  wire u2_remLo_373_;
  wire u2_remLo_373__FF_INPUT;
  wire u2_remLo_374_;
  wire u2_remLo_374__FF_INPUT;
  wire u2_remLo_375_;
  wire u2_remLo_375__FF_INPUT;
  wire u2_remLo_376_;
  wire u2_remLo_376__FF_INPUT;
  wire u2_remLo_377_;
  wire u2_remLo_377__FF_INPUT;
  wire u2_remLo_378_;
  wire u2_remLo_378__FF_INPUT;
  wire u2_remLo_379_;
  wire u2_remLo_379__FF_INPUT;
  wire u2_remLo_37_;
  wire u2_remLo_37__FF_INPUT;
  wire u2_remLo_380_;
  wire u2_remLo_380__FF_INPUT;
  wire u2_remLo_381_;
  wire u2_remLo_381__FF_INPUT;
  wire u2_remLo_382_;
  wire u2_remLo_382__FF_INPUT;
  wire u2_remLo_383_;
  wire u2_remLo_383__FF_INPUT;
  wire u2_remLo_384_;
  wire u2_remLo_384__FF_INPUT;
  wire u2_remLo_385_;
  wire u2_remLo_385__FF_INPUT;
  wire u2_remLo_386_;
  wire u2_remLo_386__FF_INPUT;
  wire u2_remLo_387_;
  wire u2_remLo_387__FF_INPUT;
  wire u2_remLo_388_;
  wire u2_remLo_388__FF_INPUT;
  wire u2_remLo_389_;
  wire u2_remLo_389__FF_INPUT;
  wire u2_remLo_38_;
  wire u2_remLo_38__FF_INPUT;
  wire u2_remLo_390_;
  wire u2_remLo_390__FF_INPUT;
  wire u2_remLo_391_;
  wire u2_remLo_391__FF_INPUT;
  wire u2_remLo_392_;
  wire u2_remLo_392__FF_INPUT;
  wire u2_remLo_393_;
  wire u2_remLo_393__FF_INPUT;
  wire u2_remLo_394_;
  wire u2_remLo_394__FF_INPUT;
  wire u2_remLo_395_;
  wire u2_remLo_395__FF_INPUT;
  wire u2_remLo_396_;
  wire u2_remLo_396__FF_INPUT;
  wire u2_remLo_397_;
  wire u2_remLo_397__FF_INPUT;
  wire u2_remLo_398_;
  wire u2_remLo_398__FF_INPUT;
  wire u2_remLo_399_;
  wire u2_remLo_399__FF_INPUT;
  wire u2_remLo_39_;
  wire u2_remLo_39__FF_INPUT;
  wire u2_remLo_3_;
  wire u2_remLo_3__FF_INPUT;
  wire u2_remLo_400_;
  wire u2_remLo_400__FF_INPUT;
  wire u2_remLo_401_;
  wire u2_remLo_401__FF_INPUT;
  wire u2_remLo_402_;
  wire u2_remLo_402__FF_INPUT;
  wire u2_remLo_403_;
  wire u2_remLo_403__FF_INPUT;
  wire u2_remLo_404_;
  wire u2_remLo_404__FF_INPUT;
  wire u2_remLo_405_;
  wire u2_remLo_405__FF_INPUT;
  wire u2_remLo_406_;
  wire u2_remLo_406__FF_INPUT;
  wire u2_remLo_407_;
  wire u2_remLo_407__FF_INPUT;
  wire u2_remLo_408_;
  wire u2_remLo_408__FF_INPUT;
  wire u2_remLo_409_;
  wire u2_remLo_409__FF_INPUT;
  wire u2_remLo_40_;
  wire u2_remLo_40__FF_INPUT;
  wire u2_remLo_410_;
  wire u2_remLo_410__FF_INPUT;
  wire u2_remLo_411_;
  wire u2_remLo_411__FF_INPUT;
  wire u2_remLo_412_;
  wire u2_remLo_412__FF_INPUT;
  wire u2_remLo_413_;
  wire u2_remLo_413__FF_INPUT;
  wire u2_remLo_414_;
  wire u2_remLo_414__FF_INPUT;
  wire u2_remLo_415_;
  wire u2_remLo_415__FF_INPUT;
  wire u2_remLo_416_;
  wire u2_remLo_416__FF_INPUT;
  wire u2_remLo_417_;
  wire u2_remLo_417__FF_INPUT;
  wire u2_remLo_418_;
  wire u2_remLo_418__FF_INPUT;
  wire u2_remLo_419_;
  wire u2_remLo_419__FF_INPUT;
  wire u2_remLo_41_;
  wire u2_remLo_41__FF_INPUT;
  wire u2_remLo_420_;
  wire u2_remLo_420__FF_INPUT;
  wire u2_remLo_421_;
  wire u2_remLo_421__FF_INPUT;
  wire u2_remLo_422_;
  wire u2_remLo_422__FF_INPUT;
  wire u2_remLo_423_;
  wire u2_remLo_423__FF_INPUT;
  wire u2_remLo_424_;
  wire u2_remLo_424__FF_INPUT;
  wire u2_remLo_425_;
  wire u2_remLo_425__FF_INPUT;
  wire u2_remLo_426_;
  wire u2_remLo_426__FF_INPUT;
  wire u2_remLo_427_;
  wire u2_remLo_427__FF_INPUT;
  wire u2_remLo_428_;
  wire u2_remLo_428__FF_INPUT;
  wire u2_remLo_429_;
  wire u2_remLo_429__FF_INPUT;
  wire u2_remLo_42_;
  wire u2_remLo_42__FF_INPUT;
  wire u2_remLo_430_;
  wire u2_remLo_430__FF_INPUT;
  wire u2_remLo_431_;
  wire u2_remLo_431__FF_INPUT;
  wire u2_remLo_432_;
  wire u2_remLo_432__FF_INPUT;
  wire u2_remLo_433_;
  wire u2_remLo_433__FF_INPUT;
  wire u2_remLo_434_;
  wire u2_remLo_434__FF_INPUT;
  wire u2_remLo_435_;
  wire u2_remLo_435__FF_INPUT;
  wire u2_remLo_436_;
  wire u2_remLo_436__FF_INPUT;
  wire u2_remLo_437_;
  wire u2_remLo_437__FF_INPUT;
  wire u2_remLo_438_;
  wire u2_remLo_438__FF_INPUT;
  wire u2_remLo_439_;
  wire u2_remLo_439__FF_INPUT;
  wire u2_remLo_43_;
  wire u2_remLo_43__FF_INPUT;
  wire u2_remLo_440_;
  wire u2_remLo_440__FF_INPUT;
  wire u2_remLo_441_;
  wire u2_remLo_441__FF_INPUT;
  wire u2_remLo_442_;
  wire u2_remLo_442__FF_INPUT;
  wire u2_remLo_443_;
  wire u2_remLo_443__FF_INPUT;
  wire u2_remLo_444_;
  wire u2_remLo_444__FF_INPUT;
  wire u2_remLo_445_;
  wire u2_remLo_445__FF_INPUT;
  wire u2_remLo_446_;
  wire u2_remLo_446__FF_INPUT;
  wire u2_remLo_447_;
  wire u2_remLo_447__FF_INPUT;
  wire u2_remLo_448_;
  wire u2_remLo_448__FF_INPUT;
  wire u2_remLo_449_;
  wire u2_remLo_449__FF_INPUT;
  wire u2_remLo_44_;
  wire u2_remLo_44__FF_INPUT;
  wire u2_remLo_450__FF_INPUT;
  wire u2_remLo_451__FF_INPUT;
  wire u2_remLo_45_;
  wire u2_remLo_45__FF_INPUT;
  wire u2_remLo_46_;
  wire u2_remLo_46__FF_INPUT;
  wire u2_remLo_47_;
  wire u2_remLo_47__FF_INPUT;
  wire u2_remLo_48_;
  wire u2_remLo_48__FF_INPUT;
  wire u2_remLo_49_;
  wire u2_remLo_49__FF_INPUT;
  wire u2_remLo_4_;
  wire u2_remLo_4__FF_INPUT;
  wire u2_remLo_50_;
  wire u2_remLo_50__FF_INPUT;
  wire u2_remLo_51_;
  wire u2_remLo_51__FF_INPUT;
  wire u2_remLo_52_;
  wire u2_remLo_52__FF_INPUT;
  wire u2_remLo_53_;
  wire u2_remLo_53__FF_INPUT;
  wire u2_remLo_54_;
  wire u2_remLo_54__FF_INPUT;
  wire u2_remLo_55_;
  wire u2_remLo_55__FF_INPUT;
  wire u2_remLo_56_;
  wire u2_remLo_56__FF_INPUT;
  wire u2_remLo_57_;
  wire u2_remLo_57__FF_INPUT;
  wire u2_remLo_58_;
  wire u2_remLo_58__FF_INPUT;
  wire u2_remLo_59_;
  wire u2_remLo_59__FF_INPUT;
  wire u2_remLo_5_;
  wire u2_remLo_5__FF_INPUT;
  wire u2_remLo_60_;
  wire u2_remLo_60__FF_INPUT;
  wire u2_remLo_61_;
  wire u2_remLo_61__FF_INPUT;
  wire u2_remLo_62_;
  wire u2_remLo_62__FF_INPUT;
  wire u2_remLo_63_;
  wire u2_remLo_63__FF_INPUT;
  wire u2_remLo_64_;
  wire u2_remLo_64__FF_INPUT;
  wire u2_remLo_65_;
  wire u2_remLo_65__FF_INPUT;
  wire u2_remLo_66_;
  wire u2_remLo_66__FF_INPUT;
  wire u2_remLo_67_;
  wire u2_remLo_67__FF_INPUT;
  wire u2_remLo_68_;
  wire u2_remLo_68__FF_INPUT;
  wire u2_remLo_69_;
  wire u2_remLo_69__FF_INPUT;
  wire u2_remLo_6_;
  wire u2_remLo_6__FF_INPUT;
  wire u2_remLo_70_;
  wire u2_remLo_70__FF_INPUT;
  wire u2_remLo_71_;
  wire u2_remLo_71__FF_INPUT;
  wire u2_remLo_72_;
  wire u2_remLo_72__FF_INPUT;
  wire u2_remLo_73_;
  wire u2_remLo_73__FF_INPUT;
  wire u2_remLo_74_;
  wire u2_remLo_74__FF_INPUT;
  wire u2_remLo_75_;
  wire u2_remLo_75__FF_INPUT;
  wire u2_remLo_76_;
  wire u2_remLo_76__FF_INPUT;
  wire u2_remLo_77_;
  wire u2_remLo_77__FF_INPUT;
  wire u2_remLo_78_;
  wire u2_remLo_78__FF_INPUT;
  wire u2_remLo_79_;
  wire u2_remLo_79__FF_INPUT;
  wire u2_remLo_7_;
  wire u2_remLo_7__FF_INPUT;
  wire u2_remLo_80_;
  wire u2_remLo_80__FF_INPUT;
  wire u2_remLo_81_;
  wire u2_remLo_81__FF_INPUT;
  wire u2_remLo_82_;
  wire u2_remLo_82__FF_INPUT;
  wire u2_remLo_83_;
  wire u2_remLo_83__FF_INPUT;
  wire u2_remLo_84_;
  wire u2_remLo_84__FF_INPUT;
  wire u2_remLo_85_;
  wire u2_remLo_85__FF_INPUT;
  wire u2_remLo_86_;
  wire u2_remLo_86__FF_INPUT;
  wire u2_remLo_87_;
  wire u2_remLo_87__FF_INPUT;
  wire u2_remLo_88_;
  wire u2_remLo_88__FF_INPUT;
  wire u2_remLo_89_;
  wire u2_remLo_89__FF_INPUT;
  wire u2_remLo_8_;
  wire u2_remLo_8__FF_INPUT;
  wire u2_remLo_90_;
  wire u2_remLo_90__FF_INPUT;
  wire u2_remLo_91_;
  wire u2_remLo_91__FF_INPUT;
  wire u2_remLo_92_;
  wire u2_remLo_92__FF_INPUT;
  wire u2_remLo_93_;
  wire u2_remLo_93__FF_INPUT;
  wire u2_remLo_94_;
  wire u2_remLo_94__FF_INPUT;
  wire u2_remLo_95_;
  wire u2_remLo_95__FF_INPUT;
  wire u2_remLo_96_;
  wire u2_remLo_96__FF_INPUT;
  wire u2_remLo_97_;
  wire u2_remLo_97__FF_INPUT;
  wire u2_remLo_98_;
  wire u2_remLo_98__FF_INPUT;
  wire u2_remLo_99_;
  wire u2_remLo_99__FF_INPUT;
  wire u2_remLo_9_;
  wire u2_remLo_9__FF_INPUT;
  wire u2_root_0_;
  wire u2_root_0__FF_INPUT;
  wire u2_root_100__FF_INPUT;
  wire u2_root_101__FF_INPUT;
  wire u2_root_102__FF_INPUT;
  wire u2_root_103__FF_INPUT;
  wire u2_root_104__FF_INPUT;
  wire u2_root_105__FF_INPUT;
  wire u2_root_106__FF_INPUT;
  wire u2_root_107__FF_INPUT;
  wire u2_root_108__FF_INPUT;
  wire u2_root_109__FF_INPUT;
  wire u2_root_10__FF_INPUT;
  wire u2_root_110__FF_INPUT;
  wire u2_root_111__FF_INPUT;
  wire u2_root_112__FF_INPUT;
  wire u2_root_113__FF_INPUT;
  wire u2_root_114__FF_INPUT;
  wire u2_root_115__FF_INPUT;
  wire u2_root_116__FF_INPUT;
  wire u2_root_117__FF_INPUT;
  wire u2_root_118__FF_INPUT;
  wire u2_root_119__FF_INPUT;
  wire u2_root_11__FF_INPUT;
  wire u2_root_120__FF_INPUT;
  wire u2_root_121__FF_INPUT;
  wire u2_root_122__FF_INPUT;
  wire u2_root_123__FF_INPUT;
  wire u2_root_124__FF_INPUT;
  wire u2_root_125__FF_INPUT;
  wire u2_root_126__FF_INPUT;
  wire u2_root_127__FF_INPUT;
  wire u2_root_128__FF_INPUT;
  wire u2_root_129__FF_INPUT;
  wire u2_root_12__FF_INPUT;
  wire u2_root_130__FF_INPUT;
  wire u2_root_131__FF_INPUT;
  wire u2_root_132__FF_INPUT;
  wire u2_root_133__FF_INPUT;
  wire u2_root_134__FF_INPUT;
  wire u2_root_135__FF_INPUT;
  wire u2_root_136__FF_INPUT;
  wire u2_root_137__FF_INPUT;
  wire u2_root_138__FF_INPUT;
  wire u2_root_139__FF_INPUT;
  wire u2_root_13__FF_INPUT;
  wire u2_root_140__FF_INPUT;
  wire u2_root_141__FF_INPUT;
  wire u2_root_142__FF_INPUT;
  wire u2_root_143__FF_INPUT;
  wire u2_root_144__FF_INPUT;
  wire u2_root_145__FF_INPUT;
  wire u2_root_146__FF_INPUT;
  wire u2_root_147__FF_INPUT;
  wire u2_root_148__FF_INPUT;
  wire u2_root_149__FF_INPUT;
  wire u2_root_14__FF_INPUT;
  wire u2_root_150__FF_INPUT;
  wire u2_root_151__FF_INPUT;
  wire u2_root_152__FF_INPUT;
  wire u2_root_153__FF_INPUT;
  wire u2_root_154__FF_INPUT;
  wire u2_root_155__FF_INPUT;
  wire u2_root_156__FF_INPUT;
  wire u2_root_157__FF_INPUT;
  wire u2_root_158__FF_INPUT;
  wire u2_root_159__FF_INPUT;
  wire u2_root_15__FF_INPUT;
  wire u2_root_160__FF_INPUT;
  wire u2_root_161__FF_INPUT;
  wire u2_root_162__FF_INPUT;
  wire u2_root_163__FF_INPUT;
  wire u2_root_164__FF_INPUT;
  wire u2_root_165__FF_INPUT;
  wire u2_root_166__FF_INPUT;
  wire u2_root_167__FF_INPUT;
  wire u2_root_168__FF_INPUT;
  wire u2_root_169__FF_INPUT;
  wire u2_root_16__FF_INPUT;
  wire u2_root_170__FF_INPUT;
  wire u2_root_171__FF_INPUT;
  wire u2_root_172__FF_INPUT;
  wire u2_root_173__FF_INPUT;
  wire u2_root_174__FF_INPUT;
  wire u2_root_175__FF_INPUT;
  wire u2_root_176__FF_INPUT;
  wire u2_root_177__FF_INPUT;
  wire u2_root_178__FF_INPUT;
  wire u2_root_179__FF_INPUT;
  wire u2_root_17__FF_INPUT;
  wire u2_root_180__FF_INPUT;
  wire u2_root_181__FF_INPUT;
  wire u2_root_182__FF_INPUT;
  wire u2_root_183__FF_INPUT;
  wire u2_root_184__FF_INPUT;
  wire u2_root_185__FF_INPUT;
  wire u2_root_186__FF_INPUT;
  wire u2_root_187__FF_INPUT;
  wire u2_root_188__FF_INPUT;
  wire u2_root_189__FF_INPUT;
  wire u2_root_18__FF_INPUT;
  wire u2_root_190__FF_INPUT;
  wire u2_root_191__FF_INPUT;
  wire u2_root_192__FF_INPUT;
  wire u2_root_193__FF_INPUT;
  wire u2_root_194__FF_INPUT;
  wire u2_root_195__FF_INPUT;
  wire u2_root_196__FF_INPUT;
  wire u2_root_197__FF_INPUT;
  wire u2_root_198__FF_INPUT;
  wire u2_root_199__FF_INPUT;
  wire u2_root_19__FF_INPUT;
  wire u2_root_1__FF_INPUT;
  wire u2_root_200__FF_INPUT;
  wire u2_root_201__FF_INPUT;
  wire u2_root_202__FF_INPUT;
  wire u2_root_203__FF_INPUT;
  wire u2_root_204__FF_INPUT;
  wire u2_root_205__FF_INPUT;
  wire u2_root_206__FF_INPUT;
  wire u2_root_207__FF_INPUT;
  wire u2_root_208__FF_INPUT;
  wire u2_root_209__FF_INPUT;
  wire u2_root_20__FF_INPUT;
  wire u2_root_210__FF_INPUT;
  wire u2_root_211__FF_INPUT;
  wire u2_root_212__FF_INPUT;
  wire u2_root_213__FF_INPUT;
  wire u2_root_214__FF_INPUT;
  wire u2_root_215__FF_INPUT;
  wire u2_root_216__FF_INPUT;
  wire u2_root_217__FF_INPUT;
  wire u2_root_218__FF_INPUT;
  wire u2_root_219__FF_INPUT;
  wire u2_root_21__FF_INPUT;
  wire u2_root_220__FF_INPUT;
  wire u2_root_221__FF_INPUT;
  wire u2_root_222__FF_INPUT;
  wire u2_root_223__FF_INPUT;
  wire u2_root_224__FF_INPUT;
  wire u2_root_225__FF_INPUT;
  wire u2_root_226__FF_INPUT;
  wire u2_root_227__FF_INPUT;
  wire u2_root_228__FF_INPUT;
  wire u2_root_229__FF_INPUT;
  wire u2_root_22__FF_INPUT;
  wire u2_root_230__FF_INPUT;
  wire u2_root_231__FF_INPUT;
  wire u2_root_232__FF_INPUT;
  wire u2_root_233__FF_INPUT;
  wire u2_root_234__FF_INPUT;
  wire u2_root_235__FF_INPUT;
  wire u2_root_236__FF_INPUT;
  wire u2_root_237__FF_INPUT;
  wire u2_root_238__FF_INPUT;
  wire u2_root_239__FF_INPUT;
  wire u2_root_23__FF_INPUT;
  wire u2_root_240__FF_INPUT;
  wire u2_root_241__FF_INPUT;
  wire u2_root_242__FF_INPUT;
  wire u2_root_243__FF_INPUT;
  wire u2_root_244__FF_INPUT;
  wire u2_root_245__FF_INPUT;
  wire u2_root_246__FF_INPUT;
  wire u2_root_247__FF_INPUT;
  wire u2_root_248__FF_INPUT;
  wire u2_root_249__FF_INPUT;
  wire u2_root_24__FF_INPUT;
  wire u2_root_250__FF_INPUT;
  wire u2_root_251__FF_INPUT;
  wire u2_root_252__FF_INPUT;
  wire u2_root_253__FF_INPUT;
  wire u2_root_254__FF_INPUT;
  wire u2_root_255__FF_INPUT;
  wire u2_root_256__FF_INPUT;
  wire u2_root_257__FF_INPUT;
  wire u2_root_258__FF_INPUT;
  wire u2_root_259__FF_INPUT;
  wire u2_root_25__FF_INPUT;
  wire u2_root_260__FF_INPUT;
  wire u2_root_261__FF_INPUT;
  wire u2_root_262__FF_INPUT;
  wire u2_root_263__FF_INPUT;
  wire u2_root_264__FF_INPUT;
  wire u2_root_265__FF_INPUT;
  wire u2_root_266__FF_INPUT;
  wire u2_root_267__FF_INPUT;
  wire u2_root_268__FF_INPUT;
  wire u2_root_269__FF_INPUT;
  wire u2_root_26__FF_INPUT;
  wire u2_root_270__FF_INPUT;
  wire u2_root_271__FF_INPUT;
  wire u2_root_272__FF_INPUT;
  wire u2_root_273__FF_INPUT;
  wire u2_root_274__FF_INPUT;
  wire u2_root_275__FF_INPUT;
  wire u2_root_276__FF_INPUT;
  wire u2_root_277__FF_INPUT;
  wire u2_root_278__FF_INPUT;
  wire u2_root_279__FF_INPUT;
  wire u2_root_27__FF_INPUT;
  wire u2_root_280__FF_INPUT;
  wire u2_root_281__FF_INPUT;
  wire u2_root_282__FF_INPUT;
  wire u2_root_283__FF_INPUT;
  wire u2_root_284__FF_INPUT;
  wire u2_root_285__FF_INPUT;
  wire u2_root_286__FF_INPUT;
  wire u2_root_287__FF_INPUT;
  wire u2_root_288__FF_INPUT;
  wire u2_root_289__FF_INPUT;
  wire u2_root_28__FF_INPUT;
  wire u2_root_290__FF_INPUT;
  wire u2_root_291__FF_INPUT;
  wire u2_root_292__FF_INPUT;
  wire u2_root_293__FF_INPUT;
  wire u2_root_294__FF_INPUT;
  wire u2_root_295__FF_INPUT;
  wire u2_root_296__FF_INPUT;
  wire u2_root_297__FF_INPUT;
  wire u2_root_298__FF_INPUT;
  wire u2_root_299__FF_INPUT;
  wire u2_root_29__FF_INPUT;
  wire u2_root_2__FF_INPUT;
  wire u2_root_300__FF_INPUT;
  wire u2_root_301__FF_INPUT;
  wire u2_root_302__FF_INPUT;
  wire u2_root_303__FF_INPUT;
  wire u2_root_304__FF_INPUT;
  wire u2_root_305__FF_INPUT;
  wire u2_root_306__FF_INPUT;
  wire u2_root_307__FF_INPUT;
  wire u2_root_308__FF_INPUT;
  wire u2_root_309__FF_INPUT;
  wire u2_root_30__FF_INPUT;
  wire u2_root_310__FF_INPUT;
  wire u2_root_311__FF_INPUT;
  wire u2_root_312__FF_INPUT;
  wire u2_root_313__FF_INPUT;
  wire u2_root_314__FF_INPUT;
  wire u2_root_315__FF_INPUT;
  wire u2_root_316__FF_INPUT;
  wire u2_root_317__FF_INPUT;
  wire u2_root_318__FF_INPUT;
  wire u2_root_319__FF_INPUT;
  wire u2_root_31__FF_INPUT;
  wire u2_root_320__FF_INPUT;
  wire u2_root_321__FF_INPUT;
  wire u2_root_322__FF_INPUT;
  wire u2_root_323__FF_INPUT;
  wire u2_root_324__FF_INPUT;
  wire u2_root_325__FF_INPUT;
  wire u2_root_326__FF_INPUT;
  wire u2_root_327__FF_INPUT;
  wire u2_root_328__FF_INPUT;
  wire u2_root_329__FF_INPUT;
  wire u2_root_32__FF_INPUT;
  wire u2_root_330__FF_INPUT;
  wire u2_root_331__FF_INPUT;
  wire u2_root_332__FF_INPUT;
  wire u2_root_333__FF_INPUT;
  wire u2_root_334__FF_INPUT;
  wire u2_root_335__FF_INPUT;
  wire u2_root_336__FF_INPUT;
  wire u2_root_337__FF_INPUT;
  wire u2_root_338__FF_INPUT;
  wire u2_root_339__FF_INPUT;
  wire u2_root_33__FF_INPUT;
  wire u2_root_340__FF_INPUT;
  wire u2_root_341__FF_INPUT;
  wire u2_root_342__FF_INPUT;
  wire u2_root_343__FF_INPUT;
  wire u2_root_344__FF_INPUT;
  wire u2_root_345__FF_INPUT;
  wire u2_root_346__FF_INPUT;
  wire u2_root_347__FF_INPUT;
  wire u2_root_348__FF_INPUT;
  wire u2_root_349__FF_INPUT;
  wire u2_root_34__FF_INPUT;
  wire u2_root_350__FF_INPUT;
  wire u2_root_351__FF_INPUT;
  wire u2_root_352__FF_INPUT;
  wire u2_root_353__FF_INPUT;
  wire u2_root_354__FF_INPUT;
  wire u2_root_355__FF_INPUT;
  wire u2_root_356__FF_INPUT;
  wire u2_root_357__FF_INPUT;
  wire u2_root_358__FF_INPUT;
  wire u2_root_359__FF_INPUT;
  wire u2_root_35__FF_INPUT;
  wire u2_root_360__FF_INPUT;
  wire u2_root_361__FF_INPUT;
  wire u2_root_362__FF_INPUT;
  wire u2_root_363__FF_INPUT;
  wire u2_root_364__FF_INPUT;
  wire u2_root_365__FF_INPUT;
  wire u2_root_366__FF_INPUT;
  wire u2_root_367__FF_INPUT;
  wire u2_root_368__FF_INPUT;
  wire u2_root_369__FF_INPUT;
  wire u2_root_36__FF_INPUT;
  wire u2_root_370__FF_INPUT;
  wire u2_root_371__FF_INPUT;
  wire u2_root_372__FF_INPUT;
  wire u2_root_373__FF_INPUT;
  wire u2_root_374__FF_INPUT;
  wire u2_root_375__FF_INPUT;
  wire u2_root_376__FF_INPUT;
  wire u2_root_377__FF_INPUT;
  wire u2_root_378__FF_INPUT;
  wire u2_root_379__FF_INPUT;
  wire u2_root_37__FF_INPUT;
  wire u2_root_380__FF_INPUT;
  wire u2_root_381__FF_INPUT;
  wire u2_root_382__FF_INPUT;
  wire u2_root_383__FF_INPUT;
  wire u2_root_384__FF_INPUT;
  wire u2_root_385__FF_INPUT;
  wire u2_root_386__FF_INPUT;
  wire u2_root_387__FF_INPUT;
  wire u2_root_388__FF_INPUT;
  wire u2_root_389__FF_INPUT;
  wire u2_root_38__FF_INPUT;
  wire u2_root_390__FF_INPUT;
  wire u2_root_391__FF_INPUT;
  wire u2_root_392__FF_INPUT;
  wire u2_root_393__FF_INPUT;
  wire u2_root_394__FF_INPUT;
  wire u2_root_395__FF_INPUT;
  wire u2_root_396__FF_INPUT;
  wire u2_root_397__FF_INPUT;
  wire u2_root_398__FF_INPUT;
  wire u2_root_399__FF_INPUT;
  wire u2_root_39__FF_INPUT;
  wire u2_root_3__FF_INPUT;
  wire u2_root_400__FF_INPUT;
  wire u2_root_401__FF_INPUT;
  wire u2_root_402__FF_INPUT;
  wire u2_root_403__FF_INPUT;
  wire u2_root_404__FF_INPUT;
  wire u2_root_405__FF_INPUT;
  wire u2_root_406__FF_INPUT;
  wire u2_root_407__FF_INPUT;
  wire u2_root_408__FF_INPUT;
  wire u2_root_409__FF_INPUT;
  wire u2_root_40__FF_INPUT;
  wire u2_root_410__FF_INPUT;
  wire u2_root_411__FF_INPUT;
  wire u2_root_412__FF_INPUT;
  wire u2_root_413__FF_INPUT;
  wire u2_root_414__FF_INPUT;
  wire u2_root_415__FF_INPUT;
  wire u2_root_416__FF_INPUT;
  wire u2_root_417__FF_INPUT;
  wire u2_root_418__FF_INPUT;
  wire u2_root_419__FF_INPUT;
  wire u2_root_41__FF_INPUT;
  wire u2_root_420__FF_INPUT;
  wire u2_root_421__FF_INPUT;
  wire u2_root_422__FF_INPUT;
  wire u2_root_423__FF_INPUT;
  wire u2_root_424__FF_INPUT;
  wire u2_root_425__FF_INPUT;
  wire u2_root_426__FF_INPUT;
  wire u2_root_427__FF_INPUT;
  wire u2_root_428__FF_INPUT;
  wire u2_root_429__FF_INPUT;
  wire u2_root_42__FF_INPUT;
  wire u2_root_430__FF_INPUT;
  wire u2_root_431__FF_INPUT;
  wire u2_root_432__FF_INPUT;
  wire u2_root_433__FF_INPUT;
  wire u2_root_434__FF_INPUT;
  wire u2_root_435__FF_INPUT;
  wire u2_root_436__FF_INPUT;
  wire u2_root_437__FF_INPUT;
  wire u2_root_438__FF_INPUT;
  wire u2_root_439__FF_INPUT;
  wire u2_root_43__FF_INPUT;
  wire u2_root_440__FF_INPUT;
  wire u2_root_441__FF_INPUT;
  wire u2_root_442__FF_INPUT;
  wire u2_root_443__FF_INPUT;
  wire u2_root_444__FF_INPUT;
  wire u2_root_445__FF_INPUT;
  wire u2_root_446__FF_INPUT;
  wire u2_root_447__FF_INPUT;
  wire u2_root_448__FF_INPUT;
  wire u2_root_449__FF_INPUT;
  wire u2_root_44__FF_INPUT;
  wire u2_root_450__FF_INPUT;
  wire u2_root_45__FF_INPUT;
  wire u2_root_46__FF_INPUT;
  wire u2_root_47__FF_INPUT;
  wire u2_root_48__FF_INPUT;
  wire u2_root_49__FF_INPUT;
  wire u2_root_4__FF_INPUT;
  wire u2_root_50__FF_INPUT;
  wire u2_root_51__FF_INPUT;
  wire u2_root_52__FF_INPUT;
  wire u2_root_53__FF_INPUT;
  wire u2_root_54__FF_INPUT;
  wire u2_root_55__FF_INPUT;
  wire u2_root_56__FF_INPUT;
  wire u2_root_57__FF_INPUT;
  wire u2_root_58__FF_INPUT;
  wire u2_root_59__FF_INPUT;
  wire u2_root_5__FF_INPUT;
  wire u2_root_60__FF_INPUT;
  wire u2_root_61__FF_INPUT;
  wire u2_root_62__FF_INPUT;
  wire u2_root_63__FF_INPUT;
  wire u2_root_64__FF_INPUT;
  wire u2_root_65__FF_INPUT;
  wire u2_root_66__FF_INPUT;
  wire u2_root_67__FF_INPUT;
  wire u2_root_68__FF_INPUT;
  wire u2_root_69__FF_INPUT;
  wire u2_root_6__FF_INPUT;
  wire u2_root_70__FF_INPUT;
  wire u2_root_71__FF_INPUT;
  wire u2_root_72__FF_INPUT;
  wire u2_root_73__FF_INPUT;
  wire u2_root_74__FF_INPUT;
  wire u2_root_75__FF_INPUT;
  wire u2_root_76__FF_INPUT;
  wire u2_root_77__FF_INPUT;
  wire u2_root_78__FF_INPUT;
  wire u2_root_79__FF_INPUT;
  wire u2_root_7__FF_INPUT;
  wire u2_root_80__FF_INPUT;
  wire u2_root_81__FF_INPUT;
  wire u2_root_82__FF_INPUT;
  wire u2_root_83__FF_INPUT;
  wire u2_root_84__FF_INPUT;
  wire u2_root_85__FF_INPUT;
  wire u2_root_86__FF_INPUT;
  wire u2_root_87__FF_INPUT;
  wire u2_root_88__FF_INPUT;
  wire u2_root_89__FF_INPUT;
  wire u2_root_8__FF_INPUT;
  wire u2_root_90__FF_INPUT;
  wire u2_root_91__FF_INPUT;
  wire u2_root_92__FF_INPUT;
  wire u2_root_93__FF_INPUT;
  wire u2_root_94__FF_INPUT;
  wire u2_root_95__FF_INPUT;
  wire u2_root_96__FF_INPUT;
  wire u2_root_97__FF_INPUT;
  wire u2_root_98__FF_INPUT;
  wire u2_root_99__FF_INPUT;
  wire u2_root_9__FF_INPUT;
  wire u2_state_0_;
  wire u2_state_2_;
  AND2X2 AND2X2_1 ( .A(_abc_64468_n753_bF_buf13), .B(sqrto_0_), .Y(_auto_iopadmap_cc_313_execute_65414_36_) );
  AND2X2 AND2X2_10 ( .A(_abc_64468_n753_bF_buf4), .B(sqrto_9_), .Y(_auto_iopadmap_cc_313_execute_65414_45_) );
  AND2X2 AND2X2_100 ( .A(_abc_64468_n900), .B(_abc_64468_n899), .Y(_auto_iopadmap_cc_313_execute_65414_135_) );
  AND2X2 AND2X2_1000 ( .A(u2__abc_44228_n4004), .B(u2__abc_44228_n3998), .Y(u2__abc_44228_n4005_1) );
  AND2X2 AND2X2_10000 ( .A(u2__abc_44228_n20168), .B(u2__abc_44228_n20171), .Y(u2__abc_44228_n20172) );
  AND2X2 AND2X2_10001 ( .A(u2__abc_44228_n20173), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_root_200__FF_INPUT) );
  AND2X2 AND2X2_10002 ( .A(u2__abc_44228_n3062_bF_buf92), .B(sqrto_200_), .Y(u2__abc_44228_n20175) );
  AND2X2 AND2X2_10003 ( .A(u2__abc_44228_n20165), .B(sqrto_199_), .Y(u2__abc_44228_n20177) );
  AND2X2 AND2X2_10004 ( .A(u2__abc_44228_n20178), .B(u2__abc_44228_n20176), .Y(u2__abc_44228_n20179) );
  AND2X2 AND2X2_10005 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n4695_1), .Y(u2__abc_44228_n20181) );
  AND2X2 AND2X2_10006 ( .A(u2__abc_44228_n20182), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n20183) );
  AND2X2 AND2X2_10007 ( .A(u2__abc_44228_n20180), .B(u2__abc_44228_n20183), .Y(u2__abc_44228_n20184) );
  AND2X2 AND2X2_10008 ( .A(u2__abc_44228_n20185), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_root_201__FF_INPUT) );
  AND2X2 AND2X2_10009 ( .A(u2__abc_44228_n3062_bF_buf91), .B(sqrto_201_), .Y(u2__abc_44228_n20187) );
  AND2X2 AND2X2_1001 ( .A(u2__abc_44228_n4006), .B(u2_remHi_78_), .Y(u2__abc_44228_n4007) );
  AND2X2 AND2X2_10010 ( .A(u2__abc_44228_n20177), .B(sqrto_200_), .Y(u2__abc_44228_n20189) );
  AND2X2 AND2X2_10011 ( .A(u2__abc_44228_n20190), .B(u2__abc_44228_n20188), .Y(u2__abc_44228_n20191) );
  AND2X2 AND2X2_10012 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n4688), .Y(u2__abc_44228_n20193) );
  AND2X2 AND2X2_10013 ( .A(u2__abc_44228_n20194), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n20195) );
  AND2X2 AND2X2_10014 ( .A(u2__abc_44228_n20192), .B(u2__abc_44228_n20195), .Y(u2__abc_44228_n20196) );
  AND2X2 AND2X2_10015 ( .A(u2__abc_44228_n20197), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_root_202__FF_INPUT) );
  AND2X2 AND2X2_10016 ( .A(u2__abc_44228_n3062_bF_buf90), .B(sqrto_202_), .Y(u2__abc_44228_n20199) );
  AND2X2 AND2X2_10017 ( .A(u2__abc_44228_n20189), .B(sqrto_201_), .Y(u2__abc_44228_n20201) );
  AND2X2 AND2X2_10018 ( .A(u2__abc_44228_n20202), .B(u2__abc_44228_n20200), .Y(u2__abc_44228_n20203) );
  AND2X2 AND2X2_10019 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n4680), .Y(u2__abc_44228_n20205) );
  AND2X2 AND2X2_1002 ( .A(u2__abc_44228_n4008), .B(sqrto_78_), .Y(u2__abc_44228_n4009) );
  AND2X2 AND2X2_10020 ( .A(u2__abc_44228_n20206), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n20207) );
  AND2X2 AND2X2_10021 ( .A(u2__abc_44228_n20204), .B(u2__abc_44228_n20207), .Y(u2__abc_44228_n20208) );
  AND2X2 AND2X2_10022 ( .A(u2__abc_44228_n20209), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_root_203__FF_INPUT) );
  AND2X2 AND2X2_10023 ( .A(u2__abc_44228_n3062_bF_buf89), .B(sqrto_203_), .Y(u2__abc_44228_n20211) );
  AND2X2 AND2X2_10024 ( .A(u2__abc_44228_n20201), .B(sqrto_202_), .Y(u2__abc_44228_n20213) );
  AND2X2 AND2X2_10025 ( .A(u2__abc_44228_n20214), .B(u2__abc_44228_n20212), .Y(u2__abc_44228_n20215) );
  AND2X2 AND2X2_10026 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n4673), .Y(u2__abc_44228_n20217) );
  AND2X2 AND2X2_10027 ( .A(u2__abc_44228_n20218), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n20219) );
  AND2X2 AND2X2_10028 ( .A(u2__abc_44228_n20216), .B(u2__abc_44228_n20219), .Y(u2__abc_44228_n20220) );
  AND2X2 AND2X2_10029 ( .A(u2__abc_44228_n20221), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_root_204__FF_INPUT) );
  AND2X2 AND2X2_1003 ( .A(u2__abc_44228_n4012), .B(u2_remHi_79_), .Y(u2__abc_44228_n4013) );
  AND2X2 AND2X2_10030 ( .A(u2__abc_44228_n3062_bF_buf88), .B(sqrto_204_), .Y(u2__abc_44228_n20223) );
  AND2X2 AND2X2_10031 ( .A(u2__abc_44228_n20213), .B(sqrto_203_), .Y(u2__abc_44228_n20225) );
  AND2X2 AND2X2_10032 ( .A(u2__abc_44228_n20226), .B(u2__abc_44228_n20224), .Y(u2__abc_44228_n20227) );
  AND2X2 AND2X2_10033 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n4666), .Y(u2__abc_44228_n20229) );
  AND2X2 AND2X2_10034 ( .A(u2__abc_44228_n20230), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n20231) );
  AND2X2 AND2X2_10035 ( .A(u2__abc_44228_n20228), .B(u2__abc_44228_n20231), .Y(u2__abc_44228_n20232) );
  AND2X2 AND2X2_10036 ( .A(u2__abc_44228_n20233), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_root_205__FF_INPUT) );
  AND2X2 AND2X2_10037 ( .A(u2__abc_44228_n3062_bF_buf87), .B(sqrto_205_), .Y(u2__abc_44228_n20235) );
  AND2X2 AND2X2_10038 ( .A(u2__abc_44228_n20225), .B(sqrto_204_), .Y(u2__abc_44228_n20237) );
  AND2X2 AND2X2_10039 ( .A(u2__abc_44228_n20238), .B(u2__abc_44228_n20236), .Y(u2__abc_44228_n20239) );
  AND2X2 AND2X2_1004 ( .A(u2__abc_44228_n4015_1), .B(sqrto_79_), .Y(u2__abc_44228_n4016) );
  AND2X2 AND2X2_10040 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n4659), .Y(u2__abc_44228_n20241) );
  AND2X2 AND2X2_10041 ( .A(u2__abc_44228_n20242), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n20243) );
  AND2X2 AND2X2_10042 ( .A(u2__abc_44228_n20240), .B(u2__abc_44228_n20243), .Y(u2__abc_44228_n20244) );
  AND2X2 AND2X2_10043 ( .A(u2__abc_44228_n20245), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_root_206__FF_INPUT) );
  AND2X2 AND2X2_10044 ( .A(u2__abc_44228_n3062_bF_buf86), .B(sqrto_206_), .Y(u2__abc_44228_n20247) );
  AND2X2 AND2X2_10045 ( .A(u2__abc_44228_n20237), .B(sqrto_205_), .Y(u2__abc_44228_n20249) );
  AND2X2 AND2X2_10046 ( .A(u2__abc_44228_n20250), .B(u2__abc_44228_n20248), .Y(u2__abc_44228_n20251) );
  AND2X2 AND2X2_10047 ( .A(u2__abc_44228_n2983_bF_buf62), .B(u2__abc_44228_n4649), .Y(u2__abc_44228_n20253) );
  AND2X2 AND2X2_10048 ( .A(u2__abc_44228_n20254), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n20255) );
  AND2X2 AND2X2_10049 ( .A(u2__abc_44228_n20252), .B(u2__abc_44228_n20255), .Y(u2__abc_44228_n20256) );
  AND2X2 AND2X2_1005 ( .A(u2__abc_44228_n4014), .B(u2__abc_44228_n4017), .Y(u2__abc_44228_n4018) );
  AND2X2 AND2X2_10050 ( .A(u2__abc_44228_n20257), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_root_207__FF_INPUT) );
  AND2X2 AND2X2_10051 ( .A(u2__abc_44228_n3062_bF_buf85), .B(sqrto_207_), .Y(u2__abc_44228_n20259) );
  AND2X2 AND2X2_10052 ( .A(u2__abc_44228_n20249), .B(sqrto_206_), .Y(u2__abc_44228_n20261) );
  AND2X2 AND2X2_10053 ( .A(u2__abc_44228_n20262), .B(u2__abc_44228_n20260), .Y(u2__abc_44228_n20263) );
  AND2X2 AND2X2_10054 ( .A(u2__abc_44228_n2983_bF_buf60), .B(u2__abc_44228_n4642), .Y(u2__abc_44228_n20265) );
  AND2X2 AND2X2_10055 ( .A(u2__abc_44228_n20266), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n20267) );
  AND2X2 AND2X2_10056 ( .A(u2__abc_44228_n20264), .B(u2__abc_44228_n20267), .Y(u2__abc_44228_n20268) );
  AND2X2 AND2X2_10057 ( .A(u2__abc_44228_n20269), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_root_208__FF_INPUT) );
  AND2X2 AND2X2_10058 ( .A(u2__abc_44228_n3062_bF_buf84), .B(sqrto_208_), .Y(u2__abc_44228_n20271) );
  AND2X2 AND2X2_10059 ( .A(u2__abc_44228_n20261), .B(sqrto_207_), .Y(u2__abc_44228_n20273) );
  AND2X2 AND2X2_1006 ( .A(u2__abc_44228_n4011), .B(u2__abc_44228_n4018), .Y(u2__abc_44228_n4019) );
  AND2X2 AND2X2_10060 ( .A(u2__abc_44228_n20274), .B(u2__abc_44228_n20272), .Y(u2__abc_44228_n20275) );
  AND2X2 AND2X2_10061 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n4635), .Y(u2__abc_44228_n20277) );
  AND2X2 AND2X2_10062 ( .A(u2__abc_44228_n20278), .B(u2__abc_44228_n2972_bF_buf87), .Y(u2__abc_44228_n20279) );
  AND2X2 AND2X2_10063 ( .A(u2__abc_44228_n20276), .B(u2__abc_44228_n20279), .Y(u2__abc_44228_n20280) );
  AND2X2 AND2X2_10064 ( .A(u2__abc_44228_n20281), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_root_209__FF_INPUT) );
  AND2X2 AND2X2_10065 ( .A(u2__abc_44228_n3062_bF_buf83), .B(sqrto_209_), .Y(u2__abc_44228_n20283) );
  AND2X2 AND2X2_10066 ( .A(u2__abc_44228_n20273), .B(sqrto_208_), .Y(u2__abc_44228_n20285) );
  AND2X2 AND2X2_10067 ( .A(u2__abc_44228_n20286), .B(u2__abc_44228_n20284), .Y(u2__abc_44228_n20287) );
  AND2X2 AND2X2_10068 ( .A(u2__abc_44228_n2983_bF_buf56), .B(u2__abc_44228_n4628), .Y(u2__abc_44228_n20289) );
  AND2X2 AND2X2_10069 ( .A(u2__abc_44228_n20290), .B(u2__abc_44228_n2972_bF_buf86), .Y(u2__abc_44228_n20291) );
  AND2X2 AND2X2_1007 ( .A(u2__abc_44228_n4005_1), .B(u2__abc_44228_n4019), .Y(u2__abc_44228_n4020) );
  AND2X2 AND2X2_10070 ( .A(u2__abc_44228_n20288), .B(u2__abc_44228_n20291), .Y(u2__abc_44228_n20292) );
  AND2X2 AND2X2_10071 ( .A(u2__abc_44228_n20293), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_root_210__FF_INPUT) );
  AND2X2 AND2X2_10072 ( .A(u2__abc_44228_n3062_bF_buf82), .B(sqrto_210_), .Y(u2__abc_44228_n20295) );
  AND2X2 AND2X2_10073 ( .A(u2__abc_44228_n20285), .B(sqrto_209_), .Y(u2__abc_44228_n20297) );
  AND2X2 AND2X2_10074 ( .A(u2__abc_44228_n20298), .B(u2__abc_44228_n20296), .Y(u2__abc_44228_n20299) );
  AND2X2 AND2X2_10075 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n4613), .Y(u2__abc_44228_n20301) );
  AND2X2 AND2X2_10076 ( .A(u2__abc_44228_n20302), .B(u2__abc_44228_n2972_bF_buf85), .Y(u2__abc_44228_n20303) );
  AND2X2 AND2X2_10077 ( .A(u2__abc_44228_n20300), .B(u2__abc_44228_n20303), .Y(u2__abc_44228_n20304) );
  AND2X2 AND2X2_10078 ( .A(u2__abc_44228_n20305), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_root_211__FF_INPUT) );
  AND2X2 AND2X2_10079 ( .A(u2__abc_44228_n3062_bF_buf81), .B(sqrto_211_), .Y(u2__abc_44228_n20307) );
  AND2X2 AND2X2_1008 ( .A(u2__abc_44228_n3991), .B(u2__abc_44228_n4020), .Y(u2__abc_44228_n4021) );
  AND2X2 AND2X2_10080 ( .A(u2__abc_44228_n20297), .B(sqrto_210_), .Y(u2__abc_44228_n20309) );
  AND2X2 AND2X2_10081 ( .A(u2__abc_44228_n20310), .B(u2__abc_44228_n20308), .Y(u2__abc_44228_n20311) );
  AND2X2 AND2X2_10082 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n4619), .Y(u2__abc_44228_n20313) );
  AND2X2 AND2X2_10083 ( .A(u2__abc_44228_n20314), .B(u2__abc_44228_n2972_bF_buf84), .Y(u2__abc_44228_n20315) );
  AND2X2 AND2X2_10084 ( .A(u2__abc_44228_n20312), .B(u2__abc_44228_n20315), .Y(u2__abc_44228_n20316) );
  AND2X2 AND2X2_10085 ( .A(u2__abc_44228_n20317), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_root_212__FF_INPUT) );
  AND2X2 AND2X2_10086 ( .A(u2__abc_44228_n3062_bF_buf80), .B(sqrto_212_), .Y(u2__abc_44228_n20319) );
  AND2X2 AND2X2_10087 ( .A(u2__abc_44228_n20309), .B(sqrto_211_), .Y(u2__abc_44228_n20321) );
  AND2X2 AND2X2_10088 ( .A(u2__abc_44228_n20322), .B(u2__abc_44228_n20320), .Y(u2__abc_44228_n20323) );
  AND2X2 AND2X2_10089 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2__abc_44228_n4606), .Y(u2__abc_44228_n20325) );
  AND2X2 AND2X2_1009 ( .A(u2__abc_44228_n3962), .B(u2__abc_44228_n4021), .Y(u2__abc_44228_n4022) );
  AND2X2 AND2X2_10090 ( .A(u2__abc_44228_n20326), .B(u2__abc_44228_n2972_bF_buf83), .Y(u2__abc_44228_n20327) );
  AND2X2 AND2X2_10091 ( .A(u2__abc_44228_n20324), .B(u2__abc_44228_n20327), .Y(u2__abc_44228_n20328) );
  AND2X2 AND2X2_10092 ( .A(u2__abc_44228_n20329), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_root_213__FF_INPUT) );
  AND2X2 AND2X2_10093 ( .A(u2__abc_44228_n3062_bF_buf79), .B(sqrto_213_), .Y(u2__abc_44228_n20331) );
  AND2X2 AND2X2_10094 ( .A(u2__abc_44228_n20321), .B(sqrto_212_), .Y(u2__abc_44228_n20333) );
  AND2X2 AND2X2_10095 ( .A(u2__abc_44228_n20334), .B(u2__abc_44228_n20332), .Y(u2__abc_44228_n20335) );
  AND2X2 AND2X2_10096 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n4599), .Y(u2__abc_44228_n20337) );
  AND2X2 AND2X2_10097 ( .A(u2__abc_44228_n20338), .B(u2__abc_44228_n2972_bF_buf82), .Y(u2__abc_44228_n20339) );
  AND2X2 AND2X2_10098 ( .A(u2__abc_44228_n20336), .B(u2__abc_44228_n20339), .Y(u2__abc_44228_n20340) );
  AND2X2 AND2X2_10099 ( .A(u2__abc_44228_n20341), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_root_214__FF_INPUT) );
  AND2X2 AND2X2_101 ( .A(_abc_64468_n903), .B(_abc_64468_n902), .Y(_auto_iopadmap_cc_313_execute_65414_136_) );
  AND2X2 AND2X2_1010 ( .A(u2__abc_44228_n4023), .B(u2_remHi_77_), .Y(u2__abc_44228_n4024_1) );
  AND2X2 AND2X2_10100 ( .A(u2__abc_44228_n3062_bF_buf78), .B(sqrto_214_), .Y(u2__abc_44228_n20343) );
  AND2X2 AND2X2_10101 ( .A(u2__abc_44228_n20333), .B(sqrto_213_), .Y(u2__abc_44228_n20345) );
  AND2X2 AND2X2_10102 ( .A(u2__abc_44228_n20346), .B(u2__abc_44228_n20344), .Y(u2__abc_44228_n20347) );
  AND2X2 AND2X2_10103 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n4583), .Y(u2__abc_44228_n20349) );
  AND2X2 AND2X2_10104 ( .A(u2__abc_44228_n20350), .B(u2__abc_44228_n2972_bF_buf81), .Y(u2__abc_44228_n20351) );
  AND2X2 AND2X2_10105 ( .A(u2__abc_44228_n20348), .B(u2__abc_44228_n20351), .Y(u2__abc_44228_n20352) );
  AND2X2 AND2X2_10106 ( .A(u2__abc_44228_n20353), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_root_215__FF_INPUT) );
  AND2X2 AND2X2_10107 ( .A(u2__abc_44228_n3062_bF_buf77), .B(sqrto_215_), .Y(u2__abc_44228_n20355) );
  AND2X2 AND2X2_10108 ( .A(u2__abc_44228_n20345), .B(sqrto_214_), .Y(u2__abc_44228_n20357) );
  AND2X2 AND2X2_10109 ( .A(u2__abc_44228_n20358), .B(u2__abc_44228_n20356), .Y(u2__abc_44228_n20359) );
  AND2X2 AND2X2_1011 ( .A(u2__abc_44228_n4026), .B(sqrto_77_), .Y(u2__abc_44228_n4027) );
  AND2X2 AND2X2_10110 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n4589), .Y(u2__abc_44228_n20361) );
  AND2X2 AND2X2_10111 ( .A(u2__abc_44228_n20362), .B(u2__abc_44228_n2972_bF_buf80), .Y(u2__abc_44228_n20363) );
  AND2X2 AND2X2_10112 ( .A(u2__abc_44228_n20360), .B(u2__abc_44228_n20363), .Y(u2__abc_44228_n20364) );
  AND2X2 AND2X2_10113 ( .A(u2__abc_44228_n20365), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_root_216__FF_INPUT) );
  AND2X2 AND2X2_10114 ( .A(u2__abc_44228_n3062_bF_buf76), .B(sqrto_216_), .Y(u2__abc_44228_n20367) );
  AND2X2 AND2X2_10115 ( .A(u2__abc_44228_n20357), .B(sqrto_215_), .Y(u2__abc_44228_n20369) );
  AND2X2 AND2X2_10116 ( .A(u2__abc_44228_n20370), .B(u2__abc_44228_n20368), .Y(u2__abc_44228_n20371) );
  AND2X2 AND2X2_10117 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n4576), .Y(u2__abc_44228_n20373) );
  AND2X2 AND2X2_10118 ( .A(u2__abc_44228_n20374), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n20375) );
  AND2X2 AND2X2_10119 ( .A(u2__abc_44228_n20372), .B(u2__abc_44228_n20375), .Y(u2__abc_44228_n20376) );
  AND2X2 AND2X2_1012 ( .A(u2__abc_44228_n4025), .B(u2__abc_44228_n4028), .Y(u2__abc_44228_n4029) );
  AND2X2 AND2X2_10120 ( .A(u2__abc_44228_n20377), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_root_217__FF_INPUT) );
  AND2X2 AND2X2_10121 ( .A(u2__abc_44228_n3062_bF_buf75), .B(sqrto_217_), .Y(u2__abc_44228_n20379) );
  AND2X2 AND2X2_10122 ( .A(u2__abc_44228_n20369), .B(sqrto_216_), .Y(u2__abc_44228_n20381) );
  AND2X2 AND2X2_10123 ( .A(u2__abc_44228_n20382), .B(u2__abc_44228_n20380), .Y(u2__abc_44228_n20383) );
  AND2X2 AND2X2_10124 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n4569), .Y(u2__abc_44228_n20385) );
  AND2X2 AND2X2_10125 ( .A(u2__abc_44228_n20386), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n20387) );
  AND2X2 AND2X2_10126 ( .A(u2__abc_44228_n20384), .B(u2__abc_44228_n20387), .Y(u2__abc_44228_n20388) );
  AND2X2 AND2X2_10127 ( .A(u2__abc_44228_n20389), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_root_218__FF_INPUT) );
  AND2X2 AND2X2_10128 ( .A(u2__abc_44228_n3062_bF_buf74), .B(sqrto_218_), .Y(u2__abc_44228_n20391) );
  AND2X2 AND2X2_10129 ( .A(u2__abc_44228_n20381), .B(sqrto_217_), .Y(u2__abc_44228_n20393) );
  AND2X2 AND2X2_1013 ( .A(u2__abc_44228_n4030), .B(u2_remHi_76_), .Y(u2__abc_44228_n4031) );
  AND2X2 AND2X2_10130 ( .A(u2__abc_44228_n20394), .B(u2__abc_44228_n20392), .Y(u2__abc_44228_n20395) );
  AND2X2 AND2X2_10131 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n4554_1), .Y(u2__abc_44228_n20397) );
  AND2X2 AND2X2_10132 ( .A(u2__abc_44228_n20398), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n20399) );
  AND2X2 AND2X2_10133 ( .A(u2__abc_44228_n20396), .B(u2__abc_44228_n20399), .Y(u2__abc_44228_n20400) );
  AND2X2 AND2X2_10134 ( .A(u2__abc_44228_n20401), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_root_219__FF_INPUT) );
  AND2X2 AND2X2_10135 ( .A(u2__abc_44228_n3062_bF_buf73), .B(sqrto_219_), .Y(u2__abc_44228_n20403) );
  AND2X2 AND2X2_10136 ( .A(u2__abc_44228_n20393), .B(sqrto_218_), .Y(u2__abc_44228_n20405) );
  AND2X2 AND2X2_10137 ( .A(u2__abc_44228_n20406), .B(u2__abc_44228_n20404), .Y(u2__abc_44228_n20407) );
  AND2X2 AND2X2_10138 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n4560), .Y(u2__abc_44228_n20409) );
  AND2X2 AND2X2_10139 ( .A(u2__abc_44228_n20410), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n20411) );
  AND2X2 AND2X2_1014 ( .A(u2__abc_44228_n4032), .B(sqrto_76_), .Y(u2__abc_44228_n4033_1) );
  AND2X2 AND2X2_10140 ( .A(u2__abc_44228_n20408), .B(u2__abc_44228_n20411), .Y(u2__abc_44228_n20412) );
  AND2X2 AND2X2_10141 ( .A(u2__abc_44228_n20413), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_root_220__FF_INPUT) );
  AND2X2 AND2X2_10142 ( .A(u2__abc_44228_n3062_bF_buf72), .B(sqrto_220_), .Y(u2__abc_44228_n20415) );
  AND2X2 AND2X2_10143 ( .A(u2__abc_44228_n20405), .B(sqrto_219_), .Y(u2__abc_44228_n20417) );
  AND2X2 AND2X2_10144 ( .A(u2__abc_44228_n20418), .B(u2__abc_44228_n20416), .Y(u2__abc_44228_n20419) );
  AND2X2 AND2X2_10145 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n4547), .Y(u2__abc_44228_n20421) );
  AND2X2 AND2X2_10146 ( .A(u2__abc_44228_n20422), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n20423) );
  AND2X2 AND2X2_10147 ( .A(u2__abc_44228_n20420), .B(u2__abc_44228_n20423), .Y(u2__abc_44228_n20424) );
  AND2X2 AND2X2_10148 ( .A(u2__abc_44228_n20425), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_root_221__FF_INPUT) );
  AND2X2 AND2X2_10149 ( .A(u2__abc_44228_n3062_bF_buf71), .B(sqrto_221_), .Y(u2__abc_44228_n20427) );
  AND2X2 AND2X2_1015 ( .A(u2__abc_44228_n4035), .B(u2__abc_44228_n4029), .Y(u2__abc_44228_n4036) );
  AND2X2 AND2X2_10150 ( .A(u2__abc_44228_n20417), .B(sqrto_220_), .Y(u2__abc_44228_n20429) );
  AND2X2 AND2X2_10151 ( .A(u2__abc_44228_n20430), .B(u2__abc_44228_n20428), .Y(u2__abc_44228_n20431) );
  AND2X2 AND2X2_10152 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n4540), .Y(u2__abc_44228_n20433) );
  AND2X2 AND2X2_10153 ( .A(u2__abc_44228_n20434), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n20435) );
  AND2X2 AND2X2_10154 ( .A(u2__abc_44228_n20432), .B(u2__abc_44228_n20435), .Y(u2__abc_44228_n20436) );
  AND2X2 AND2X2_10155 ( .A(u2__abc_44228_n20437), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_root_222__FF_INPUT) );
  AND2X2 AND2X2_10156 ( .A(u2__abc_44228_n3062_bF_buf70), .B(sqrto_222_), .Y(u2__abc_44228_n20439) );
  AND2X2 AND2X2_10157 ( .A(u2__abc_44228_n20429), .B(sqrto_221_), .Y(u2__abc_44228_n20441) );
  AND2X2 AND2X2_10158 ( .A(u2__abc_44228_n20442), .B(u2__abc_44228_n20440), .Y(u2__abc_44228_n20443) );
  AND2X2 AND2X2_10159 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n4522), .Y(u2__abc_44228_n20445) );
  AND2X2 AND2X2_1016 ( .A(u2__abc_44228_n4037), .B(u2_remHi_74_), .Y(u2__abc_44228_n4038) );
  AND2X2 AND2X2_10160 ( .A(u2__abc_44228_n20446), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n20447) );
  AND2X2 AND2X2_10161 ( .A(u2__abc_44228_n20444), .B(u2__abc_44228_n20447), .Y(u2__abc_44228_n20448) );
  AND2X2 AND2X2_10162 ( .A(u2__abc_44228_n20449), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_root_223__FF_INPUT) );
  AND2X2 AND2X2_10163 ( .A(u2__abc_44228_n3062_bF_buf69), .B(sqrto_223_), .Y(u2__abc_44228_n20451) );
  AND2X2 AND2X2_10164 ( .A(u2__abc_44228_n20441), .B(sqrto_222_), .Y(u2__abc_44228_n20453) );
  AND2X2 AND2X2_10165 ( .A(u2__abc_44228_n20454), .B(u2__abc_44228_n20452), .Y(u2__abc_44228_n20455) );
  AND2X2 AND2X2_10166 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n4528), .Y(u2__abc_44228_n20457) );
  AND2X2 AND2X2_10167 ( .A(u2__abc_44228_n20458), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n20459) );
  AND2X2 AND2X2_10168 ( .A(u2__abc_44228_n20456), .B(u2__abc_44228_n20459), .Y(u2__abc_44228_n20460) );
  AND2X2 AND2X2_10169 ( .A(u2__abc_44228_n20461), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_root_224__FF_INPUT) );
  AND2X2 AND2X2_1017 ( .A(u2__abc_44228_n4039), .B(sqrto_74_), .Y(u2__abc_44228_n4040) );
  AND2X2 AND2X2_10170 ( .A(u2__abc_44228_n3062_bF_buf68), .B(sqrto_224_), .Y(u2__abc_44228_n20463) );
  AND2X2 AND2X2_10171 ( .A(u2__abc_44228_n20453), .B(sqrto_223_), .Y(u2__abc_44228_n20465) );
  AND2X2 AND2X2_10172 ( .A(u2__abc_44228_n20466), .B(u2__abc_44228_n20464), .Y(u2__abc_44228_n20467) );
  AND2X2 AND2X2_10173 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n4515), .Y(u2__abc_44228_n20469) );
  AND2X2 AND2X2_10174 ( .A(u2__abc_44228_n20470), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n20471) );
  AND2X2 AND2X2_10175 ( .A(u2__abc_44228_n20468), .B(u2__abc_44228_n20471), .Y(u2__abc_44228_n20472) );
  AND2X2 AND2X2_10176 ( .A(u2__abc_44228_n20473), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_root_225__FF_INPUT) );
  AND2X2 AND2X2_10177 ( .A(u2__abc_44228_n3062_bF_buf67), .B(sqrto_225_), .Y(u2__abc_44228_n20475) );
  AND2X2 AND2X2_10178 ( .A(u2__abc_44228_n20465), .B(sqrto_224_), .Y(u2__abc_44228_n20477) );
  AND2X2 AND2X2_10179 ( .A(u2__abc_44228_n20478), .B(u2__abc_44228_n20476), .Y(u2__abc_44228_n20479) );
  AND2X2 AND2X2_1018 ( .A(u2__abc_44228_n4043), .B(u2_remHi_75_), .Y(u2__abc_44228_n4044) );
  AND2X2 AND2X2_10180 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n4508_1), .Y(u2__abc_44228_n20481) );
  AND2X2 AND2X2_10181 ( .A(u2__abc_44228_n20482), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n20483) );
  AND2X2 AND2X2_10182 ( .A(u2__abc_44228_n20480), .B(u2__abc_44228_n20483), .Y(u2__abc_44228_n20484) );
  AND2X2 AND2X2_10183 ( .A(u2__abc_44228_n20485), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_root_226__FF_INPUT) );
  AND2X2 AND2X2_10184 ( .A(u2__abc_44228_n3062_bF_buf66), .B(u2_o_226_), .Y(u2__abc_44228_n20487) );
  AND2X2 AND2X2_10185 ( .A(u2__abc_44228_n20477), .B(sqrto_225_), .Y(u2__abc_44228_n20489) );
  AND2X2 AND2X2_10186 ( .A(u2__abc_44228_n20490), .B(u2__abc_44228_n20488), .Y(u2__abc_44228_n20491) );
  AND2X2 AND2X2_10187 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n4493), .Y(u2__abc_44228_n20493) );
  AND2X2 AND2X2_10188 ( .A(u2__abc_44228_n20494), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n20495) );
  AND2X2 AND2X2_10189 ( .A(u2__abc_44228_n20492), .B(u2__abc_44228_n20495), .Y(u2__abc_44228_n20496) );
  AND2X2 AND2X2_1019 ( .A(u2__abc_44228_n4046), .B(sqrto_75_), .Y(u2__abc_44228_n4047) );
  AND2X2 AND2X2_10190 ( .A(u2__abc_44228_n20497), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_root_227__FF_INPUT) );
  AND2X2 AND2X2_10191 ( .A(u2__abc_44228_n3062_bF_buf65), .B(u2_o_227_), .Y(u2__abc_44228_n20499) );
  AND2X2 AND2X2_10192 ( .A(u2__abc_44228_n20489), .B(u2_o_226_), .Y(u2__abc_44228_n20501) );
  AND2X2 AND2X2_10193 ( .A(u2__abc_44228_n20502), .B(u2__abc_44228_n20500), .Y(u2__abc_44228_n20503) );
  AND2X2 AND2X2_10194 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n4499), .Y(u2__abc_44228_n20505) );
  AND2X2 AND2X2_10195 ( .A(u2__abc_44228_n20506), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n20507) );
  AND2X2 AND2X2_10196 ( .A(u2__abc_44228_n20504), .B(u2__abc_44228_n20507), .Y(u2__abc_44228_n20508) );
  AND2X2 AND2X2_10197 ( .A(u2__abc_44228_n20509), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_root_228__FF_INPUT) );
  AND2X2 AND2X2_10198 ( .A(u2__abc_44228_n3062_bF_buf64), .B(u2_o_228_), .Y(u2__abc_44228_n20511) );
  AND2X2 AND2X2_10199 ( .A(u2__abc_44228_n20501), .B(u2_o_227_), .Y(u2__abc_44228_n20513) );
  AND2X2 AND2X2_102 ( .A(_abc_64468_n906), .B(_abc_64468_n905), .Y(_auto_iopadmap_cc_313_execute_65414_137_) );
  AND2X2 AND2X2_1020 ( .A(u2__abc_44228_n4045), .B(u2__abc_44228_n4048), .Y(u2__abc_44228_n4049) );
  AND2X2 AND2X2_10200 ( .A(u2__abc_44228_n20514), .B(u2__abc_44228_n20512), .Y(u2__abc_44228_n20515) );
  AND2X2 AND2X2_10201 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n4486), .Y(u2__abc_44228_n20517) );
  AND2X2 AND2X2_10202 ( .A(u2__abc_44228_n20518), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n20519) );
  AND2X2 AND2X2_10203 ( .A(u2__abc_44228_n20516), .B(u2__abc_44228_n20519), .Y(u2__abc_44228_n20520) );
  AND2X2 AND2X2_10204 ( .A(u2__abc_44228_n20521), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_root_229__FF_INPUT) );
  AND2X2 AND2X2_10205 ( .A(u2__abc_44228_n3062_bF_buf63), .B(u2_o_229_), .Y(u2__abc_44228_n20523) );
  AND2X2 AND2X2_10206 ( .A(u2__abc_44228_n20513), .B(u2_o_228_), .Y(u2__abc_44228_n20525) );
  AND2X2 AND2X2_10207 ( .A(u2__abc_44228_n20526), .B(u2__abc_44228_n20524), .Y(u2__abc_44228_n20527) );
  AND2X2 AND2X2_10208 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n4479), .Y(u2__abc_44228_n20529) );
  AND2X2 AND2X2_10209 ( .A(u2__abc_44228_n20530), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n20531) );
  AND2X2 AND2X2_1021 ( .A(u2__abc_44228_n4042), .B(u2__abc_44228_n4049), .Y(u2__abc_44228_n4050_1) );
  AND2X2 AND2X2_10210 ( .A(u2__abc_44228_n20528), .B(u2__abc_44228_n20531), .Y(u2__abc_44228_n20532) );
  AND2X2 AND2X2_10211 ( .A(u2__abc_44228_n20533), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_root_230__FF_INPUT) );
  AND2X2 AND2X2_10212 ( .A(u2__abc_44228_n3062_bF_buf62), .B(u2_o_230_), .Y(u2__abc_44228_n20535) );
  AND2X2 AND2X2_10213 ( .A(u2__abc_44228_n20525), .B(u2_o_229_), .Y(u2__abc_44228_n20537) );
  AND2X2 AND2X2_10214 ( .A(u2__abc_44228_n20538), .B(u2__abc_44228_n20536), .Y(u2__abc_44228_n20539) );
  AND2X2 AND2X2_10215 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n4456), .Y(u2__abc_44228_n20541) );
  AND2X2 AND2X2_10216 ( .A(u2__abc_44228_n20542), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n20543) );
  AND2X2 AND2X2_10217 ( .A(u2__abc_44228_n20540), .B(u2__abc_44228_n20543), .Y(u2__abc_44228_n20544) );
  AND2X2 AND2X2_10218 ( .A(u2__abc_44228_n20545), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_root_231__FF_INPUT) );
  AND2X2 AND2X2_10219 ( .A(u2__abc_44228_n3062_bF_buf61), .B(u2_o_231_), .Y(u2__abc_44228_n20547) );
  AND2X2 AND2X2_1022 ( .A(u2__abc_44228_n4036), .B(u2__abc_44228_n4050_1), .Y(u2__abc_44228_n4051) );
  AND2X2 AND2X2_10220 ( .A(u2__abc_44228_n20537), .B(u2_o_230_), .Y(u2__abc_44228_n20549) );
  AND2X2 AND2X2_10221 ( .A(u2__abc_44228_n20550), .B(u2__abc_44228_n20548), .Y(u2__abc_44228_n20551) );
  AND2X2 AND2X2_10222 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n4449), .Y(u2__abc_44228_n20553) );
  AND2X2 AND2X2_10223 ( .A(u2__abc_44228_n20554), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n20555) );
  AND2X2 AND2X2_10224 ( .A(u2__abc_44228_n20552), .B(u2__abc_44228_n20555), .Y(u2__abc_44228_n20556) );
  AND2X2 AND2X2_10225 ( .A(u2__abc_44228_n20557), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_root_232__FF_INPUT) );
  AND2X2 AND2X2_10226 ( .A(u2__abc_44228_n3062_bF_buf60), .B(u2_o_232_), .Y(u2__abc_44228_n20559) );
  AND2X2 AND2X2_10227 ( .A(u2__abc_44228_n20549), .B(u2_o_231_), .Y(u2__abc_44228_n20561) );
  AND2X2 AND2X2_10228 ( .A(u2__abc_44228_n20562), .B(u2__abc_44228_n20560), .Y(u2__abc_44228_n20563) );
  AND2X2 AND2X2_10229 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n4470), .Y(u2__abc_44228_n20565) );
  AND2X2 AND2X2_1023 ( .A(u2__abc_44228_n4052), .B(u2_remHi_71_), .Y(u2__abc_44228_n4053) );
  AND2X2 AND2X2_10230 ( .A(u2__abc_44228_n20566), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n20567) );
  AND2X2 AND2X2_10231 ( .A(u2__abc_44228_n20564), .B(u2__abc_44228_n20567), .Y(u2__abc_44228_n20568) );
  AND2X2 AND2X2_10232 ( .A(u2__abc_44228_n20569), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_root_233__FF_INPUT) );
  AND2X2 AND2X2_10233 ( .A(u2__abc_44228_n3062_bF_buf59), .B(u2_o_233_), .Y(u2__abc_44228_n20571) );
  AND2X2 AND2X2_10234 ( .A(u2__abc_44228_n20561), .B(u2_o_232_), .Y(u2__abc_44228_n20573) );
  AND2X2 AND2X2_10235 ( .A(u2__abc_44228_n20574), .B(u2__abc_44228_n20572), .Y(u2__abc_44228_n20575) );
  AND2X2 AND2X2_10236 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n4463), .Y(u2__abc_44228_n20577) );
  AND2X2 AND2X2_10237 ( .A(u2__abc_44228_n20578), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n20579) );
  AND2X2 AND2X2_10238 ( .A(u2__abc_44228_n20576), .B(u2__abc_44228_n20579), .Y(u2__abc_44228_n20580) );
  AND2X2 AND2X2_10239 ( .A(u2__abc_44228_n20581), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_root_234__FF_INPUT) );
  AND2X2 AND2X2_1024 ( .A(u2__abc_44228_n4055), .B(sqrto_71_), .Y(u2__abc_44228_n4056) );
  AND2X2 AND2X2_10240 ( .A(u2__abc_44228_n3062_bF_buf58), .B(u2_o_234_), .Y(u2__abc_44228_n20583) );
  AND2X2 AND2X2_10241 ( .A(u2__abc_44228_n20573), .B(u2_o_233_), .Y(u2__abc_44228_n20585) );
  AND2X2 AND2X2_10242 ( .A(u2__abc_44228_n20586), .B(u2__abc_44228_n20584), .Y(u2__abc_44228_n20587) );
  AND2X2 AND2X2_10243 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n4434), .Y(u2__abc_44228_n20589) );
  AND2X2 AND2X2_10244 ( .A(u2__abc_44228_n20590), .B(u2__abc_44228_n2972_bF_buf61), .Y(u2__abc_44228_n20591) );
  AND2X2 AND2X2_10245 ( .A(u2__abc_44228_n20588), .B(u2__abc_44228_n20591), .Y(u2__abc_44228_n20592) );
  AND2X2 AND2X2_10246 ( .A(u2__abc_44228_n20593), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_root_235__FF_INPUT) );
  AND2X2 AND2X2_10247 ( .A(u2__abc_44228_n3062_bF_buf57), .B(u2_o_235_), .Y(u2__abc_44228_n20595) );
  AND2X2 AND2X2_10248 ( .A(u2__abc_44228_n20585), .B(u2_o_234_), .Y(u2__abc_44228_n20597) );
  AND2X2 AND2X2_10249 ( .A(u2__abc_44228_n20598), .B(u2__abc_44228_n20596), .Y(u2__abc_44228_n20599) );
  AND2X2 AND2X2_1025 ( .A(u2__abc_44228_n4054), .B(u2__abc_44228_n4057), .Y(u2__abc_44228_n4058) );
  AND2X2 AND2X2_10250 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n4440), .Y(u2__abc_44228_n20601) );
  AND2X2 AND2X2_10251 ( .A(u2__abc_44228_n20602), .B(u2__abc_44228_n2972_bF_buf60), .Y(u2__abc_44228_n20603) );
  AND2X2 AND2X2_10252 ( .A(u2__abc_44228_n20600), .B(u2__abc_44228_n20603), .Y(u2__abc_44228_n20604) );
  AND2X2 AND2X2_10253 ( .A(u2__abc_44228_n20605), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_root_236__FF_INPUT) );
  AND2X2 AND2X2_10254 ( .A(u2__abc_44228_n3062_bF_buf56), .B(u2_o_236_), .Y(u2__abc_44228_n20607) );
  AND2X2 AND2X2_10255 ( .A(u2__abc_44228_n20597), .B(u2_o_235_), .Y(u2__abc_44228_n20609) );
  AND2X2 AND2X2_10256 ( .A(u2__abc_44228_n20610), .B(u2__abc_44228_n20608), .Y(u2__abc_44228_n20611) );
  AND2X2 AND2X2_10257 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n4427), .Y(u2__abc_44228_n20613) );
  AND2X2 AND2X2_10258 ( .A(u2__abc_44228_n20614), .B(u2__abc_44228_n2972_bF_buf59), .Y(u2__abc_44228_n20615) );
  AND2X2 AND2X2_10259 ( .A(u2__abc_44228_n20612), .B(u2__abc_44228_n20615), .Y(u2__abc_44228_n20616) );
  AND2X2 AND2X2_1026 ( .A(u2__abc_44228_n4059), .B(u2_remHi_70_), .Y(u2__abc_44228_n4060) );
  AND2X2 AND2X2_10260 ( .A(u2__abc_44228_n20617), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_root_237__FF_INPUT) );
  AND2X2 AND2X2_10261 ( .A(u2__abc_44228_n3062_bF_buf55), .B(u2_o_237_), .Y(u2__abc_44228_n20619) );
  AND2X2 AND2X2_10262 ( .A(u2__abc_44228_n20609), .B(u2_o_236_), .Y(u2__abc_44228_n20621) );
  AND2X2 AND2X2_10263 ( .A(u2__abc_44228_n20622), .B(u2__abc_44228_n20620), .Y(u2__abc_44228_n20623) );
  AND2X2 AND2X2_10264 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n4420), .Y(u2__abc_44228_n20625) );
  AND2X2 AND2X2_10265 ( .A(u2__abc_44228_n20626), .B(u2__abc_44228_n2972_bF_buf58), .Y(u2__abc_44228_n20627) );
  AND2X2 AND2X2_10266 ( .A(u2__abc_44228_n20624), .B(u2__abc_44228_n20627), .Y(u2__abc_44228_n20628) );
  AND2X2 AND2X2_10267 ( .A(u2__abc_44228_n20629), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_root_238__FF_INPUT) );
  AND2X2 AND2X2_10268 ( .A(u2__abc_44228_n3062_bF_buf54), .B(u2_o_238_), .Y(u2__abc_44228_n20631) );
  AND2X2 AND2X2_10269 ( .A(u2__abc_44228_n20621), .B(u2_o_237_), .Y(u2__abc_44228_n20633) );
  AND2X2 AND2X2_1027 ( .A(u2__abc_44228_n4061_1), .B(sqrto_70_), .Y(u2__abc_44228_n4062) );
  AND2X2 AND2X2_10270 ( .A(u2__abc_44228_n20634), .B(u2__abc_44228_n20632), .Y(u2__abc_44228_n20635) );
  AND2X2 AND2X2_10271 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n4403), .Y(u2__abc_44228_n20637) );
  AND2X2 AND2X2_10272 ( .A(u2__abc_44228_n20638), .B(u2__abc_44228_n2972_bF_buf57), .Y(u2__abc_44228_n20639) );
  AND2X2 AND2X2_10273 ( .A(u2__abc_44228_n20636), .B(u2__abc_44228_n20639), .Y(u2__abc_44228_n20640) );
  AND2X2 AND2X2_10274 ( .A(u2__abc_44228_n20641), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_root_239__FF_INPUT) );
  AND2X2 AND2X2_10275 ( .A(u2__abc_44228_n3062_bF_buf53), .B(u2_o_239_), .Y(u2__abc_44228_n20643) );
  AND2X2 AND2X2_10276 ( .A(u2__abc_44228_n20633), .B(u2_o_238_), .Y(u2__abc_44228_n20645) );
  AND2X2 AND2X2_10277 ( .A(u2__abc_44228_n20646), .B(u2__abc_44228_n20644), .Y(u2__abc_44228_n20647) );
  AND2X2 AND2X2_10278 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n4409), .Y(u2__abc_44228_n20649) );
  AND2X2 AND2X2_10279 ( .A(u2__abc_44228_n20650), .B(u2__abc_44228_n2972_bF_buf56), .Y(u2__abc_44228_n20651) );
  AND2X2 AND2X2_1028 ( .A(u2__abc_44228_n4064), .B(u2__abc_44228_n4058), .Y(u2__abc_44228_n4065) );
  AND2X2 AND2X2_10280 ( .A(u2__abc_44228_n20648), .B(u2__abc_44228_n20651), .Y(u2__abc_44228_n20652) );
  AND2X2 AND2X2_10281 ( .A(u2__abc_44228_n20653), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_root_240__FF_INPUT) );
  AND2X2 AND2X2_10282 ( .A(u2__abc_44228_n3062_bF_buf52), .B(u2_o_240_), .Y(u2__abc_44228_n20655) );
  AND2X2 AND2X2_10283 ( .A(u2__abc_44228_n20645), .B(u2_o_239_), .Y(u2__abc_44228_n20657) );
  AND2X2 AND2X2_10284 ( .A(u2__abc_44228_n20658), .B(u2__abc_44228_n20656), .Y(u2__abc_44228_n20659) );
  AND2X2 AND2X2_10285 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n4396_1), .Y(u2__abc_44228_n20661) );
  AND2X2 AND2X2_10286 ( .A(u2__abc_44228_n20662), .B(u2__abc_44228_n2972_bF_buf55), .Y(u2__abc_44228_n20663) );
  AND2X2 AND2X2_10287 ( .A(u2__abc_44228_n20660), .B(u2__abc_44228_n20663), .Y(u2__abc_44228_n20664) );
  AND2X2 AND2X2_10288 ( .A(u2__abc_44228_n20665), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_root_241__FF_INPUT) );
  AND2X2 AND2X2_10289 ( .A(u2__abc_44228_n3062_bF_buf51), .B(u2_o_241_), .Y(u2__abc_44228_n20667) );
  AND2X2 AND2X2_1029 ( .A(u2__abc_44228_n4066), .B(u2_remHi_73_), .Y(u2__abc_44228_n4067) );
  AND2X2 AND2X2_10290 ( .A(u2__abc_44228_n20657), .B(u2_o_240_), .Y(u2__abc_44228_n20669) );
  AND2X2 AND2X2_10291 ( .A(u2__abc_44228_n20670), .B(u2__abc_44228_n20668), .Y(u2__abc_44228_n20671) );
  AND2X2 AND2X2_10292 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n4389), .Y(u2__abc_44228_n20673) );
  AND2X2 AND2X2_10293 ( .A(u2__abc_44228_n20674), .B(u2__abc_44228_n2972_bF_buf54), .Y(u2__abc_44228_n20675) );
  AND2X2 AND2X2_10294 ( .A(u2__abc_44228_n20672), .B(u2__abc_44228_n20675), .Y(u2__abc_44228_n20676) );
  AND2X2 AND2X2_10295 ( .A(u2__abc_44228_n20677), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_root_242__FF_INPUT) );
  AND2X2 AND2X2_10296 ( .A(u2__abc_44228_n3062_bF_buf50), .B(u2_o_242_), .Y(u2__abc_44228_n20679) );
  AND2X2 AND2X2_10297 ( .A(u2__abc_44228_n20669), .B(u2_o_241_), .Y(u2__abc_44228_n20681) );
  AND2X2 AND2X2_10298 ( .A(u2__abc_44228_n20682), .B(u2__abc_44228_n20680), .Y(u2__abc_44228_n20683) );
  AND2X2 AND2X2_10299 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n4374), .Y(u2__abc_44228_n20685) );
  AND2X2 AND2X2_103 ( .A(_abc_64468_n909), .B(_abc_64468_n908), .Y(_auto_iopadmap_cc_313_execute_65414_138_) );
  AND2X2 AND2X2_1030 ( .A(u2__abc_44228_n4069), .B(sqrto_73_), .Y(u2__abc_44228_n4070_1) );
  AND2X2 AND2X2_10300 ( .A(u2__abc_44228_n20686), .B(u2__abc_44228_n2972_bF_buf53), .Y(u2__abc_44228_n20687) );
  AND2X2 AND2X2_10301 ( .A(u2__abc_44228_n20684), .B(u2__abc_44228_n20687), .Y(u2__abc_44228_n20688) );
  AND2X2 AND2X2_10302 ( .A(u2__abc_44228_n20689), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_root_243__FF_INPUT) );
  AND2X2 AND2X2_10303 ( .A(u2__abc_44228_n3062_bF_buf49), .B(u2_o_243_), .Y(u2__abc_44228_n20691) );
  AND2X2 AND2X2_10304 ( .A(u2__abc_44228_n20681), .B(u2_o_242_), .Y(u2__abc_44228_n20693) );
  AND2X2 AND2X2_10305 ( .A(u2__abc_44228_n20694), .B(u2__abc_44228_n20692), .Y(u2__abc_44228_n20695) );
  AND2X2 AND2X2_10306 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n4380), .Y(u2__abc_44228_n20697) );
  AND2X2 AND2X2_10307 ( .A(u2__abc_44228_n20698), .B(u2__abc_44228_n2972_bF_buf52), .Y(u2__abc_44228_n20699) );
  AND2X2 AND2X2_10308 ( .A(u2__abc_44228_n20696), .B(u2__abc_44228_n20699), .Y(u2__abc_44228_n20700) );
  AND2X2 AND2X2_10309 ( .A(u2__abc_44228_n20701), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_root_244__FF_INPUT) );
  AND2X2 AND2X2_1031 ( .A(u2__abc_44228_n4068), .B(u2__abc_44228_n4071), .Y(u2__abc_44228_n4072) );
  AND2X2 AND2X2_10310 ( .A(u2__abc_44228_n3062_bF_buf48), .B(u2_o_244_), .Y(u2__abc_44228_n20703) );
  AND2X2 AND2X2_10311 ( .A(u2__abc_44228_n20693), .B(u2_o_243_), .Y(u2__abc_44228_n20705) );
  AND2X2 AND2X2_10312 ( .A(u2__abc_44228_n20706), .B(u2__abc_44228_n20704), .Y(u2__abc_44228_n20707) );
  AND2X2 AND2X2_10313 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n4367), .Y(u2__abc_44228_n20709) );
  AND2X2 AND2X2_10314 ( .A(u2__abc_44228_n20710), .B(u2__abc_44228_n2972_bF_buf51), .Y(u2__abc_44228_n20711) );
  AND2X2 AND2X2_10315 ( .A(u2__abc_44228_n20708), .B(u2__abc_44228_n20711), .Y(u2__abc_44228_n20712) );
  AND2X2 AND2X2_10316 ( .A(u2__abc_44228_n20713), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_root_245__FF_INPUT) );
  AND2X2 AND2X2_10317 ( .A(u2__abc_44228_n3062_bF_buf47), .B(u2_o_245_), .Y(u2__abc_44228_n20715) );
  AND2X2 AND2X2_10318 ( .A(u2__abc_44228_n20705), .B(u2_o_244_), .Y(u2__abc_44228_n20717) );
  AND2X2 AND2X2_10319 ( .A(u2__abc_44228_n20718), .B(u2__abc_44228_n20716), .Y(u2__abc_44228_n20719) );
  AND2X2 AND2X2_1032 ( .A(u2__abc_44228_n4073), .B(u2_remHi_72_), .Y(u2__abc_44228_n4074) );
  AND2X2 AND2X2_10320 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n4360), .Y(u2__abc_44228_n20721) );
  AND2X2 AND2X2_10321 ( .A(u2__abc_44228_n20722), .B(u2__abc_44228_n2972_bF_buf50), .Y(u2__abc_44228_n20723) );
  AND2X2 AND2X2_10322 ( .A(u2__abc_44228_n20720), .B(u2__abc_44228_n20723), .Y(u2__abc_44228_n20724) );
  AND2X2 AND2X2_10323 ( .A(u2__abc_44228_n20725), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_root_246__FF_INPUT) );
  AND2X2 AND2X2_10324 ( .A(u2__abc_44228_n3062_bF_buf46), .B(u2_o_246_), .Y(u2__abc_44228_n20727) );
  AND2X2 AND2X2_10325 ( .A(u2__abc_44228_n20717), .B(u2_o_245_), .Y(u2__abc_44228_n20729) );
  AND2X2 AND2X2_10326 ( .A(u2__abc_44228_n20730), .B(u2__abc_44228_n20728), .Y(u2__abc_44228_n20731) );
  AND2X2 AND2X2_10327 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n4344), .Y(u2__abc_44228_n20733) );
  AND2X2 AND2X2_10328 ( .A(u2__abc_44228_n20734), .B(u2__abc_44228_n2972_bF_buf49), .Y(u2__abc_44228_n20735) );
  AND2X2 AND2X2_10329 ( .A(u2__abc_44228_n20732), .B(u2__abc_44228_n20735), .Y(u2__abc_44228_n20736) );
  AND2X2 AND2X2_1033 ( .A(u2__abc_44228_n4075), .B(sqrto_72_), .Y(u2__abc_44228_n4076) );
  AND2X2 AND2X2_10330 ( .A(u2__abc_44228_n20737), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_root_247__FF_INPUT) );
  AND2X2 AND2X2_10331 ( .A(u2__abc_44228_n3062_bF_buf45), .B(u2_o_247_), .Y(u2__abc_44228_n20739) );
  AND2X2 AND2X2_10332 ( .A(u2__abc_44228_n20729), .B(u2_o_246_), .Y(u2__abc_44228_n20741) );
  AND2X2 AND2X2_10333 ( .A(u2__abc_44228_n20742), .B(u2__abc_44228_n20740), .Y(u2__abc_44228_n20743) );
  AND2X2 AND2X2_10334 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n4350), .Y(u2__abc_44228_n20745) );
  AND2X2 AND2X2_10335 ( .A(u2__abc_44228_n20746), .B(u2__abc_44228_n2972_bF_buf48), .Y(u2__abc_44228_n20747) );
  AND2X2 AND2X2_10336 ( .A(u2__abc_44228_n20744), .B(u2__abc_44228_n20747), .Y(u2__abc_44228_n20748) );
  AND2X2 AND2X2_10337 ( .A(u2__abc_44228_n20749), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_root_248__FF_INPUT) );
  AND2X2 AND2X2_10338 ( .A(u2__abc_44228_n3062_bF_buf44), .B(u2_o_248_), .Y(u2__abc_44228_n20751) );
  AND2X2 AND2X2_10339 ( .A(u2__abc_44228_n20741), .B(u2_o_247_), .Y(u2__abc_44228_n20753) );
  AND2X2 AND2X2_1034 ( .A(u2__abc_44228_n4078), .B(u2__abc_44228_n4072), .Y(u2__abc_44228_n4079) );
  AND2X2 AND2X2_10340 ( .A(u2__abc_44228_n20754), .B(u2__abc_44228_n20752), .Y(u2__abc_44228_n20755) );
  AND2X2 AND2X2_10341 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n4337), .Y(u2__abc_44228_n20757) );
  AND2X2 AND2X2_10342 ( .A(u2__abc_44228_n20758), .B(u2__abc_44228_n2972_bF_buf47), .Y(u2__abc_44228_n20759) );
  AND2X2 AND2X2_10343 ( .A(u2__abc_44228_n20756), .B(u2__abc_44228_n20759), .Y(u2__abc_44228_n20760) );
  AND2X2 AND2X2_10344 ( .A(u2__abc_44228_n20761), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_root_249__FF_INPUT) );
  AND2X2 AND2X2_10345 ( .A(u2__abc_44228_n3062_bF_buf43), .B(u2_o_249_), .Y(u2__abc_44228_n20763) );
  AND2X2 AND2X2_10346 ( .A(u2__abc_44228_n20753), .B(u2_o_248_), .Y(u2__abc_44228_n20765) );
  AND2X2 AND2X2_10347 ( .A(u2__abc_44228_n20766), .B(u2__abc_44228_n20764), .Y(u2__abc_44228_n20767) );
  AND2X2 AND2X2_10348 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n4330), .Y(u2__abc_44228_n20769) );
  AND2X2 AND2X2_10349 ( .A(u2__abc_44228_n20770), .B(u2__abc_44228_n2972_bF_buf46), .Y(u2__abc_44228_n20771) );
  AND2X2 AND2X2_1035 ( .A(u2__abc_44228_n4065), .B(u2__abc_44228_n4079), .Y(u2__abc_44228_n4080_1) );
  AND2X2 AND2X2_10350 ( .A(u2__abc_44228_n20768), .B(u2__abc_44228_n20771), .Y(u2__abc_44228_n20772) );
  AND2X2 AND2X2_10351 ( .A(u2__abc_44228_n20773), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_root_250__FF_INPUT) );
  AND2X2 AND2X2_10352 ( .A(u2__abc_44228_n3062_bF_buf42), .B(u2_o_250_), .Y(u2__abc_44228_n20775) );
  AND2X2 AND2X2_10353 ( .A(u2__abc_44228_n20765), .B(u2_o_249_), .Y(u2__abc_44228_n20777) );
  AND2X2 AND2X2_10354 ( .A(u2__abc_44228_n20778), .B(u2__abc_44228_n20776), .Y(u2__abc_44228_n20779) );
  AND2X2 AND2X2_10355 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n4315), .Y(u2__abc_44228_n20781) );
  AND2X2 AND2X2_10356 ( .A(u2__abc_44228_n20782), .B(u2__abc_44228_n2972_bF_buf45), .Y(u2__abc_44228_n20783) );
  AND2X2 AND2X2_10357 ( .A(u2__abc_44228_n20780), .B(u2__abc_44228_n20783), .Y(u2__abc_44228_n20784) );
  AND2X2 AND2X2_10358 ( .A(u2__abc_44228_n20785), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_root_251__FF_INPUT) );
  AND2X2 AND2X2_10359 ( .A(u2__abc_44228_n3062_bF_buf41), .B(u2_o_251_), .Y(u2__abc_44228_n20787) );
  AND2X2 AND2X2_1036 ( .A(u2__abc_44228_n4051), .B(u2__abc_44228_n4080_1), .Y(u2__abc_44228_n4081) );
  AND2X2 AND2X2_10360 ( .A(u2__abc_44228_n20777), .B(u2_o_250_), .Y(u2__abc_44228_n20789) );
  AND2X2 AND2X2_10361 ( .A(u2__abc_44228_n20790), .B(u2__abc_44228_n20788), .Y(u2__abc_44228_n20791) );
  AND2X2 AND2X2_10362 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n4321), .Y(u2__abc_44228_n20793) );
  AND2X2 AND2X2_10363 ( .A(u2__abc_44228_n20794), .B(u2__abc_44228_n2972_bF_buf44), .Y(u2__abc_44228_n20795) );
  AND2X2 AND2X2_10364 ( .A(u2__abc_44228_n20792), .B(u2__abc_44228_n20795), .Y(u2__abc_44228_n20796) );
  AND2X2 AND2X2_10365 ( .A(u2__abc_44228_n20797), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_root_252__FF_INPUT) );
  AND2X2 AND2X2_10366 ( .A(u2__abc_44228_n3062_bF_buf40), .B(u2_o_252_), .Y(u2__abc_44228_n20799) );
  AND2X2 AND2X2_10367 ( .A(u2__abc_44228_n20789), .B(u2_o_251_), .Y(u2__abc_44228_n20801) );
  AND2X2 AND2X2_10368 ( .A(u2__abc_44228_n20802), .B(u2__abc_44228_n20800), .Y(u2__abc_44228_n20803) );
  AND2X2 AND2X2_10369 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n4308), .Y(u2__abc_44228_n20805) );
  AND2X2 AND2X2_1037 ( .A(u2__abc_44228_n4082), .B(u2_remHi_69_), .Y(u2__abc_44228_n4083) );
  AND2X2 AND2X2_10370 ( .A(u2__abc_44228_n20806), .B(u2__abc_44228_n2972_bF_buf43), .Y(u2__abc_44228_n20807) );
  AND2X2 AND2X2_10371 ( .A(u2__abc_44228_n20804), .B(u2__abc_44228_n20807), .Y(u2__abc_44228_n20808) );
  AND2X2 AND2X2_10372 ( .A(u2__abc_44228_n20809), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_root_253__FF_INPUT) );
  AND2X2 AND2X2_10373 ( .A(u2__abc_44228_n3062_bF_buf39), .B(u2_o_253_), .Y(u2__abc_44228_n20811) );
  AND2X2 AND2X2_10374 ( .A(u2__abc_44228_n20801), .B(u2_o_252_), .Y(u2__abc_44228_n20813) );
  AND2X2 AND2X2_10375 ( .A(u2__abc_44228_n20814), .B(u2__abc_44228_n20812), .Y(u2__abc_44228_n20815) );
  AND2X2 AND2X2_10376 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n4301), .Y(u2__abc_44228_n20817) );
  AND2X2 AND2X2_10377 ( .A(u2__abc_44228_n20818), .B(u2__abc_44228_n2972_bF_buf42), .Y(u2__abc_44228_n20819) );
  AND2X2 AND2X2_10378 ( .A(u2__abc_44228_n20816), .B(u2__abc_44228_n20819), .Y(u2__abc_44228_n20820) );
  AND2X2 AND2X2_10379 ( .A(u2__abc_44228_n20821), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_root_254__FF_INPUT) );
  AND2X2 AND2X2_1038 ( .A(u2__abc_44228_n4085), .B(sqrto_69_), .Y(u2__abc_44228_n4086) );
  AND2X2 AND2X2_10380 ( .A(u2__abc_44228_n3062_bF_buf38), .B(u2_o_254_), .Y(u2__abc_44228_n20823) );
  AND2X2 AND2X2_10381 ( .A(u2__abc_44228_n20813), .B(u2_o_253_), .Y(u2__abc_44228_n20825) );
  AND2X2 AND2X2_10382 ( .A(u2__abc_44228_n20826), .B(u2__abc_44228_n20824), .Y(u2__abc_44228_n20827) );
  AND2X2 AND2X2_10383 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n6519), .Y(u2__abc_44228_n20829) );
  AND2X2 AND2X2_10384 ( .A(u2__abc_44228_n20830), .B(u2__abc_44228_n2972_bF_buf41), .Y(u2__abc_44228_n20831) );
  AND2X2 AND2X2_10385 ( .A(u2__abc_44228_n20828), .B(u2__abc_44228_n20831), .Y(u2__abc_44228_n20832) );
  AND2X2 AND2X2_10386 ( .A(u2__abc_44228_n20833), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_root_255__FF_INPUT) );
  AND2X2 AND2X2_10387 ( .A(u2__abc_44228_n3062_bF_buf37), .B(u2_o_255_), .Y(u2__abc_44228_n20835) );
  AND2X2 AND2X2_10388 ( .A(u2__abc_44228_n20825), .B(u2_o_254_), .Y(u2__abc_44228_n20837) );
  AND2X2 AND2X2_10389 ( .A(u2__abc_44228_n20838), .B(u2__abc_44228_n20836), .Y(u2__abc_44228_n20839) );
  AND2X2 AND2X2_1039 ( .A(u2__abc_44228_n4084), .B(u2__abc_44228_n4087), .Y(u2__abc_44228_n4088) );
  AND2X2 AND2X2_10390 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n6512), .Y(u2__abc_44228_n20841) );
  AND2X2 AND2X2_10391 ( .A(u2__abc_44228_n20842), .B(u2__abc_44228_n2972_bF_buf40), .Y(u2__abc_44228_n20843) );
  AND2X2 AND2X2_10392 ( .A(u2__abc_44228_n20840), .B(u2__abc_44228_n20843), .Y(u2__abc_44228_n20844) );
  AND2X2 AND2X2_10393 ( .A(u2__abc_44228_n20845), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_root_256__FF_INPUT) );
  AND2X2 AND2X2_10394 ( .A(u2__abc_44228_n3062_bF_buf36), .B(u2_o_256_), .Y(u2__abc_44228_n20847) );
  AND2X2 AND2X2_10395 ( .A(u2__abc_44228_n20837), .B(u2_o_255_), .Y(u2__abc_44228_n20849) );
  AND2X2 AND2X2_10396 ( .A(u2__abc_44228_n20850), .B(u2__abc_44228_n20848), .Y(u2__abc_44228_n20851) );
  AND2X2 AND2X2_10397 ( .A(u2__abc_44228_n2983_bF_buf104), .B(u2__abc_44228_n6505), .Y(u2__abc_44228_n20853) );
  AND2X2 AND2X2_10398 ( .A(u2__abc_44228_n20854), .B(u2__abc_44228_n2972_bF_buf39), .Y(u2__abc_44228_n20855) );
  AND2X2 AND2X2_10399 ( .A(u2__abc_44228_n20852), .B(u2__abc_44228_n20855), .Y(u2__abc_44228_n20856) );
  AND2X2 AND2X2_104 ( .A(_abc_64468_n912), .B(_abc_64468_n911), .Y(_auto_iopadmap_cc_313_execute_65414_139_) );
  AND2X2 AND2X2_1040 ( .A(u2__abc_44228_n4089), .B(u2_remHi_68_), .Y(u2__abc_44228_n4090_1) );
  AND2X2 AND2X2_10400 ( .A(u2__abc_44228_n20857), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_root_257__FF_INPUT) );
  AND2X2 AND2X2_10401 ( .A(u2__abc_44228_n3062_bF_buf35), .B(u2_o_257_), .Y(u2__abc_44228_n20859) );
  AND2X2 AND2X2_10402 ( .A(u2__abc_44228_n20849), .B(u2_o_256_), .Y(u2__abc_44228_n20861) );
  AND2X2 AND2X2_10403 ( .A(u2__abc_44228_n20862), .B(u2__abc_44228_n20860), .Y(u2__abc_44228_n20863) );
  AND2X2 AND2X2_10404 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n6498), .Y(u2__abc_44228_n20865) );
  AND2X2 AND2X2_10405 ( .A(u2__abc_44228_n20866), .B(u2__abc_44228_n2972_bF_buf38), .Y(u2__abc_44228_n20867) );
  AND2X2 AND2X2_10406 ( .A(u2__abc_44228_n20864), .B(u2__abc_44228_n20867), .Y(u2__abc_44228_n20868) );
  AND2X2 AND2X2_10407 ( .A(u2__abc_44228_n20869), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_root_258__FF_INPUT) );
  AND2X2 AND2X2_10408 ( .A(u2__abc_44228_n3062_bF_buf34), .B(u2_o_258_), .Y(u2__abc_44228_n20871) );
  AND2X2 AND2X2_10409 ( .A(u2__abc_44228_n20861), .B(u2_o_257_), .Y(u2__abc_44228_n20873) );
  AND2X2 AND2X2_1041 ( .A(u2__abc_44228_n4091), .B(sqrto_68_), .Y(u2__abc_44228_n4092) );
  AND2X2 AND2X2_10410 ( .A(u2__abc_44228_n20874), .B(u2__abc_44228_n20872), .Y(u2__abc_44228_n20875) );
  AND2X2 AND2X2_10411 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n6490), .Y(u2__abc_44228_n20877) );
  AND2X2 AND2X2_10412 ( .A(u2__abc_44228_n20878), .B(u2__abc_44228_n2972_bF_buf37), .Y(u2__abc_44228_n20879) );
  AND2X2 AND2X2_10413 ( .A(u2__abc_44228_n20876), .B(u2__abc_44228_n20879), .Y(u2__abc_44228_n20880) );
  AND2X2 AND2X2_10414 ( .A(u2__abc_44228_n20881), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_root_259__FF_INPUT) );
  AND2X2 AND2X2_10415 ( .A(u2__abc_44228_n3062_bF_buf33), .B(u2_o_259_), .Y(u2__abc_44228_n20883) );
  AND2X2 AND2X2_10416 ( .A(u2__abc_44228_n20873), .B(u2_o_258_), .Y(u2__abc_44228_n20885) );
  AND2X2 AND2X2_10417 ( .A(u2__abc_44228_n20886), .B(u2__abc_44228_n20884), .Y(u2__abc_44228_n20887) );
  AND2X2 AND2X2_10418 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n6483), .Y(u2__abc_44228_n20889) );
  AND2X2 AND2X2_10419 ( .A(u2__abc_44228_n20890), .B(u2__abc_44228_n2972_bF_buf36), .Y(u2__abc_44228_n20891) );
  AND2X2 AND2X2_1042 ( .A(u2__abc_44228_n4094), .B(u2__abc_44228_n4088), .Y(u2__abc_44228_n4095) );
  AND2X2 AND2X2_10420 ( .A(u2__abc_44228_n20888), .B(u2__abc_44228_n20891), .Y(u2__abc_44228_n20892) );
  AND2X2 AND2X2_10421 ( .A(u2__abc_44228_n20893), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_root_260__FF_INPUT) );
  AND2X2 AND2X2_10422 ( .A(u2__abc_44228_n3062_bF_buf32), .B(u2_o_260_), .Y(u2__abc_44228_n20895) );
  AND2X2 AND2X2_10423 ( .A(u2__abc_44228_n20885), .B(u2_o_259_), .Y(u2__abc_44228_n20897) );
  AND2X2 AND2X2_10424 ( .A(u2__abc_44228_n20898), .B(u2__abc_44228_n20896), .Y(u2__abc_44228_n20899) );
  AND2X2 AND2X2_10425 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n6476), .Y(u2__abc_44228_n20901) );
  AND2X2 AND2X2_10426 ( .A(u2__abc_44228_n20902), .B(u2__abc_44228_n2972_bF_buf35), .Y(u2__abc_44228_n20903) );
  AND2X2 AND2X2_10427 ( .A(u2__abc_44228_n20900), .B(u2__abc_44228_n20903), .Y(u2__abc_44228_n20904) );
  AND2X2 AND2X2_10428 ( .A(u2__abc_44228_n20905), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_root_261__FF_INPUT) );
  AND2X2 AND2X2_10429 ( .A(u2__abc_44228_n3062_bF_buf31), .B(u2_o_261_), .Y(u2__abc_44228_n20907) );
  AND2X2 AND2X2_1043 ( .A(u2__abc_44228_n4096), .B(u2_remHi_67_), .Y(u2__abc_44228_n4097) );
  AND2X2 AND2X2_10430 ( .A(u2__abc_44228_n20897), .B(u2_o_260_), .Y(u2__abc_44228_n20909) );
  AND2X2 AND2X2_10431 ( .A(u2__abc_44228_n20910), .B(u2__abc_44228_n20908), .Y(u2__abc_44228_n20911) );
  AND2X2 AND2X2_10432 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n6469), .Y(u2__abc_44228_n20913) );
  AND2X2 AND2X2_10433 ( .A(u2__abc_44228_n20914), .B(u2__abc_44228_n2972_bF_buf34), .Y(u2__abc_44228_n20915) );
  AND2X2 AND2X2_10434 ( .A(u2__abc_44228_n20912), .B(u2__abc_44228_n20915), .Y(u2__abc_44228_n20916) );
  AND2X2 AND2X2_10435 ( .A(u2__abc_44228_n20917), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_root_262__FF_INPUT) );
  AND2X2 AND2X2_10436 ( .A(u2__abc_44228_n3062_bF_buf30), .B(u2_o_262_), .Y(u2__abc_44228_n20919) );
  AND2X2 AND2X2_10437 ( .A(u2__abc_44228_n20909), .B(u2_o_261_), .Y(u2__abc_44228_n20921) );
  AND2X2 AND2X2_10438 ( .A(u2__abc_44228_n20922), .B(u2__abc_44228_n20920), .Y(u2__abc_44228_n20923) );
  AND2X2 AND2X2_10439 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n6460), .Y(u2__abc_44228_n20925) );
  AND2X2 AND2X2_1044 ( .A(u2__abc_44228_n4099), .B(sqrto_67_), .Y(u2__abc_44228_n4100_1) );
  AND2X2 AND2X2_10440 ( .A(u2__abc_44228_n20926), .B(u2__abc_44228_n2972_bF_buf33), .Y(u2__abc_44228_n20927) );
  AND2X2 AND2X2_10441 ( .A(u2__abc_44228_n20924), .B(u2__abc_44228_n20927), .Y(u2__abc_44228_n20928) );
  AND2X2 AND2X2_10442 ( .A(u2__abc_44228_n20929), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_root_263__FF_INPUT) );
  AND2X2 AND2X2_10443 ( .A(u2__abc_44228_n3062_bF_buf29), .B(u2_o_263_), .Y(u2__abc_44228_n20931) );
  AND2X2 AND2X2_10444 ( .A(u2__abc_44228_n20921), .B(u2_o_262_), .Y(u2__abc_44228_n20933) );
  AND2X2 AND2X2_10445 ( .A(u2__abc_44228_n20934), .B(u2__abc_44228_n20932), .Y(u2__abc_44228_n20935) );
  AND2X2 AND2X2_10446 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n6453_1), .Y(u2__abc_44228_n20937) );
  AND2X2 AND2X2_10447 ( .A(u2__abc_44228_n20938), .B(u2__abc_44228_n2972_bF_buf32), .Y(u2__abc_44228_n20939) );
  AND2X2 AND2X2_10448 ( .A(u2__abc_44228_n20936), .B(u2__abc_44228_n20939), .Y(u2__abc_44228_n20940) );
  AND2X2 AND2X2_10449 ( .A(u2__abc_44228_n20941), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_root_264__FF_INPUT) );
  AND2X2 AND2X2_1045 ( .A(u2__abc_44228_n4098), .B(u2__abc_44228_n4101), .Y(u2__abc_44228_n4102) );
  AND2X2 AND2X2_10450 ( .A(u2__abc_44228_n3062_bF_buf28), .B(u2_o_264_), .Y(u2__abc_44228_n20943) );
  AND2X2 AND2X2_10451 ( .A(u2__abc_44228_n20933), .B(u2_o_263_), .Y(u2__abc_44228_n20945) );
  AND2X2 AND2X2_10452 ( .A(u2__abc_44228_n20946), .B(u2__abc_44228_n20944), .Y(u2__abc_44228_n20947) );
  AND2X2 AND2X2_10453 ( .A(u2__abc_44228_n2983_bF_buf88), .B(u2__abc_44228_n6446), .Y(u2__abc_44228_n20949) );
  AND2X2 AND2X2_10454 ( .A(u2__abc_44228_n20950), .B(u2__abc_44228_n2972_bF_buf31), .Y(u2__abc_44228_n20951) );
  AND2X2 AND2X2_10455 ( .A(u2__abc_44228_n20948), .B(u2__abc_44228_n20951), .Y(u2__abc_44228_n20952) );
  AND2X2 AND2X2_10456 ( .A(u2__abc_44228_n20953), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_root_265__FF_INPUT) );
  AND2X2 AND2X2_10457 ( .A(u2__abc_44228_n3062_bF_buf27), .B(u2_o_265_), .Y(u2__abc_44228_n20955) );
  AND2X2 AND2X2_10458 ( .A(u2__abc_44228_n20945), .B(u2_o_264_), .Y(u2__abc_44228_n20957) );
  AND2X2 AND2X2_10459 ( .A(u2__abc_44228_n20958), .B(u2__abc_44228_n20956), .Y(u2__abc_44228_n20959) );
  AND2X2 AND2X2_1046 ( .A(u2__abc_44228_n4103), .B(u2_remHi_66_), .Y(u2__abc_44228_n4104) );
  AND2X2 AND2X2_10460 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n6439), .Y(u2__abc_44228_n20961) );
  AND2X2 AND2X2_10461 ( .A(u2__abc_44228_n20962), .B(u2__abc_44228_n2972_bF_buf30), .Y(u2__abc_44228_n20963) );
  AND2X2 AND2X2_10462 ( .A(u2__abc_44228_n20960), .B(u2__abc_44228_n20963), .Y(u2__abc_44228_n20964) );
  AND2X2 AND2X2_10463 ( .A(u2__abc_44228_n20965), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_root_266__FF_INPUT) );
  AND2X2 AND2X2_10464 ( .A(u2__abc_44228_n3062_bF_buf26), .B(u2_o_266_), .Y(u2__abc_44228_n20967) );
  AND2X2 AND2X2_10465 ( .A(u2__abc_44228_n20957), .B(u2_o_265_), .Y(u2__abc_44228_n20969) );
  AND2X2 AND2X2_10466 ( .A(u2__abc_44228_n20970), .B(u2__abc_44228_n20968), .Y(u2__abc_44228_n20971) );
  AND2X2 AND2X2_10467 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n6431), .Y(u2__abc_44228_n20973) );
  AND2X2 AND2X2_10468 ( .A(u2__abc_44228_n20974), .B(u2__abc_44228_n2972_bF_buf29), .Y(u2__abc_44228_n20975) );
  AND2X2 AND2X2_10469 ( .A(u2__abc_44228_n20972), .B(u2__abc_44228_n20975), .Y(u2__abc_44228_n20976) );
  AND2X2 AND2X2_1047 ( .A(u2__abc_44228_n4105), .B(sqrto_66_), .Y(u2__abc_44228_n4106) );
  AND2X2 AND2X2_10470 ( .A(u2__abc_44228_n20977), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_root_267__FF_INPUT) );
  AND2X2 AND2X2_10471 ( .A(u2__abc_44228_n3062_bF_buf25), .B(u2_o_267_), .Y(u2__abc_44228_n20979) );
  AND2X2 AND2X2_10472 ( .A(u2__abc_44228_n20969), .B(u2_o_266_), .Y(u2__abc_44228_n20981) );
  AND2X2 AND2X2_10473 ( .A(u2__abc_44228_n20982), .B(u2__abc_44228_n20980), .Y(u2__abc_44228_n20983) );
  AND2X2 AND2X2_10474 ( .A(u2__abc_44228_n2983_bF_buf82), .B(u2__abc_44228_n6424), .Y(u2__abc_44228_n20985) );
  AND2X2 AND2X2_10475 ( .A(u2__abc_44228_n20986), .B(u2__abc_44228_n2972_bF_buf28), .Y(u2__abc_44228_n20987) );
  AND2X2 AND2X2_10476 ( .A(u2__abc_44228_n20984), .B(u2__abc_44228_n20987), .Y(u2__abc_44228_n20988) );
  AND2X2 AND2X2_10477 ( .A(u2__abc_44228_n20989), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_root_268__FF_INPUT) );
  AND2X2 AND2X2_10478 ( .A(u2__abc_44228_n3062_bF_buf24), .B(u2_o_268_), .Y(u2__abc_44228_n20991) );
  AND2X2 AND2X2_10479 ( .A(u2__abc_44228_n20981), .B(u2_o_267_), .Y(u2__abc_44228_n20993) );
  AND2X2 AND2X2_1048 ( .A(u2__abc_44228_n4108), .B(u2__abc_44228_n4102), .Y(u2__abc_44228_n4109_1) );
  AND2X2 AND2X2_10480 ( .A(u2__abc_44228_n20994), .B(u2__abc_44228_n20992), .Y(u2__abc_44228_n20995) );
  AND2X2 AND2X2_10481 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n6417), .Y(u2__abc_44228_n20997) );
  AND2X2 AND2X2_10482 ( .A(u2__abc_44228_n20998), .B(u2__abc_44228_n2972_bF_buf27), .Y(u2__abc_44228_n20999) );
  AND2X2 AND2X2_10483 ( .A(u2__abc_44228_n20996), .B(u2__abc_44228_n20999), .Y(u2__abc_44228_n21000) );
  AND2X2 AND2X2_10484 ( .A(u2__abc_44228_n21001), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_root_269__FF_INPUT) );
  AND2X2 AND2X2_10485 ( .A(u2__abc_44228_n3062_bF_buf23), .B(u2_o_269_), .Y(u2__abc_44228_n21003) );
  AND2X2 AND2X2_10486 ( .A(u2__abc_44228_n20993), .B(u2_o_268_), .Y(u2__abc_44228_n21005) );
  AND2X2 AND2X2_10487 ( .A(u2__abc_44228_n21006), .B(u2__abc_44228_n21004), .Y(u2__abc_44228_n21007) );
  AND2X2 AND2X2_10488 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n6410), .Y(u2__abc_44228_n21009) );
  AND2X2 AND2X2_10489 ( .A(u2__abc_44228_n21010), .B(u2__abc_44228_n2972_bF_buf26), .Y(u2__abc_44228_n21011) );
  AND2X2 AND2X2_1049 ( .A(u2__abc_44228_n4095), .B(u2__abc_44228_n4109_1), .Y(u2__abc_44228_n4110) );
  AND2X2 AND2X2_10490 ( .A(u2__abc_44228_n21008), .B(u2__abc_44228_n21011), .Y(u2__abc_44228_n21012) );
  AND2X2 AND2X2_10491 ( .A(u2__abc_44228_n21013), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_root_270__FF_INPUT) );
  AND2X2 AND2X2_10492 ( .A(u2__abc_44228_n3062_bF_buf22), .B(u2_o_270_), .Y(u2__abc_44228_n21015) );
  AND2X2 AND2X2_10493 ( .A(u2__abc_44228_n21005), .B(u2_o_269_), .Y(u2__abc_44228_n21017) );
  AND2X2 AND2X2_10494 ( .A(u2__abc_44228_n21018), .B(u2__abc_44228_n21016), .Y(u2__abc_44228_n21019) );
  AND2X2 AND2X2_10495 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n6393), .Y(u2__abc_44228_n21021) );
  AND2X2 AND2X2_10496 ( .A(u2__abc_44228_n21022), .B(u2__abc_44228_n2972_bF_buf25), .Y(u2__abc_44228_n21023) );
  AND2X2 AND2X2_10497 ( .A(u2__abc_44228_n21020), .B(u2__abc_44228_n21023), .Y(u2__abc_44228_n21024) );
  AND2X2 AND2X2_10498 ( .A(u2__abc_44228_n21025), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_root_271__FF_INPUT) );
  AND2X2 AND2X2_10499 ( .A(u2__abc_44228_n3062_bF_buf21), .B(u2_o_271_), .Y(u2__abc_44228_n21027) );
  AND2X2 AND2X2_105 ( .A(_abc_64468_n915), .B(_abc_64468_n914), .Y(_auto_iopadmap_cc_313_execute_65414_140_) );
  AND2X2 AND2X2_1050 ( .A(u2__abc_44228_n4112), .B(u2__abc_44228_n4114), .Y(u2__abc_44228_n4115) );
  AND2X2 AND2X2_10500 ( .A(u2__abc_44228_n21017), .B(u2_o_270_), .Y(u2__abc_44228_n21029) );
  AND2X2 AND2X2_10501 ( .A(u2__abc_44228_n21030), .B(u2__abc_44228_n21028), .Y(u2__abc_44228_n21031) );
  AND2X2 AND2X2_10502 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n6399), .Y(u2__abc_44228_n21033) );
  AND2X2 AND2X2_10503 ( .A(u2__abc_44228_n21034), .B(u2__abc_44228_n2972_bF_buf24), .Y(u2__abc_44228_n21035) );
  AND2X2 AND2X2_10504 ( .A(u2__abc_44228_n21032), .B(u2__abc_44228_n21035), .Y(u2__abc_44228_n21036) );
  AND2X2 AND2X2_10505 ( .A(u2__abc_44228_n21037), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_root_272__FF_INPUT) );
  AND2X2 AND2X2_10506 ( .A(u2__abc_44228_n3062_bF_buf20), .B(u2_o_272_), .Y(u2__abc_44228_n21039) );
  AND2X2 AND2X2_10507 ( .A(u2__abc_44228_n21029), .B(u2_o_271_), .Y(u2__abc_44228_n21041) );
  AND2X2 AND2X2_10508 ( .A(u2__abc_44228_n21042), .B(u2__abc_44228_n21040), .Y(u2__abc_44228_n21043) );
  AND2X2 AND2X2_10509 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n6386), .Y(u2__abc_44228_n21045) );
  AND2X2 AND2X2_1051 ( .A(u2__abc_44228_n4117), .B(u2__abc_44228_n4119_1), .Y(u2__abc_44228_n4120) );
  AND2X2 AND2X2_10510 ( .A(u2__abc_44228_n21046), .B(u2__abc_44228_n2972_bF_buf23), .Y(u2__abc_44228_n21047) );
  AND2X2 AND2X2_10511 ( .A(u2__abc_44228_n21044), .B(u2__abc_44228_n21047), .Y(u2__abc_44228_n21048) );
  AND2X2 AND2X2_10512 ( .A(u2__abc_44228_n21049), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_root_273__FF_INPUT) );
  AND2X2 AND2X2_10513 ( .A(u2__abc_44228_n3062_bF_buf19), .B(u2_o_273_), .Y(u2__abc_44228_n21051) );
  AND2X2 AND2X2_10514 ( .A(u2__abc_44228_n21041), .B(u2_o_272_), .Y(u2__abc_44228_n21053) );
  AND2X2 AND2X2_10515 ( .A(u2__abc_44228_n21054), .B(u2__abc_44228_n21052), .Y(u2__abc_44228_n21055) );
  AND2X2 AND2X2_10516 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n6379_1), .Y(u2__abc_44228_n21057) );
  AND2X2 AND2X2_10517 ( .A(u2__abc_44228_n21058), .B(u2__abc_44228_n2972_bF_buf22), .Y(u2__abc_44228_n21059) );
  AND2X2 AND2X2_10518 ( .A(u2__abc_44228_n21056), .B(u2__abc_44228_n21059), .Y(u2__abc_44228_n21060) );
  AND2X2 AND2X2_10519 ( .A(u2__abc_44228_n21061), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_root_274__FF_INPUT) );
  AND2X2 AND2X2_1052 ( .A(u2__abc_44228_n4115), .B(u2__abc_44228_n4120), .Y(u2__abc_44228_n4121) );
  AND2X2 AND2X2_10520 ( .A(u2__abc_44228_n3062_bF_buf18), .B(u2_o_274_), .Y(u2__abc_44228_n21063) );
  AND2X2 AND2X2_10521 ( .A(u2__abc_44228_n21053), .B(u2_o_273_), .Y(u2__abc_44228_n21065) );
  AND2X2 AND2X2_10522 ( .A(u2__abc_44228_n21066), .B(u2__abc_44228_n21064), .Y(u2__abc_44228_n21067) );
  AND2X2 AND2X2_10523 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n6371_1), .Y(u2__abc_44228_n21069) );
  AND2X2 AND2X2_10524 ( .A(u2__abc_44228_n21070), .B(u2__abc_44228_n2972_bF_buf21), .Y(u2__abc_44228_n21071) );
  AND2X2 AND2X2_10525 ( .A(u2__abc_44228_n21068), .B(u2__abc_44228_n21071), .Y(u2__abc_44228_n21072) );
  AND2X2 AND2X2_10526 ( .A(u2__abc_44228_n21073), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_root_275__FF_INPUT) );
  AND2X2 AND2X2_10527 ( .A(u2__abc_44228_n3062_bF_buf17), .B(u2_o_275_), .Y(u2__abc_44228_n21075) );
  AND2X2 AND2X2_10528 ( .A(u2__abc_44228_n21065), .B(u2_o_274_), .Y(u2__abc_44228_n21077) );
  AND2X2 AND2X2_10529 ( .A(u2__abc_44228_n21078), .B(u2__abc_44228_n21076), .Y(u2__abc_44228_n21079) );
  AND2X2 AND2X2_1053 ( .A(u2__abc_44228_n4122), .B(u2_remHi_63_), .Y(u2__abc_44228_n4123) );
  AND2X2 AND2X2_10530 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n6364), .Y(u2__abc_44228_n21081) );
  AND2X2 AND2X2_10531 ( .A(u2__abc_44228_n21082), .B(u2__abc_44228_n2972_bF_buf20), .Y(u2__abc_44228_n21083) );
  AND2X2 AND2X2_10532 ( .A(u2__abc_44228_n21080), .B(u2__abc_44228_n21083), .Y(u2__abc_44228_n21084) );
  AND2X2 AND2X2_10533 ( .A(u2__abc_44228_n21085), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_root_276__FF_INPUT) );
  AND2X2 AND2X2_10534 ( .A(u2__abc_44228_n3062_bF_buf16), .B(u2_o_276_), .Y(u2__abc_44228_n21087) );
  AND2X2 AND2X2_10535 ( .A(u2__abc_44228_n21077), .B(u2_o_275_), .Y(u2__abc_44228_n21089) );
  AND2X2 AND2X2_10536 ( .A(u2__abc_44228_n21090), .B(u2__abc_44228_n21088), .Y(u2__abc_44228_n21091) );
  AND2X2 AND2X2_10537 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n6357), .Y(u2__abc_44228_n21093) );
  AND2X2 AND2X2_10538 ( .A(u2__abc_44228_n21094), .B(u2__abc_44228_n2972_bF_buf19), .Y(u2__abc_44228_n21095) );
  AND2X2 AND2X2_10539 ( .A(u2__abc_44228_n21092), .B(u2__abc_44228_n21095), .Y(u2__abc_44228_n21096) );
  AND2X2 AND2X2_1054 ( .A(u2__abc_44228_n4125), .B(sqrto_63_), .Y(u2__abc_44228_n4126) );
  AND2X2 AND2X2_10540 ( .A(u2__abc_44228_n21097), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_root_277__FF_INPUT) );
  AND2X2 AND2X2_10541 ( .A(u2__abc_44228_n3062_bF_buf15), .B(u2_o_277_), .Y(u2__abc_44228_n21099) );
  AND2X2 AND2X2_10542 ( .A(u2__abc_44228_n21089), .B(u2_o_276_), .Y(u2__abc_44228_n21101) );
  AND2X2 AND2X2_10543 ( .A(u2__abc_44228_n21102), .B(u2__abc_44228_n21100), .Y(u2__abc_44228_n21103) );
  AND2X2 AND2X2_10544 ( .A(u2__abc_44228_n2983_bF_buf62), .B(u2__abc_44228_n6350), .Y(u2__abc_44228_n21105) );
  AND2X2 AND2X2_10545 ( .A(u2__abc_44228_n21106), .B(u2__abc_44228_n2972_bF_buf18), .Y(u2__abc_44228_n21107) );
  AND2X2 AND2X2_10546 ( .A(u2__abc_44228_n21104), .B(u2__abc_44228_n21107), .Y(u2__abc_44228_n21108) );
  AND2X2 AND2X2_10547 ( .A(u2__abc_44228_n21109), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_root_278__FF_INPUT) );
  AND2X2 AND2X2_10548 ( .A(u2__abc_44228_n3062_bF_buf14), .B(u2_o_278_), .Y(u2__abc_44228_n21111) );
  AND2X2 AND2X2_10549 ( .A(u2__abc_44228_n21101), .B(u2_o_277_), .Y(u2__abc_44228_n21113) );
  AND2X2 AND2X2_1055 ( .A(u2__abc_44228_n4124), .B(u2__abc_44228_n4127), .Y(u2__abc_44228_n4128_1) );
  AND2X2 AND2X2_10550 ( .A(u2__abc_44228_n21114), .B(u2__abc_44228_n21112), .Y(u2__abc_44228_n21115) );
  AND2X2 AND2X2_10551 ( .A(u2__abc_44228_n2983_bF_buf60), .B(u2__abc_44228_n6327), .Y(u2__abc_44228_n21117) );
  AND2X2 AND2X2_10552 ( .A(u2__abc_44228_n21118), .B(u2__abc_44228_n2972_bF_buf17), .Y(u2__abc_44228_n21119) );
  AND2X2 AND2X2_10553 ( .A(u2__abc_44228_n21116), .B(u2__abc_44228_n21119), .Y(u2__abc_44228_n21120) );
  AND2X2 AND2X2_10554 ( .A(u2__abc_44228_n21121), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_root_279__FF_INPUT) );
  AND2X2 AND2X2_10555 ( .A(u2__abc_44228_n3062_bF_buf13), .B(u2_o_279_), .Y(u2__abc_44228_n21123) );
  AND2X2 AND2X2_10556 ( .A(u2__abc_44228_n21113), .B(u2_o_278_), .Y(u2__abc_44228_n21125) );
  AND2X2 AND2X2_10557 ( .A(u2__abc_44228_n21126), .B(u2__abc_44228_n21124), .Y(u2__abc_44228_n21127) );
  AND2X2 AND2X2_10558 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n6320), .Y(u2__abc_44228_n21129) );
  AND2X2 AND2X2_10559 ( .A(u2__abc_44228_n21130), .B(u2__abc_44228_n2972_bF_buf16), .Y(u2__abc_44228_n21131) );
  AND2X2 AND2X2_1056 ( .A(u2__abc_44228_n4129), .B(u2_remHi_62_), .Y(u2__abc_44228_n4130) );
  AND2X2 AND2X2_10560 ( .A(u2__abc_44228_n21128), .B(u2__abc_44228_n21131), .Y(u2__abc_44228_n21132) );
  AND2X2 AND2X2_10561 ( .A(u2__abc_44228_n21133), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_root_280__FF_INPUT) );
  AND2X2 AND2X2_10562 ( .A(u2__abc_44228_n3062_bF_buf12), .B(u2_o_280_), .Y(u2__abc_44228_n21135) );
  AND2X2 AND2X2_10563 ( .A(u2__abc_44228_n21125), .B(u2_o_279_), .Y(u2__abc_44228_n21137) );
  AND2X2 AND2X2_10564 ( .A(u2__abc_44228_n21138), .B(u2__abc_44228_n21136), .Y(u2__abc_44228_n21139) );
  AND2X2 AND2X2_10565 ( .A(u2__abc_44228_n2983_bF_buf56), .B(u2__abc_44228_n6341), .Y(u2__abc_44228_n21141) );
  AND2X2 AND2X2_10566 ( .A(u2__abc_44228_n21142), .B(u2__abc_44228_n2972_bF_buf15), .Y(u2__abc_44228_n21143) );
  AND2X2 AND2X2_10567 ( .A(u2__abc_44228_n21140), .B(u2__abc_44228_n21143), .Y(u2__abc_44228_n21144) );
  AND2X2 AND2X2_10568 ( .A(u2__abc_44228_n21145), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_root_281__FF_INPUT) );
  AND2X2 AND2X2_10569 ( .A(u2__abc_44228_n3062_bF_buf11), .B(u2_o_281_), .Y(u2__abc_44228_n21147) );
  AND2X2 AND2X2_1057 ( .A(u2__abc_44228_n4131), .B(sqrto_62_), .Y(u2__abc_44228_n4132) );
  AND2X2 AND2X2_10570 ( .A(u2__abc_44228_n21137), .B(u2_o_280_), .Y(u2__abc_44228_n21149) );
  AND2X2 AND2X2_10571 ( .A(u2__abc_44228_n21150), .B(u2__abc_44228_n21148), .Y(u2__abc_44228_n21151) );
  AND2X2 AND2X2_10572 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n6334), .Y(u2__abc_44228_n21153) );
  AND2X2 AND2X2_10573 ( .A(u2__abc_44228_n21154), .B(u2__abc_44228_n2972_bF_buf14), .Y(u2__abc_44228_n21155) );
  AND2X2 AND2X2_10574 ( .A(u2__abc_44228_n21152), .B(u2__abc_44228_n21155), .Y(u2__abc_44228_n21156) );
  AND2X2 AND2X2_10575 ( .A(u2__abc_44228_n21157), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_root_282__FF_INPUT) );
  AND2X2 AND2X2_10576 ( .A(u2__abc_44228_n3062_bF_buf10), .B(u2_o_282_), .Y(u2__abc_44228_n21159) );
  AND2X2 AND2X2_10577 ( .A(u2__abc_44228_n21149), .B(u2_o_281_), .Y(u2__abc_44228_n21161) );
  AND2X2 AND2X2_10578 ( .A(u2__abc_44228_n21162), .B(u2__abc_44228_n21160), .Y(u2__abc_44228_n21163) );
  AND2X2 AND2X2_10579 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n6312), .Y(u2__abc_44228_n21165) );
  AND2X2 AND2X2_1058 ( .A(u2__abc_44228_n4134), .B(u2__abc_44228_n4128_1), .Y(u2__abc_44228_n4135) );
  AND2X2 AND2X2_10580 ( .A(u2__abc_44228_n21166), .B(u2__abc_44228_n2972_bF_buf13), .Y(u2__abc_44228_n21167) );
  AND2X2 AND2X2_10581 ( .A(u2__abc_44228_n21164), .B(u2__abc_44228_n21167), .Y(u2__abc_44228_n21168) );
  AND2X2 AND2X2_10582 ( .A(u2__abc_44228_n21169), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_root_283__FF_INPUT) );
  AND2X2 AND2X2_10583 ( .A(u2__abc_44228_n3062_bF_buf9), .B(u2_o_283_), .Y(u2__abc_44228_n21171) );
  AND2X2 AND2X2_10584 ( .A(u2__abc_44228_n21161), .B(u2_o_282_), .Y(u2__abc_44228_n21173) );
  AND2X2 AND2X2_10585 ( .A(u2__abc_44228_n21174), .B(u2__abc_44228_n21172), .Y(u2__abc_44228_n21175) );
  AND2X2 AND2X2_10586 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2__abc_44228_n6305_1), .Y(u2__abc_44228_n21177) );
  AND2X2 AND2X2_10587 ( .A(u2__abc_44228_n21178), .B(u2__abc_44228_n2972_bF_buf12), .Y(u2__abc_44228_n21179) );
  AND2X2 AND2X2_10588 ( .A(u2__abc_44228_n21176), .B(u2__abc_44228_n21179), .Y(u2__abc_44228_n21180) );
  AND2X2 AND2X2_10589 ( .A(u2__abc_44228_n21181), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_root_284__FF_INPUT) );
  AND2X2 AND2X2_1059 ( .A(u2__abc_44228_n4135), .B(u2__abc_44228_n4121), .Y(u2__abc_44228_n4136) );
  AND2X2 AND2X2_10590 ( .A(u2__abc_44228_n3062_bF_buf8), .B(u2_o_284_), .Y(u2__abc_44228_n21183) );
  AND2X2 AND2X2_10591 ( .A(u2__abc_44228_n21173), .B(u2_o_283_), .Y(u2__abc_44228_n21185) );
  AND2X2 AND2X2_10592 ( .A(u2__abc_44228_n21186), .B(u2__abc_44228_n21184), .Y(u2__abc_44228_n21187) );
  AND2X2 AND2X2_10593 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n6298), .Y(u2__abc_44228_n21189) );
  AND2X2 AND2X2_10594 ( .A(u2__abc_44228_n21190), .B(u2__abc_44228_n2972_bF_buf11), .Y(u2__abc_44228_n21191) );
  AND2X2 AND2X2_10595 ( .A(u2__abc_44228_n21188), .B(u2__abc_44228_n21191), .Y(u2__abc_44228_n21192) );
  AND2X2 AND2X2_10596 ( .A(u2__abc_44228_n21193), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_root_285__FF_INPUT) );
  AND2X2 AND2X2_10597 ( .A(u2__abc_44228_n3062_bF_buf7), .B(u2_o_285_), .Y(u2__abc_44228_n21195) );
  AND2X2 AND2X2_10598 ( .A(u2__abc_44228_n21185), .B(u2_o_284_), .Y(u2__abc_44228_n21197) );
  AND2X2 AND2X2_10599 ( .A(u2__abc_44228_n21198), .B(u2__abc_44228_n21196), .Y(u2__abc_44228_n21199) );
  AND2X2 AND2X2_106 ( .A(_abc_64468_n918), .B(_abc_64468_n917), .Y(_auto_iopadmap_cc_313_execute_65414_141_) );
  AND2X2 AND2X2_1060 ( .A(u2__abc_44228_n4110), .B(u2__abc_44228_n4136), .Y(u2__abc_44228_n4137) );
  AND2X2 AND2X2_10600 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n6291), .Y(u2__abc_44228_n21201) );
  AND2X2 AND2X2_10601 ( .A(u2__abc_44228_n21202), .B(u2__abc_44228_n2972_bF_buf10), .Y(u2__abc_44228_n21203) );
  AND2X2 AND2X2_10602 ( .A(u2__abc_44228_n21200), .B(u2__abc_44228_n21203), .Y(u2__abc_44228_n21204) );
  AND2X2 AND2X2_10603 ( .A(u2__abc_44228_n21205), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_root_286__FF_INPUT) );
  AND2X2 AND2X2_10604 ( .A(u2__abc_44228_n3062_bF_buf6), .B(u2_o_286_), .Y(u2__abc_44228_n21207) );
  AND2X2 AND2X2_10605 ( .A(u2__abc_44228_n21197), .B(u2_o_285_), .Y(u2__abc_44228_n21209) );
  AND2X2 AND2X2_10606 ( .A(u2__abc_44228_n21210), .B(u2__abc_44228_n21208), .Y(u2__abc_44228_n21211) );
  AND2X2 AND2X2_10607 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n6280), .Y(u2__abc_44228_n21213) );
  AND2X2 AND2X2_10608 ( .A(u2__abc_44228_n21214), .B(u2__abc_44228_n2972_bF_buf9), .Y(u2__abc_44228_n21215) );
  AND2X2 AND2X2_10609 ( .A(u2__abc_44228_n21212), .B(u2__abc_44228_n21215), .Y(u2__abc_44228_n21216) );
  AND2X2 AND2X2_1061 ( .A(u2__abc_44228_n4081), .B(u2__abc_44228_n4137), .Y(u2__abc_44228_n4138_1) );
  AND2X2 AND2X2_10610 ( .A(u2__abc_44228_n21217), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_root_287__FF_INPUT) );
  AND2X2 AND2X2_10611 ( .A(u2__abc_44228_n3062_bF_buf5), .B(u2_o_287_), .Y(u2__abc_44228_n21219) );
  AND2X2 AND2X2_10612 ( .A(u2__abc_44228_n21209), .B(u2_o_286_), .Y(u2__abc_44228_n21221) );
  AND2X2 AND2X2_10613 ( .A(u2__abc_44228_n21222), .B(u2__abc_44228_n21220), .Y(u2__abc_44228_n21223) );
  AND2X2 AND2X2_10614 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n6273), .Y(u2__abc_44228_n21225) );
  AND2X2 AND2X2_10615 ( .A(u2__abc_44228_n21226), .B(u2__abc_44228_n2972_bF_buf8), .Y(u2__abc_44228_n21227) );
  AND2X2 AND2X2_10616 ( .A(u2__abc_44228_n21224), .B(u2__abc_44228_n21227), .Y(u2__abc_44228_n21228) );
  AND2X2 AND2X2_10617 ( .A(u2__abc_44228_n21229), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_root_288__FF_INPUT) );
  AND2X2 AND2X2_10618 ( .A(u2__abc_44228_n3062_bF_buf4), .B(u2_o_288_), .Y(u2__abc_44228_n21231) );
  AND2X2 AND2X2_10619 ( .A(u2__abc_44228_n21221), .B(u2_o_287_), .Y(u2__abc_44228_n21233) );
  AND2X2 AND2X2_1062 ( .A(u2__abc_44228_n4022), .B(u2__abc_44228_n4138_1), .Y(u2__abc_44228_n4139) );
  AND2X2 AND2X2_10620 ( .A(u2__abc_44228_n21234), .B(u2__abc_44228_n21232), .Y(u2__abc_44228_n21235) );
  AND2X2 AND2X2_10621 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n6266), .Y(u2__abc_44228_n21237) );
  AND2X2 AND2X2_10622 ( .A(u2__abc_44228_n21238), .B(u2__abc_44228_n2972_bF_buf7), .Y(u2__abc_44228_n21239) );
  AND2X2 AND2X2_10623 ( .A(u2__abc_44228_n21236), .B(u2__abc_44228_n21239), .Y(u2__abc_44228_n21240) );
  AND2X2 AND2X2_10624 ( .A(u2__abc_44228_n21241), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_root_289__FF_INPUT) );
  AND2X2 AND2X2_10625 ( .A(u2__abc_44228_n3062_bF_buf3), .B(u2_o_289_), .Y(u2__abc_44228_n21243) );
  AND2X2 AND2X2_10626 ( .A(u2__abc_44228_n21233), .B(u2_o_288_), .Y(u2__abc_44228_n21245) );
  AND2X2 AND2X2_10627 ( .A(u2__abc_44228_n21246), .B(u2__abc_44228_n21244), .Y(u2__abc_44228_n21247) );
  AND2X2 AND2X2_10628 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n6259), .Y(u2__abc_44228_n21249) );
  AND2X2 AND2X2_10629 ( .A(u2__abc_44228_n21250), .B(u2__abc_44228_n2972_bF_buf6), .Y(u2__abc_44228_n21251) );
  AND2X2 AND2X2_1063 ( .A(u2__abc_44228_n3903_1), .B(u2__abc_44228_n4139), .Y(u2__abc_44228_n4140) );
  AND2X2 AND2X2_10630 ( .A(u2__abc_44228_n21248), .B(u2__abc_44228_n21251), .Y(u2__abc_44228_n21252) );
  AND2X2 AND2X2_10631 ( .A(u2__abc_44228_n21253), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_root_290__FF_INPUT) );
  AND2X2 AND2X2_10632 ( .A(u2__abc_44228_n3062_bF_buf2), .B(u2_o_290_), .Y(u2__abc_44228_n21255) );
  AND2X2 AND2X2_10633 ( .A(u2__abc_44228_n21245), .B(u2_o_289_), .Y(u2__abc_44228_n21257) );
  AND2X2 AND2X2_10634 ( .A(u2__abc_44228_n21258), .B(u2__abc_44228_n21256), .Y(u2__abc_44228_n21259) );
  AND2X2 AND2X2_10635 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n6251_1), .Y(u2__abc_44228_n21261) );
  AND2X2 AND2X2_10636 ( .A(u2__abc_44228_n21262), .B(u2__abc_44228_n2972_bF_buf5), .Y(u2__abc_44228_n21263) );
  AND2X2 AND2X2_10637 ( .A(u2__abc_44228_n21260), .B(u2__abc_44228_n21263), .Y(u2__abc_44228_n21264) );
  AND2X2 AND2X2_10638 ( .A(u2__abc_44228_n21265), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_root_291__FF_INPUT) );
  AND2X2 AND2X2_10639 ( .A(u2__abc_44228_n3062_bF_buf1), .B(u2_o_291_), .Y(u2__abc_44228_n21267) );
  AND2X2 AND2X2_1064 ( .A(u2__abc_44228_n3664), .B(u2__abc_44228_n4140), .Y(u2__abc_44228_n4141) );
  AND2X2 AND2X2_10640 ( .A(u2__abc_44228_n21257), .B(u2_o_290_), .Y(u2__abc_44228_n21269) );
  AND2X2 AND2X2_10641 ( .A(u2__abc_44228_n21270), .B(u2__abc_44228_n21268), .Y(u2__abc_44228_n21271) );
  AND2X2 AND2X2_10642 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n6244), .Y(u2__abc_44228_n21273) );
  AND2X2 AND2X2_10643 ( .A(u2__abc_44228_n21274), .B(u2__abc_44228_n2972_bF_buf4), .Y(u2__abc_44228_n21275) );
  AND2X2 AND2X2_10644 ( .A(u2__abc_44228_n21272), .B(u2__abc_44228_n21275), .Y(u2__abc_44228_n21276) );
  AND2X2 AND2X2_10645 ( .A(u2__abc_44228_n21277), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_root_292__FF_INPUT) );
  AND2X2 AND2X2_10646 ( .A(u2__abc_44228_n3062_bF_buf0), .B(u2_o_292_), .Y(u2__abc_44228_n21279) );
  AND2X2 AND2X2_10647 ( .A(u2__abc_44228_n21269), .B(u2_o_291_), .Y(u2__abc_44228_n21281) );
  AND2X2 AND2X2_10648 ( .A(u2__abc_44228_n21282), .B(u2__abc_44228_n21280), .Y(u2__abc_44228_n21283) );
  AND2X2 AND2X2_10649 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n6237), .Y(u2__abc_44228_n21285) );
  AND2X2 AND2X2_1065 ( .A(u2__abc_44228_n4142), .B(u2__abc_44228_n4127), .Y(u2__abc_44228_n4143) );
  AND2X2 AND2X2_10650 ( .A(u2__abc_44228_n21286), .B(u2__abc_44228_n2972_bF_buf3), .Y(u2__abc_44228_n21287) );
  AND2X2 AND2X2_10651 ( .A(u2__abc_44228_n21284), .B(u2__abc_44228_n21287), .Y(u2__abc_44228_n21288) );
  AND2X2 AND2X2_10652 ( .A(u2__abc_44228_n21289), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_root_293__FF_INPUT) );
  AND2X2 AND2X2_10653 ( .A(u2__abc_44228_n3062_bF_buf92), .B(u2_o_293_), .Y(u2__abc_44228_n21291) );
  AND2X2 AND2X2_10654 ( .A(u2__abc_44228_n21281), .B(u2_o_292_), .Y(u2__abc_44228_n21293) );
  AND2X2 AND2X2_10655 ( .A(u2__abc_44228_n21294), .B(u2__abc_44228_n21292), .Y(u2__abc_44228_n21295) );
  AND2X2 AND2X2_10656 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n6230), .Y(u2__abc_44228_n21297) );
  AND2X2 AND2X2_10657 ( .A(u2__abc_44228_n21298), .B(u2__abc_44228_n2972_bF_buf2), .Y(u2__abc_44228_n21299) );
  AND2X2 AND2X2_10658 ( .A(u2__abc_44228_n21296), .B(u2__abc_44228_n21299), .Y(u2__abc_44228_n21300) );
  AND2X2 AND2X2_10659 ( .A(u2__abc_44228_n21301), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_root_294__FF_INPUT) );
  AND2X2 AND2X2_1066 ( .A(u2__abc_44228_n4143), .B(u2__abc_44228_n4121), .Y(u2__abc_44228_n4144) );
  AND2X2 AND2X2_10660 ( .A(u2__abc_44228_n3062_bF_buf91), .B(u2_o_294_), .Y(u2__abc_44228_n21303) );
  AND2X2 AND2X2_10661 ( .A(u2__abc_44228_n21293), .B(u2_o_293_), .Y(u2__abc_44228_n21305) );
  AND2X2 AND2X2_10662 ( .A(u2__abc_44228_n21306), .B(u2__abc_44228_n21304), .Y(u2__abc_44228_n21307) );
  AND2X2 AND2X2_10663 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n6207), .Y(u2__abc_44228_n21309) );
  AND2X2 AND2X2_10664 ( .A(u2__abc_44228_n21310), .B(u2__abc_44228_n2972_bF_buf1), .Y(u2__abc_44228_n21311) );
  AND2X2 AND2X2_10665 ( .A(u2__abc_44228_n21308), .B(u2__abc_44228_n21311), .Y(u2__abc_44228_n21312) );
  AND2X2 AND2X2_10666 ( .A(u2__abc_44228_n21313), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_root_295__FF_INPUT) );
  AND2X2 AND2X2_10667 ( .A(u2__abc_44228_n3062_bF_buf90), .B(u2_o_295_), .Y(u2__abc_44228_n21315) );
  AND2X2 AND2X2_10668 ( .A(u2__abc_44228_n21305), .B(u2_o_294_), .Y(u2__abc_44228_n21317) );
  AND2X2 AND2X2_10669 ( .A(u2__abc_44228_n21318), .B(u2__abc_44228_n21316), .Y(u2__abc_44228_n21319) );
  AND2X2 AND2X2_1067 ( .A(u2__abc_44228_n4146), .B(u2__abc_44228_n4114), .Y(u2__abc_44228_n4147_1) );
  AND2X2 AND2X2_10670 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n6200), .Y(u2__abc_44228_n21321) );
  AND2X2 AND2X2_10671 ( .A(u2__abc_44228_n21322), .B(u2__abc_44228_n2972_bF_buf0), .Y(u2__abc_44228_n21323) );
  AND2X2 AND2X2_10672 ( .A(u2__abc_44228_n21320), .B(u2__abc_44228_n21323), .Y(u2__abc_44228_n21324) );
  AND2X2 AND2X2_10673 ( .A(u2__abc_44228_n21325), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_root_296__FF_INPUT) );
  AND2X2 AND2X2_10674 ( .A(u2__abc_44228_n3062_bF_buf89), .B(u2_o_296_), .Y(u2__abc_44228_n21327) );
  AND2X2 AND2X2_10675 ( .A(u2__abc_44228_n21317), .B(u2_o_295_), .Y(u2__abc_44228_n21329) );
  AND2X2 AND2X2_10676 ( .A(u2__abc_44228_n21330), .B(u2__abc_44228_n21328), .Y(u2__abc_44228_n21331) );
  AND2X2 AND2X2_10677 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n6221), .Y(u2__abc_44228_n21333) );
  AND2X2 AND2X2_10678 ( .A(u2__abc_44228_n21334), .B(u2__abc_44228_n2972_bF_buf107), .Y(u2__abc_44228_n21335) );
  AND2X2 AND2X2_10679 ( .A(u2__abc_44228_n21332), .B(u2__abc_44228_n21335), .Y(u2__abc_44228_n21336) );
  AND2X2 AND2X2_1068 ( .A(u2__abc_44228_n4149), .B(u2__abc_44228_n4110), .Y(u2__abc_44228_n4150) );
  AND2X2 AND2X2_10680 ( .A(u2__abc_44228_n21337), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_root_297__FF_INPUT) );
  AND2X2 AND2X2_10681 ( .A(u2__abc_44228_n3062_bF_buf88), .B(u2_o_297_), .Y(u2__abc_44228_n21339) );
  AND2X2 AND2X2_10682 ( .A(u2__abc_44228_n21329), .B(u2_o_296_), .Y(u2__abc_44228_n21341) );
  AND2X2 AND2X2_10683 ( .A(u2__abc_44228_n21342), .B(u2__abc_44228_n21340), .Y(u2__abc_44228_n21343) );
  AND2X2 AND2X2_10684 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n6214_1), .Y(u2__abc_44228_n21345) );
  AND2X2 AND2X2_10685 ( .A(u2__abc_44228_n21346), .B(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n21347) );
  AND2X2 AND2X2_10686 ( .A(u2__abc_44228_n21344), .B(u2__abc_44228_n21347), .Y(u2__abc_44228_n21348) );
  AND2X2 AND2X2_10687 ( .A(u2__abc_44228_n21349), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_root_298__FF_INPUT) );
  AND2X2 AND2X2_10688 ( .A(u2__abc_44228_n3062_bF_buf87), .B(u2_o_298_), .Y(u2__abc_44228_n21351) );
  AND2X2 AND2X2_10689 ( .A(u2__abc_44228_n21341), .B(u2_o_297_), .Y(u2__abc_44228_n21353) );
  AND2X2 AND2X2_1069 ( .A(u2__abc_44228_n4151), .B(u2__abc_44228_n4101), .Y(u2__abc_44228_n4152) );
  AND2X2 AND2X2_10690 ( .A(u2__abc_44228_n21354), .B(u2__abc_44228_n21352), .Y(u2__abc_44228_n21355) );
  AND2X2 AND2X2_10691 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n6192), .Y(u2__abc_44228_n21357) );
  AND2X2 AND2X2_10692 ( .A(u2__abc_44228_n21358), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n21359) );
  AND2X2 AND2X2_10693 ( .A(u2__abc_44228_n21356), .B(u2__abc_44228_n21359), .Y(u2__abc_44228_n21360) );
  AND2X2 AND2X2_10694 ( .A(u2__abc_44228_n21361), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_root_299__FF_INPUT) );
  AND2X2 AND2X2_10695 ( .A(u2__abc_44228_n3062_bF_buf86), .B(u2_o_299_), .Y(u2__abc_44228_n21363) );
  AND2X2 AND2X2_10696 ( .A(u2__abc_44228_n21353), .B(u2_o_298_), .Y(u2__abc_44228_n21365) );
  AND2X2 AND2X2_10697 ( .A(u2__abc_44228_n21366), .B(u2__abc_44228_n21364), .Y(u2__abc_44228_n21367) );
  AND2X2 AND2X2_10698 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n6185), .Y(u2__abc_44228_n21369) );
  AND2X2 AND2X2_10699 ( .A(u2__abc_44228_n21370), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n21371) );
  AND2X2 AND2X2_107 ( .A(_abc_64468_n921), .B(_abc_64468_n920), .Y(_auto_iopadmap_cc_313_execute_65414_142_) );
  AND2X2 AND2X2_1070 ( .A(u2__abc_44228_n4095), .B(u2__abc_44228_n4152), .Y(u2__abc_44228_n4153) );
  AND2X2 AND2X2_10700 ( .A(u2__abc_44228_n21368), .B(u2__abc_44228_n21371), .Y(u2__abc_44228_n21372) );
  AND2X2 AND2X2_10701 ( .A(u2__abc_44228_n21373), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_root_300__FF_INPUT) );
  AND2X2 AND2X2_10702 ( .A(u2__abc_44228_n3062_bF_buf85), .B(u2_o_300_), .Y(u2__abc_44228_n21375) );
  AND2X2 AND2X2_10703 ( .A(u2__abc_44228_n21365), .B(u2_o_299_), .Y(u2__abc_44228_n21377) );
  AND2X2 AND2X2_10704 ( .A(u2__abc_44228_n21378), .B(u2__abc_44228_n21376), .Y(u2__abc_44228_n21379) );
  AND2X2 AND2X2_10705 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n6178_1), .Y(u2__abc_44228_n21381) );
  AND2X2 AND2X2_10706 ( .A(u2__abc_44228_n21382), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n21383) );
  AND2X2 AND2X2_10707 ( .A(u2__abc_44228_n21380), .B(u2__abc_44228_n21383), .Y(u2__abc_44228_n21384) );
  AND2X2 AND2X2_10708 ( .A(u2__abc_44228_n21385), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_root_301__FF_INPUT) );
  AND2X2 AND2X2_10709 ( .A(u2__abc_44228_n3062_bF_buf84), .B(u2_o_301_), .Y(u2__abc_44228_n21387) );
  AND2X2 AND2X2_1071 ( .A(u2__abc_44228_n4087), .B(u2__abc_44228_n4090_1), .Y(u2__abc_44228_n4154) );
  AND2X2 AND2X2_10710 ( .A(u2__abc_44228_n21377), .B(u2_o_300_), .Y(u2__abc_44228_n21389) );
  AND2X2 AND2X2_10711 ( .A(u2__abc_44228_n21390), .B(u2__abc_44228_n21388), .Y(u2__abc_44228_n21391) );
  AND2X2 AND2X2_10712 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n6171), .Y(u2__abc_44228_n21393) );
  AND2X2 AND2X2_10713 ( .A(u2__abc_44228_n21394), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n21395) );
  AND2X2 AND2X2_10714 ( .A(u2__abc_44228_n21392), .B(u2__abc_44228_n21395), .Y(u2__abc_44228_n21396) );
  AND2X2 AND2X2_10715 ( .A(u2__abc_44228_n21397), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_root_302__FF_INPUT) );
  AND2X2 AND2X2_10716 ( .A(u2__abc_44228_n3062_bF_buf83), .B(u2_o_302_), .Y(u2__abc_44228_n21399) );
  AND2X2 AND2X2_10717 ( .A(u2__abc_44228_n21389), .B(u2_o_301_), .Y(u2__abc_44228_n21401) );
  AND2X2 AND2X2_10718 ( .A(u2__abc_44228_n21402), .B(u2__abc_44228_n21400), .Y(u2__abc_44228_n21403) );
  AND2X2 AND2X2_10719 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n6154), .Y(u2__abc_44228_n21405) );
  AND2X2 AND2X2_1072 ( .A(u2__abc_44228_n4157_1), .B(u2__abc_44228_n4081), .Y(u2__abc_44228_n4158) );
  AND2X2 AND2X2_10720 ( .A(u2__abc_44228_n21406), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n21407) );
  AND2X2 AND2X2_10721 ( .A(u2__abc_44228_n21404), .B(u2__abc_44228_n21407), .Y(u2__abc_44228_n21408) );
  AND2X2 AND2X2_10722 ( .A(u2__abc_44228_n21409), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_root_303__FF_INPUT) );
  AND2X2 AND2X2_10723 ( .A(u2__abc_44228_n3062_bF_buf82), .B(u2_o_303_), .Y(u2__abc_44228_n21411) );
  AND2X2 AND2X2_10724 ( .A(u2__abc_44228_n21401), .B(u2_o_302_), .Y(u2__abc_44228_n21413) );
  AND2X2 AND2X2_10725 ( .A(u2__abc_44228_n21414), .B(u2__abc_44228_n21412), .Y(u2__abc_44228_n21415) );
  AND2X2 AND2X2_10726 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n6160), .Y(u2__abc_44228_n21417) );
  AND2X2 AND2X2_10727 ( .A(u2__abc_44228_n21418), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n21419) );
  AND2X2 AND2X2_10728 ( .A(u2__abc_44228_n21416), .B(u2__abc_44228_n21419), .Y(u2__abc_44228_n21420) );
  AND2X2 AND2X2_10729 ( .A(u2__abc_44228_n21421), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_root_304__FF_INPUT) );
  AND2X2 AND2X2_1073 ( .A(u2__abc_44228_n4159), .B(u2__abc_44228_n4057), .Y(u2__abc_44228_n4160) );
  AND2X2 AND2X2_10730 ( .A(u2__abc_44228_n3062_bF_buf81), .B(u2_o_304_), .Y(u2__abc_44228_n21423) );
  AND2X2 AND2X2_10731 ( .A(u2__abc_44228_n21413), .B(u2_o_303_), .Y(u2__abc_44228_n21425) );
  AND2X2 AND2X2_10732 ( .A(u2__abc_44228_n21426), .B(u2__abc_44228_n21424), .Y(u2__abc_44228_n21427) );
  AND2X2 AND2X2_10733 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n6147), .Y(u2__abc_44228_n21429) );
  AND2X2 AND2X2_10734 ( .A(u2__abc_44228_n21430), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n21431) );
  AND2X2 AND2X2_10735 ( .A(u2__abc_44228_n21428), .B(u2__abc_44228_n21431), .Y(u2__abc_44228_n21432) );
  AND2X2 AND2X2_10736 ( .A(u2__abc_44228_n21433), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_root_305__FF_INPUT) );
  AND2X2 AND2X2_10737 ( .A(u2__abc_44228_n3062_bF_buf80), .B(u2_o_305_), .Y(u2__abc_44228_n21435) );
  AND2X2 AND2X2_10738 ( .A(u2__abc_44228_n21425), .B(u2_o_304_), .Y(u2__abc_44228_n21437) );
  AND2X2 AND2X2_10739 ( .A(u2__abc_44228_n21438), .B(u2__abc_44228_n21436), .Y(u2__abc_44228_n21439) );
  AND2X2 AND2X2_1074 ( .A(u2__abc_44228_n4079), .B(u2__abc_44228_n4160), .Y(u2__abc_44228_n4161) );
  AND2X2 AND2X2_10740 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n6140), .Y(u2__abc_44228_n21441) );
  AND2X2 AND2X2_10741 ( .A(u2__abc_44228_n21442), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n21443) );
  AND2X2 AND2X2_10742 ( .A(u2__abc_44228_n21440), .B(u2__abc_44228_n21443), .Y(u2__abc_44228_n21444) );
  AND2X2 AND2X2_10743 ( .A(u2__abc_44228_n21445), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_root_306__FF_INPUT) );
  AND2X2 AND2X2_10744 ( .A(u2__abc_44228_n3062_bF_buf79), .B(u2_o_306_), .Y(u2__abc_44228_n21447) );
  AND2X2 AND2X2_10745 ( .A(u2__abc_44228_n21437), .B(u2_o_305_), .Y(u2__abc_44228_n21449) );
  AND2X2 AND2X2_10746 ( .A(u2__abc_44228_n21450), .B(u2__abc_44228_n21448), .Y(u2__abc_44228_n21451) );
  AND2X2 AND2X2_10747 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n6125), .Y(u2__abc_44228_n21453) );
  AND2X2 AND2X2_10748 ( .A(u2__abc_44228_n21454), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n21455) );
  AND2X2 AND2X2_10749 ( .A(u2__abc_44228_n21452), .B(u2__abc_44228_n21455), .Y(u2__abc_44228_n21456) );
  AND2X2 AND2X2_1075 ( .A(u2__abc_44228_n4068), .B(u2__abc_44228_n4162), .Y(u2__abc_44228_n4163) );
  AND2X2 AND2X2_10750 ( .A(u2__abc_44228_n21457), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_root_307__FF_INPUT) );
  AND2X2 AND2X2_10751 ( .A(u2__abc_44228_n3062_bF_buf78), .B(u2_o_307_), .Y(u2__abc_44228_n21459) );
  AND2X2 AND2X2_10752 ( .A(u2__abc_44228_n21449), .B(u2_o_306_), .Y(u2__abc_44228_n21461) );
  AND2X2 AND2X2_10753 ( .A(u2__abc_44228_n21462), .B(u2__abc_44228_n21460), .Y(u2__abc_44228_n21463) );
  AND2X2 AND2X2_10754 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n6131), .Y(u2__abc_44228_n21465) );
  AND2X2 AND2X2_10755 ( .A(u2__abc_44228_n21466), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n21467) );
  AND2X2 AND2X2_10756 ( .A(u2__abc_44228_n21464), .B(u2__abc_44228_n21467), .Y(u2__abc_44228_n21468) );
  AND2X2 AND2X2_10757 ( .A(u2__abc_44228_n21469), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_root_308__FF_INPUT) );
  AND2X2 AND2X2_10758 ( .A(u2__abc_44228_n3062_bF_buf77), .B(u2_o_308_), .Y(u2__abc_44228_n21471) );
  AND2X2 AND2X2_10759 ( .A(u2__abc_44228_n21461), .B(u2_o_307_), .Y(u2__abc_44228_n21473) );
  AND2X2 AND2X2_1076 ( .A(u2__abc_44228_n4164), .B(u2__abc_44228_n4071), .Y(u2__abc_44228_n4165) );
  AND2X2 AND2X2_10760 ( .A(u2__abc_44228_n21474), .B(u2__abc_44228_n21472), .Y(u2__abc_44228_n21475) );
  AND2X2 AND2X2_10761 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n6118), .Y(u2__abc_44228_n21477) );
  AND2X2 AND2X2_10762 ( .A(u2__abc_44228_n21478), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n21479) );
  AND2X2 AND2X2_10763 ( .A(u2__abc_44228_n21476), .B(u2__abc_44228_n21479), .Y(u2__abc_44228_n21480) );
  AND2X2 AND2X2_10764 ( .A(u2__abc_44228_n21481), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_root_309__FF_INPUT) );
  AND2X2 AND2X2_10765 ( .A(u2__abc_44228_n3062_bF_buf76), .B(u2_o_309_), .Y(u2__abc_44228_n21483) );
  AND2X2 AND2X2_10766 ( .A(u2__abc_44228_n21473), .B(u2_o_308_), .Y(u2__abc_44228_n21485) );
  AND2X2 AND2X2_10767 ( .A(u2__abc_44228_n21486), .B(u2__abc_44228_n21484), .Y(u2__abc_44228_n21487) );
  AND2X2 AND2X2_10768 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n6111), .Y(u2__abc_44228_n21489) );
  AND2X2 AND2X2_10769 ( .A(u2__abc_44228_n21490), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n21491) );
  AND2X2 AND2X2_1077 ( .A(u2__abc_44228_n4166), .B(u2__abc_44228_n4051), .Y(u2__abc_44228_n4167_1) );
  AND2X2 AND2X2_10770 ( .A(u2__abc_44228_n21488), .B(u2__abc_44228_n21491), .Y(u2__abc_44228_n21492) );
  AND2X2 AND2X2_10771 ( .A(u2__abc_44228_n21493), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_root_310__FF_INPUT) );
  AND2X2 AND2X2_10772 ( .A(u2__abc_44228_n3062_bF_buf75), .B(u2_o_310_), .Y(u2__abc_44228_n21495) );
  AND2X2 AND2X2_10773 ( .A(u2__abc_44228_n21485), .B(u2_o_309_), .Y(u2__abc_44228_n21497) );
  AND2X2 AND2X2_10774 ( .A(u2__abc_44228_n21498), .B(u2__abc_44228_n21496), .Y(u2__abc_44228_n21499) );
  AND2X2 AND2X2_10775 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n6102), .Y(u2__abc_44228_n21501) );
  AND2X2 AND2X2_10776 ( .A(u2__abc_44228_n21502), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n21503) );
  AND2X2 AND2X2_10777 ( .A(u2__abc_44228_n21500), .B(u2__abc_44228_n21503), .Y(u2__abc_44228_n21504) );
  AND2X2 AND2X2_10778 ( .A(u2__abc_44228_n21505), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_root_311__FF_INPUT) );
  AND2X2 AND2X2_10779 ( .A(u2__abc_44228_n3062_bF_buf74), .B(u2_o_311_), .Y(u2__abc_44228_n21507) );
  AND2X2 AND2X2_1078 ( .A(u2__abc_44228_n4028), .B(u2__abc_44228_n4031), .Y(u2__abc_44228_n4168) );
  AND2X2 AND2X2_10780 ( .A(u2__abc_44228_n21497), .B(u2_o_310_), .Y(u2__abc_44228_n21509) );
  AND2X2 AND2X2_10781 ( .A(u2__abc_44228_n21510), .B(u2__abc_44228_n21508), .Y(u2__abc_44228_n21511) );
  AND2X2 AND2X2_10782 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n6095), .Y(u2__abc_44228_n21513) );
  AND2X2 AND2X2_10783 ( .A(u2__abc_44228_n21514), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n21515) );
  AND2X2 AND2X2_10784 ( .A(u2__abc_44228_n21512), .B(u2__abc_44228_n21515), .Y(u2__abc_44228_n21516) );
  AND2X2 AND2X2_10785 ( .A(u2__abc_44228_n21517), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_root_312__FF_INPUT) );
  AND2X2 AND2X2_10786 ( .A(u2__abc_44228_n3062_bF_buf73), .B(u2_o_312_), .Y(u2__abc_44228_n21519) );
  AND2X2 AND2X2_10787 ( .A(u2__abc_44228_n21509), .B(u2_o_311_), .Y(u2__abc_44228_n21521) );
  AND2X2 AND2X2_10788 ( .A(u2__abc_44228_n21522), .B(u2__abc_44228_n21520), .Y(u2__abc_44228_n21523) );
  AND2X2 AND2X2_10789 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n6088), .Y(u2__abc_44228_n21525) );
  AND2X2 AND2X2_1079 ( .A(u2__abc_44228_n4169), .B(u2__abc_44228_n4045), .Y(u2__abc_44228_n4170) );
  AND2X2 AND2X2_10790 ( .A(u2__abc_44228_n21526), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n21527) );
  AND2X2 AND2X2_10791 ( .A(u2__abc_44228_n21524), .B(u2__abc_44228_n21527), .Y(u2__abc_44228_n21528) );
  AND2X2 AND2X2_10792 ( .A(u2__abc_44228_n21529), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_root_313__FF_INPUT) );
  AND2X2 AND2X2_10793 ( .A(u2__abc_44228_n3062_bF_buf72), .B(u2_o_313_), .Y(u2__abc_44228_n21531) );
  AND2X2 AND2X2_10794 ( .A(u2__abc_44228_n21521), .B(u2_o_312_), .Y(u2__abc_44228_n21533) );
  AND2X2 AND2X2_10795 ( .A(u2__abc_44228_n21534), .B(u2__abc_44228_n21532), .Y(u2__abc_44228_n21535) );
  AND2X2 AND2X2_10796 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n6081), .Y(u2__abc_44228_n21537) );
  AND2X2 AND2X2_10797 ( .A(u2__abc_44228_n21538), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n21539) );
  AND2X2 AND2X2_10798 ( .A(u2__abc_44228_n21536), .B(u2__abc_44228_n21539), .Y(u2__abc_44228_n21540) );
  AND2X2 AND2X2_10799 ( .A(u2__abc_44228_n21541), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_root_314__FF_INPUT) );
  AND2X2 AND2X2_108 ( .A(_abc_64468_n924), .B(_abc_64468_n923), .Y(_auto_iopadmap_cc_313_execute_65414_143_) );
  AND2X2 AND2X2_1080 ( .A(u2__abc_44228_n4171), .B(u2__abc_44228_n4048), .Y(u2__abc_44228_n4172) );
  AND2X2 AND2X2_10800 ( .A(u2__abc_44228_n3062_bF_buf71), .B(u2_o_314_), .Y(u2__abc_44228_n21543) );
  AND2X2 AND2X2_10801 ( .A(u2__abc_44228_n21533), .B(u2_o_313_), .Y(u2__abc_44228_n21545) );
  AND2X2 AND2X2_10802 ( .A(u2__abc_44228_n21546), .B(u2__abc_44228_n21544), .Y(u2__abc_44228_n21547) );
  AND2X2 AND2X2_10803 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n6073), .Y(u2__abc_44228_n21549) );
  AND2X2 AND2X2_10804 ( .A(u2__abc_44228_n21550), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n21551) );
  AND2X2 AND2X2_10805 ( .A(u2__abc_44228_n21548), .B(u2__abc_44228_n21551), .Y(u2__abc_44228_n21552) );
  AND2X2 AND2X2_10806 ( .A(u2__abc_44228_n21553), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_root_315__FF_INPUT) );
  AND2X2 AND2X2_10807 ( .A(u2__abc_44228_n3062_bF_buf70), .B(u2_o_315_), .Y(u2__abc_44228_n21555) );
  AND2X2 AND2X2_10808 ( .A(u2__abc_44228_n21545), .B(u2_o_314_), .Y(u2__abc_44228_n21557) );
  AND2X2 AND2X2_10809 ( .A(u2__abc_44228_n21558), .B(u2__abc_44228_n21556), .Y(u2__abc_44228_n21559) );
  AND2X2 AND2X2_1081 ( .A(u2__abc_44228_n4172), .B(u2__abc_44228_n4036), .Y(u2__abc_44228_n4173) );
  AND2X2 AND2X2_10810 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n6066), .Y(u2__abc_44228_n21561) );
  AND2X2 AND2X2_10811 ( .A(u2__abc_44228_n21562), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n21563) );
  AND2X2 AND2X2_10812 ( .A(u2__abc_44228_n21560), .B(u2__abc_44228_n21563), .Y(u2__abc_44228_n21564) );
  AND2X2 AND2X2_10813 ( .A(u2__abc_44228_n21565), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_root_316__FF_INPUT) );
  AND2X2 AND2X2_10814 ( .A(u2__abc_44228_n3062_bF_buf69), .B(u2_o_316_), .Y(u2__abc_44228_n21567) );
  AND2X2 AND2X2_10815 ( .A(u2__abc_44228_n21557), .B(u2_o_315_), .Y(u2__abc_44228_n21569) );
  AND2X2 AND2X2_10816 ( .A(u2__abc_44228_n21570), .B(u2__abc_44228_n21568), .Y(u2__abc_44228_n21571) );
  AND2X2 AND2X2_10817 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n6059_1), .Y(u2__abc_44228_n21573) );
  AND2X2 AND2X2_10818 ( .A(u2__abc_44228_n21574), .B(u2__abc_44228_n2972_bF_buf87), .Y(u2__abc_44228_n21575) );
  AND2X2 AND2X2_10819 ( .A(u2__abc_44228_n21572), .B(u2__abc_44228_n21575), .Y(u2__abc_44228_n21576) );
  AND2X2 AND2X2_1082 ( .A(u2__abc_44228_n4177), .B(u2__abc_44228_n4022), .Y(u2__abc_44228_n4178) );
  AND2X2 AND2X2_10820 ( .A(u2__abc_44228_n21577), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_root_317__FF_INPUT) );
  AND2X2 AND2X2_10821 ( .A(u2__abc_44228_n3062_bF_buf68), .B(u2_o_317_), .Y(u2__abc_44228_n21579) );
  AND2X2 AND2X2_10822 ( .A(u2__abc_44228_n21569), .B(u2_o_316_), .Y(u2__abc_44228_n21581) );
  AND2X2 AND2X2_10823 ( .A(u2__abc_44228_n21582), .B(u2__abc_44228_n21580), .Y(u2__abc_44228_n21583) );
  AND2X2 AND2X2_10824 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n6052), .Y(u2__abc_44228_n21585) );
  AND2X2 AND2X2_10825 ( .A(u2__abc_44228_n21586), .B(u2__abc_44228_n2972_bF_buf86), .Y(u2__abc_44228_n21587) );
  AND2X2 AND2X2_10826 ( .A(u2__abc_44228_n21584), .B(u2__abc_44228_n21587), .Y(u2__abc_44228_n21588) );
  AND2X2 AND2X2_10827 ( .A(u2__abc_44228_n21589), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_root_318__FF_INPUT) );
  AND2X2 AND2X2_10828 ( .A(u2__abc_44228_n3062_bF_buf67), .B(u2_o_318_), .Y(u2__abc_44228_n21591) );
  AND2X2 AND2X2_10829 ( .A(u2__abc_44228_n21581), .B(u2_o_317_), .Y(u2__abc_44228_n21593) );
  AND2X2 AND2X2_1083 ( .A(u2__abc_44228_n4179), .B(u2__abc_44228_n4014), .Y(u2__abc_44228_n4180) );
  AND2X2 AND2X2_10830 ( .A(u2__abc_44228_n21594), .B(u2__abc_44228_n21592), .Y(u2__abc_44228_n21595) );
  AND2X2 AND2X2_10831 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n6033), .Y(u2__abc_44228_n21597) );
  AND2X2 AND2X2_10832 ( .A(u2__abc_44228_n21598), .B(u2__abc_44228_n2972_bF_buf85), .Y(u2__abc_44228_n21599) );
  AND2X2 AND2X2_10833 ( .A(u2__abc_44228_n21596), .B(u2__abc_44228_n21599), .Y(u2__abc_44228_n21600) );
  AND2X2 AND2X2_10834 ( .A(u2__abc_44228_n21601), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_root_319__FF_INPUT) );
  AND2X2 AND2X2_10835 ( .A(u2__abc_44228_n3062_bF_buf66), .B(u2_o_319_), .Y(u2__abc_44228_n21603) );
  AND2X2 AND2X2_10836 ( .A(u2__abc_44228_n21593), .B(u2_o_318_), .Y(u2__abc_44228_n21605) );
  AND2X2 AND2X2_10837 ( .A(u2__abc_44228_n21606), .B(u2__abc_44228_n21604), .Y(u2__abc_44228_n21607) );
  AND2X2 AND2X2_10838 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n6039), .Y(u2__abc_44228_n21609) );
  AND2X2 AND2X2_10839 ( .A(u2__abc_44228_n21610), .B(u2__abc_44228_n2972_bF_buf84), .Y(u2__abc_44228_n21611) );
  AND2X2 AND2X2_1084 ( .A(u2__abc_44228_n4181), .B(u2__abc_44228_n4017), .Y(u2__abc_44228_n4182) );
  AND2X2 AND2X2_10840 ( .A(u2__abc_44228_n21608), .B(u2__abc_44228_n21611), .Y(u2__abc_44228_n21612) );
  AND2X2 AND2X2_10841 ( .A(u2__abc_44228_n21613), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_root_320__FF_INPUT) );
  AND2X2 AND2X2_10842 ( .A(u2__abc_44228_n3062_bF_buf65), .B(u2_o_320_), .Y(u2__abc_44228_n21615) );
  AND2X2 AND2X2_10843 ( .A(u2__abc_44228_n21605), .B(u2_o_319_), .Y(u2__abc_44228_n21617) );
  AND2X2 AND2X2_10844 ( .A(u2__abc_44228_n21618), .B(u2__abc_44228_n21616), .Y(u2__abc_44228_n21619) );
  AND2X2 AND2X2_10845 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n6026), .Y(u2__abc_44228_n21621) );
  AND2X2 AND2X2_10846 ( .A(u2__abc_44228_n21622), .B(u2__abc_44228_n2972_bF_buf83), .Y(u2__abc_44228_n21623) );
  AND2X2 AND2X2_10847 ( .A(u2__abc_44228_n21620), .B(u2__abc_44228_n21623), .Y(u2__abc_44228_n21624) );
  AND2X2 AND2X2_10848 ( .A(u2__abc_44228_n21625), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_root_321__FF_INPUT) );
  AND2X2 AND2X2_10849 ( .A(u2__abc_44228_n3062_bF_buf64), .B(u2_o_321_), .Y(u2__abc_44228_n21627) );
  AND2X2 AND2X2_1085 ( .A(u2__abc_44228_n4182), .B(u2__abc_44228_n4005_1), .Y(u2__abc_44228_n4183) );
  AND2X2 AND2X2_10850 ( .A(u2__abc_44228_n21617), .B(u2_o_320_), .Y(u2__abc_44228_n21629) );
  AND2X2 AND2X2_10851 ( .A(u2__abc_44228_n21630), .B(u2__abc_44228_n21628), .Y(u2__abc_44228_n21631) );
  AND2X2 AND2X2_10852 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n6019), .Y(u2__abc_44228_n21633) );
  AND2X2 AND2X2_10853 ( .A(u2__abc_44228_n21634), .B(u2__abc_44228_n2972_bF_buf82), .Y(u2__abc_44228_n21635) );
  AND2X2 AND2X2_10854 ( .A(u2__abc_44228_n21632), .B(u2__abc_44228_n21635), .Y(u2__abc_44228_n21636) );
  AND2X2 AND2X2_10855 ( .A(u2__abc_44228_n21637), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_root_322__FF_INPUT) );
  AND2X2 AND2X2_10856 ( .A(u2__abc_44228_n3062_bF_buf63), .B(u2_o_322_), .Y(u2__abc_44228_n21639) );
  AND2X2 AND2X2_10857 ( .A(u2__abc_44228_n21629), .B(u2_o_321_), .Y(u2__abc_44228_n21641) );
  AND2X2 AND2X2_10858 ( .A(u2__abc_44228_n21642), .B(u2__abc_44228_n21640), .Y(u2__abc_44228_n21643) );
  AND2X2 AND2X2_10859 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n6004), .Y(u2__abc_44228_n21645) );
  AND2X2 AND2X2_1086 ( .A(u2__abc_44228_n3997), .B(u2__abc_44228_n4000), .Y(u2__abc_44228_n4184) );
  AND2X2 AND2X2_10860 ( .A(u2__abc_44228_n21646), .B(u2__abc_44228_n2972_bF_buf81), .Y(u2__abc_44228_n21647) );
  AND2X2 AND2X2_10861 ( .A(u2__abc_44228_n21644), .B(u2__abc_44228_n21647), .Y(u2__abc_44228_n21648) );
  AND2X2 AND2X2_10862 ( .A(u2__abc_44228_n21649), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_root_323__FF_INPUT) );
  AND2X2 AND2X2_10863 ( .A(u2__abc_44228_n3062_bF_buf62), .B(u2_o_323_), .Y(u2__abc_44228_n21651) );
  AND2X2 AND2X2_10864 ( .A(u2__abc_44228_n21641), .B(u2_o_322_), .Y(u2__abc_44228_n21653) );
  AND2X2 AND2X2_10865 ( .A(u2__abc_44228_n21654), .B(u2__abc_44228_n21652), .Y(u2__abc_44228_n21655) );
  AND2X2 AND2X2_10866 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n6010), .Y(u2__abc_44228_n21657) );
  AND2X2 AND2X2_10867 ( .A(u2__abc_44228_n21658), .B(u2__abc_44228_n2972_bF_buf80), .Y(u2__abc_44228_n21659) );
  AND2X2 AND2X2_10868 ( .A(u2__abc_44228_n21656), .B(u2__abc_44228_n21659), .Y(u2__abc_44228_n21660) );
  AND2X2 AND2X2_10869 ( .A(u2__abc_44228_n21661), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_root_324__FF_INPUT) );
  AND2X2 AND2X2_1087 ( .A(u2__abc_44228_n4186), .B(u2__abc_44228_n3991), .Y(u2__abc_44228_n4187) );
  AND2X2 AND2X2_10870 ( .A(u2__abc_44228_n3062_bF_buf61), .B(u2_o_324_), .Y(u2__abc_44228_n21663) );
  AND2X2 AND2X2_10871 ( .A(u2__abc_44228_n21653), .B(u2_o_323_), .Y(u2__abc_44228_n21665) );
  AND2X2 AND2X2_10872 ( .A(u2__abc_44228_n21666), .B(u2__abc_44228_n21664), .Y(u2__abc_44228_n21667) );
  AND2X2 AND2X2_10873 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n5997), .Y(u2__abc_44228_n21669) );
  AND2X2 AND2X2_10874 ( .A(u2__abc_44228_n21670), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n21671) );
  AND2X2 AND2X2_10875 ( .A(u2__abc_44228_n21668), .B(u2__abc_44228_n21671), .Y(u2__abc_44228_n21672) );
  AND2X2 AND2X2_10876 ( .A(u2__abc_44228_n21673), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_root_325__FF_INPUT) );
  AND2X2 AND2X2_10877 ( .A(u2__abc_44228_n3062_bF_buf60), .B(u2_o_325_), .Y(u2__abc_44228_n21675) );
  AND2X2 AND2X2_10878 ( .A(u2__abc_44228_n21665), .B(u2_o_324_), .Y(u2__abc_44228_n21677) );
  AND2X2 AND2X2_10879 ( .A(u2__abc_44228_n21678), .B(u2__abc_44228_n21676), .Y(u2__abc_44228_n21679) );
  AND2X2 AND2X2_1088 ( .A(u2__abc_44228_n4189), .B(u2__abc_44228_n3985), .Y(u2__abc_44228_n4190) );
  AND2X2 AND2X2_10880 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n5990), .Y(u2__abc_44228_n21681) );
  AND2X2 AND2X2_10881 ( .A(u2__abc_44228_n21682), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n21683) );
  AND2X2 AND2X2_10882 ( .A(u2__abc_44228_n21680), .B(u2__abc_44228_n21683), .Y(u2__abc_44228_n21684) );
  AND2X2 AND2X2_10883 ( .A(u2__abc_44228_n21685), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_root_326__FF_INPUT) );
  AND2X2 AND2X2_10884 ( .A(u2__abc_44228_n3062_bF_buf59), .B(u2_o_326_), .Y(u2__abc_44228_n21687) );
  AND2X2 AND2X2_10885 ( .A(u2__abc_44228_n21677), .B(u2_o_325_), .Y(u2__abc_44228_n21689) );
  AND2X2 AND2X2_10886 ( .A(u2__abc_44228_n21690), .B(u2__abc_44228_n21688), .Y(u2__abc_44228_n21691) );
  AND2X2 AND2X2_10887 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n5981), .Y(u2__abc_44228_n21693) );
  AND2X2 AND2X2_10888 ( .A(u2__abc_44228_n21694), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n21695) );
  AND2X2 AND2X2_10889 ( .A(u2__abc_44228_n21692), .B(u2__abc_44228_n21695), .Y(u2__abc_44228_n21696) );
  AND2X2 AND2X2_1089 ( .A(u2__abc_44228_n4191), .B(u2__abc_44228_n3976_1), .Y(u2__abc_44228_n4192) );
  AND2X2 AND2X2_10890 ( .A(u2__abc_44228_n21697), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_root_327__FF_INPUT) );
  AND2X2 AND2X2_10891 ( .A(u2__abc_44228_n3062_bF_buf58), .B(u2_o_327_), .Y(u2__abc_44228_n21699) );
  AND2X2 AND2X2_10892 ( .A(u2__abc_44228_n21689), .B(u2_o_326_), .Y(u2__abc_44228_n21701) );
  AND2X2 AND2X2_10893 ( .A(u2__abc_44228_n21702), .B(u2__abc_44228_n21700), .Y(u2__abc_44228_n21703) );
  AND2X2 AND2X2_10894 ( .A(u2__abc_44228_n2983_bF_buf104), .B(u2__abc_44228_n5974), .Y(u2__abc_44228_n21705) );
  AND2X2 AND2X2_10895 ( .A(u2__abc_44228_n21706), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n21707) );
  AND2X2 AND2X2_10896 ( .A(u2__abc_44228_n21704), .B(u2__abc_44228_n21707), .Y(u2__abc_44228_n21708) );
  AND2X2 AND2X2_10897 ( .A(u2__abc_44228_n21709), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_root_328__FF_INPUT) );
  AND2X2 AND2X2_10898 ( .A(u2__abc_44228_n3062_bF_buf57), .B(u2_o_328_), .Y(u2__abc_44228_n21711) );
  AND2X2 AND2X2_10899 ( .A(u2__abc_44228_n21701), .B(u2_o_327_), .Y(u2__abc_44228_n21713) );
  AND2X2 AND2X2_109 ( .A(_abc_64468_n927), .B(_abc_64468_n926), .Y(_auto_iopadmap_cc_313_execute_65414_144_) );
  AND2X2 AND2X2_1090 ( .A(u2__abc_44228_n3968), .B(u2__abc_44228_n3971), .Y(u2__abc_44228_n4193) );
  AND2X2 AND2X2_10900 ( .A(u2__abc_44228_n21714), .B(u2__abc_44228_n21712), .Y(u2__abc_44228_n21715) );
  AND2X2 AND2X2_10901 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n5967), .Y(u2__abc_44228_n21717) );
  AND2X2 AND2X2_10902 ( .A(u2__abc_44228_n21718), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n21719) );
  AND2X2 AND2X2_10903 ( .A(u2__abc_44228_n21716), .B(u2__abc_44228_n21719), .Y(u2__abc_44228_n21720) );
  AND2X2 AND2X2_10904 ( .A(u2__abc_44228_n21721), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_root_329__FF_INPUT) );
  AND2X2 AND2X2_10905 ( .A(u2__abc_44228_n3062_bF_buf56), .B(u2_o_329_), .Y(u2__abc_44228_n21723) );
  AND2X2 AND2X2_10906 ( .A(u2__abc_44228_n21713), .B(u2_o_328_), .Y(u2__abc_44228_n21725) );
  AND2X2 AND2X2_10907 ( .A(u2__abc_44228_n21726), .B(u2__abc_44228_n21724), .Y(u2__abc_44228_n21727) );
  AND2X2 AND2X2_10908 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n5960), .Y(u2__abc_44228_n21729) );
  AND2X2 AND2X2_10909 ( .A(u2__abc_44228_n21730), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n21731) );
  AND2X2 AND2X2_1091 ( .A(u2__abc_44228_n4196), .B(u2__abc_44228_n3962), .Y(u2__abc_44228_n4197) );
  AND2X2 AND2X2_10910 ( .A(u2__abc_44228_n21728), .B(u2__abc_44228_n21731), .Y(u2__abc_44228_n21732) );
  AND2X2 AND2X2_10911 ( .A(u2__abc_44228_n21733), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_root_330__FF_INPUT) );
  AND2X2 AND2X2_10912 ( .A(u2__abc_44228_n3062_bF_buf55), .B(u2_o_330_), .Y(u2__abc_44228_n21735) );
  AND2X2 AND2X2_10913 ( .A(u2__abc_44228_n21725), .B(u2_o_329_), .Y(u2__abc_44228_n21737) );
  AND2X2 AND2X2_10914 ( .A(u2__abc_44228_n21738), .B(u2__abc_44228_n21736), .Y(u2__abc_44228_n21739) );
  AND2X2 AND2X2_10915 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n5952), .Y(u2__abc_44228_n21741) );
  AND2X2 AND2X2_10916 ( .A(u2__abc_44228_n21742), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n21743) );
  AND2X2 AND2X2_10917 ( .A(u2__abc_44228_n21740), .B(u2__abc_44228_n21743), .Y(u2__abc_44228_n21744) );
  AND2X2 AND2X2_10918 ( .A(u2__abc_44228_n21745), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_root_331__FF_INPUT) );
  AND2X2 AND2X2_10919 ( .A(u2__abc_44228_n3062_bF_buf54), .B(u2_o_331_), .Y(u2__abc_44228_n21747) );
  AND2X2 AND2X2_1092 ( .A(u2__abc_44228_n4198), .B(u2__abc_44228_n3955), .Y(u2__abc_44228_n4199) );
  AND2X2 AND2X2_10920 ( .A(u2__abc_44228_n21737), .B(u2_o_330_), .Y(u2__abc_44228_n21749) );
  AND2X2 AND2X2_10921 ( .A(u2__abc_44228_n21750), .B(u2__abc_44228_n21748), .Y(u2__abc_44228_n21751) );
  AND2X2 AND2X2_10922 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n5945), .Y(u2__abc_44228_n21753) );
  AND2X2 AND2X2_10923 ( .A(u2__abc_44228_n21754), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n21755) );
  AND2X2 AND2X2_10924 ( .A(u2__abc_44228_n21752), .B(u2__abc_44228_n21755), .Y(u2__abc_44228_n21756) );
  AND2X2 AND2X2_10925 ( .A(u2__abc_44228_n21757), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_root_332__FF_INPUT) );
  AND2X2 AND2X2_10926 ( .A(u2__abc_44228_n3062_bF_buf53), .B(u2_o_332_), .Y(u2__abc_44228_n21759) );
  AND2X2 AND2X2_10927 ( .A(u2__abc_44228_n21749), .B(u2_o_331_), .Y(u2__abc_44228_n21761) );
  AND2X2 AND2X2_10928 ( .A(u2__abc_44228_n21762), .B(u2__abc_44228_n21760), .Y(u2__abc_44228_n21763) );
  AND2X2 AND2X2_10929 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n5938_1), .Y(u2__abc_44228_n21765) );
  AND2X2 AND2X2_1093 ( .A(u2__abc_44228_n4200), .B(u2__abc_44228_n3958_1), .Y(u2__abc_44228_n4201) );
  AND2X2 AND2X2_10930 ( .A(u2__abc_44228_n21766), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n21767) );
  AND2X2 AND2X2_10931 ( .A(u2__abc_44228_n21764), .B(u2__abc_44228_n21767), .Y(u2__abc_44228_n21768) );
  AND2X2 AND2X2_10932 ( .A(u2__abc_44228_n21769), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_root_333__FF_INPUT) );
  AND2X2 AND2X2_10933 ( .A(u2__abc_44228_n3062_bF_buf52), .B(u2_o_333_), .Y(u2__abc_44228_n21771) );
  AND2X2 AND2X2_10934 ( .A(u2__abc_44228_n21761), .B(u2_o_332_), .Y(u2__abc_44228_n21773) );
  AND2X2 AND2X2_10935 ( .A(u2__abc_44228_n21774), .B(u2__abc_44228_n21772), .Y(u2__abc_44228_n21775) );
  AND2X2 AND2X2_10936 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n5931), .Y(u2__abc_44228_n21777) );
  AND2X2 AND2X2_10937 ( .A(u2__abc_44228_n21778), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n21779) );
  AND2X2 AND2X2_10938 ( .A(u2__abc_44228_n21776), .B(u2__abc_44228_n21779), .Y(u2__abc_44228_n21780) );
  AND2X2 AND2X2_10939 ( .A(u2__abc_44228_n21781), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_root_334__FF_INPUT) );
  AND2X2 AND2X2_1094 ( .A(u2__abc_44228_n4201), .B(u2__abc_44228_n3946), .Y(u2__abc_44228_n4202) );
  AND2X2 AND2X2_10940 ( .A(u2__abc_44228_n3062_bF_buf51), .B(u2_o_334_), .Y(u2__abc_44228_n21783) );
  AND2X2 AND2X2_10941 ( .A(u2__abc_44228_n21773), .B(u2_o_333_), .Y(u2__abc_44228_n21785) );
  AND2X2 AND2X2_10942 ( .A(u2__abc_44228_n21786), .B(u2__abc_44228_n21784), .Y(u2__abc_44228_n21787) );
  AND2X2 AND2X2_10943 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n5921), .Y(u2__abc_44228_n21789) );
  AND2X2 AND2X2_10944 ( .A(u2__abc_44228_n21790), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n21791) );
  AND2X2 AND2X2_10945 ( .A(u2__abc_44228_n21788), .B(u2__abc_44228_n21791), .Y(u2__abc_44228_n21792) );
  AND2X2 AND2X2_10946 ( .A(u2__abc_44228_n21793), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_root_335__FF_INPUT) );
  AND2X2 AND2X2_10947 ( .A(u2__abc_44228_n3062_bF_buf50), .B(u2_o_335_), .Y(u2__abc_44228_n21795) );
  AND2X2 AND2X2_10948 ( .A(u2__abc_44228_n21785), .B(u2_o_334_), .Y(u2__abc_44228_n21797) );
  AND2X2 AND2X2_10949 ( .A(u2__abc_44228_n21798), .B(u2__abc_44228_n21796), .Y(u2__abc_44228_n21799) );
  AND2X2 AND2X2_1095 ( .A(u2__abc_44228_n3938), .B(u2__abc_44228_n3941), .Y(u2__abc_44228_n4203) );
  AND2X2 AND2X2_10950 ( .A(u2__abc_44228_n2983_bF_buf88), .B(u2__abc_44228_n5914), .Y(u2__abc_44228_n21801) );
  AND2X2 AND2X2_10951 ( .A(u2__abc_44228_n21802), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n21803) );
  AND2X2 AND2X2_10952 ( .A(u2__abc_44228_n21800), .B(u2__abc_44228_n21803), .Y(u2__abc_44228_n21804) );
  AND2X2 AND2X2_10953 ( .A(u2__abc_44228_n21805), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_root_336__FF_INPUT) );
  AND2X2 AND2X2_10954 ( .A(u2__abc_44228_n3062_bF_buf49), .B(u2_o_336_), .Y(u2__abc_44228_n21807) );
  AND2X2 AND2X2_10955 ( .A(u2__abc_44228_n21797), .B(u2_o_335_), .Y(u2__abc_44228_n21809) );
  AND2X2 AND2X2_10956 ( .A(u2__abc_44228_n21810), .B(u2__abc_44228_n21808), .Y(u2__abc_44228_n21811) );
  AND2X2 AND2X2_10957 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n5907), .Y(u2__abc_44228_n21813) );
  AND2X2 AND2X2_10958 ( .A(u2__abc_44228_n21814), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n21815) );
  AND2X2 AND2X2_10959 ( .A(u2__abc_44228_n21812), .B(u2__abc_44228_n21815), .Y(u2__abc_44228_n21816) );
  AND2X2 AND2X2_1096 ( .A(u2__abc_44228_n4205_1), .B(u2__abc_44228_n3932), .Y(u2__abc_44228_n4206) );
  AND2X2 AND2X2_10960 ( .A(u2__abc_44228_n21817), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_root_337__FF_INPUT) );
  AND2X2 AND2X2_10961 ( .A(u2__abc_44228_n3062_bF_buf48), .B(u2_o_337_), .Y(u2__abc_44228_n21819) );
  AND2X2 AND2X2_10962 ( .A(u2__abc_44228_n21809), .B(u2_o_336_), .Y(u2__abc_44228_n21821) );
  AND2X2 AND2X2_10963 ( .A(u2__abc_44228_n21822), .B(u2__abc_44228_n21820), .Y(u2__abc_44228_n21823) );
  AND2X2 AND2X2_10964 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n5900), .Y(u2__abc_44228_n21825) );
  AND2X2 AND2X2_10965 ( .A(u2__abc_44228_n21826), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n21827) );
  AND2X2 AND2X2_10966 ( .A(u2__abc_44228_n21824), .B(u2__abc_44228_n21827), .Y(u2__abc_44228_n21828) );
  AND2X2 AND2X2_10967 ( .A(u2__abc_44228_n21829), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_root_338__FF_INPUT) );
  AND2X2 AND2X2_10968 ( .A(u2__abc_44228_n3062_bF_buf47), .B(u2_o_338_), .Y(u2__abc_44228_n21831) );
  AND2X2 AND2X2_10969 ( .A(u2__abc_44228_n21821), .B(u2_o_337_), .Y(u2__abc_44228_n21833) );
  AND2X2 AND2X2_1097 ( .A(u2__abc_44228_n4207), .B(u2__abc_44228_n3926), .Y(u2__abc_44228_n4208) );
  AND2X2 AND2X2_10970 ( .A(u2__abc_44228_n21834), .B(u2__abc_44228_n21832), .Y(u2__abc_44228_n21835) );
  AND2X2 AND2X2_10971 ( .A(u2__abc_44228_n2983_bF_buf82), .B(u2__abc_44228_n5885), .Y(u2__abc_44228_n21837) );
  AND2X2 AND2X2_10972 ( .A(u2__abc_44228_n21838), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n21839) );
  AND2X2 AND2X2_10973 ( .A(u2__abc_44228_n21836), .B(u2__abc_44228_n21839), .Y(u2__abc_44228_n21840) );
  AND2X2 AND2X2_10974 ( .A(u2__abc_44228_n21841), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_root_339__FF_INPUT) );
  AND2X2 AND2X2_10975 ( .A(u2__abc_44228_n3062_bF_buf46), .B(u2_o_339_), .Y(u2__abc_44228_n21843) );
  AND2X2 AND2X2_10976 ( .A(u2__abc_44228_n21833), .B(u2_o_338_), .Y(u2__abc_44228_n21845) );
  AND2X2 AND2X2_10977 ( .A(u2__abc_44228_n21846), .B(u2__abc_44228_n21844), .Y(u2__abc_44228_n21847) );
  AND2X2 AND2X2_10978 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n5891), .Y(u2__abc_44228_n21849) );
  AND2X2 AND2X2_10979 ( .A(u2__abc_44228_n21850), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n21851) );
  AND2X2 AND2X2_1098 ( .A(u2__abc_44228_n4209), .B(u2__abc_44228_n3929), .Y(u2__abc_44228_n4210) );
  AND2X2 AND2X2_10980 ( .A(u2__abc_44228_n21848), .B(u2__abc_44228_n21851), .Y(u2__abc_44228_n21852) );
  AND2X2 AND2X2_10981 ( .A(u2__abc_44228_n21853), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_root_340__FF_INPUT) );
  AND2X2 AND2X2_10982 ( .A(u2__abc_44228_n3062_bF_buf45), .B(u2_o_340_), .Y(u2__abc_44228_n21855) );
  AND2X2 AND2X2_10983 ( .A(u2__abc_44228_n21845), .B(u2_o_339_), .Y(u2__abc_44228_n21857) );
  AND2X2 AND2X2_10984 ( .A(u2__abc_44228_n21858), .B(u2__abc_44228_n21856), .Y(u2__abc_44228_n21859) );
  AND2X2 AND2X2_10985 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n5878), .Y(u2__abc_44228_n21861) );
  AND2X2 AND2X2_10986 ( .A(u2__abc_44228_n21862), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n21863) );
  AND2X2 AND2X2_10987 ( .A(u2__abc_44228_n21860), .B(u2__abc_44228_n21863), .Y(u2__abc_44228_n21864) );
  AND2X2 AND2X2_10988 ( .A(u2__abc_44228_n21865), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_root_341__FF_INPUT) );
  AND2X2 AND2X2_10989 ( .A(u2__abc_44228_n3062_bF_buf44), .B(u2_o_341_), .Y(u2__abc_44228_n21867) );
  AND2X2 AND2X2_1099 ( .A(u2__abc_44228_n4210), .B(u2__abc_44228_n3917), .Y(u2__abc_44228_n4211) );
  AND2X2 AND2X2_10990 ( .A(u2__abc_44228_n21857), .B(u2_o_340_), .Y(u2__abc_44228_n21869) );
  AND2X2 AND2X2_10991 ( .A(u2__abc_44228_n21870), .B(u2__abc_44228_n21868), .Y(u2__abc_44228_n21871) );
  AND2X2 AND2X2_10992 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n5871), .Y(u2__abc_44228_n21873) );
  AND2X2 AND2X2_10993 ( .A(u2__abc_44228_n21874), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n21875) );
  AND2X2 AND2X2_10994 ( .A(u2__abc_44228_n21872), .B(u2__abc_44228_n21875), .Y(u2__abc_44228_n21876) );
  AND2X2 AND2X2_10995 ( .A(u2__abc_44228_n21877), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_root_342__FF_INPUT) );
  AND2X2 AND2X2_10996 ( .A(u2__abc_44228_n3062_bF_buf43), .B(u2_o_342_), .Y(u2__abc_44228_n21879) );
  AND2X2 AND2X2_10997 ( .A(u2__abc_44228_n21869), .B(u2_o_341_), .Y(u2__abc_44228_n21881) );
  AND2X2 AND2X2_10998 ( .A(u2__abc_44228_n21882), .B(u2__abc_44228_n21880), .Y(u2__abc_44228_n21883) );
  AND2X2 AND2X2_10999 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n5848), .Y(u2__abc_44228_n21885) );
  AND2X2 AND2X2_11 ( .A(_abc_64468_n753_bF_buf3), .B(sqrto_10_), .Y(_auto_iopadmap_cc_313_execute_65414_46_) );
  AND2X2 AND2X2_110 ( .A(_abc_64468_n930), .B(_abc_64468_n929), .Y(_auto_iopadmap_cc_313_execute_65414_145_) );
  AND2X2 AND2X2_1100 ( .A(u2__abc_44228_n3909), .B(u2__abc_44228_n3912_1), .Y(u2__abc_44228_n4212) );
  AND2X2 AND2X2_11000 ( .A(u2__abc_44228_n21886), .B(u2__abc_44228_n2972_bF_buf61), .Y(u2__abc_44228_n21887) );
  AND2X2 AND2X2_11001 ( .A(u2__abc_44228_n21884), .B(u2__abc_44228_n21887), .Y(u2__abc_44228_n21888) );
  AND2X2 AND2X2_11002 ( .A(u2__abc_44228_n21889), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_root_343__FF_INPUT) );
  AND2X2 AND2X2_11003 ( .A(u2__abc_44228_n3062_bF_buf42), .B(u2_o_343_), .Y(u2__abc_44228_n21891) );
  AND2X2 AND2X2_11004 ( .A(u2__abc_44228_n21881), .B(u2_o_342_), .Y(u2__abc_44228_n21893) );
  AND2X2 AND2X2_11005 ( .A(u2__abc_44228_n21894), .B(u2__abc_44228_n21892), .Y(u2__abc_44228_n21895) );
  AND2X2 AND2X2_11006 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n5841), .Y(u2__abc_44228_n21897) );
  AND2X2 AND2X2_11007 ( .A(u2__abc_44228_n21898), .B(u2__abc_44228_n2972_bF_buf60), .Y(u2__abc_44228_n21899) );
  AND2X2 AND2X2_11008 ( .A(u2__abc_44228_n21896), .B(u2__abc_44228_n21899), .Y(u2__abc_44228_n21900) );
  AND2X2 AND2X2_11009 ( .A(u2__abc_44228_n21901), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_root_344__FF_INPUT) );
  AND2X2 AND2X2_1101 ( .A(u2__abc_44228_n4217), .B(u2__abc_44228_n3903_1), .Y(u2__abc_44228_n4218) );
  AND2X2 AND2X2_11010 ( .A(u2__abc_44228_n3062_bF_buf41), .B(u2_o_344_), .Y(u2__abc_44228_n21903) );
  AND2X2 AND2X2_11011 ( .A(u2__abc_44228_n21893), .B(u2_o_343_), .Y(u2__abc_44228_n21905) );
  AND2X2 AND2X2_11012 ( .A(u2__abc_44228_n21906), .B(u2__abc_44228_n21904), .Y(u2__abc_44228_n21907) );
  AND2X2 AND2X2_11013 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n5862), .Y(u2__abc_44228_n21909) );
  AND2X2 AND2X2_11014 ( .A(u2__abc_44228_n21910), .B(u2__abc_44228_n2972_bF_buf59), .Y(u2__abc_44228_n21911) );
  AND2X2 AND2X2_11015 ( .A(u2__abc_44228_n21908), .B(u2__abc_44228_n21911), .Y(u2__abc_44228_n21912) );
  AND2X2 AND2X2_11016 ( .A(u2__abc_44228_n21913), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_root_345__FF_INPUT) );
  AND2X2 AND2X2_11017 ( .A(u2__abc_44228_n3062_bF_buf40), .B(u2_o_345_), .Y(u2__abc_44228_n21915) );
  AND2X2 AND2X2_11018 ( .A(u2__abc_44228_n21905), .B(u2_o_344_), .Y(u2__abc_44228_n21917) );
  AND2X2 AND2X2_11019 ( .A(u2__abc_44228_n21918), .B(u2__abc_44228_n21916), .Y(u2__abc_44228_n21919) );
  AND2X2 AND2X2_1102 ( .A(u2__abc_44228_n4219), .B(u2__abc_44228_n3894), .Y(u2__abc_44228_n4220) );
  AND2X2 AND2X2_11020 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n5855), .Y(u2__abc_44228_n21921) );
  AND2X2 AND2X2_11021 ( .A(u2__abc_44228_n21922), .B(u2__abc_44228_n2972_bF_buf58), .Y(u2__abc_44228_n21923) );
  AND2X2 AND2X2_11022 ( .A(u2__abc_44228_n21920), .B(u2__abc_44228_n21923), .Y(u2__abc_44228_n21924) );
  AND2X2 AND2X2_11023 ( .A(u2__abc_44228_n21925), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_root_346__FF_INPUT) );
  AND2X2 AND2X2_11024 ( .A(u2__abc_44228_n3062_bF_buf39), .B(u2_o_346_), .Y(u2__abc_44228_n21927) );
  AND2X2 AND2X2_11025 ( .A(u2__abc_44228_n21917), .B(u2_o_345_), .Y(u2__abc_44228_n21929) );
  AND2X2 AND2X2_11026 ( .A(u2__abc_44228_n21930), .B(u2__abc_44228_n21928), .Y(u2__abc_44228_n21931) );
  AND2X2 AND2X2_11027 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n5826), .Y(u2__abc_44228_n21933) );
  AND2X2 AND2X2_11028 ( .A(u2__abc_44228_n21934), .B(u2__abc_44228_n2972_bF_buf57), .Y(u2__abc_44228_n21935) );
  AND2X2 AND2X2_11029 ( .A(u2__abc_44228_n21932), .B(u2__abc_44228_n21935), .Y(u2__abc_44228_n21936) );
  AND2X2 AND2X2_1103 ( .A(u2__abc_44228_n4221), .B(u2__abc_44228_n3897), .Y(u2__abc_44228_n4222) );
  AND2X2 AND2X2_11030 ( .A(u2__abc_44228_n21937), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_root_347__FF_INPUT) );
  AND2X2 AND2X2_11031 ( .A(u2__abc_44228_n3062_bF_buf38), .B(u2_o_347_), .Y(u2__abc_44228_n21939) );
  AND2X2 AND2X2_11032 ( .A(u2__abc_44228_n21929), .B(u2_o_346_), .Y(u2__abc_44228_n21941) );
  AND2X2 AND2X2_11033 ( .A(u2__abc_44228_n21942), .B(u2__abc_44228_n21940), .Y(u2__abc_44228_n21943) );
  AND2X2 AND2X2_11034 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n5832), .Y(u2__abc_44228_n21945) );
  AND2X2 AND2X2_11035 ( .A(u2__abc_44228_n21946), .B(u2__abc_44228_n2972_bF_buf56), .Y(u2__abc_44228_n21947) );
  AND2X2 AND2X2_11036 ( .A(u2__abc_44228_n21944), .B(u2__abc_44228_n21947), .Y(u2__abc_44228_n21948) );
  AND2X2 AND2X2_11037 ( .A(u2__abc_44228_n21949), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_root_348__FF_INPUT) );
  AND2X2 AND2X2_11038 ( .A(u2__abc_44228_n3062_bF_buf37), .B(u2_o_348_), .Y(u2__abc_44228_n21951) );
  AND2X2 AND2X2_11039 ( .A(u2__abc_44228_n21941), .B(u2_o_347_), .Y(u2__abc_44228_n21953) );
  AND2X2 AND2X2_1104 ( .A(u2__abc_44228_n4222), .B(u2__abc_44228_n3885), .Y(u2__abc_44228_n4223) );
  AND2X2 AND2X2_11040 ( .A(u2__abc_44228_n21954), .B(u2__abc_44228_n21952), .Y(u2__abc_44228_n21955) );
  AND2X2 AND2X2_11041 ( .A(u2__abc_44228_n2983_bF_buf62), .B(u2__abc_44228_n5819), .Y(u2__abc_44228_n21957) );
  AND2X2 AND2X2_11042 ( .A(u2__abc_44228_n21958), .B(u2__abc_44228_n2972_bF_buf55), .Y(u2__abc_44228_n21959) );
  AND2X2 AND2X2_11043 ( .A(u2__abc_44228_n21956), .B(u2__abc_44228_n21959), .Y(u2__abc_44228_n21960) );
  AND2X2 AND2X2_11044 ( .A(u2__abc_44228_n21961), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_root_349__FF_INPUT) );
  AND2X2 AND2X2_11045 ( .A(u2__abc_44228_n3062_bF_buf36), .B(u2_o_349_), .Y(u2__abc_44228_n21963) );
  AND2X2 AND2X2_11046 ( .A(u2__abc_44228_n21953), .B(u2_o_348_), .Y(u2__abc_44228_n21965) );
  AND2X2 AND2X2_11047 ( .A(u2__abc_44228_n21966), .B(u2__abc_44228_n21964), .Y(u2__abc_44228_n21967) );
  AND2X2 AND2X2_11048 ( .A(u2__abc_44228_n2983_bF_buf60), .B(u2__abc_44228_n5812_1), .Y(u2__abc_44228_n21969) );
  AND2X2 AND2X2_11049 ( .A(u2__abc_44228_n21970), .B(u2__abc_44228_n2972_bF_buf54), .Y(u2__abc_44228_n21971) );
  AND2X2 AND2X2_1105 ( .A(u2__abc_44228_n3877), .B(u2__abc_44228_n3880), .Y(u2__abc_44228_n4224_1) );
  AND2X2 AND2X2_11050 ( .A(u2__abc_44228_n21968), .B(u2__abc_44228_n21971), .Y(u2__abc_44228_n21972) );
  AND2X2 AND2X2_11051 ( .A(u2__abc_44228_n21973), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_root_350__FF_INPUT) );
  AND2X2 AND2X2_11052 ( .A(u2__abc_44228_n3062_bF_buf35), .B(u2_o_350_), .Y(u2__abc_44228_n21975) );
  AND2X2 AND2X2_11053 ( .A(u2__abc_44228_n21965), .B(u2_o_349_), .Y(u2__abc_44228_n21977) );
  AND2X2 AND2X2_11054 ( .A(u2__abc_44228_n21978), .B(u2__abc_44228_n21976), .Y(u2__abc_44228_n21979) );
  AND2X2 AND2X2_11055 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n5801), .Y(u2__abc_44228_n21981) );
  AND2X2 AND2X2_11056 ( .A(u2__abc_44228_n21982), .B(u2__abc_44228_n2972_bF_buf53), .Y(u2__abc_44228_n21983) );
  AND2X2 AND2X2_11057 ( .A(u2__abc_44228_n21980), .B(u2__abc_44228_n21983), .Y(u2__abc_44228_n21984) );
  AND2X2 AND2X2_11058 ( .A(u2__abc_44228_n21985), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_root_351__FF_INPUT) );
  AND2X2 AND2X2_11059 ( .A(u2__abc_44228_n3062_bF_buf34), .B(u2_o_351_), .Y(u2__abc_44228_n21987) );
  AND2X2 AND2X2_1106 ( .A(u2__abc_44228_n4226), .B(u2__abc_44228_n3871), .Y(u2__abc_44228_n4227) );
  AND2X2 AND2X2_11060 ( .A(u2__abc_44228_n21977), .B(u2_o_350_), .Y(u2__abc_44228_n21989) );
  AND2X2 AND2X2_11061 ( .A(u2__abc_44228_n21990), .B(u2__abc_44228_n21988), .Y(u2__abc_44228_n21991) );
  AND2X2 AND2X2_11062 ( .A(u2__abc_44228_n2983_bF_buf56), .B(u2__abc_44228_n5794), .Y(u2__abc_44228_n21993) );
  AND2X2 AND2X2_11063 ( .A(u2__abc_44228_n21994), .B(u2__abc_44228_n2972_bF_buf52), .Y(u2__abc_44228_n21995) );
  AND2X2 AND2X2_11064 ( .A(u2__abc_44228_n21992), .B(u2__abc_44228_n21995), .Y(u2__abc_44228_n21996) );
  AND2X2 AND2X2_11065 ( .A(u2__abc_44228_n21997), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_root_352__FF_INPUT) );
  AND2X2 AND2X2_11066 ( .A(u2__abc_44228_n3062_bF_buf33), .B(u2_o_352_), .Y(u2__abc_44228_n21999) );
  AND2X2 AND2X2_11067 ( .A(u2__abc_44228_n21989), .B(u2_o_351_), .Y(u2__abc_44228_n22001) );
  AND2X2 AND2X2_11068 ( .A(u2__abc_44228_n22002), .B(u2__abc_44228_n22000), .Y(u2__abc_44228_n22003) );
  AND2X2 AND2X2_11069 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n5787), .Y(u2__abc_44228_n22005) );
  AND2X2 AND2X2_1107 ( .A(u2__abc_44228_n4229), .B(u2__abc_44228_n3865), .Y(u2__abc_44228_n4230) );
  AND2X2 AND2X2_11070 ( .A(u2__abc_44228_n22006), .B(u2__abc_44228_n2972_bF_buf51), .Y(u2__abc_44228_n22007) );
  AND2X2 AND2X2_11071 ( .A(u2__abc_44228_n22004), .B(u2__abc_44228_n22007), .Y(u2__abc_44228_n22008) );
  AND2X2 AND2X2_11072 ( .A(u2__abc_44228_n22009), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_root_353__FF_INPUT) );
  AND2X2 AND2X2_11073 ( .A(u2__abc_44228_n3062_bF_buf32), .B(u2_o_353_), .Y(u2__abc_44228_n22011) );
  AND2X2 AND2X2_11074 ( .A(u2__abc_44228_n22001), .B(u2_o_352_), .Y(u2__abc_44228_n22013) );
  AND2X2 AND2X2_11075 ( .A(u2__abc_44228_n22014), .B(u2__abc_44228_n22012), .Y(u2__abc_44228_n22015) );
  AND2X2 AND2X2_11076 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n5780), .Y(u2__abc_44228_n22017) );
  AND2X2 AND2X2_11077 ( .A(u2__abc_44228_n22018), .B(u2__abc_44228_n2972_bF_buf50), .Y(u2__abc_44228_n22019) );
  AND2X2 AND2X2_11078 ( .A(u2__abc_44228_n22016), .B(u2__abc_44228_n22019), .Y(u2__abc_44228_n22020) );
  AND2X2 AND2X2_11079 ( .A(u2__abc_44228_n22021), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_root_354__FF_INPUT) );
  AND2X2 AND2X2_1108 ( .A(u2__abc_44228_n4231), .B(u2__abc_44228_n3856), .Y(u2__abc_44228_n4232) );
  AND2X2 AND2X2_11080 ( .A(u2__abc_44228_n3062_bF_buf31), .B(u2_o_354_), .Y(u2__abc_44228_n22023) );
  AND2X2 AND2X2_11081 ( .A(u2__abc_44228_n22013), .B(u2_o_353_), .Y(u2__abc_44228_n22025) );
  AND2X2 AND2X2_11082 ( .A(u2__abc_44228_n22026), .B(u2__abc_44228_n22024), .Y(u2__abc_44228_n22027) );
  AND2X2 AND2X2_11083 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2__abc_44228_n5765_1), .Y(u2__abc_44228_n22029) );
  AND2X2 AND2X2_11084 ( .A(u2__abc_44228_n22030), .B(u2__abc_44228_n2972_bF_buf49), .Y(u2__abc_44228_n22031) );
  AND2X2 AND2X2_11085 ( .A(u2__abc_44228_n22028), .B(u2__abc_44228_n22031), .Y(u2__abc_44228_n22032) );
  AND2X2 AND2X2_11086 ( .A(u2__abc_44228_n22033), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_root_355__FF_INPUT) );
  AND2X2 AND2X2_11087 ( .A(u2__abc_44228_n3062_bF_buf30), .B(u2_o_355_), .Y(u2__abc_44228_n22035) );
  AND2X2 AND2X2_11088 ( .A(u2__abc_44228_n22025), .B(u2_o_354_), .Y(u2__abc_44228_n22037) );
  AND2X2 AND2X2_11089 ( .A(u2__abc_44228_n22038), .B(u2__abc_44228_n22036), .Y(u2__abc_44228_n22039) );
  AND2X2 AND2X2_1109 ( .A(u2__abc_44228_n3848), .B(u2__abc_44228_n3851), .Y(u2__abc_44228_n4233_1) );
  AND2X2 AND2X2_11090 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n5771), .Y(u2__abc_44228_n22041) );
  AND2X2 AND2X2_11091 ( .A(u2__abc_44228_n22042), .B(u2__abc_44228_n2972_bF_buf48), .Y(u2__abc_44228_n22043) );
  AND2X2 AND2X2_11092 ( .A(u2__abc_44228_n22040), .B(u2__abc_44228_n22043), .Y(u2__abc_44228_n22044) );
  AND2X2 AND2X2_11093 ( .A(u2__abc_44228_n22045), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_root_356__FF_INPUT) );
  AND2X2 AND2X2_11094 ( .A(u2__abc_44228_n3062_bF_buf29), .B(u2_o_356_), .Y(u2__abc_44228_n22047) );
  AND2X2 AND2X2_11095 ( .A(u2__abc_44228_n22037), .B(u2_o_355_), .Y(u2__abc_44228_n22049) );
  AND2X2 AND2X2_11096 ( .A(u2__abc_44228_n22050), .B(u2__abc_44228_n22048), .Y(u2__abc_44228_n22051) );
  AND2X2 AND2X2_11097 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n5758), .Y(u2__abc_44228_n22053) );
  AND2X2 AND2X2_11098 ( .A(u2__abc_44228_n22054), .B(u2__abc_44228_n2972_bF_buf47), .Y(u2__abc_44228_n22055) );
  AND2X2 AND2X2_11099 ( .A(u2__abc_44228_n22052), .B(u2__abc_44228_n22055), .Y(u2__abc_44228_n22056) );
  AND2X2 AND2X2_111 ( .A(_abc_64468_n933), .B(_abc_64468_n932), .Y(_auto_iopadmap_cc_313_execute_65414_146_) );
  AND2X2 AND2X2_1110 ( .A(u2__abc_44228_n4236), .B(u2__abc_44228_n3842), .Y(u2__abc_44228_n4237) );
  AND2X2 AND2X2_11100 ( .A(u2__abc_44228_n22057), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_root_357__FF_INPUT) );
  AND2X2 AND2X2_11101 ( .A(u2__abc_44228_n3062_bF_buf28), .B(u2_o_357_), .Y(u2__abc_44228_n22059) );
  AND2X2 AND2X2_11102 ( .A(u2__abc_44228_n22049), .B(u2_o_356_), .Y(u2__abc_44228_n22061) );
  AND2X2 AND2X2_11103 ( .A(u2__abc_44228_n22062), .B(u2__abc_44228_n22060), .Y(u2__abc_44228_n22063) );
  AND2X2 AND2X2_11104 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n5751), .Y(u2__abc_44228_n22065) );
  AND2X2 AND2X2_11105 ( .A(u2__abc_44228_n22066), .B(u2__abc_44228_n2972_bF_buf46), .Y(u2__abc_44228_n22067) );
  AND2X2 AND2X2_11106 ( .A(u2__abc_44228_n22064), .B(u2__abc_44228_n22067), .Y(u2__abc_44228_n22068) );
  AND2X2 AND2X2_11107 ( .A(u2__abc_44228_n22069), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_root_358__FF_INPUT) );
  AND2X2 AND2X2_11108 ( .A(u2__abc_44228_n3062_bF_buf27), .B(u2_o_358_), .Y(u2__abc_44228_n22071) );
  AND2X2 AND2X2_11109 ( .A(u2__abc_44228_n22061), .B(u2_o_357_), .Y(u2__abc_44228_n22073) );
  AND2X2 AND2X2_1111 ( .A(u2__abc_44228_n4239), .B(u2__abc_44228_n3815), .Y(u2__abc_44228_n4240) );
  AND2X2 AND2X2_11110 ( .A(u2__abc_44228_n22074), .B(u2__abc_44228_n22072), .Y(u2__abc_44228_n22075) );
  AND2X2 AND2X2_11111 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n5728_1), .Y(u2__abc_44228_n22077) );
  AND2X2 AND2X2_11112 ( .A(u2__abc_44228_n22078), .B(u2__abc_44228_n2972_bF_buf45), .Y(u2__abc_44228_n22079) );
  AND2X2 AND2X2_11113 ( .A(u2__abc_44228_n22076), .B(u2__abc_44228_n22079), .Y(u2__abc_44228_n22080) );
  AND2X2 AND2X2_11114 ( .A(u2__abc_44228_n22081), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_root_359__FF_INPUT) );
  AND2X2 AND2X2_11115 ( .A(u2__abc_44228_n3062_bF_buf26), .B(u2_o_359_), .Y(u2__abc_44228_n22083) );
  AND2X2 AND2X2_11116 ( .A(u2__abc_44228_n22073), .B(u2_o_358_), .Y(u2__abc_44228_n22085) );
  AND2X2 AND2X2_11117 ( .A(u2__abc_44228_n22086), .B(u2__abc_44228_n22084), .Y(u2__abc_44228_n22087) );
  AND2X2 AND2X2_11118 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n5721), .Y(u2__abc_44228_n22089) );
  AND2X2 AND2X2_11119 ( .A(u2__abc_44228_n22090), .B(u2__abc_44228_n2972_bF_buf44), .Y(u2__abc_44228_n22091) );
  AND2X2 AND2X2_1112 ( .A(u2__abc_44228_n4241), .B(u2__abc_44228_n3840), .Y(u2__abc_44228_n4242) );
  AND2X2 AND2X2_11120 ( .A(u2__abc_44228_n22088), .B(u2__abc_44228_n22091), .Y(u2__abc_44228_n22092) );
  AND2X2 AND2X2_11121 ( .A(u2__abc_44228_n22093), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_root_360__FF_INPUT) );
  AND2X2 AND2X2_11122 ( .A(u2__abc_44228_n3062_bF_buf25), .B(u2_o_360_), .Y(u2__abc_44228_n22095) );
  AND2X2 AND2X2_11123 ( .A(u2__abc_44228_n22085), .B(u2_o_359_), .Y(u2__abc_44228_n22097) );
  AND2X2 AND2X2_11124 ( .A(u2__abc_44228_n22098), .B(u2__abc_44228_n22096), .Y(u2__abc_44228_n22099) );
  AND2X2 AND2X2_11125 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n5742), .Y(u2__abc_44228_n22101) );
  AND2X2 AND2X2_11126 ( .A(u2__abc_44228_n22102), .B(u2__abc_44228_n2972_bF_buf43), .Y(u2__abc_44228_n22103) );
  AND2X2 AND2X2_11127 ( .A(u2__abc_44228_n22100), .B(u2__abc_44228_n22103), .Y(u2__abc_44228_n22104) );
  AND2X2 AND2X2_11128 ( .A(u2__abc_44228_n22105), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_root_361__FF_INPUT) );
  AND2X2 AND2X2_11129 ( .A(u2__abc_44228_n3062_bF_buf24), .B(u2_o_361_), .Y(u2__abc_44228_n22107) );
  AND2X2 AND2X2_1113 ( .A(u2__abc_44228_n3829), .B(u2__abc_44228_n4243_1), .Y(u2__abc_44228_n4244) );
  AND2X2 AND2X2_11130 ( .A(u2__abc_44228_n22097), .B(u2_o_360_), .Y(u2__abc_44228_n22109) );
  AND2X2 AND2X2_11131 ( .A(u2__abc_44228_n22110), .B(u2__abc_44228_n22108), .Y(u2__abc_44228_n22111) );
  AND2X2 AND2X2_11132 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n5735), .Y(u2__abc_44228_n22113) );
  AND2X2 AND2X2_11133 ( .A(u2__abc_44228_n22114), .B(u2__abc_44228_n2972_bF_buf42), .Y(u2__abc_44228_n22115) );
  AND2X2 AND2X2_11134 ( .A(u2__abc_44228_n22112), .B(u2__abc_44228_n22115), .Y(u2__abc_44228_n22116) );
  AND2X2 AND2X2_11135 ( .A(u2__abc_44228_n22117), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_root_362__FF_INPUT) );
  AND2X2 AND2X2_11136 ( .A(u2__abc_44228_n3062_bF_buf23), .B(u2_o_362_), .Y(u2__abc_44228_n22119) );
  AND2X2 AND2X2_11137 ( .A(u2__abc_44228_n22109), .B(u2_o_361_), .Y(u2__abc_44228_n22121) );
  AND2X2 AND2X2_11138 ( .A(u2__abc_44228_n22122), .B(u2__abc_44228_n22120), .Y(u2__abc_44228_n22123) );
  AND2X2 AND2X2_11139 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n5713), .Y(u2__abc_44228_n22125) );
  AND2X2 AND2X2_1114 ( .A(u2__abc_44228_n4245), .B(u2__abc_44228_n3832), .Y(u2__abc_44228_n4246) );
  AND2X2 AND2X2_11140 ( .A(u2__abc_44228_n22126), .B(u2__abc_44228_n2972_bF_buf41), .Y(u2__abc_44228_n22127) );
  AND2X2 AND2X2_11141 ( .A(u2__abc_44228_n22124), .B(u2__abc_44228_n22127), .Y(u2__abc_44228_n22128) );
  AND2X2 AND2X2_11142 ( .A(u2__abc_44228_n22129), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_root_363__FF_INPUT) );
  AND2X2 AND2X2_11143 ( .A(u2__abc_44228_n3062_bF_buf22), .B(u2_o_363_), .Y(u2__abc_44228_n22131) );
  AND2X2 AND2X2_11144 ( .A(u2__abc_44228_n22121), .B(u2_o_362_), .Y(u2__abc_44228_n22133) );
  AND2X2 AND2X2_11145 ( .A(u2__abc_44228_n22134), .B(u2__abc_44228_n22132), .Y(u2__abc_44228_n22135) );
  AND2X2 AND2X2_11146 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n5706), .Y(u2__abc_44228_n22137) );
  AND2X2 AND2X2_11147 ( .A(u2__abc_44228_n22138), .B(u2__abc_44228_n2972_bF_buf40), .Y(u2__abc_44228_n22139) );
  AND2X2 AND2X2_11148 ( .A(u2__abc_44228_n22136), .B(u2__abc_44228_n22139), .Y(u2__abc_44228_n22140) );
  AND2X2 AND2X2_11149 ( .A(u2__abc_44228_n22141), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_root_364__FF_INPUT) );
  AND2X2 AND2X2_1115 ( .A(u2__abc_44228_n4247), .B(u2__abc_44228_n3812), .Y(u2__abc_44228_n4248) );
  AND2X2 AND2X2_11150 ( .A(u2__abc_44228_n3062_bF_buf21), .B(u2_o_364_), .Y(u2__abc_44228_n22143) );
  AND2X2 AND2X2_11151 ( .A(u2__abc_44228_n22133), .B(u2_o_363_), .Y(u2__abc_44228_n22145) );
  AND2X2 AND2X2_11152 ( .A(u2__abc_44228_n22146), .B(u2__abc_44228_n22144), .Y(u2__abc_44228_n22147) );
  AND2X2 AND2X2_11153 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n5699), .Y(u2__abc_44228_n22149) );
  AND2X2 AND2X2_11154 ( .A(u2__abc_44228_n22150), .B(u2__abc_44228_n2972_bF_buf39), .Y(u2__abc_44228_n22151) );
  AND2X2 AND2X2_11155 ( .A(u2__abc_44228_n22148), .B(u2__abc_44228_n22151), .Y(u2__abc_44228_n22152) );
  AND2X2 AND2X2_11156 ( .A(u2__abc_44228_n22153), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_root_365__FF_INPUT) );
  AND2X2 AND2X2_11157 ( .A(u2__abc_44228_n3062_bF_buf20), .B(u2_o_365_), .Y(u2__abc_44228_n22155) );
  AND2X2 AND2X2_11158 ( .A(u2__abc_44228_n22145), .B(u2_o_364_), .Y(u2__abc_44228_n22157) );
  AND2X2 AND2X2_11159 ( .A(u2__abc_44228_n22158), .B(u2__abc_44228_n22156), .Y(u2__abc_44228_n22159) );
  AND2X2 AND2X2_1116 ( .A(u2__abc_44228_n4249), .B(u2__abc_44228_n3806), .Y(u2__abc_44228_n4250) );
  AND2X2 AND2X2_11160 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n5692), .Y(u2__abc_44228_n22161) );
  AND2X2 AND2X2_11161 ( .A(u2__abc_44228_n22162), .B(u2__abc_44228_n2972_bF_buf38), .Y(u2__abc_44228_n22163) );
  AND2X2 AND2X2_11162 ( .A(u2__abc_44228_n22160), .B(u2__abc_44228_n22163), .Y(u2__abc_44228_n22164) );
  AND2X2 AND2X2_11163 ( .A(u2__abc_44228_n22165), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_root_366__FF_INPUT) );
  AND2X2 AND2X2_11164 ( .A(u2__abc_44228_n3062_bF_buf19), .B(u2_o_366_), .Y(u2__abc_44228_n22167) );
  AND2X2 AND2X2_11165 ( .A(u2__abc_44228_n22157), .B(u2_o_365_), .Y(u2__abc_44228_n22169) );
  AND2X2 AND2X2_11166 ( .A(u2__abc_44228_n22170), .B(u2__abc_44228_n22168), .Y(u2__abc_44228_n22171) );
  AND2X2 AND2X2_11167 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n5668), .Y(u2__abc_44228_n22173) );
  AND2X2 AND2X2_11168 ( .A(u2__abc_44228_n22174), .B(u2__abc_44228_n2972_bF_buf37), .Y(u2__abc_44228_n22175) );
  AND2X2 AND2X2_11169 ( .A(u2__abc_44228_n22172), .B(u2__abc_44228_n22175), .Y(u2__abc_44228_n22176) );
  AND2X2 AND2X2_1117 ( .A(u2__abc_44228_n4251), .B(u2__abc_44228_n3809), .Y(u2__abc_44228_n4252) );
  AND2X2 AND2X2_11170 ( .A(u2__abc_44228_n22177), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_root_367__FF_INPUT) );
  AND2X2 AND2X2_11171 ( .A(u2__abc_44228_n3062_bF_buf18), .B(u2_o_367_), .Y(u2__abc_44228_n22179) );
  AND2X2 AND2X2_11172 ( .A(u2__abc_44228_n22169), .B(u2_o_366_), .Y(u2__abc_44228_n22181) );
  AND2X2 AND2X2_11173 ( .A(u2__abc_44228_n22182), .B(u2__abc_44228_n22180), .Y(u2__abc_44228_n22183) );
  AND2X2 AND2X2_11174 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n5661), .Y(u2__abc_44228_n22185) );
  AND2X2 AND2X2_11175 ( .A(u2__abc_44228_n22186), .B(u2__abc_44228_n2972_bF_buf36), .Y(u2__abc_44228_n22187) );
  AND2X2 AND2X2_11176 ( .A(u2__abc_44228_n22184), .B(u2__abc_44228_n22187), .Y(u2__abc_44228_n22188) );
  AND2X2 AND2X2_11177 ( .A(u2__abc_44228_n22189), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_root_368__FF_INPUT) );
  AND2X2 AND2X2_11178 ( .A(u2__abc_44228_n3062_bF_buf17), .B(u2_o_368_), .Y(u2__abc_44228_n22191) );
  AND2X2 AND2X2_11179 ( .A(u2__abc_44228_n22181), .B(u2_o_367_), .Y(u2__abc_44228_n22193) );
  AND2X2 AND2X2_1118 ( .A(u2__abc_44228_n4252), .B(u2__abc_44228_n3797), .Y(u2__abc_44228_n4253_1) );
  AND2X2 AND2X2_11180 ( .A(u2__abc_44228_n22194), .B(u2__abc_44228_n22192), .Y(u2__abc_44228_n22195) );
  AND2X2 AND2X2_11181 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n5682), .Y(u2__abc_44228_n22197) );
  AND2X2 AND2X2_11182 ( .A(u2__abc_44228_n22198), .B(u2__abc_44228_n2972_bF_buf35), .Y(u2__abc_44228_n22199) );
  AND2X2 AND2X2_11183 ( .A(u2__abc_44228_n22196), .B(u2__abc_44228_n22199), .Y(u2__abc_44228_n22200) );
  AND2X2 AND2X2_11184 ( .A(u2__abc_44228_n22201), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_root_369__FF_INPUT) );
  AND2X2 AND2X2_11185 ( .A(u2__abc_44228_n3062_bF_buf16), .B(u2_o_369_), .Y(u2__abc_44228_n22203) );
  AND2X2 AND2X2_11186 ( .A(u2__abc_44228_n22193), .B(u2_o_368_), .Y(u2__abc_44228_n22205) );
  AND2X2 AND2X2_11187 ( .A(u2__abc_44228_n22206), .B(u2__abc_44228_n22204), .Y(u2__abc_44228_n22207) );
  AND2X2 AND2X2_11188 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n5675), .Y(u2__abc_44228_n22209) );
  AND2X2 AND2X2_11189 ( .A(u2__abc_44228_n22210), .B(u2__abc_44228_n2972_bF_buf34), .Y(u2__abc_44228_n22211) );
  AND2X2 AND2X2_1119 ( .A(u2__abc_44228_n3789_1), .B(u2__abc_44228_n3792), .Y(u2__abc_44228_n4254) );
  AND2X2 AND2X2_11190 ( .A(u2__abc_44228_n22208), .B(u2__abc_44228_n22211), .Y(u2__abc_44228_n22212) );
  AND2X2 AND2X2_11191 ( .A(u2__abc_44228_n22213), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_root_370__FF_INPUT) );
  AND2X2 AND2X2_11192 ( .A(u2__abc_44228_n3062_bF_buf15), .B(u2_o_370_), .Y(u2__abc_44228_n22215) );
  AND2X2 AND2X2_11193 ( .A(u2__abc_44228_n22205), .B(u2_o_369_), .Y(u2__abc_44228_n22217) );
  AND2X2 AND2X2_11194 ( .A(u2__abc_44228_n22218), .B(u2__abc_44228_n22216), .Y(u2__abc_44228_n22219) );
  AND2X2 AND2X2_11195 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n5646), .Y(u2__abc_44228_n22221) );
  AND2X2 AND2X2_11196 ( .A(u2__abc_44228_n22222), .B(u2__abc_44228_n2972_bF_buf33), .Y(u2__abc_44228_n22223) );
  AND2X2 AND2X2_11197 ( .A(u2__abc_44228_n22220), .B(u2__abc_44228_n22223), .Y(u2__abc_44228_n22224) );
  AND2X2 AND2X2_11198 ( .A(u2__abc_44228_n22225), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_root_371__FF_INPUT) );
  AND2X2 AND2X2_11199 ( .A(u2__abc_44228_n3062_bF_buf14), .B(u2_o_371_), .Y(u2__abc_44228_n22227) );
  AND2X2 AND2X2_112 ( .A(_abc_64468_n936), .B(_abc_64468_n935), .Y(_auto_iopadmap_cc_313_execute_65414_147_) );
  AND2X2 AND2X2_1120 ( .A(u2__abc_44228_n4258), .B(u2__abc_44228_n3783), .Y(u2__abc_44228_n4259) );
  AND2X2 AND2X2_11200 ( .A(u2__abc_44228_n22217), .B(u2_o_370_), .Y(u2__abc_44228_n22229) );
  AND2X2 AND2X2_11201 ( .A(u2__abc_44228_n22230), .B(u2__abc_44228_n22228), .Y(u2__abc_44228_n22231) );
  AND2X2 AND2X2_11202 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n5652_1), .Y(u2__abc_44228_n22233) );
  AND2X2 AND2X2_11203 ( .A(u2__abc_44228_n22234), .B(u2__abc_44228_n2972_bF_buf32), .Y(u2__abc_44228_n22235) );
  AND2X2 AND2X2_11204 ( .A(u2__abc_44228_n22232), .B(u2__abc_44228_n22235), .Y(u2__abc_44228_n22236) );
  AND2X2 AND2X2_11205 ( .A(u2__abc_44228_n22237), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_root_372__FF_INPUT) );
  AND2X2 AND2X2_11206 ( .A(u2__abc_44228_n3062_bF_buf13), .B(u2_o_372_), .Y(u2__abc_44228_n22239) );
  AND2X2 AND2X2_11207 ( .A(u2__abc_44228_n22229), .B(u2_o_371_), .Y(u2__abc_44228_n22241) );
  AND2X2 AND2X2_11208 ( .A(u2__abc_44228_n22242), .B(u2__abc_44228_n22240), .Y(u2__abc_44228_n22243) );
  AND2X2 AND2X2_11209 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n5639), .Y(u2__abc_44228_n22245) );
  AND2X2 AND2X2_1121 ( .A(u2__abc_44228_n4261), .B(u2__abc_44228_n3696), .Y(u2__abc_44228_n4262_1) );
  AND2X2 AND2X2_11210 ( .A(u2__abc_44228_n22246), .B(u2__abc_44228_n2972_bF_buf31), .Y(u2__abc_44228_n22247) );
  AND2X2 AND2X2_11211 ( .A(u2__abc_44228_n22244), .B(u2__abc_44228_n22247), .Y(u2__abc_44228_n22248) );
  AND2X2 AND2X2_11212 ( .A(u2__abc_44228_n22249), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_root_373__FF_INPUT) );
  AND2X2 AND2X2_11213 ( .A(u2__abc_44228_n3062_bF_buf12), .B(u2_o_373_), .Y(u2__abc_44228_n22251) );
  AND2X2 AND2X2_11214 ( .A(u2__abc_44228_n22241), .B(u2_o_372_), .Y(u2__abc_44228_n22253) );
  AND2X2 AND2X2_11215 ( .A(u2__abc_44228_n22254), .B(u2__abc_44228_n22252), .Y(u2__abc_44228_n22255) );
  AND2X2 AND2X2_11216 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n5632), .Y(u2__abc_44228_n22257) );
  AND2X2 AND2X2_11217 ( .A(u2__abc_44228_n22258), .B(u2__abc_44228_n2972_bF_buf30), .Y(u2__abc_44228_n22259) );
  AND2X2 AND2X2_11218 ( .A(u2__abc_44228_n22256), .B(u2__abc_44228_n22259), .Y(u2__abc_44228_n22260) );
  AND2X2 AND2X2_11219 ( .A(u2__abc_44228_n22261), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_root_374__FF_INPUT) );
  AND2X2 AND2X2_1122 ( .A(u2__abc_44228_n4263), .B(u2__abc_44228_n3721), .Y(u2__abc_44228_n4264) );
  AND2X2 AND2X2_11220 ( .A(u2__abc_44228_n3062_bF_buf11), .B(u2_o_374_), .Y(u2__abc_44228_n22263) );
  AND2X2 AND2X2_11221 ( .A(u2__abc_44228_n22253), .B(u2_o_373_), .Y(u2__abc_44228_n22265) );
  AND2X2 AND2X2_11222 ( .A(u2__abc_44228_n22266), .B(u2__abc_44228_n22264), .Y(u2__abc_44228_n22267) );
  AND2X2 AND2X2_11223 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n5609), .Y(u2__abc_44228_n22269) );
  AND2X2 AND2X2_11224 ( .A(u2__abc_44228_n22270), .B(u2__abc_44228_n2972_bF_buf29), .Y(u2__abc_44228_n22271) );
  AND2X2 AND2X2_11225 ( .A(u2__abc_44228_n22268), .B(u2__abc_44228_n22271), .Y(u2__abc_44228_n22272) );
  AND2X2 AND2X2_11226 ( .A(u2__abc_44228_n22273), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_root_375__FF_INPUT) );
  AND2X2 AND2X2_11227 ( .A(u2__abc_44228_n3062_bF_buf10), .B(u2_o_375_), .Y(u2__abc_44228_n22275) );
  AND2X2 AND2X2_11228 ( .A(u2__abc_44228_n22265), .B(u2_o_374_), .Y(u2__abc_44228_n22277) );
  AND2X2 AND2X2_11229 ( .A(u2__abc_44228_n22278), .B(u2__abc_44228_n22276), .Y(u2__abc_44228_n22279) );
  AND2X2 AND2X2_1123 ( .A(u2__abc_44228_n4265), .B(u2__abc_44228_n3713), .Y(u2__abc_44228_n4266) );
  AND2X2 AND2X2_11230 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n5602), .Y(u2__abc_44228_n22281) );
  AND2X2 AND2X2_11231 ( .A(u2__abc_44228_n22282), .B(u2__abc_44228_n2972_bF_buf28), .Y(u2__abc_44228_n22283) );
  AND2X2 AND2X2_11232 ( .A(u2__abc_44228_n22280), .B(u2__abc_44228_n22283), .Y(u2__abc_44228_n22284) );
  AND2X2 AND2X2_11233 ( .A(u2__abc_44228_n22285), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_root_376__FF_INPUT) );
  AND2X2 AND2X2_11234 ( .A(u2__abc_44228_n3062_bF_buf9), .B(u2_o_376_), .Y(u2__abc_44228_n22287) );
  AND2X2 AND2X2_11235 ( .A(u2__abc_44228_n22277), .B(u2_o_375_), .Y(u2__abc_44228_n22289) );
  AND2X2 AND2X2_11236 ( .A(u2__abc_44228_n22290), .B(u2__abc_44228_n22288), .Y(u2__abc_44228_n22291) );
  AND2X2 AND2X2_11237 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n5623), .Y(u2__abc_44228_n22293) );
  AND2X2 AND2X2_11238 ( .A(u2__abc_44228_n22294), .B(u2__abc_44228_n2972_bF_buf27), .Y(u2__abc_44228_n22295) );
  AND2X2 AND2X2_11239 ( .A(u2__abc_44228_n22292), .B(u2__abc_44228_n22295), .Y(u2__abc_44228_n22296) );
  AND2X2 AND2X2_1124 ( .A(u2__abc_44228_n4267), .B(u2__abc_44228_n3693), .Y(u2__abc_44228_n4268) );
  AND2X2 AND2X2_11240 ( .A(u2__abc_44228_n22297), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_root_377__FF_INPUT) );
  AND2X2 AND2X2_11241 ( .A(u2__abc_44228_n3062_bF_buf8), .B(u2_o_377_), .Y(u2__abc_44228_n22299) );
  AND2X2 AND2X2_11242 ( .A(u2__abc_44228_n22289), .B(u2_o_376_), .Y(u2__abc_44228_n22301) );
  AND2X2 AND2X2_11243 ( .A(u2__abc_44228_n22302), .B(u2__abc_44228_n22300), .Y(u2__abc_44228_n22303) );
  AND2X2 AND2X2_11244 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n5616), .Y(u2__abc_44228_n22305) );
  AND2X2 AND2X2_11245 ( .A(u2__abc_44228_n22306), .B(u2__abc_44228_n2972_bF_buf26), .Y(u2__abc_44228_n22307) );
  AND2X2 AND2X2_11246 ( .A(u2__abc_44228_n22304), .B(u2__abc_44228_n22307), .Y(u2__abc_44228_n22308) );
  AND2X2 AND2X2_11247 ( .A(u2__abc_44228_n22309), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_root_378__FF_INPUT) );
  AND2X2 AND2X2_11248 ( .A(u2__abc_44228_n3062_bF_buf7), .B(u2_o_378_), .Y(u2__abc_44228_n22311) );
  AND2X2 AND2X2_11249 ( .A(u2__abc_44228_n22301), .B(u2_o_377_), .Y(u2__abc_44228_n22313) );
  AND2X2 AND2X2_1125 ( .A(u2__abc_44228_n4269), .B(u2__abc_44228_n3687), .Y(u2__abc_44228_n4270) );
  AND2X2 AND2X2_11250 ( .A(u2__abc_44228_n22314), .B(u2__abc_44228_n22312), .Y(u2__abc_44228_n22315) );
  AND2X2 AND2X2_11251 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n5594), .Y(u2__abc_44228_n22317) );
  AND2X2 AND2X2_11252 ( .A(u2__abc_44228_n22318), .B(u2__abc_44228_n2972_bF_buf25), .Y(u2__abc_44228_n22319) );
  AND2X2 AND2X2_11253 ( .A(u2__abc_44228_n22316), .B(u2__abc_44228_n22319), .Y(u2__abc_44228_n22320) );
  AND2X2 AND2X2_11254 ( .A(u2__abc_44228_n22321), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_root_379__FF_INPUT) );
  AND2X2 AND2X2_11255 ( .A(u2__abc_44228_n3062_bF_buf6), .B(u2_o_379_), .Y(u2__abc_44228_n22323) );
  AND2X2 AND2X2_11256 ( .A(u2__abc_44228_n22313), .B(u2_o_378_), .Y(u2__abc_44228_n22325) );
  AND2X2 AND2X2_11257 ( .A(u2__abc_44228_n22326), .B(u2__abc_44228_n22324), .Y(u2__abc_44228_n22327) );
  AND2X2 AND2X2_11258 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n5587_1), .Y(u2__abc_44228_n22329) );
  AND2X2 AND2X2_11259 ( .A(u2__abc_44228_n22330), .B(u2__abc_44228_n2972_bF_buf24), .Y(u2__abc_44228_n22331) );
  AND2X2 AND2X2_1126 ( .A(u2__abc_44228_n4271), .B(u2__abc_44228_n3690), .Y(u2__abc_44228_n4272_1) );
  AND2X2 AND2X2_11260 ( .A(u2__abc_44228_n22328), .B(u2__abc_44228_n22331), .Y(u2__abc_44228_n22332) );
  AND2X2 AND2X2_11261 ( .A(u2__abc_44228_n22333), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_root_380__FF_INPUT) );
  AND2X2 AND2X2_11262 ( .A(u2__abc_44228_n3062_bF_buf5), .B(u2_o_380_), .Y(u2__abc_44228_n22335) );
  AND2X2 AND2X2_11263 ( .A(u2__abc_44228_n22325), .B(u2_o_379_), .Y(u2__abc_44228_n22337) );
  AND2X2 AND2X2_11264 ( .A(u2__abc_44228_n22338), .B(u2__abc_44228_n22336), .Y(u2__abc_44228_n22339) );
  AND2X2 AND2X2_11265 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n5580), .Y(u2__abc_44228_n22341) );
  AND2X2 AND2X2_11266 ( .A(u2__abc_44228_n22342), .B(u2__abc_44228_n2972_bF_buf23), .Y(u2__abc_44228_n22343) );
  AND2X2 AND2X2_11267 ( .A(u2__abc_44228_n22340), .B(u2__abc_44228_n22343), .Y(u2__abc_44228_n22344) );
  AND2X2 AND2X2_11268 ( .A(u2__abc_44228_n22345), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_root_381__FF_INPUT) );
  AND2X2 AND2X2_11269 ( .A(u2__abc_44228_n3062_bF_buf4), .B(u2_o_381_), .Y(u2__abc_44228_n22347) );
  AND2X2 AND2X2_1127 ( .A(u2__abc_44228_n4272_1), .B(u2__abc_44228_n3678), .Y(u2__abc_44228_n4273) );
  AND2X2 AND2X2_11270 ( .A(u2__abc_44228_n22337), .B(u2_o_380_), .Y(u2__abc_44228_n22349) );
  AND2X2 AND2X2_11271 ( .A(u2__abc_44228_n22350), .B(u2__abc_44228_n22348), .Y(u2__abc_44228_n22351) );
  AND2X2 AND2X2_11272 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n5573), .Y(u2__abc_44228_n22353) );
  AND2X2 AND2X2_11273 ( .A(u2__abc_44228_n22354), .B(u2__abc_44228_n2972_bF_buf22), .Y(u2__abc_44228_n22355) );
  AND2X2 AND2X2_11274 ( .A(u2__abc_44228_n22352), .B(u2__abc_44228_n22355), .Y(u2__abc_44228_n22356) );
  AND2X2 AND2X2_11275 ( .A(u2__abc_44228_n22357), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_root_382__FF_INPUT) );
  AND2X2 AND2X2_11276 ( .A(u2__abc_44228_n3062_bF_buf3), .B(u2_o_382_), .Y(u2__abc_44228_n22359) );
  AND2X2 AND2X2_11277 ( .A(u2__abc_44228_n22349), .B(u2_o_381_), .Y(u2__abc_44228_n22361) );
  AND2X2 AND2X2_11278 ( .A(u2__abc_44228_n22362), .B(u2__abc_44228_n22360), .Y(u2__abc_44228_n22363) );
  AND2X2 AND2X2_11279 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n7333), .Y(u2__abc_44228_n22365) );
  AND2X2 AND2X2_1128 ( .A(u2__abc_44228_n3670), .B(u2__abc_44228_n3673), .Y(u2__abc_44228_n4274) );
  AND2X2 AND2X2_11280 ( .A(u2__abc_44228_n22366), .B(u2__abc_44228_n2972_bF_buf21), .Y(u2__abc_44228_n22367) );
  AND2X2 AND2X2_11281 ( .A(u2__abc_44228_n22364), .B(u2__abc_44228_n22367), .Y(u2__abc_44228_n22368) );
  AND2X2 AND2X2_11282 ( .A(u2__abc_44228_n22369), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_root_383__FF_INPUT) );
  AND2X2 AND2X2_11283 ( .A(u2__abc_44228_n3062_bF_buf2), .B(u2_o_383_), .Y(u2__abc_44228_n22371) );
  AND2X2 AND2X2_11284 ( .A(u2__abc_44228_n22361), .B(u2_o_382_), .Y(u2__abc_44228_n22373) );
  AND2X2 AND2X2_11285 ( .A(u2__abc_44228_n22374), .B(u2__abc_44228_n22372), .Y(u2__abc_44228_n22375) );
  AND2X2 AND2X2_11286 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n7326), .Y(u2__abc_44228_n22377) );
  AND2X2 AND2X2_11287 ( .A(u2__abc_44228_n22378), .B(u2__abc_44228_n2972_bF_buf20), .Y(u2__abc_44228_n22379) );
  AND2X2 AND2X2_11288 ( .A(u2__abc_44228_n22376), .B(u2__abc_44228_n22379), .Y(u2__abc_44228_n22380) );
  AND2X2 AND2X2_11289 ( .A(u2__abc_44228_n22381), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_root_384__FF_INPUT) );
  AND2X2 AND2X2_1129 ( .A(u2__abc_44228_n4278), .B(u2__abc_44228_n3775), .Y(u2__abc_44228_n4279) );
  AND2X2 AND2X2_11290 ( .A(u2__abc_44228_n3062_bF_buf1), .B(u2_o_384_), .Y(u2__abc_44228_n22383) );
  AND2X2 AND2X2_11291 ( .A(u2__abc_44228_n22373), .B(u2_o_383_), .Y(u2__abc_44228_n22385) );
  AND2X2 AND2X2_11292 ( .A(u2__abc_44228_n22386), .B(u2__abc_44228_n22384), .Y(u2__abc_44228_n22387) );
  AND2X2 AND2X2_11293 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n7319_1), .Y(u2__abc_44228_n22389) );
  AND2X2 AND2X2_11294 ( .A(u2__abc_44228_n22390), .B(u2__abc_44228_n2972_bF_buf19), .Y(u2__abc_44228_n22391) );
  AND2X2 AND2X2_11295 ( .A(u2__abc_44228_n22388), .B(u2__abc_44228_n22391), .Y(u2__abc_44228_n22392) );
  AND2X2 AND2X2_11296 ( .A(u2__abc_44228_n22393), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_root_385__FF_INPUT) );
  AND2X2 AND2X2_11297 ( .A(u2__abc_44228_n3062_bF_buf0), .B(u2_o_385_), .Y(u2__abc_44228_n22395) );
  AND2X2 AND2X2_11298 ( .A(u2__abc_44228_n22385), .B(u2_o_384_), .Y(u2__abc_44228_n22397) );
  AND2X2 AND2X2_11299 ( .A(u2__abc_44228_n22398), .B(u2__abc_44228_n22396), .Y(u2__abc_44228_n22399) );
  AND2X2 AND2X2_113 ( .A(_abc_64468_n939), .B(_abc_64468_n938), .Y(_auto_iopadmap_cc_313_execute_65414_148_) );
  AND2X2 AND2X2_1130 ( .A(u2__abc_44228_n4280), .B(u2__abc_44228_n3778), .Y(u2__abc_44228_n4281_1) );
  AND2X2 AND2X2_11300 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n7312), .Y(u2__abc_44228_n22401) );
  AND2X2 AND2X2_11301 ( .A(u2__abc_44228_n22402), .B(u2__abc_44228_n2972_bF_buf18), .Y(u2__abc_44228_n22403) );
  AND2X2 AND2X2_11302 ( .A(u2__abc_44228_n22400), .B(u2__abc_44228_n22403), .Y(u2__abc_44228_n22404) );
  AND2X2 AND2X2_11303 ( .A(u2__abc_44228_n22405), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_root_386__FF_INPUT) );
  AND2X2 AND2X2_11304 ( .A(u2__abc_44228_n3062_bF_buf92), .B(u2_o_386_), .Y(u2__abc_44228_n22407) );
  AND2X2 AND2X2_11305 ( .A(u2__abc_44228_n22397), .B(u2_o_385_), .Y(u2__abc_44228_n22409) );
  AND2X2 AND2X2_11306 ( .A(u2__abc_44228_n22410), .B(u2__abc_44228_n22408), .Y(u2__abc_44228_n22411) );
  AND2X2 AND2X2_11307 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n7297), .Y(u2__abc_44228_n22413) );
  AND2X2 AND2X2_11308 ( .A(u2__abc_44228_n22414), .B(u2__abc_44228_n2972_bF_buf17), .Y(u2__abc_44228_n22415) );
  AND2X2 AND2X2_11309 ( .A(u2__abc_44228_n22412), .B(u2__abc_44228_n22415), .Y(u2__abc_44228_n22416) );
  AND2X2 AND2X2_1131 ( .A(u2__abc_44228_n4281_1), .B(u2__abc_44228_n3766), .Y(u2__abc_44228_n4282) );
  AND2X2 AND2X2_11310 ( .A(u2__abc_44228_n22417), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_root_387__FF_INPUT) );
  AND2X2 AND2X2_11311 ( .A(u2__abc_44228_n3062_bF_buf91), .B(u2_o_387_), .Y(u2__abc_44228_n22419) );
  AND2X2 AND2X2_11312 ( .A(u2__abc_44228_n22409), .B(u2_o_386_), .Y(u2__abc_44228_n22421) );
  AND2X2 AND2X2_11313 ( .A(u2__abc_44228_n22422), .B(u2__abc_44228_n22420), .Y(u2__abc_44228_n22423) );
  AND2X2 AND2X2_11314 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n7303), .Y(u2__abc_44228_n22425) );
  AND2X2 AND2X2_11315 ( .A(u2__abc_44228_n22426), .B(u2__abc_44228_n2972_bF_buf16), .Y(u2__abc_44228_n22427) );
  AND2X2 AND2X2_11316 ( .A(u2__abc_44228_n22424), .B(u2__abc_44228_n22427), .Y(u2__abc_44228_n22428) );
  AND2X2 AND2X2_11317 ( .A(u2__abc_44228_n22429), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_root_388__FF_INPUT) );
  AND2X2 AND2X2_11318 ( .A(u2__abc_44228_n3062_bF_buf90), .B(u2_o_388_), .Y(u2__abc_44228_n22431) );
  AND2X2 AND2X2_11319 ( .A(u2__abc_44228_n22421), .B(u2_o_387_), .Y(u2__abc_44228_n22433) );
  AND2X2 AND2X2_1132 ( .A(u2__abc_44228_n3758), .B(u2__abc_44228_n3761), .Y(u2__abc_44228_n4283) );
  AND2X2 AND2X2_11320 ( .A(u2__abc_44228_n22434), .B(u2__abc_44228_n22432), .Y(u2__abc_44228_n22435) );
  AND2X2 AND2X2_11321 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n7290), .Y(u2__abc_44228_n22437) );
  AND2X2 AND2X2_11322 ( .A(u2__abc_44228_n22438), .B(u2__abc_44228_n2972_bF_buf15), .Y(u2__abc_44228_n22439) );
  AND2X2 AND2X2_11323 ( .A(u2__abc_44228_n22436), .B(u2__abc_44228_n22439), .Y(u2__abc_44228_n22440) );
  AND2X2 AND2X2_11324 ( .A(u2__abc_44228_n22441), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_root_389__FF_INPUT) );
  AND2X2 AND2X2_11325 ( .A(u2__abc_44228_n3062_bF_buf89), .B(u2_o_389_), .Y(u2__abc_44228_n22443) );
  AND2X2 AND2X2_11326 ( .A(u2__abc_44228_n22433), .B(u2_o_388_), .Y(u2__abc_44228_n22445) );
  AND2X2 AND2X2_11327 ( .A(u2__abc_44228_n22446), .B(u2__abc_44228_n22444), .Y(u2__abc_44228_n22447) );
  AND2X2 AND2X2_11328 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n7283), .Y(u2__abc_44228_n22449) );
  AND2X2 AND2X2_11329 ( .A(u2__abc_44228_n22450), .B(u2__abc_44228_n2972_bF_buf14), .Y(u2__abc_44228_n22451) );
  AND2X2 AND2X2_1133 ( .A(u2__abc_44228_n4285), .B(u2__abc_44228_n3752), .Y(u2__abc_44228_n4286) );
  AND2X2 AND2X2_11330 ( .A(u2__abc_44228_n22448), .B(u2__abc_44228_n22451), .Y(u2__abc_44228_n22452) );
  AND2X2 AND2X2_11331 ( .A(u2__abc_44228_n22453), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_root_390__FF_INPUT) );
  AND2X2 AND2X2_11332 ( .A(u2__abc_44228_n3062_bF_buf88), .B(u2_o_390_), .Y(u2__abc_44228_n22455) );
  AND2X2 AND2X2_11333 ( .A(u2__abc_44228_n22445), .B(u2_o_389_), .Y(u2__abc_44228_n22457) );
  AND2X2 AND2X2_11334 ( .A(u2__abc_44228_n22458), .B(u2__abc_44228_n22456), .Y(u2__abc_44228_n22459) );
  AND2X2 AND2X2_11335 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n7267), .Y(u2__abc_44228_n22461) );
  AND2X2 AND2X2_11336 ( .A(u2__abc_44228_n22462), .B(u2__abc_44228_n2972_bF_buf13), .Y(u2__abc_44228_n22463) );
  AND2X2 AND2X2_11337 ( .A(u2__abc_44228_n22460), .B(u2__abc_44228_n22463), .Y(u2__abc_44228_n22464) );
  AND2X2 AND2X2_11338 ( .A(u2__abc_44228_n22465), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_root_391__FF_INPUT) );
  AND2X2 AND2X2_11339 ( .A(u2__abc_44228_n3062_bF_buf87), .B(u2_o_391_), .Y(u2__abc_44228_n22467) );
  AND2X2 AND2X2_1134 ( .A(u2__abc_44228_n4288), .B(u2__abc_44228_n3740_1), .Y(u2__abc_44228_n4289) );
  AND2X2 AND2X2_11340 ( .A(u2__abc_44228_n22457), .B(u2_o_390_), .Y(u2__abc_44228_n22469) );
  AND2X2 AND2X2_11341 ( .A(u2__abc_44228_n22470), .B(u2__abc_44228_n22468), .Y(u2__abc_44228_n22471) );
  AND2X2 AND2X2_11342 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n7273), .Y(u2__abc_44228_n22473) );
  AND2X2 AND2X2_11343 ( .A(u2__abc_44228_n22474), .B(u2__abc_44228_n2972_bF_buf12), .Y(u2__abc_44228_n22475) );
  AND2X2 AND2X2_11344 ( .A(u2__abc_44228_n22472), .B(u2__abc_44228_n22475), .Y(u2__abc_44228_n22476) );
  AND2X2 AND2X2_11345 ( .A(u2__abc_44228_n22477), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_root_392__FF_INPUT) );
  AND2X2 AND2X2_11346 ( .A(u2__abc_44228_n3062_bF_buf86), .B(u2_o_392_), .Y(u2__abc_44228_n22479) );
  AND2X2 AND2X2_11347 ( .A(u2__abc_44228_n22469), .B(u2_o_391_), .Y(u2__abc_44228_n22481) );
  AND2X2 AND2X2_11348 ( .A(u2__abc_44228_n22482), .B(u2__abc_44228_n22480), .Y(u2__abc_44228_n22483) );
  AND2X2 AND2X2_11349 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n7260), .Y(u2__abc_44228_n22485) );
  AND2X2 AND2X2_1135 ( .A(u2__abc_44228_n4290), .B(u2__abc_44228_n3737), .Y(u2__abc_44228_n4291_1) );
  AND2X2 AND2X2_11350 ( .A(u2__abc_44228_n22486), .B(u2__abc_44228_n2972_bF_buf11), .Y(u2__abc_44228_n22487) );
  AND2X2 AND2X2_11351 ( .A(u2__abc_44228_n22484), .B(u2__abc_44228_n22487), .Y(u2__abc_44228_n22488) );
  AND2X2 AND2X2_11352 ( .A(u2__abc_44228_n22489), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_root_393__FF_INPUT) );
  AND2X2 AND2X2_11353 ( .A(u2__abc_44228_n3062_bF_buf85), .B(u2_o_393_), .Y(u2__abc_44228_n22491) );
  AND2X2 AND2X2_11354 ( .A(u2__abc_44228_n22481), .B(u2_o_392_), .Y(u2__abc_44228_n22493) );
  AND2X2 AND2X2_11355 ( .A(u2__abc_44228_n22494), .B(u2__abc_44228_n22492), .Y(u2__abc_44228_n22495) );
  AND2X2 AND2X2_11356 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n7253), .Y(u2__abc_44228_n22497) );
  AND2X2 AND2X2_11357 ( .A(u2__abc_44228_n22498), .B(u2__abc_44228_n2972_bF_buf10), .Y(u2__abc_44228_n22499) );
  AND2X2 AND2X2_11358 ( .A(u2__abc_44228_n22496), .B(u2__abc_44228_n22499), .Y(u2__abc_44228_n22500) );
  AND2X2 AND2X2_11359 ( .A(u2__abc_44228_n22501), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_root_394__FF_INPUT) );
  AND2X2 AND2X2_1136 ( .A(u2__abc_44228_n3729), .B(u2__abc_44228_n3732_1), .Y(u2__abc_44228_n4292) );
  AND2X2 AND2X2_11360 ( .A(u2__abc_44228_n3062_bF_buf84), .B(u2_o_394_), .Y(u2__abc_44228_n22503) );
  AND2X2 AND2X2_11361 ( .A(u2__abc_44228_n22493), .B(u2_o_393_), .Y(u2__abc_44228_n22505) );
  AND2X2 AND2X2_11362 ( .A(u2__abc_44228_n22506), .B(u2__abc_44228_n22504), .Y(u2__abc_44228_n22507) );
  AND2X2 AND2X2_11363 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n7238), .Y(u2__abc_44228_n22509) );
  AND2X2 AND2X2_11364 ( .A(u2__abc_44228_n22510), .B(u2__abc_44228_n2972_bF_buf9), .Y(u2__abc_44228_n22511) );
  AND2X2 AND2X2_11365 ( .A(u2__abc_44228_n22508), .B(u2__abc_44228_n22511), .Y(u2__abc_44228_n22512) );
  AND2X2 AND2X2_11366 ( .A(u2__abc_44228_n22513), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_root_395__FF_INPUT) );
  AND2X2 AND2X2_11367 ( .A(u2__abc_44228_n3062_bF_buf83), .B(u2_o_395_), .Y(u2__abc_44228_n22515) );
  AND2X2 AND2X2_11368 ( .A(u2__abc_44228_n22505), .B(u2_o_394_), .Y(u2__abc_44228_n22517) );
  AND2X2 AND2X2_11369 ( .A(u2__abc_44228_n22518), .B(u2__abc_44228_n22516), .Y(u2__abc_44228_n22519) );
  AND2X2 AND2X2_1137 ( .A(u2__abc_44228_n4295), .B(u2__abc_44228_n3723_1), .Y(u2__abc_44228_n4296) );
  AND2X2 AND2X2_11370 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n7244_1), .Y(u2__abc_44228_n22521) );
  AND2X2 AND2X2_11371 ( .A(u2__abc_44228_n22522), .B(u2__abc_44228_n2972_bF_buf8), .Y(u2__abc_44228_n22523) );
  AND2X2 AND2X2_11372 ( .A(u2__abc_44228_n22520), .B(u2__abc_44228_n22523), .Y(u2__abc_44228_n22524) );
  AND2X2 AND2X2_11373 ( .A(u2__abc_44228_n22525), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_root_396__FF_INPUT) );
  AND2X2 AND2X2_11374 ( .A(u2__abc_44228_n3062_bF_buf82), .B(u2_o_396_), .Y(u2__abc_44228_n22527) );
  AND2X2 AND2X2_11375 ( .A(u2__abc_44228_n22517), .B(u2_o_395_), .Y(u2__abc_44228_n22529) );
  AND2X2 AND2X2_11376 ( .A(u2__abc_44228_n22530), .B(u2__abc_44228_n22528), .Y(u2__abc_44228_n22531) );
  AND2X2 AND2X2_11377 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n7231), .Y(u2__abc_44228_n22533) );
  AND2X2 AND2X2_11378 ( .A(u2__abc_44228_n22534), .B(u2__abc_44228_n2972_bF_buf7), .Y(u2__abc_44228_n22535) );
  AND2X2 AND2X2_11379 ( .A(u2__abc_44228_n22532), .B(u2__abc_44228_n22535), .Y(u2__abc_44228_n22536) );
  AND2X2 AND2X2_1138 ( .A(u2__abc_44228_n4301), .B(u2_remHi_253_), .Y(u2__abc_44228_n4302) );
  AND2X2 AND2X2_11380 ( .A(u2__abc_44228_n22537), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_root_397__FF_INPUT) );
  AND2X2 AND2X2_11381 ( .A(u2__abc_44228_n3062_bF_buf81), .B(u2_o_397_), .Y(u2__abc_44228_n22539) );
  AND2X2 AND2X2_11382 ( .A(u2__abc_44228_n22529), .B(u2_o_396_), .Y(u2__abc_44228_n22541) );
  AND2X2 AND2X2_11383 ( .A(u2__abc_44228_n22542), .B(u2__abc_44228_n22540), .Y(u2__abc_44228_n22543) );
  AND2X2 AND2X2_11384 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n7224), .Y(u2__abc_44228_n22545) );
  AND2X2 AND2X2_11385 ( .A(u2__abc_44228_n22546), .B(u2__abc_44228_n2972_bF_buf6), .Y(u2__abc_44228_n22547) );
  AND2X2 AND2X2_11386 ( .A(u2__abc_44228_n22544), .B(u2__abc_44228_n22547), .Y(u2__abc_44228_n22548) );
  AND2X2 AND2X2_11387 ( .A(u2__abc_44228_n22549), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_root_398__FF_INPUT) );
  AND2X2 AND2X2_11388 ( .A(u2__abc_44228_n3062_bF_buf80), .B(u2_o_398_), .Y(u2__abc_44228_n22551) );
  AND2X2 AND2X2_11389 ( .A(u2__abc_44228_n22541), .B(u2_o_397_), .Y(u2__abc_44228_n22553) );
  AND2X2 AND2X2_1139 ( .A(u2__abc_44228_n4304), .B(u2_o_253_), .Y(u2__abc_44228_n4305) );
  AND2X2 AND2X2_11390 ( .A(u2__abc_44228_n22554), .B(u2__abc_44228_n22552), .Y(u2__abc_44228_n22555) );
  AND2X2 AND2X2_11391 ( .A(u2__abc_44228_n2983_bF_buf104), .B(u2__abc_44228_n7207), .Y(u2__abc_44228_n22557) );
  AND2X2 AND2X2_11392 ( .A(u2__abc_44228_n22558), .B(u2__abc_44228_n2972_bF_buf5), .Y(u2__abc_44228_n22559) );
  AND2X2 AND2X2_11393 ( .A(u2__abc_44228_n22556), .B(u2__abc_44228_n22559), .Y(u2__abc_44228_n22560) );
  AND2X2 AND2X2_11394 ( .A(u2__abc_44228_n22561), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_root_399__FF_INPUT) );
  AND2X2 AND2X2_11395 ( .A(u2__abc_44228_n3062_bF_buf79), .B(u2_o_399_), .Y(u2__abc_44228_n22563) );
  AND2X2 AND2X2_11396 ( .A(u2__abc_44228_n22553), .B(u2_o_398_), .Y(u2__abc_44228_n22565) );
  AND2X2 AND2X2_11397 ( .A(u2__abc_44228_n22566), .B(u2__abc_44228_n22564), .Y(u2__abc_44228_n22567) );
  AND2X2 AND2X2_11398 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n7213), .Y(u2__abc_44228_n22569) );
  AND2X2 AND2X2_11399 ( .A(u2__abc_44228_n22570), .B(u2__abc_44228_n2972_bF_buf4), .Y(u2__abc_44228_n22571) );
  AND2X2 AND2X2_114 ( .A(_abc_64468_n942), .B(_abc_64468_n941), .Y(_auto_iopadmap_cc_313_execute_65414_149_) );
  AND2X2 AND2X2_1140 ( .A(u2__abc_44228_n4303), .B(u2__abc_44228_n4306), .Y(u2__abc_44228_n4307) );
  AND2X2 AND2X2_11400 ( .A(u2__abc_44228_n22568), .B(u2__abc_44228_n22571), .Y(u2__abc_44228_n22572) );
  AND2X2 AND2X2_11401 ( .A(u2__abc_44228_n22573), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_root_400__FF_INPUT) );
  AND2X2 AND2X2_11402 ( .A(u2__abc_44228_n3062_bF_buf78), .B(u2_o_400_), .Y(u2__abc_44228_n22575) );
  AND2X2 AND2X2_11403 ( .A(u2__abc_44228_n22565), .B(u2_o_399_), .Y(u2__abc_44228_n22577) );
  AND2X2 AND2X2_11404 ( .A(u2__abc_44228_n22578), .B(u2__abc_44228_n22576), .Y(u2__abc_44228_n22579) );
  AND2X2 AND2X2_11405 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n7200), .Y(u2__abc_44228_n22581) );
  AND2X2 AND2X2_11406 ( .A(u2__abc_44228_n22582), .B(u2__abc_44228_n2972_bF_buf3), .Y(u2__abc_44228_n22583) );
  AND2X2 AND2X2_11407 ( .A(u2__abc_44228_n22580), .B(u2__abc_44228_n22583), .Y(u2__abc_44228_n22584) );
  AND2X2 AND2X2_11408 ( .A(u2__abc_44228_n22585), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_root_401__FF_INPUT) );
  AND2X2 AND2X2_11409 ( .A(u2__abc_44228_n3062_bF_buf77), .B(u2_o_401_), .Y(u2__abc_44228_n22587) );
  AND2X2 AND2X2_1141 ( .A(u2__abc_44228_n4308), .B(u2_remHi_252_), .Y(u2__abc_44228_n4309) );
  AND2X2 AND2X2_11410 ( .A(u2__abc_44228_n22577), .B(u2_o_400_), .Y(u2__abc_44228_n22589) );
  AND2X2 AND2X2_11411 ( .A(u2__abc_44228_n22590), .B(u2__abc_44228_n22588), .Y(u2__abc_44228_n22591) );
  AND2X2 AND2X2_11412 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n7193), .Y(u2__abc_44228_n22593) );
  AND2X2 AND2X2_11413 ( .A(u2__abc_44228_n22594), .B(u2__abc_44228_n2972_bF_buf2), .Y(u2__abc_44228_n22595) );
  AND2X2 AND2X2_11414 ( .A(u2__abc_44228_n22592), .B(u2__abc_44228_n22595), .Y(u2__abc_44228_n22596) );
  AND2X2 AND2X2_11415 ( .A(u2__abc_44228_n22597), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_root_402__FF_INPUT) );
  AND2X2 AND2X2_11416 ( .A(u2__abc_44228_n3062_bF_buf76), .B(u2_o_402_), .Y(u2__abc_44228_n22599) );
  AND2X2 AND2X2_11417 ( .A(u2__abc_44228_n22589), .B(u2_o_401_), .Y(u2__abc_44228_n22601) );
  AND2X2 AND2X2_11418 ( .A(u2__abc_44228_n22602), .B(u2__abc_44228_n22600), .Y(u2__abc_44228_n22603) );
  AND2X2 AND2X2_11419 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n7185), .Y(u2__abc_44228_n22605) );
  AND2X2 AND2X2_1142 ( .A(u2__abc_44228_n4310_1), .B(u2_o_252_), .Y(u2__abc_44228_n4311) );
  AND2X2 AND2X2_11420 ( .A(u2__abc_44228_n22606), .B(u2__abc_44228_n2972_bF_buf1), .Y(u2__abc_44228_n22607) );
  AND2X2 AND2X2_11421 ( .A(u2__abc_44228_n22604), .B(u2__abc_44228_n22607), .Y(u2__abc_44228_n22608) );
  AND2X2 AND2X2_11422 ( .A(u2__abc_44228_n22609), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_root_403__FF_INPUT) );
  AND2X2 AND2X2_11423 ( .A(u2__abc_44228_n3062_bF_buf75), .B(u2_o_403_), .Y(u2__abc_44228_n22611) );
  AND2X2 AND2X2_11424 ( .A(u2__abc_44228_n22601), .B(u2_o_402_), .Y(u2__abc_44228_n22613) );
  AND2X2 AND2X2_11425 ( .A(u2__abc_44228_n22614), .B(u2__abc_44228_n22612), .Y(u2__abc_44228_n22615) );
  AND2X2 AND2X2_11426 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n7178), .Y(u2__abc_44228_n22617) );
  AND2X2 AND2X2_11427 ( .A(u2__abc_44228_n22618), .B(u2__abc_44228_n2972_bF_buf0), .Y(u2__abc_44228_n22619) );
  AND2X2 AND2X2_11428 ( .A(u2__abc_44228_n22616), .B(u2__abc_44228_n22619), .Y(u2__abc_44228_n22620) );
  AND2X2 AND2X2_11429 ( .A(u2__abc_44228_n22621), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_root_404__FF_INPUT) );
  AND2X2 AND2X2_1143 ( .A(u2__abc_44228_n4313), .B(u2__abc_44228_n4307), .Y(u2__abc_44228_n4314) );
  AND2X2 AND2X2_11430 ( .A(u2__abc_44228_n3062_bF_buf74), .B(u2_o_404_), .Y(u2__abc_44228_n22623) );
  AND2X2 AND2X2_11431 ( .A(u2__abc_44228_n22613), .B(u2_o_403_), .Y(u2__abc_44228_n22625) );
  AND2X2 AND2X2_11432 ( .A(u2__abc_44228_n22626), .B(u2__abc_44228_n22624), .Y(u2__abc_44228_n22627) );
  AND2X2 AND2X2_11433 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n7171), .Y(u2__abc_44228_n22629) );
  AND2X2 AND2X2_11434 ( .A(u2__abc_44228_n22630), .B(u2__abc_44228_n2972_bF_buf107), .Y(u2__abc_44228_n22631) );
  AND2X2 AND2X2_11435 ( .A(u2__abc_44228_n22628), .B(u2__abc_44228_n22631), .Y(u2__abc_44228_n22632) );
  AND2X2 AND2X2_11436 ( .A(u2__abc_44228_n22633), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_root_405__FF_INPUT) );
  AND2X2 AND2X2_11437 ( .A(u2__abc_44228_n3062_bF_buf73), .B(u2_o_405_), .Y(u2__abc_44228_n22635) );
  AND2X2 AND2X2_11438 ( .A(u2__abc_44228_n22625), .B(u2_o_404_), .Y(u2__abc_44228_n22637) );
  AND2X2 AND2X2_11439 ( .A(u2__abc_44228_n22638), .B(u2__abc_44228_n22636), .Y(u2__abc_44228_n22639) );
  AND2X2 AND2X2_1144 ( .A(u2__abc_44228_n4315), .B(u2_remHi_250_), .Y(u2__abc_44228_n4316) );
  AND2X2 AND2X2_11440 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n7164), .Y(u2__abc_44228_n22641) );
  AND2X2 AND2X2_11441 ( .A(u2__abc_44228_n22642), .B(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n22643) );
  AND2X2 AND2X2_11442 ( .A(u2__abc_44228_n22640), .B(u2__abc_44228_n22643), .Y(u2__abc_44228_n22644) );
  AND2X2 AND2X2_11443 ( .A(u2__abc_44228_n22645), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_root_406__FF_INPUT) );
  AND2X2 AND2X2_11444 ( .A(u2__abc_44228_n3062_bF_buf72), .B(u2_o_406_), .Y(u2__abc_44228_n22647) );
  AND2X2 AND2X2_11445 ( .A(u2__abc_44228_n22637), .B(u2_o_405_), .Y(u2__abc_44228_n22649) );
  AND2X2 AND2X2_11446 ( .A(u2__abc_44228_n22650), .B(u2__abc_44228_n22648), .Y(u2__abc_44228_n22651) );
  AND2X2 AND2X2_11447 ( .A(u2__abc_44228_n2983_bF_buf88), .B(u2__abc_44228_n7155), .Y(u2__abc_44228_n22653) );
  AND2X2 AND2X2_11448 ( .A(u2__abc_44228_n22654), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n22655) );
  AND2X2 AND2X2_11449 ( .A(u2__abc_44228_n22652), .B(u2__abc_44228_n22655), .Y(u2__abc_44228_n22656) );
  AND2X2 AND2X2_1145 ( .A(u2__abc_44228_n4317), .B(u2_o_250_), .Y(u2__abc_44228_n4318) );
  AND2X2 AND2X2_11450 ( .A(u2__abc_44228_n22657), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_root_407__FF_INPUT) );
  AND2X2 AND2X2_11451 ( .A(u2__abc_44228_n3062_bF_buf71), .B(u2_o_407_), .Y(u2__abc_44228_n22659) );
  AND2X2 AND2X2_11452 ( .A(u2__abc_44228_n22649), .B(u2_o_406_), .Y(u2__abc_44228_n22661) );
  AND2X2 AND2X2_11453 ( .A(u2__abc_44228_n22662), .B(u2__abc_44228_n22660), .Y(u2__abc_44228_n22663) );
  AND2X2 AND2X2_11454 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n7148), .Y(u2__abc_44228_n22665) );
  AND2X2 AND2X2_11455 ( .A(u2__abc_44228_n22666), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n22667) );
  AND2X2 AND2X2_11456 ( .A(u2__abc_44228_n22664), .B(u2__abc_44228_n22667), .Y(u2__abc_44228_n22668) );
  AND2X2 AND2X2_11457 ( .A(u2__abc_44228_n22669), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_root_408__FF_INPUT) );
  AND2X2 AND2X2_11458 ( .A(u2__abc_44228_n3062_bF_buf70), .B(u2_o_408_), .Y(u2__abc_44228_n22671) );
  AND2X2 AND2X2_11459 ( .A(u2__abc_44228_n22661), .B(u2_o_407_), .Y(u2__abc_44228_n22673) );
  AND2X2 AND2X2_1146 ( .A(u2__abc_44228_n4321), .B(u2_remHi_251_), .Y(u2__abc_44228_n4322) );
  AND2X2 AND2X2_11460 ( .A(u2__abc_44228_n22674), .B(u2__abc_44228_n22672), .Y(u2__abc_44228_n22675) );
  AND2X2 AND2X2_11461 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n7141), .Y(u2__abc_44228_n22677) );
  AND2X2 AND2X2_11462 ( .A(u2__abc_44228_n22678), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n22679) );
  AND2X2 AND2X2_11463 ( .A(u2__abc_44228_n22676), .B(u2__abc_44228_n22679), .Y(u2__abc_44228_n22680) );
  AND2X2 AND2X2_11464 ( .A(u2__abc_44228_n22681), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_root_409__FF_INPUT) );
  AND2X2 AND2X2_11465 ( .A(u2__abc_44228_n3062_bF_buf69), .B(u2_o_409_), .Y(u2__abc_44228_n22683) );
  AND2X2 AND2X2_11466 ( .A(u2__abc_44228_n22673), .B(u2_o_408_), .Y(u2__abc_44228_n22685) );
  AND2X2 AND2X2_11467 ( .A(u2__abc_44228_n22686), .B(u2__abc_44228_n22684), .Y(u2__abc_44228_n22687) );
  AND2X2 AND2X2_11468 ( .A(u2__abc_44228_n2983_bF_buf82), .B(u2__abc_44228_n7134_1), .Y(u2__abc_44228_n22689) );
  AND2X2 AND2X2_11469 ( .A(u2__abc_44228_n22690), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n22691) );
  AND2X2 AND2X2_1147 ( .A(u2__abc_44228_n4324), .B(u2_o_251_), .Y(u2__abc_44228_n4325) );
  AND2X2 AND2X2_11470 ( .A(u2__abc_44228_n22688), .B(u2__abc_44228_n22691), .Y(u2__abc_44228_n22692) );
  AND2X2 AND2X2_11471 ( .A(u2__abc_44228_n22693), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_root_410__FF_INPUT) );
  AND2X2 AND2X2_11472 ( .A(u2__abc_44228_n3062_bF_buf68), .B(u2_o_410_), .Y(u2__abc_44228_n22695) );
  AND2X2 AND2X2_11473 ( .A(u2__abc_44228_n22685), .B(u2_o_409_), .Y(u2__abc_44228_n22697) );
  AND2X2 AND2X2_11474 ( .A(u2__abc_44228_n22698), .B(u2__abc_44228_n22696), .Y(u2__abc_44228_n22699) );
  AND2X2 AND2X2_11475 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n7126), .Y(u2__abc_44228_n22701) );
  AND2X2 AND2X2_11476 ( .A(u2__abc_44228_n22702), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n22703) );
  AND2X2 AND2X2_11477 ( .A(u2__abc_44228_n22700), .B(u2__abc_44228_n22703), .Y(u2__abc_44228_n22704) );
  AND2X2 AND2X2_11478 ( .A(u2__abc_44228_n22705), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_root_411__FF_INPUT) );
  AND2X2 AND2X2_11479 ( .A(u2__abc_44228_n3062_bF_buf67), .B(u2_o_411_), .Y(u2__abc_44228_n22707) );
  AND2X2 AND2X2_1148 ( .A(u2__abc_44228_n4323), .B(u2__abc_44228_n4326), .Y(u2__abc_44228_n4327) );
  AND2X2 AND2X2_11480 ( .A(u2__abc_44228_n22697), .B(u2_o_410_), .Y(u2__abc_44228_n22709) );
  AND2X2 AND2X2_11481 ( .A(u2__abc_44228_n22710), .B(u2__abc_44228_n22708), .Y(u2__abc_44228_n22711) );
  AND2X2 AND2X2_11482 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n7119), .Y(u2__abc_44228_n22713) );
  AND2X2 AND2X2_11483 ( .A(u2__abc_44228_n22714), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n22715) );
  AND2X2 AND2X2_11484 ( .A(u2__abc_44228_n22712), .B(u2__abc_44228_n22715), .Y(u2__abc_44228_n22716) );
  AND2X2 AND2X2_11485 ( .A(u2__abc_44228_n22717), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_root_412__FF_INPUT) );
  AND2X2 AND2X2_11486 ( .A(u2__abc_44228_n3062_bF_buf66), .B(u2_o_412_), .Y(u2__abc_44228_n22719) );
  AND2X2 AND2X2_11487 ( .A(u2__abc_44228_n22709), .B(u2_o_411_), .Y(u2__abc_44228_n22721) );
  AND2X2 AND2X2_11488 ( .A(u2__abc_44228_n22722), .B(u2__abc_44228_n22720), .Y(u2__abc_44228_n22723) );
  AND2X2 AND2X2_11489 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n7112), .Y(u2__abc_44228_n22725) );
  AND2X2 AND2X2_1149 ( .A(u2__abc_44228_n4320_1), .B(u2__abc_44228_n4327), .Y(u2__abc_44228_n4328) );
  AND2X2 AND2X2_11490 ( .A(u2__abc_44228_n22726), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n22727) );
  AND2X2 AND2X2_11491 ( .A(u2__abc_44228_n22724), .B(u2__abc_44228_n22727), .Y(u2__abc_44228_n22728) );
  AND2X2 AND2X2_11492 ( .A(u2__abc_44228_n22729), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_root_413__FF_INPUT) );
  AND2X2 AND2X2_11493 ( .A(u2__abc_44228_n3062_bF_buf65), .B(u2_o_413_), .Y(u2__abc_44228_n22731) );
  AND2X2 AND2X2_11494 ( .A(u2__abc_44228_n22721), .B(u2_o_412_), .Y(u2__abc_44228_n22733) );
  AND2X2 AND2X2_11495 ( .A(u2__abc_44228_n22734), .B(u2__abc_44228_n22732), .Y(u2__abc_44228_n22735) );
  AND2X2 AND2X2_11496 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n7105), .Y(u2__abc_44228_n22737) );
  AND2X2 AND2X2_11497 ( .A(u2__abc_44228_n22738), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n22739) );
  AND2X2 AND2X2_11498 ( .A(u2__abc_44228_n22736), .B(u2__abc_44228_n22739), .Y(u2__abc_44228_n22740) );
  AND2X2 AND2X2_11499 ( .A(u2__abc_44228_n22741), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_root_414__FF_INPUT) );
  AND2X2 AND2X2_115 ( .A(_abc_64468_n945), .B(_abc_64468_n944), .Y(_auto_iopadmap_cc_313_execute_65414_150_) );
  AND2X2 AND2X2_1150 ( .A(u2__abc_44228_n4314), .B(u2__abc_44228_n4328), .Y(u2__abc_44228_n4329_1) );
  AND2X2 AND2X2_11500 ( .A(u2__abc_44228_n3062_bF_buf64), .B(u2_o_414_), .Y(u2__abc_44228_n22743) );
  AND2X2 AND2X2_11501 ( .A(u2__abc_44228_n22733), .B(u2_o_413_), .Y(u2__abc_44228_n22745) );
  AND2X2 AND2X2_11502 ( .A(u2__abc_44228_n22746), .B(u2__abc_44228_n22744), .Y(u2__abc_44228_n22747) );
  AND2X2 AND2X2_11503 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n7087), .Y(u2__abc_44228_n22749) );
  AND2X2 AND2X2_11504 ( .A(u2__abc_44228_n22750), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n22751) );
  AND2X2 AND2X2_11505 ( .A(u2__abc_44228_n22748), .B(u2__abc_44228_n22751), .Y(u2__abc_44228_n22752) );
  AND2X2 AND2X2_11506 ( .A(u2__abc_44228_n22753), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_root_415__FF_INPUT) );
  AND2X2 AND2X2_11507 ( .A(u2__abc_44228_n3062_bF_buf63), .B(u2_o_415_), .Y(u2__abc_44228_n22755) );
  AND2X2 AND2X2_11508 ( .A(u2__abc_44228_n22745), .B(u2_o_414_), .Y(u2__abc_44228_n22757) );
  AND2X2 AND2X2_11509 ( .A(u2__abc_44228_n22758), .B(u2__abc_44228_n22756), .Y(u2__abc_44228_n22759) );
  AND2X2 AND2X2_1151 ( .A(u2__abc_44228_n4330), .B(u2_remHi_249_), .Y(u2__abc_44228_n4331) );
  AND2X2 AND2X2_11510 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n7093), .Y(u2__abc_44228_n22761) );
  AND2X2 AND2X2_11511 ( .A(u2__abc_44228_n22762), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n22763) );
  AND2X2 AND2X2_11512 ( .A(u2__abc_44228_n22760), .B(u2__abc_44228_n22763), .Y(u2__abc_44228_n22764) );
  AND2X2 AND2X2_11513 ( .A(u2__abc_44228_n22765), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_root_416__FF_INPUT) );
  AND2X2 AND2X2_11514 ( .A(u2__abc_44228_n3062_bF_buf62), .B(u2_o_416_), .Y(u2__abc_44228_n22767) );
  AND2X2 AND2X2_11515 ( .A(u2__abc_44228_n22757), .B(u2_o_415_), .Y(u2__abc_44228_n22769) );
  AND2X2 AND2X2_11516 ( .A(u2__abc_44228_n22770), .B(u2__abc_44228_n22768), .Y(u2__abc_44228_n22771) );
  AND2X2 AND2X2_11517 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n7080), .Y(u2__abc_44228_n22773) );
  AND2X2 AND2X2_11518 ( .A(u2__abc_44228_n22774), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n22775) );
  AND2X2 AND2X2_11519 ( .A(u2__abc_44228_n22772), .B(u2__abc_44228_n22775), .Y(u2__abc_44228_n22776) );
  AND2X2 AND2X2_1152 ( .A(u2__abc_44228_n4333), .B(u2_o_249_), .Y(u2__abc_44228_n4334) );
  AND2X2 AND2X2_11520 ( .A(u2__abc_44228_n22777), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_root_417__FF_INPUT) );
  AND2X2 AND2X2_11521 ( .A(u2__abc_44228_n3062_bF_buf61), .B(u2_o_417_), .Y(u2__abc_44228_n22779) );
  AND2X2 AND2X2_11522 ( .A(u2__abc_44228_n22769), .B(u2_o_416_), .Y(u2__abc_44228_n22781) );
  AND2X2 AND2X2_11523 ( .A(u2__abc_44228_n22782), .B(u2__abc_44228_n22780), .Y(u2__abc_44228_n22783) );
  AND2X2 AND2X2_11524 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n7073), .Y(u2__abc_44228_n22785) );
  AND2X2 AND2X2_11525 ( .A(u2__abc_44228_n22786), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n22787) );
  AND2X2 AND2X2_11526 ( .A(u2__abc_44228_n22784), .B(u2__abc_44228_n22787), .Y(u2__abc_44228_n22788) );
  AND2X2 AND2X2_11527 ( .A(u2__abc_44228_n22789), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_root_418__FF_INPUT) );
  AND2X2 AND2X2_11528 ( .A(u2__abc_44228_n3062_bF_buf60), .B(u2_o_418_), .Y(u2__abc_44228_n22791) );
  AND2X2 AND2X2_11529 ( .A(u2__abc_44228_n22781), .B(u2_o_417_), .Y(u2__abc_44228_n22793) );
  AND2X2 AND2X2_1153 ( .A(u2__abc_44228_n4332), .B(u2__abc_44228_n4335), .Y(u2__abc_44228_n4336) );
  AND2X2 AND2X2_11530 ( .A(u2__abc_44228_n22794), .B(u2__abc_44228_n22792), .Y(u2__abc_44228_n22795) );
  AND2X2 AND2X2_11531 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n7065), .Y(u2__abc_44228_n22797) );
  AND2X2 AND2X2_11532 ( .A(u2__abc_44228_n22798), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n22799) );
  AND2X2 AND2X2_11533 ( .A(u2__abc_44228_n22796), .B(u2__abc_44228_n22799), .Y(u2__abc_44228_n22800) );
  AND2X2 AND2X2_11534 ( .A(u2__abc_44228_n22801), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_root_419__FF_INPUT) );
  AND2X2 AND2X2_11535 ( .A(u2__abc_44228_n3062_bF_buf59), .B(u2_o_419_), .Y(u2__abc_44228_n22803) );
  AND2X2 AND2X2_11536 ( .A(u2__abc_44228_n22793), .B(u2_o_418_), .Y(u2__abc_44228_n22805) );
  AND2X2 AND2X2_11537 ( .A(u2__abc_44228_n22806), .B(u2__abc_44228_n22804), .Y(u2__abc_44228_n22807) );
  AND2X2 AND2X2_11538 ( .A(u2__abc_44228_n2983_bF_buf62), .B(u2__abc_44228_n7058), .Y(u2__abc_44228_n22809) );
  AND2X2 AND2X2_11539 ( .A(u2__abc_44228_n22810), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n22811) );
  AND2X2 AND2X2_1154 ( .A(u2__abc_44228_n4337), .B(u2_remHi_248_), .Y(u2__abc_44228_n4338_1) );
  AND2X2 AND2X2_11540 ( .A(u2__abc_44228_n22808), .B(u2__abc_44228_n22811), .Y(u2__abc_44228_n22812) );
  AND2X2 AND2X2_11541 ( .A(u2__abc_44228_n22813), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_root_420__FF_INPUT) );
  AND2X2 AND2X2_11542 ( .A(u2__abc_44228_n3062_bF_buf58), .B(u2_o_420_), .Y(u2__abc_44228_n22815) );
  AND2X2 AND2X2_11543 ( .A(u2__abc_44228_n22805), .B(u2_o_419_), .Y(u2__abc_44228_n22817) );
  AND2X2 AND2X2_11544 ( .A(u2__abc_44228_n22818), .B(u2__abc_44228_n22816), .Y(u2__abc_44228_n22819) );
  AND2X2 AND2X2_11545 ( .A(u2__abc_44228_n2983_bF_buf60), .B(u2__abc_44228_n7051), .Y(u2__abc_44228_n22821) );
  AND2X2 AND2X2_11546 ( .A(u2__abc_44228_n22822), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n22823) );
  AND2X2 AND2X2_11547 ( .A(u2__abc_44228_n22820), .B(u2__abc_44228_n22823), .Y(u2__abc_44228_n22824) );
  AND2X2 AND2X2_11548 ( .A(u2__abc_44228_n22825), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_root_421__FF_INPUT) );
  AND2X2 AND2X2_11549 ( .A(u2__abc_44228_n3062_bF_buf57), .B(u2_o_421_), .Y(u2__abc_44228_n22827) );
  AND2X2 AND2X2_1155 ( .A(u2__abc_44228_n4339), .B(u2_o_248_), .Y(u2__abc_44228_n4340) );
  AND2X2 AND2X2_11550 ( .A(u2__abc_44228_n22817), .B(u2_o_420_), .Y(u2__abc_44228_n22829) );
  AND2X2 AND2X2_11551 ( .A(u2__abc_44228_n22830), .B(u2__abc_44228_n22828), .Y(u2__abc_44228_n22831) );
  AND2X2 AND2X2_11552 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n7044), .Y(u2__abc_44228_n22833) );
  AND2X2 AND2X2_11553 ( .A(u2__abc_44228_n22834), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n22835) );
  AND2X2 AND2X2_11554 ( .A(u2__abc_44228_n22832), .B(u2__abc_44228_n22835), .Y(u2__abc_44228_n22836) );
  AND2X2 AND2X2_11555 ( .A(u2__abc_44228_n22837), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_root_422__FF_INPUT) );
  AND2X2 AND2X2_11556 ( .A(u2__abc_44228_n3062_bF_buf56), .B(u2_o_422_), .Y(u2__abc_44228_n22839) );
  AND2X2 AND2X2_11557 ( .A(u2__abc_44228_n22829), .B(u2_o_421_), .Y(u2__abc_44228_n22841) );
  AND2X2 AND2X2_11558 ( .A(u2__abc_44228_n22842), .B(u2__abc_44228_n22840), .Y(u2__abc_44228_n22843) );
  AND2X2 AND2X2_11559 ( .A(u2__abc_44228_n2983_bF_buf56), .B(u2__abc_44228_n7035), .Y(u2__abc_44228_n22845) );
  AND2X2 AND2X2_1156 ( .A(u2__abc_44228_n4342), .B(u2__abc_44228_n4336), .Y(u2__abc_44228_n4343) );
  AND2X2 AND2X2_11560 ( .A(u2__abc_44228_n22846), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n22847) );
  AND2X2 AND2X2_11561 ( .A(u2__abc_44228_n22844), .B(u2__abc_44228_n22847), .Y(u2__abc_44228_n22848) );
  AND2X2 AND2X2_11562 ( .A(u2__abc_44228_n22849), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_root_423__FF_INPUT) );
  AND2X2 AND2X2_11563 ( .A(u2__abc_44228_n3062_bF_buf55), .B(u2_o_423_), .Y(u2__abc_44228_n22851) );
  AND2X2 AND2X2_11564 ( .A(u2__abc_44228_n22841), .B(u2_o_422_), .Y(u2__abc_44228_n22853) );
  AND2X2 AND2X2_11565 ( .A(u2__abc_44228_n22854), .B(u2__abc_44228_n22852), .Y(u2__abc_44228_n22855) );
  AND2X2 AND2X2_11566 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n7028), .Y(u2__abc_44228_n22857) );
  AND2X2 AND2X2_11567 ( .A(u2__abc_44228_n22858), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n22859) );
  AND2X2 AND2X2_11568 ( .A(u2__abc_44228_n22856), .B(u2__abc_44228_n22859), .Y(u2__abc_44228_n22860) );
  AND2X2 AND2X2_11569 ( .A(u2__abc_44228_n22861), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_root_424__FF_INPUT) );
  AND2X2 AND2X2_1157 ( .A(u2__abc_44228_n4344), .B(u2_remHi_246_), .Y(u2__abc_44228_n4345) );
  AND2X2 AND2X2_11570 ( .A(u2__abc_44228_n3062_bF_buf54), .B(u2_o_424_), .Y(u2__abc_44228_n22863) );
  AND2X2 AND2X2_11571 ( .A(u2__abc_44228_n22853), .B(u2_o_423_), .Y(u2__abc_44228_n22865) );
  AND2X2 AND2X2_11572 ( .A(u2__abc_44228_n22866), .B(u2__abc_44228_n22864), .Y(u2__abc_44228_n22867) );
  AND2X2 AND2X2_11573 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n7021), .Y(u2__abc_44228_n22869) );
  AND2X2 AND2X2_11574 ( .A(u2__abc_44228_n22870), .B(u2__abc_44228_n2972_bF_buf87), .Y(u2__abc_44228_n22871) );
  AND2X2 AND2X2_11575 ( .A(u2__abc_44228_n22868), .B(u2__abc_44228_n22871), .Y(u2__abc_44228_n22872) );
  AND2X2 AND2X2_11576 ( .A(u2__abc_44228_n22873), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_root_425__FF_INPUT) );
  AND2X2 AND2X2_11577 ( .A(u2__abc_44228_n3062_bF_buf53), .B(u2_o_425_), .Y(u2__abc_44228_n22875) );
  AND2X2 AND2X2_11578 ( .A(u2__abc_44228_n22865), .B(u2_o_424_), .Y(u2__abc_44228_n22877) );
  AND2X2 AND2X2_11579 ( .A(u2__abc_44228_n22878), .B(u2__abc_44228_n22876), .Y(u2__abc_44228_n22879) );
  AND2X2 AND2X2_1158 ( .A(u2__abc_44228_n4346), .B(u2_o_246_), .Y(u2__abc_44228_n4347) );
  AND2X2 AND2X2_11580 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2__abc_44228_n7014_1), .Y(u2__abc_44228_n22881) );
  AND2X2 AND2X2_11581 ( .A(u2__abc_44228_n22882), .B(u2__abc_44228_n2972_bF_buf86), .Y(u2__abc_44228_n22883) );
  AND2X2 AND2X2_11582 ( .A(u2__abc_44228_n22880), .B(u2__abc_44228_n22883), .Y(u2__abc_44228_n22884) );
  AND2X2 AND2X2_11583 ( .A(u2__abc_44228_n22885), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_root_426__FF_INPUT) );
  AND2X2 AND2X2_11584 ( .A(u2__abc_44228_n3062_bF_buf52), .B(u2_o_426_), .Y(u2__abc_44228_n22887) );
  AND2X2 AND2X2_11585 ( .A(u2__abc_44228_n22877), .B(u2_o_425_), .Y(u2__abc_44228_n22889) );
  AND2X2 AND2X2_11586 ( .A(u2__abc_44228_n22890), .B(u2__abc_44228_n22888), .Y(u2__abc_44228_n22891) );
  AND2X2 AND2X2_11587 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n7006), .Y(u2__abc_44228_n22893) );
  AND2X2 AND2X2_11588 ( .A(u2__abc_44228_n22894), .B(u2__abc_44228_n2972_bF_buf85), .Y(u2__abc_44228_n22895) );
  AND2X2 AND2X2_11589 ( .A(u2__abc_44228_n22892), .B(u2__abc_44228_n22895), .Y(u2__abc_44228_n22896) );
  AND2X2 AND2X2_1159 ( .A(u2__abc_44228_n4350), .B(u2_remHi_247_), .Y(u2__abc_44228_n4351) );
  AND2X2 AND2X2_11590 ( .A(u2__abc_44228_n22897), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_root_427__FF_INPUT) );
  AND2X2 AND2X2_11591 ( .A(u2__abc_44228_n3062_bF_buf51), .B(u2_o_427_), .Y(u2__abc_44228_n22899) );
  AND2X2 AND2X2_11592 ( .A(u2__abc_44228_n22889), .B(u2_o_426_), .Y(u2__abc_44228_n22901) );
  AND2X2 AND2X2_11593 ( .A(u2__abc_44228_n22902), .B(u2__abc_44228_n22900), .Y(u2__abc_44228_n22903) );
  AND2X2 AND2X2_11594 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n6999), .Y(u2__abc_44228_n22905) );
  AND2X2 AND2X2_11595 ( .A(u2__abc_44228_n22906), .B(u2__abc_44228_n2972_bF_buf84), .Y(u2__abc_44228_n22907) );
  AND2X2 AND2X2_11596 ( .A(u2__abc_44228_n22904), .B(u2__abc_44228_n22907), .Y(u2__abc_44228_n22908) );
  AND2X2 AND2X2_11597 ( .A(u2__abc_44228_n22909), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_root_428__FF_INPUT) );
  AND2X2 AND2X2_11598 ( .A(u2__abc_44228_n3062_bF_buf50), .B(u2_o_428_), .Y(u2__abc_44228_n22911) );
  AND2X2 AND2X2_11599 ( .A(u2__abc_44228_n22901), .B(u2_o_427_), .Y(u2__abc_44228_n22913) );
  AND2X2 AND2X2_116 ( .A(_abc_64468_n948), .B(_abc_64468_n947), .Y(_auto_iopadmap_cc_313_execute_65414_151_) );
  AND2X2 AND2X2_1160 ( .A(u2__abc_44228_n4353), .B(u2_o_247_), .Y(u2__abc_44228_n4354) );
  AND2X2 AND2X2_11600 ( .A(u2__abc_44228_n22914), .B(u2__abc_44228_n22912), .Y(u2__abc_44228_n22915) );
  AND2X2 AND2X2_11601 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n6992), .Y(u2__abc_44228_n22917) );
  AND2X2 AND2X2_11602 ( .A(u2__abc_44228_n22918), .B(u2__abc_44228_n2972_bF_buf83), .Y(u2__abc_44228_n22919) );
  AND2X2 AND2X2_11603 ( .A(u2__abc_44228_n22916), .B(u2__abc_44228_n22919), .Y(u2__abc_44228_n22920) );
  AND2X2 AND2X2_11604 ( .A(u2__abc_44228_n22921), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_root_429__FF_INPUT) );
  AND2X2 AND2X2_11605 ( .A(u2__abc_44228_n3062_bF_buf49), .B(u2_o_429_), .Y(u2__abc_44228_n22923) );
  AND2X2 AND2X2_11606 ( .A(u2__abc_44228_n22913), .B(u2_o_428_), .Y(u2__abc_44228_n22925) );
  AND2X2 AND2X2_11607 ( .A(u2__abc_44228_n22926), .B(u2__abc_44228_n22924), .Y(u2__abc_44228_n22927) );
  AND2X2 AND2X2_11608 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n6985), .Y(u2__abc_44228_n22929) );
  AND2X2 AND2X2_11609 ( .A(u2__abc_44228_n22930), .B(u2__abc_44228_n2972_bF_buf82), .Y(u2__abc_44228_n22931) );
  AND2X2 AND2X2_1161 ( .A(u2__abc_44228_n4352), .B(u2__abc_44228_n4355), .Y(u2__abc_44228_n4356) );
  AND2X2 AND2X2_11610 ( .A(u2__abc_44228_n22928), .B(u2__abc_44228_n22931), .Y(u2__abc_44228_n22932) );
  AND2X2 AND2X2_11611 ( .A(u2__abc_44228_n22933), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_root_430__FF_INPUT) );
  AND2X2 AND2X2_11612 ( .A(u2__abc_44228_n3062_bF_buf48), .B(u2_o_430_), .Y(u2__abc_44228_n22935) );
  AND2X2 AND2X2_11613 ( .A(u2__abc_44228_n22925), .B(u2_o_429_), .Y(u2__abc_44228_n22937) );
  AND2X2 AND2X2_11614 ( .A(u2__abc_44228_n22938), .B(u2__abc_44228_n22936), .Y(u2__abc_44228_n22939) );
  AND2X2 AND2X2_11615 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n6961_1), .Y(u2__abc_44228_n22941) );
  AND2X2 AND2X2_11616 ( .A(u2__abc_44228_n22942), .B(u2__abc_44228_n2972_bF_buf81), .Y(u2__abc_44228_n22943) );
  AND2X2 AND2X2_11617 ( .A(u2__abc_44228_n22940), .B(u2__abc_44228_n22943), .Y(u2__abc_44228_n22944) );
  AND2X2 AND2X2_11618 ( .A(u2__abc_44228_n22945), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_root_431__FF_INPUT) );
  AND2X2 AND2X2_11619 ( .A(u2__abc_44228_n3062_bF_buf47), .B(u2_o_431_), .Y(u2__abc_44228_n22947) );
  AND2X2 AND2X2_1162 ( .A(u2__abc_44228_n4349_1), .B(u2__abc_44228_n4356), .Y(u2__abc_44228_n4357) );
  AND2X2 AND2X2_11620 ( .A(u2__abc_44228_n22937), .B(u2_o_430_), .Y(u2__abc_44228_n22949) );
  AND2X2 AND2X2_11621 ( .A(u2__abc_44228_n22950), .B(u2__abc_44228_n22948), .Y(u2__abc_44228_n22951) );
  AND2X2 AND2X2_11622 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n6954), .Y(u2__abc_44228_n22953) );
  AND2X2 AND2X2_11623 ( .A(u2__abc_44228_n22954), .B(u2__abc_44228_n2972_bF_buf80), .Y(u2__abc_44228_n22955) );
  AND2X2 AND2X2_11624 ( .A(u2__abc_44228_n22952), .B(u2__abc_44228_n22955), .Y(u2__abc_44228_n22956) );
  AND2X2 AND2X2_11625 ( .A(u2__abc_44228_n22957), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_root_432__FF_INPUT) );
  AND2X2 AND2X2_11626 ( .A(u2__abc_44228_n3062_bF_buf46), .B(u2_o_432_), .Y(u2__abc_44228_n22959) );
  AND2X2 AND2X2_11627 ( .A(u2__abc_44228_n22949), .B(u2_o_431_), .Y(u2__abc_44228_n22961) );
  AND2X2 AND2X2_11628 ( .A(u2__abc_44228_n22962), .B(u2__abc_44228_n22960), .Y(u2__abc_44228_n22963) );
  AND2X2 AND2X2_11629 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n6975), .Y(u2__abc_44228_n22965) );
  AND2X2 AND2X2_1163 ( .A(u2__abc_44228_n4343), .B(u2__abc_44228_n4357), .Y(u2__abc_44228_n4358) );
  AND2X2 AND2X2_11630 ( .A(u2__abc_44228_n22966), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n22967) );
  AND2X2 AND2X2_11631 ( .A(u2__abc_44228_n22964), .B(u2__abc_44228_n22967), .Y(u2__abc_44228_n22968) );
  AND2X2 AND2X2_11632 ( .A(u2__abc_44228_n22969), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_root_433__FF_INPUT) );
  AND2X2 AND2X2_11633 ( .A(u2__abc_44228_n3062_bF_buf45), .B(u2_o_433_), .Y(u2__abc_44228_n22971) );
  AND2X2 AND2X2_11634 ( .A(u2__abc_44228_n22961), .B(u2_o_432_), .Y(u2__abc_44228_n22973) );
  AND2X2 AND2X2_11635 ( .A(u2__abc_44228_n22974), .B(u2__abc_44228_n22972), .Y(u2__abc_44228_n22975) );
  AND2X2 AND2X2_11636 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n6968), .Y(u2__abc_44228_n22977) );
  AND2X2 AND2X2_11637 ( .A(u2__abc_44228_n22978), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n22979) );
  AND2X2 AND2X2_11638 ( .A(u2__abc_44228_n22976), .B(u2__abc_44228_n22979), .Y(u2__abc_44228_n22980) );
  AND2X2 AND2X2_11639 ( .A(u2__abc_44228_n22981), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_root_434__FF_INPUT) );
  AND2X2 AND2X2_1164 ( .A(u2__abc_44228_n4329_1), .B(u2__abc_44228_n4358), .Y(u2__abc_44228_n4359_1) );
  AND2X2 AND2X2_11640 ( .A(u2__abc_44228_n3062_bF_buf44), .B(u2_o_434_), .Y(u2__abc_44228_n22983) );
  AND2X2 AND2X2_11641 ( .A(u2__abc_44228_n22973), .B(u2_o_433_), .Y(u2__abc_44228_n22985) );
  AND2X2 AND2X2_11642 ( .A(u2__abc_44228_n22986), .B(u2__abc_44228_n22984), .Y(u2__abc_44228_n22987) );
  AND2X2 AND2X2_11643 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n6939), .Y(u2__abc_44228_n22989) );
  AND2X2 AND2X2_11644 ( .A(u2__abc_44228_n22990), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n22991) );
  AND2X2 AND2X2_11645 ( .A(u2__abc_44228_n22988), .B(u2__abc_44228_n22991), .Y(u2__abc_44228_n22992) );
  AND2X2 AND2X2_11646 ( .A(u2__abc_44228_n22993), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_root_435__FF_INPUT) );
  AND2X2 AND2X2_11647 ( .A(u2__abc_44228_n3062_bF_buf43), .B(u2_o_435_), .Y(u2__abc_44228_n22995) );
  AND2X2 AND2X2_11648 ( .A(u2__abc_44228_n22985), .B(u2_o_434_), .Y(u2__abc_44228_n22997) );
  AND2X2 AND2X2_11649 ( .A(u2__abc_44228_n22998), .B(u2__abc_44228_n22996), .Y(u2__abc_44228_n22999) );
  AND2X2 AND2X2_1165 ( .A(u2__abc_44228_n4360), .B(u2_remHi_245_), .Y(u2__abc_44228_n4361) );
  AND2X2 AND2X2_11650 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n6945), .Y(u2__abc_44228_n23001) );
  AND2X2 AND2X2_11651 ( .A(u2__abc_44228_n23002), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n23003) );
  AND2X2 AND2X2_11652 ( .A(u2__abc_44228_n23000), .B(u2__abc_44228_n23003), .Y(u2__abc_44228_n23004) );
  AND2X2 AND2X2_11653 ( .A(u2__abc_44228_n23005), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_root_436__FF_INPUT) );
  AND2X2 AND2X2_11654 ( .A(u2__abc_44228_n3062_bF_buf42), .B(u2_o_436_), .Y(u2__abc_44228_n23007) );
  AND2X2 AND2X2_11655 ( .A(u2__abc_44228_n22997), .B(u2_o_435_), .Y(u2__abc_44228_n23009) );
  AND2X2 AND2X2_11656 ( .A(u2__abc_44228_n23010), .B(u2__abc_44228_n23008), .Y(u2__abc_44228_n23011) );
  AND2X2 AND2X2_11657 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n6932), .Y(u2__abc_44228_n23013) );
  AND2X2 AND2X2_11658 ( .A(u2__abc_44228_n23014), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n23015) );
  AND2X2 AND2X2_11659 ( .A(u2__abc_44228_n23012), .B(u2__abc_44228_n23015), .Y(u2__abc_44228_n23016) );
  AND2X2 AND2X2_1166 ( .A(u2__abc_44228_n4363), .B(u2_o_245_), .Y(u2__abc_44228_n4364) );
  AND2X2 AND2X2_11660 ( .A(u2__abc_44228_n23017), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_root_437__FF_INPUT) );
  AND2X2 AND2X2_11661 ( .A(u2__abc_44228_n3062_bF_buf41), .B(u2_o_437_), .Y(u2__abc_44228_n23019) );
  AND2X2 AND2X2_11662 ( .A(u2__abc_44228_n23009), .B(u2_o_436_), .Y(u2__abc_44228_n23021) );
  AND2X2 AND2X2_11663 ( .A(u2__abc_44228_n23022), .B(u2__abc_44228_n23020), .Y(u2__abc_44228_n23023) );
  AND2X2 AND2X2_11664 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n6925), .Y(u2__abc_44228_n23025) );
  AND2X2 AND2X2_11665 ( .A(u2__abc_44228_n23026), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n23027) );
  AND2X2 AND2X2_11666 ( .A(u2__abc_44228_n23024), .B(u2__abc_44228_n23027), .Y(u2__abc_44228_n23028) );
  AND2X2 AND2X2_11667 ( .A(u2__abc_44228_n23029), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_root_438__FF_INPUT) );
  AND2X2 AND2X2_11668 ( .A(u2__abc_44228_n3062_bF_buf40), .B(u2_o_438_), .Y(u2__abc_44228_n23031) );
  AND2X2 AND2X2_11669 ( .A(u2__abc_44228_n23021), .B(u2_o_437_), .Y(u2__abc_44228_n23033) );
  AND2X2 AND2X2_1167 ( .A(u2__abc_44228_n4362), .B(u2__abc_44228_n4365), .Y(u2__abc_44228_n4366) );
  AND2X2 AND2X2_11670 ( .A(u2__abc_44228_n23034), .B(u2__abc_44228_n23032), .Y(u2__abc_44228_n23035) );
  AND2X2 AND2X2_11671 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n6916), .Y(u2__abc_44228_n23037) );
  AND2X2 AND2X2_11672 ( .A(u2__abc_44228_n23038), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n23039) );
  AND2X2 AND2X2_11673 ( .A(u2__abc_44228_n23036), .B(u2__abc_44228_n23039), .Y(u2__abc_44228_n23040) );
  AND2X2 AND2X2_11674 ( .A(u2__abc_44228_n23041), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_root_439__FF_INPUT) );
  AND2X2 AND2X2_11675 ( .A(u2__abc_44228_n3062_bF_buf39), .B(u2_o_439_), .Y(u2__abc_44228_n23043) );
  AND2X2 AND2X2_11676 ( .A(u2__abc_44228_n23033), .B(u2_o_438_), .Y(u2__abc_44228_n23045) );
  AND2X2 AND2X2_11677 ( .A(u2__abc_44228_n23046), .B(u2__abc_44228_n23044), .Y(u2__abc_44228_n23047) );
  AND2X2 AND2X2_11678 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n6909), .Y(u2__abc_44228_n23049) );
  AND2X2 AND2X2_11679 ( .A(u2__abc_44228_n23050), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n23051) );
  AND2X2 AND2X2_1168 ( .A(u2__abc_44228_n4367), .B(u2_remHi_244_), .Y(u2__abc_44228_n4368_1) );
  AND2X2 AND2X2_11680 ( .A(u2__abc_44228_n23048), .B(u2__abc_44228_n23051), .Y(u2__abc_44228_n23052) );
  AND2X2 AND2X2_11681 ( .A(u2__abc_44228_n23053), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_root_440__FF_INPUT) );
  AND2X2 AND2X2_11682 ( .A(u2__abc_44228_n3062_bF_buf38), .B(u2_o_440_), .Y(u2__abc_44228_n23055) );
  AND2X2 AND2X2_11683 ( .A(u2__abc_44228_n23045), .B(u2_o_439_), .Y(u2__abc_44228_n23057) );
  AND2X2 AND2X2_11684 ( .A(u2__abc_44228_n23058), .B(u2__abc_44228_n23056), .Y(u2__abc_44228_n23059) );
  AND2X2 AND2X2_11685 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n6902), .Y(u2__abc_44228_n23061) );
  AND2X2 AND2X2_11686 ( .A(u2__abc_44228_n23062), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n23063) );
  AND2X2 AND2X2_11687 ( .A(u2__abc_44228_n23060), .B(u2__abc_44228_n23063), .Y(u2__abc_44228_n23064) );
  AND2X2 AND2X2_11688 ( .A(u2__abc_44228_n23065), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_root_441__FF_INPUT) );
  AND2X2 AND2X2_11689 ( .A(u2__abc_44228_n3062_bF_buf37), .B(u2_o_441_), .Y(u2__abc_44228_n23067) );
  AND2X2 AND2X2_1169 ( .A(u2__abc_44228_n4369), .B(u2_o_244_), .Y(u2__abc_44228_n4370) );
  AND2X2 AND2X2_11690 ( .A(u2__abc_44228_n23057), .B(u2_o_440_), .Y(u2__abc_44228_n23069) );
  AND2X2 AND2X2_11691 ( .A(u2__abc_44228_n23070), .B(u2__abc_44228_n23068), .Y(u2__abc_44228_n23071) );
  AND2X2 AND2X2_11692 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n6895), .Y(u2__abc_44228_n23073) );
  AND2X2 AND2X2_11693 ( .A(u2__abc_44228_n23074), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n23075) );
  AND2X2 AND2X2_11694 ( .A(u2__abc_44228_n23072), .B(u2__abc_44228_n23075), .Y(u2__abc_44228_n23076) );
  AND2X2 AND2X2_11695 ( .A(u2__abc_44228_n23077), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_root_442__FF_INPUT) );
  AND2X2 AND2X2_11696 ( .A(u2__abc_44228_n3062_bF_buf36), .B(u2_o_442_), .Y(u2__abc_44228_n23079) );
  AND2X2 AND2X2_11697 ( .A(u2__abc_44228_n23069), .B(u2_o_441_), .Y(u2__abc_44228_n23081) );
  AND2X2 AND2X2_11698 ( .A(u2__abc_44228_n23082), .B(u2__abc_44228_n23080), .Y(u2__abc_44228_n23083) );
  AND2X2 AND2X2_11699 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n6887_1), .Y(u2__abc_44228_n23085) );
  AND2X2 AND2X2_117 ( .A(_abc_64468_n951), .B(_abc_64468_n950), .Y(_auto_iopadmap_cc_313_execute_65414_152_) );
  AND2X2 AND2X2_1170 ( .A(u2__abc_44228_n4372), .B(u2__abc_44228_n4366), .Y(u2__abc_44228_n4373) );
  AND2X2 AND2X2_11700 ( .A(u2__abc_44228_n23086), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n23087) );
  AND2X2 AND2X2_11701 ( .A(u2__abc_44228_n23084), .B(u2__abc_44228_n23087), .Y(u2__abc_44228_n23088) );
  AND2X2 AND2X2_11702 ( .A(u2__abc_44228_n23089), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_root_443__FF_INPUT) );
  AND2X2 AND2X2_11703 ( .A(u2__abc_44228_n3062_bF_buf35), .B(u2_o_443_), .Y(u2__abc_44228_n23091) );
  AND2X2 AND2X2_11704 ( .A(u2__abc_44228_n23081), .B(u2_o_442_), .Y(u2__abc_44228_n23093) );
  AND2X2 AND2X2_11705 ( .A(u2__abc_44228_n23094), .B(u2__abc_44228_n23092), .Y(u2__abc_44228_n23095) );
  AND2X2 AND2X2_11706 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n6880), .Y(u2__abc_44228_n23097) );
  AND2X2 AND2X2_11707 ( .A(u2__abc_44228_n23098), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n23099) );
  AND2X2 AND2X2_11708 ( .A(u2__abc_44228_n23096), .B(u2__abc_44228_n23099), .Y(u2__abc_44228_n23100) );
  AND2X2 AND2X2_11709 ( .A(u2__abc_44228_n23101), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_root_444__FF_INPUT) );
  AND2X2 AND2X2_1171 ( .A(u2__abc_44228_n4374), .B(u2_remHi_242_), .Y(u2__abc_44228_n4375) );
  AND2X2 AND2X2_11710 ( .A(u2__abc_44228_n3062_bF_buf34), .B(u2_o_444_), .Y(u2__abc_44228_n23103) );
  AND2X2 AND2X2_11711 ( .A(u2__abc_44228_n23093), .B(u2_o_443_), .Y(u2__abc_44228_n23105) );
  AND2X2 AND2X2_11712 ( .A(u2__abc_44228_n23106), .B(u2__abc_44228_n23104), .Y(u2__abc_44228_n23107) );
  AND2X2 AND2X2_11713 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n6873), .Y(u2__abc_44228_n23109) );
  AND2X2 AND2X2_11714 ( .A(u2__abc_44228_n23110), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n23111) );
  AND2X2 AND2X2_11715 ( .A(u2__abc_44228_n23108), .B(u2__abc_44228_n23111), .Y(u2__abc_44228_n23112) );
  AND2X2 AND2X2_11716 ( .A(u2__abc_44228_n23113), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_root_445__FF_INPUT) );
  AND2X2 AND2X2_11717 ( .A(u2__abc_44228_n3062_bF_buf33), .B(u2_o_445_), .Y(u2__abc_44228_n23115) );
  AND2X2 AND2X2_11718 ( .A(u2__abc_44228_n23105), .B(u2_o_444_), .Y(u2__abc_44228_n23117) );
  AND2X2 AND2X2_11719 ( .A(u2__abc_44228_n23118), .B(u2__abc_44228_n23116), .Y(u2__abc_44228_n23119) );
  AND2X2 AND2X2_1172 ( .A(u2__abc_44228_n4376), .B(u2_o_242_), .Y(u2__abc_44228_n4377_1) );
  AND2X2 AND2X2_11720 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n6866), .Y(u2__abc_44228_n23121) );
  AND2X2 AND2X2_11721 ( .A(u2__abc_44228_n23122), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n23123) );
  AND2X2 AND2X2_11722 ( .A(u2__abc_44228_n23120), .B(u2__abc_44228_n23123), .Y(u2__abc_44228_n23124) );
  AND2X2 AND2X2_11723 ( .A(u2__abc_44228_n23125), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_root_446__FF_INPUT) );
  AND2X2 AND2X2_11724 ( .A(u2__abc_44228_n3062_bF_buf32), .B(u2_o_446_), .Y(u2__abc_44228_n23127) );
  AND2X2 AND2X2_11725 ( .A(u2__abc_44228_n23117), .B(u2_o_445_), .Y(u2__abc_44228_n23129) );
  AND2X2 AND2X2_11726 ( .A(u2__abc_44228_n23130), .B(u2__abc_44228_n23128), .Y(u2__abc_44228_n23131) );
  AND2X2 AND2X2_11727 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n7523), .Y(u2__abc_44228_n23133) );
  AND2X2 AND2X2_11728 ( .A(u2__abc_44228_n23134), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n23135) );
  AND2X2 AND2X2_11729 ( .A(u2__abc_44228_n23132), .B(u2__abc_44228_n23135), .Y(u2__abc_44228_n23136) );
  AND2X2 AND2X2_1173 ( .A(u2__abc_44228_n4380), .B(u2_remHi_243_), .Y(u2__abc_44228_n4381) );
  AND2X2 AND2X2_11730 ( .A(u2__abc_44228_n23137), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_root_447__FF_INPUT) );
  AND2X2 AND2X2_11731 ( .A(u2__abc_44228_n3062_bF_buf31), .B(u2_o_447_), .Y(u2__abc_44228_n23139) );
  AND2X2 AND2X2_11732 ( .A(u2__abc_44228_n23129), .B(u2_o_446_), .Y(u2__abc_44228_n23141) );
  AND2X2 AND2X2_11733 ( .A(u2__abc_44228_n23142), .B(u2__abc_44228_n23140), .Y(u2__abc_44228_n23143) );
  AND2X2 AND2X2_11734 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n7529), .Y(u2__abc_44228_n23145) );
  AND2X2 AND2X2_11735 ( .A(u2__abc_44228_n23146), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n23147) );
  AND2X2 AND2X2_11736 ( .A(u2__abc_44228_n23144), .B(u2__abc_44228_n23147), .Y(u2__abc_44228_n23148) );
  AND2X2 AND2X2_11737 ( .A(u2__abc_44228_n23149), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_root_448__FF_INPUT) );
  AND2X2 AND2X2_11738 ( .A(u2__abc_44228_n3062_bF_buf30), .B(u2_o_448_), .Y(u2__abc_44228_n23151) );
  AND2X2 AND2X2_11739 ( .A(u2__abc_44228_n23141), .B(u2_o_447_), .Y(u2__abc_44228_n23153) );
  AND2X2 AND2X2_1174 ( .A(u2__abc_44228_n4383), .B(u2_o_243_), .Y(u2__abc_44228_n4384) );
  AND2X2 AND2X2_11740 ( .A(u2__abc_44228_n23154), .B(u2__abc_44228_n23152), .Y(u2__abc_44228_n23155) );
  AND2X2 AND2X2_11741 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n7516), .Y(u2__abc_44228_n23157) );
  AND2X2 AND2X2_11742 ( .A(u2__abc_44228_n23158), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n23159) );
  AND2X2 AND2X2_11743 ( .A(u2__abc_44228_n23156), .B(u2__abc_44228_n23159), .Y(u2__abc_44228_n23160) );
  AND2X2 AND2X2_11744 ( .A(u2__abc_44228_n23161), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_root_449__FF_INPUT) );
  AND2X2 AND2X2_11745 ( .A(u2__abc_44228_n3062_bF_buf29), .B(u2_o_449_), .Y(u2__abc_44228_n23163) );
  AND2X2 AND2X2_11746 ( .A(u2__abc_44228_n23153), .B(u2_o_448_), .Y(u2__abc_44228_n23165) );
  AND2X2 AND2X2_11747 ( .A(u2__abc_44228_n23166), .B(u2__abc_44228_n23164), .Y(u2__abc_44228_n23167) );
  AND2X2 AND2X2_11748 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n7509), .Y(u2__abc_44228_n23169) );
  AND2X2 AND2X2_11749 ( .A(u2__abc_44228_n23170), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n23171) );
  AND2X2 AND2X2_1175 ( .A(u2__abc_44228_n4382), .B(u2__abc_44228_n4385), .Y(u2__abc_44228_n4386_1) );
  AND2X2 AND2X2_11750 ( .A(u2__abc_44228_n23168), .B(u2__abc_44228_n23171), .Y(u2__abc_44228_n23172) );
  AND2X2 AND2X2_11751 ( .A(u2__abc_44228_n23173), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_root_450__FF_INPUT) );
  AND2X2 AND2X2_1176 ( .A(u2__abc_44228_n4379), .B(u2__abc_44228_n4386_1), .Y(u2__abc_44228_n4387) );
  AND2X2 AND2X2_1177 ( .A(u2__abc_44228_n4373), .B(u2__abc_44228_n4387), .Y(u2__abc_44228_n4388) );
  AND2X2 AND2X2_1178 ( .A(u2__abc_44228_n4389), .B(u2_remHi_241_), .Y(u2__abc_44228_n4390) );
  AND2X2 AND2X2_1179 ( .A(u2__abc_44228_n4392), .B(u2_o_241_), .Y(u2__abc_44228_n4393) );
  AND2X2 AND2X2_118 ( .A(_abc_64468_n954), .B(_abc_64468_n953), .Y(_auto_iopadmap_cc_313_execute_65414_153_) );
  AND2X2 AND2X2_1180 ( .A(u2__abc_44228_n4391), .B(u2__abc_44228_n4394), .Y(u2__abc_44228_n4395) );
  AND2X2 AND2X2_1181 ( .A(u2__abc_44228_n4396_1), .B(u2_remHi_240_), .Y(u2__abc_44228_n4397) );
  AND2X2 AND2X2_1182 ( .A(u2__abc_44228_n4398), .B(u2_o_240_), .Y(u2__abc_44228_n4399) );
  AND2X2 AND2X2_1183 ( .A(u2__abc_44228_n4401), .B(u2__abc_44228_n4395), .Y(u2__abc_44228_n4402) );
  AND2X2 AND2X2_1184 ( .A(u2__abc_44228_n4403), .B(u2_remHi_238_), .Y(u2__abc_44228_n4404) );
  AND2X2 AND2X2_1185 ( .A(u2__abc_44228_n4405_1), .B(u2_o_238_), .Y(u2__abc_44228_n4406) );
  AND2X2 AND2X2_1186 ( .A(u2__abc_44228_n4409), .B(u2_remHi_239_), .Y(u2__abc_44228_n4410) );
  AND2X2 AND2X2_1187 ( .A(u2__abc_44228_n4412), .B(u2_o_239_), .Y(u2__abc_44228_n4413) );
  AND2X2 AND2X2_1188 ( .A(u2__abc_44228_n4411), .B(u2__abc_44228_n4414_1), .Y(u2__abc_44228_n4415) );
  AND2X2 AND2X2_1189 ( .A(u2__abc_44228_n4408), .B(u2__abc_44228_n4415), .Y(u2__abc_44228_n4416) );
  AND2X2 AND2X2_119 ( .A(_abc_64468_n957), .B(_abc_64468_n956), .Y(_auto_iopadmap_cc_313_execute_65414_154_) );
  AND2X2 AND2X2_1190 ( .A(u2__abc_44228_n4402), .B(u2__abc_44228_n4416), .Y(u2__abc_44228_n4417) );
  AND2X2 AND2X2_1191 ( .A(u2__abc_44228_n4388), .B(u2__abc_44228_n4417), .Y(u2__abc_44228_n4418) );
  AND2X2 AND2X2_1192 ( .A(u2__abc_44228_n4359_1), .B(u2__abc_44228_n4418), .Y(u2__abc_44228_n4419) );
  AND2X2 AND2X2_1193 ( .A(u2__abc_44228_n4420), .B(u2_remHi_237_), .Y(u2__abc_44228_n4421) );
  AND2X2 AND2X2_1194 ( .A(u2__abc_44228_n4423_1), .B(u2_o_237_), .Y(u2__abc_44228_n4424) );
  AND2X2 AND2X2_1195 ( .A(u2__abc_44228_n4422), .B(u2__abc_44228_n4425), .Y(u2__abc_44228_n4426) );
  AND2X2 AND2X2_1196 ( .A(u2__abc_44228_n4427), .B(u2_remHi_236_), .Y(u2__abc_44228_n4428) );
  AND2X2 AND2X2_1197 ( .A(u2__abc_44228_n4429), .B(u2_o_236_), .Y(u2__abc_44228_n4430) );
  AND2X2 AND2X2_1198 ( .A(u2__abc_44228_n4432_1), .B(u2__abc_44228_n4426), .Y(u2__abc_44228_n4433) );
  AND2X2 AND2X2_1199 ( .A(u2__abc_44228_n4434), .B(u2_remHi_234_), .Y(u2__abc_44228_n4435) );
  AND2X2 AND2X2_12 ( .A(_abc_64468_n753_bF_buf2), .B(sqrto_11_), .Y(_auto_iopadmap_cc_313_execute_65414_47_) );
  AND2X2 AND2X2_120 ( .A(_abc_64468_n960), .B(_abc_64468_n959), .Y(_auto_iopadmap_cc_313_execute_65414_155_) );
  AND2X2 AND2X2_1200 ( .A(u2__abc_44228_n4436), .B(u2_o_234_), .Y(u2__abc_44228_n4437) );
  AND2X2 AND2X2_1201 ( .A(u2__abc_44228_n4440), .B(u2_remHi_235_), .Y(u2__abc_44228_n4441) );
  AND2X2 AND2X2_1202 ( .A(u2__abc_44228_n4443), .B(u2_o_235_), .Y(u2__abc_44228_n4444) );
  AND2X2 AND2X2_1203 ( .A(u2__abc_44228_n4442_1), .B(u2__abc_44228_n4445), .Y(u2__abc_44228_n4446) );
  AND2X2 AND2X2_1204 ( .A(u2__abc_44228_n4439), .B(u2__abc_44228_n4446), .Y(u2__abc_44228_n4447) );
  AND2X2 AND2X2_1205 ( .A(u2__abc_44228_n4433), .B(u2__abc_44228_n4447), .Y(u2__abc_44228_n4448) );
  AND2X2 AND2X2_1206 ( .A(u2__abc_44228_n4449), .B(u2_remHi_231_), .Y(u2__abc_44228_n4450) );
  AND2X2 AND2X2_1207 ( .A(u2__abc_44228_n4452), .B(u2_o_231_), .Y(u2__abc_44228_n4453) );
  AND2X2 AND2X2_1208 ( .A(u2__abc_44228_n4451_1), .B(u2__abc_44228_n4454), .Y(u2__abc_44228_n4455) );
  AND2X2 AND2X2_1209 ( .A(u2__abc_44228_n4456), .B(u2_remHi_230_), .Y(u2__abc_44228_n4457) );
  AND2X2 AND2X2_121 ( .A(_abc_64468_n963), .B(_abc_64468_n962), .Y(_auto_iopadmap_cc_313_execute_65414_156_) );
  AND2X2 AND2X2_1210 ( .A(u2__abc_44228_n4458), .B(u2_o_230_), .Y(u2__abc_44228_n4459) );
  AND2X2 AND2X2_1211 ( .A(u2__abc_44228_n4461_1), .B(u2__abc_44228_n4455), .Y(u2__abc_44228_n4462) );
  AND2X2 AND2X2_1212 ( .A(u2__abc_44228_n4463), .B(u2_remHi_233_), .Y(u2__abc_44228_n4464) );
  AND2X2 AND2X2_1213 ( .A(u2__abc_44228_n4466), .B(u2_o_233_), .Y(u2__abc_44228_n4467) );
  AND2X2 AND2X2_1214 ( .A(u2__abc_44228_n4465), .B(u2__abc_44228_n4468), .Y(u2__abc_44228_n4469) );
  AND2X2 AND2X2_1215 ( .A(u2__abc_44228_n4470), .B(u2_remHi_232_), .Y(u2__abc_44228_n4471_1) );
  AND2X2 AND2X2_1216 ( .A(u2__abc_44228_n4472), .B(u2_o_232_), .Y(u2__abc_44228_n4473) );
  AND2X2 AND2X2_1217 ( .A(u2__abc_44228_n4475), .B(u2__abc_44228_n4469), .Y(u2__abc_44228_n4476) );
  AND2X2 AND2X2_1218 ( .A(u2__abc_44228_n4462), .B(u2__abc_44228_n4476), .Y(u2__abc_44228_n4477) );
  AND2X2 AND2X2_1219 ( .A(u2__abc_44228_n4448), .B(u2__abc_44228_n4477), .Y(u2__abc_44228_n4478) );
  AND2X2 AND2X2_122 ( .A(_abc_64468_n966), .B(_abc_64468_n965), .Y(_auto_iopadmap_cc_313_execute_65414_157_) );
  AND2X2 AND2X2_1220 ( .A(u2__abc_44228_n4479), .B(u2_remHi_229_), .Y(u2__abc_44228_n4480_1) );
  AND2X2 AND2X2_1221 ( .A(u2__abc_44228_n4482), .B(u2_o_229_), .Y(u2__abc_44228_n4483) );
  AND2X2 AND2X2_1222 ( .A(u2__abc_44228_n4481), .B(u2__abc_44228_n4484), .Y(u2__abc_44228_n4485) );
  AND2X2 AND2X2_1223 ( .A(u2__abc_44228_n4486), .B(u2_remHi_228_), .Y(u2__abc_44228_n4487) );
  AND2X2 AND2X2_1224 ( .A(u2__abc_44228_n4488), .B(u2_o_228_), .Y(u2__abc_44228_n4489_1) );
  AND2X2 AND2X2_1225 ( .A(u2__abc_44228_n4491), .B(u2__abc_44228_n4485), .Y(u2__abc_44228_n4492) );
  AND2X2 AND2X2_1226 ( .A(u2__abc_44228_n4493), .B(u2_remHi_226_), .Y(u2__abc_44228_n4494) );
  AND2X2 AND2X2_1227 ( .A(u2__abc_44228_n4495), .B(u2_o_226_), .Y(u2__abc_44228_n4496) );
  AND2X2 AND2X2_1228 ( .A(u2__abc_44228_n4499), .B(u2_remHi_227_), .Y(u2__abc_44228_n4500) );
  AND2X2 AND2X2_1229 ( .A(u2__abc_44228_n4502), .B(u2_o_227_), .Y(u2__abc_44228_n4503) );
  AND2X2 AND2X2_123 ( .A(_abc_64468_n969), .B(_abc_64468_n968), .Y(_auto_iopadmap_cc_313_execute_65414_158_) );
  AND2X2 AND2X2_1230 ( .A(u2__abc_44228_n4501), .B(u2__abc_44228_n4504), .Y(u2__abc_44228_n4505) );
  AND2X2 AND2X2_1231 ( .A(u2__abc_44228_n4498_1), .B(u2__abc_44228_n4505), .Y(u2__abc_44228_n4506) );
  AND2X2 AND2X2_1232 ( .A(u2__abc_44228_n4492), .B(u2__abc_44228_n4506), .Y(u2__abc_44228_n4507) );
  AND2X2 AND2X2_1233 ( .A(u2__abc_44228_n4508_1), .B(u2_remHi_225_), .Y(u2__abc_44228_n4509) );
  AND2X2 AND2X2_1234 ( .A(u2__abc_44228_n4511), .B(sqrto_225_), .Y(u2__abc_44228_n4512) );
  AND2X2 AND2X2_1235 ( .A(u2__abc_44228_n4510), .B(u2__abc_44228_n4513), .Y(u2__abc_44228_n4514) );
  AND2X2 AND2X2_1236 ( .A(u2__abc_44228_n4515), .B(u2_remHi_224_), .Y(u2__abc_44228_n4516) );
  AND2X2 AND2X2_1237 ( .A(u2__abc_44228_n4517_1), .B(sqrto_224_), .Y(u2__abc_44228_n4518) );
  AND2X2 AND2X2_1238 ( .A(u2__abc_44228_n4520), .B(u2__abc_44228_n4514), .Y(u2__abc_44228_n4521) );
  AND2X2 AND2X2_1239 ( .A(u2__abc_44228_n4522), .B(u2_remHi_222_), .Y(u2__abc_44228_n4523) );
  AND2X2 AND2X2_124 ( .A(_abc_64468_n972), .B(_abc_64468_n971), .Y(_auto_iopadmap_cc_313_execute_65414_159_) );
  AND2X2 AND2X2_1240 ( .A(u2__abc_44228_n4524), .B(sqrto_222_), .Y(u2__abc_44228_n4525) );
  AND2X2 AND2X2_1241 ( .A(u2__abc_44228_n4528), .B(u2_remHi_223_), .Y(u2__abc_44228_n4529) );
  AND2X2 AND2X2_1242 ( .A(u2__abc_44228_n4531), .B(sqrto_223_), .Y(u2__abc_44228_n4532) );
  AND2X2 AND2X2_1243 ( .A(u2__abc_44228_n4530), .B(u2__abc_44228_n4533), .Y(u2__abc_44228_n4534) );
  AND2X2 AND2X2_1244 ( .A(u2__abc_44228_n4527), .B(u2__abc_44228_n4534), .Y(u2__abc_44228_n4535_1) );
  AND2X2 AND2X2_1245 ( .A(u2__abc_44228_n4521), .B(u2__abc_44228_n4535_1), .Y(u2__abc_44228_n4536) );
  AND2X2 AND2X2_1246 ( .A(u2__abc_44228_n4507), .B(u2__abc_44228_n4536), .Y(u2__abc_44228_n4537) );
  AND2X2 AND2X2_1247 ( .A(u2__abc_44228_n4478), .B(u2__abc_44228_n4537), .Y(u2__abc_44228_n4538) );
  AND2X2 AND2X2_1248 ( .A(u2__abc_44228_n4419), .B(u2__abc_44228_n4538), .Y(u2__abc_44228_n4539) );
  AND2X2 AND2X2_1249 ( .A(u2__abc_44228_n4540), .B(u2_remHi_221_), .Y(u2__abc_44228_n4541) );
  AND2X2 AND2X2_125 ( .A(_abc_64468_n975), .B(_abc_64468_n974), .Y(_auto_iopadmap_cc_313_execute_65414_160_) );
  AND2X2 AND2X2_1250 ( .A(u2__abc_44228_n4543), .B(sqrto_221_), .Y(u2__abc_44228_n4544) );
  AND2X2 AND2X2_1251 ( .A(u2__abc_44228_n4542), .B(u2__abc_44228_n4545_1), .Y(u2__abc_44228_n4546) );
  AND2X2 AND2X2_1252 ( .A(u2__abc_44228_n4547), .B(u2_remHi_220_), .Y(u2__abc_44228_n4548) );
  AND2X2 AND2X2_1253 ( .A(u2__abc_44228_n4549), .B(sqrto_220_), .Y(u2__abc_44228_n4550) );
  AND2X2 AND2X2_1254 ( .A(u2__abc_44228_n4552), .B(u2__abc_44228_n4546), .Y(u2__abc_44228_n4553) );
  AND2X2 AND2X2_1255 ( .A(u2__abc_44228_n4554_1), .B(u2_remHi_218_), .Y(u2__abc_44228_n4555) );
  AND2X2 AND2X2_1256 ( .A(u2__abc_44228_n4556), .B(sqrto_218_), .Y(u2__abc_44228_n4557) );
  AND2X2 AND2X2_1257 ( .A(u2__abc_44228_n4560), .B(u2_remHi_219_), .Y(u2__abc_44228_n4561) );
  AND2X2 AND2X2_1258 ( .A(u2__abc_44228_n4563_1), .B(sqrto_219_), .Y(u2__abc_44228_n4564) );
  AND2X2 AND2X2_1259 ( .A(u2__abc_44228_n4562), .B(u2__abc_44228_n4565), .Y(u2__abc_44228_n4566) );
  AND2X2 AND2X2_126 ( .A(_abc_64468_n978), .B(_abc_64468_n977), .Y(_auto_iopadmap_cc_313_execute_65414_161_) );
  AND2X2 AND2X2_1260 ( .A(u2__abc_44228_n4559), .B(u2__abc_44228_n4566), .Y(u2__abc_44228_n4567) );
  AND2X2 AND2X2_1261 ( .A(u2__abc_44228_n4553), .B(u2__abc_44228_n4567), .Y(u2__abc_44228_n4568) );
  AND2X2 AND2X2_1262 ( .A(u2__abc_44228_n4569), .B(u2_remHi_217_), .Y(u2__abc_44228_n4570) );
  AND2X2 AND2X2_1263 ( .A(u2__abc_44228_n4572_1), .B(sqrto_217_), .Y(u2__abc_44228_n4573) );
  AND2X2 AND2X2_1264 ( .A(u2__abc_44228_n4571), .B(u2__abc_44228_n4574), .Y(u2__abc_44228_n4575) );
  AND2X2 AND2X2_1265 ( .A(u2__abc_44228_n4576), .B(u2_remHi_216_), .Y(u2__abc_44228_n4577) );
  AND2X2 AND2X2_1266 ( .A(u2__abc_44228_n4578), .B(sqrto_216_), .Y(u2__abc_44228_n4579) );
  AND2X2 AND2X2_1267 ( .A(u2__abc_44228_n4581_1), .B(u2__abc_44228_n4575), .Y(u2__abc_44228_n4582) );
  AND2X2 AND2X2_1268 ( .A(u2__abc_44228_n4583), .B(u2_remHi_214_), .Y(u2__abc_44228_n4584) );
  AND2X2 AND2X2_1269 ( .A(u2__abc_44228_n4585), .B(sqrto_214_), .Y(u2__abc_44228_n4586) );
  AND2X2 AND2X2_127 ( .A(_abc_64468_n981), .B(_abc_64468_n980), .Y(_auto_iopadmap_cc_313_execute_65414_162_) );
  AND2X2 AND2X2_1270 ( .A(u2__abc_44228_n4589), .B(u2_remHi_215_), .Y(u2__abc_44228_n4590) );
  AND2X2 AND2X2_1271 ( .A(u2__abc_44228_n4592), .B(sqrto_215_), .Y(u2__abc_44228_n4593) );
  AND2X2 AND2X2_1272 ( .A(u2__abc_44228_n4591_1), .B(u2__abc_44228_n4594), .Y(u2__abc_44228_n4595) );
  AND2X2 AND2X2_1273 ( .A(u2__abc_44228_n4588), .B(u2__abc_44228_n4595), .Y(u2__abc_44228_n4596) );
  AND2X2 AND2X2_1274 ( .A(u2__abc_44228_n4582), .B(u2__abc_44228_n4596), .Y(u2__abc_44228_n4597) );
  AND2X2 AND2X2_1275 ( .A(u2__abc_44228_n4568), .B(u2__abc_44228_n4597), .Y(u2__abc_44228_n4598) );
  AND2X2 AND2X2_1276 ( .A(u2__abc_44228_n4599), .B(u2_remHi_213_), .Y(u2__abc_44228_n4600_1) );
  AND2X2 AND2X2_1277 ( .A(u2__abc_44228_n4602), .B(sqrto_213_), .Y(u2__abc_44228_n4603) );
  AND2X2 AND2X2_1278 ( .A(u2__abc_44228_n4601), .B(u2__abc_44228_n4604), .Y(u2__abc_44228_n4605) );
  AND2X2 AND2X2_1279 ( .A(u2__abc_44228_n4606), .B(u2_remHi_212_), .Y(u2__abc_44228_n4607) );
  AND2X2 AND2X2_128 ( .A(_abc_64468_n984), .B(_abc_64468_n983), .Y(_auto_iopadmap_cc_313_execute_65414_163_) );
  AND2X2 AND2X2_1280 ( .A(u2__abc_44228_n4608), .B(sqrto_212_), .Y(u2__abc_44228_n4609) );
  AND2X2 AND2X2_1281 ( .A(u2__abc_44228_n4611), .B(u2__abc_44228_n4605), .Y(u2__abc_44228_n4612) );
  AND2X2 AND2X2_1282 ( .A(u2__abc_44228_n4613), .B(u2_remHi_210_), .Y(u2__abc_44228_n4614) );
  AND2X2 AND2X2_1283 ( .A(u2__abc_44228_n4615), .B(sqrto_210_), .Y(u2__abc_44228_n4616) );
  AND2X2 AND2X2_1284 ( .A(u2__abc_44228_n4619), .B(u2_remHi_211_), .Y(u2__abc_44228_n4620_1) );
  AND2X2 AND2X2_1285 ( .A(u2__abc_44228_n4622), .B(sqrto_211_), .Y(u2__abc_44228_n4623) );
  AND2X2 AND2X2_1286 ( .A(u2__abc_44228_n4621), .B(u2__abc_44228_n4624), .Y(u2__abc_44228_n4625) );
  AND2X2 AND2X2_1287 ( .A(u2__abc_44228_n4618), .B(u2__abc_44228_n4625), .Y(u2__abc_44228_n4626) );
  AND2X2 AND2X2_1288 ( .A(u2__abc_44228_n4612), .B(u2__abc_44228_n4626), .Y(u2__abc_44228_n4627) );
  AND2X2 AND2X2_1289 ( .A(u2__abc_44228_n4628), .B(u2_remHi_209_), .Y(u2__abc_44228_n4629_1) );
  AND2X2 AND2X2_129 ( .A(_abc_64468_n987), .B(_abc_64468_n986), .Y(_auto_iopadmap_cc_313_execute_65414_164_) );
  AND2X2 AND2X2_1290 ( .A(u2__abc_44228_n4631), .B(sqrto_209_), .Y(u2__abc_44228_n4632) );
  AND2X2 AND2X2_1291 ( .A(u2__abc_44228_n4630), .B(u2__abc_44228_n4633), .Y(u2__abc_44228_n4634) );
  AND2X2 AND2X2_1292 ( .A(u2__abc_44228_n4635), .B(u2_remHi_208_), .Y(u2__abc_44228_n4636) );
  AND2X2 AND2X2_1293 ( .A(u2__abc_44228_n4637), .B(sqrto_208_), .Y(u2__abc_44228_n4638_1) );
  AND2X2 AND2X2_1294 ( .A(u2__abc_44228_n4640), .B(u2__abc_44228_n4634), .Y(u2__abc_44228_n4641) );
  AND2X2 AND2X2_1295 ( .A(u2__abc_44228_n4642), .B(u2_remHi_207_), .Y(u2__abc_44228_n4643) );
  AND2X2 AND2X2_1296 ( .A(u2__abc_44228_n4645), .B(sqrto_207_), .Y(u2__abc_44228_n4646_1) );
  AND2X2 AND2X2_1297 ( .A(u2__abc_44228_n4644), .B(u2__abc_44228_n4647), .Y(u2__abc_44228_n4648) );
  AND2X2 AND2X2_1298 ( .A(u2__abc_44228_n4649), .B(u2_remHi_206_), .Y(u2__abc_44228_n4650) );
  AND2X2 AND2X2_1299 ( .A(u2__abc_44228_n4651), .B(sqrto_206_), .Y(u2__abc_44228_n4652) );
  AND2X2 AND2X2_13 ( .A(_abc_64468_n753_bF_buf1), .B(sqrto_12_), .Y(_auto_iopadmap_cc_313_execute_65414_48_) );
  AND2X2 AND2X2_130 ( .A(_abc_64468_n990), .B(_abc_64468_n989), .Y(_auto_iopadmap_cc_313_execute_65414_165_) );
  AND2X2 AND2X2_1300 ( .A(u2__abc_44228_n4654), .B(u2__abc_44228_n4648), .Y(u2__abc_44228_n4655) );
  AND2X2 AND2X2_1301 ( .A(u2__abc_44228_n4641), .B(u2__abc_44228_n4655), .Y(u2__abc_44228_n4656_1) );
  AND2X2 AND2X2_1302 ( .A(u2__abc_44228_n4627), .B(u2__abc_44228_n4656_1), .Y(u2__abc_44228_n4657) );
  AND2X2 AND2X2_1303 ( .A(u2__abc_44228_n4598), .B(u2__abc_44228_n4657), .Y(u2__abc_44228_n4658) );
  AND2X2 AND2X2_1304 ( .A(u2__abc_44228_n4659), .B(u2_remHi_205_), .Y(u2__abc_44228_n4660) );
  AND2X2 AND2X2_1305 ( .A(u2__abc_44228_n4662), .B(sqrto_205_), .Y(u2__abc_44228_n4663) );
  AND2X2 AND2X2_1306 ( .A(u2__abc_44228_n4661), .B(u2__abc_44228_n4664), .Y(u2__abc_44228_n4665_1) );
  AND2X2 AND2X2_1307 ( .A(u2__abc_44228_n4666), .B(u2_remHi_204_), .Y(u2__abc_44228_n4667) );
  AND2X2 AND2X2_1308 ( .A(u2__abc_44228_n4668), .B(sqrto_204_), .Y(u2__abc_44228_n4669) );
  AND2X2 AND2X2_1309 ( .A(u2__abc_44228_n4671), .B(u2__abc_44228_n4665_1), .Y(u2__abc_44228_n4672) );
  AND2X2 AND2X2_131 ( .A(_abc_64468_n993), .B(_abc_64468_n992), .Y(_auto_iopadmap_cc_313_execute_65414_166_) );
  AND2X2 AND2X2_1310 ( .A(u2__abc_44228_n4673), .B(u2_remHi_203_), .Y(u2__abc_44228_n4674_1) );
  AND2X2 AND2X2_1311 ( .A(u2__abc_44228_n4676), .B(sqrto_203_), .Y(u2__abc_44228_n4677) );
  AND2X2 AND2X2_1312 ( .A(u2__abc_44228_n4675), .B(u2__abc_44228_n4678), .Y(u2__abc_44228_n4679) );
  AND2X2 AND2X2_1313 ( .A(u2__abc_44228_n4680), .B(u2_remHi_202_), .Y(u2__abc_44228_n4681) );
  AND2X2 AND2X2_1314 ( .A(u2__abc_44228_n4682), .B(sqrto_202_), .Y(u2__abc_44228_n4683) );
  AND2X2 AND2X2_1315 ( .A(u2__abc_44228_n4685_1), .B(u2__abc_44228_n4679), .Y(u2__abc_44228_n4686) );
  AND2X2 AND2X2_1316 ( .A(u2__abc_44228_n4672), .B(u2__abc_44228_n4686), .Y(u2__abc_44228_n4687) );
  AND2X2 AND2X2_1317 ( .A(u2__abc_44228_n4688), .B(u2_remHi_201_), .Y(u2__abc_44228_n4689) );
  AND2X2 AND2X2_1318 ( .A(u2__abc_44228_n4691), .B(sqrto_201_), .Y(u2__abc_44228_n4692) );
  AND2X2 AND2X2_1319 ( .A(u2__abc_44228_n4690), .B(u2__abc_44228_n4693), .Y(u2__abc_44228_n4694) );
  AND2X2 AND2X2_132 ( .A(_abc_64468_n996), .B(_abc_64468_n995), .Y(_auto_iopadmap_cc_313_execute_65414_167_) );
  AND2X2 AND2X2_1320 ( .A(u2__abc_44228_n4695_1), .B(u2_remHi_200_), .Y(u2__abc_44228_n4696) );
  AND2X2 AND2X2_1321 ( .A(u2__abc_44228_n4697), .B(sqrto_200_), .Y(u2__abc_44228_n4698) );
  AND2X2 AND2X2_1322 ( .A(u2__abc_44228_n4700), .B(u2__abc_44228_n4694), .Y(u2__abc_44228_n4701) );
  AND2X2 AND2X2_1323 ( .A(u2__abc_44228_n4702), .B(u2_remHi_198_), .Y(u2__abc_44228_n4703) );
  AND2X2 AND2X2_1324 ( .A(u2__abc_44228_n4704_1), .B(sqrto_198_), .Y(u2__abc_44228_n4705) );
  AND2X2 AND2X2_1325 ( .A(u2__abc_44228_n4708), .B(u2_remHi_199_), .Y(u2__abc_44228_n4709) );
  AND2X2 AND2X2_1326 ( .A(u2__abc_44228_n4711), .B(sqrto_199_), .Y(u2__abc_44228_n4712) );
  AND2X2 AND2X2_1327 ( .A(u2__abc_44228_n4710), .B(u2__abc_44228_n4713_1), .Y(u2__abc_44228_n4714) );
  AND2X2 AND2X2_1328 ( .A(u2__abc_44228_n4707), .B(u2__abc_44228_n4714), .Y(u2__abc_44228_n4715) );
  AND2X2 AND2X2_1329 ( .A(u2__abc_44228_n4701), .B(u2__abc_44228_n4715), .Y(u2__abc_44228_n4716) );
  AND2X2 AND2X2_133 ( .A(_abc_64468_n999), .B(_abc_64468_n998), .Y(_auto_iopadmap_cc_313_execute_65414_168_) );
  AND2X2 AND2X2_1330 ( .A(u2__abc_44228_n4687), .B(u2__abc_44228_n4716), .Y(u2__abc_44228_n4717) );
  AND2X2 AND2X2_1331 ( .A(u2__abc_44228_n4718), .B(u2_remHi_197_), .Y(u2__abc_44228_n4719) );
  AND2X2 AND2X2_1332 ( .A(u2__abc_44228_n4721), .B(sqrto_197_), .Y(u2__abc_44228_n4722_1) );
  AND2X2 AND2X2_1333 ( .A(u2__abc_44228_n4720), .B(u2__abc_44228_n4723), .Y(u2__abc_44228_n4724) );
  AND2X2 AND2X2_1334 ( .A(u2__abc_44228_n4725), .B(u2_remHi_196_), .Y(u2__abc_44228_n4726) );
  AND2X2 AND2X2_1335 ( .A(u2__abc_44228_n4727), .B(sqrto_196_), .Y(u2__abc_44228_n4728) );
  AND2X2 AND2X2_1336 ( .A(u2__abc_44228_n4730), .B(u2__abc_44228_n4724), .Y(u2__abc_44228_n4731_1) );
  AND2X2 AND2X2_1337 ( .A(u2__abc_44228_n4732), .B(u2_remHi_195_), .Y(u2__abc_44228_n4733) );
  AND2X2 AND2X2_1338 ( .A(u2__abc_44228_n4735), .B(sqrto_195_), .Y(u2__abc_44228_n4736) );
  AND2X2 AND2X2_1339 ( .A(u2__abc_44228_n4734), .B(u2__abc_44228_n4737), .Y(u2__abc_44228_n4738) );
  AND2X2 AND2X2_134 ( .A(_abc_64468_n1002), .B(_abc_64468_n1001), .Y(_auto_iopadmap_cc_313_execute_65414_169_) );
  AND2X2 AND2X2_1340 ( .A(u2__abc_44228_n4739), .B(u2_remHi_194_), .Y(u2__abc_44228_n4740) );
  AND2X2 AND2X2_1341 ( .A(u2__abc_44228_n4741_1), .B(sqrto_194_), .Y(u2__abc_44228_n4742) );
  AND2X2 AND2X2_1342 ( .A(u2__abc_44228_n4744), .B(u2__abc_44228_n4738), .Y(u2__abc_44228_n4745) );
  AND2X2 AND2X2_1343 ( .A(u2__abc_44228_n4731_1), .B(u2__abc_44228_n4745), .Y(u2__abc_44228_n4746) );
  AND2X2 AND2X2_1344 ( .A(u2__abc_44228_n4747), .B(u2_remHi_193_), .Y(u2__abc_44228_n4748) );
  AND2X2 AND2X2_1345 ( .A(u2__abc_44228_n4750_1), .B(sqrto_193_), .Y(u2__abc_44228_n4751) );
  AND2X2 AND2X2_1346 ( .A(u2__abc_44228_n4749), .B(u2__abc_44228_n4752), .Y(u2__abc_44228_n4753) );
  AND2X2 AND2X2_1347 ( .A(u2__abc_44228_n4754), .B(u2_remHi_192_), .Y(u2__abc_44228_n4755) );
  AND2X2 AND2X2_1348 ( .A(u2__abc_44228_n4756), .B(sqrto_192_), .Y(u2__abc_44228_n4757) );
  AND2X2 AND2X2_1349 ( .A(u2__abc_44228_n4759), .B(u2__abc_44228_n4753), .Y(u2__abc_44228_n4760_1) );
  AND2X2 AND2X2_135 ( .A(_abc_64468_n1005), .B(_abc_64468_n1004), .Y(_auto_iopadmap_cc_313_execute_65414_170_) );
  AND2X2 AND2X2_1350 ( .A(u2__abc_44228_n4761), .B(u2_remHi_190_), .Y(u2__abc_44228_n4762) );
  AND2X2 AND2X2_1351 ( .A(u2__abc_44228_n4763), .B(sqrto_190_), .Y(u2__abc_44228_n4764) );
  AND2X2 AND2X2_1352 ( .A(u2__abc_44228_n4767), .B(u2_remHi_191_), .Y(u2__abc_44228_n4768) );
  AND2X2 AND2X2_1353 ( .A(u2__abc_44228_n4770_1), .B(sqrto_191_), .Y(u2__abc_44228_n4771) );
  AND2X2 AND2X2_1354 ( .A(u2__abc_44228_n4769), .B(u2__abc_44228_n4772), .Y(u2__abc_44228_n4773) );
  AND2X2 AND2X2_1355 ( .A(u2__abc_44228_n4766), .B(u2__abc_44228_n4773), .Y(u2__abc_44228_n4774) );
  AND2X2 AND2X2_1356 ( .A(u2__abc_44228_n4760_1), .B(u2__abc_44228_n4774), .Y(u2__abc_44228_n4775) );
  AND2X2 AND2X2_1357 ( .A(u2__abc_44228_n4746), .B(u2__abc_44228_n4775), .Y(u2__abc_44228_n4776) );
  AND2X2 AND2X2_1358 ( .A(u2__abc_44228_n4717), .B(u2__abc_44228_n4776), .Y(u2__abc_44228_n4777) );
  AND2X2 AND2X2_1359 ( .A(u2__abc_44228_n4658), .B(u2__abc_44228_n4777), .Y(u2__abc_44228_n4778) );
  AND2X2 AND2X2_136 ( .A(_abc_64468_n1008), .B(_abc_64468_n1007), .Y(_auto_iopadmap_cc_313_execute_65414_171_) );
  AND2X2 AND2X2_1360 ( .A(u2__abc_44228_n4539), .B(u2__abc_44228_n4778), .Y(u2__abc_44228_n4779_1) );
  AND2X2 AND2X2_1361 ( .A(u2__abc_44228_n4780), .B(u2_remHi_189_), .Y(u2__abc_44228_n4781) );
  AND2X2 AND2X2_1362 ( .A(u2__abc_44228_n4783), .B(sqrto_189_), .Y(u2__abc_44228_n4784) );
  AND2X2 AND2X2_1363 ( .A(u2__abc_44228_n4782), .B(u2__abc_44228_n4785), .Y(u2__abc_44228_n4786) );
  AND2X2 AND2X2_1364 ( .A(u2__abc_44228_n4787), .B(u2_remHi_188_), .Y(u2__abc_44228_n4788_1) );
  AND2X2 AND2X2_1365 ( .A(u2__abc_44228_n4789), .B(sqrto_188_), .Y(u2__abc_44228_n4790) );
  AND2X2 AND2X2_1366 ( .A(u2__abc_44228_n4792), .B(u2__abc_44228_n4786), .Y(u2__abc_44228_n4793) );
  AND2X2 AND2X2_1367 ( .A(u2__abc_44228_n4794), .B(u2_remHi_187_), .Y(u2__abc_44228_n4795) );
  AND2X2 AND2X2_1368 ( .A(u2__abc_44228_n4797), .B(sqrto_187_), .Y(u2__abc_44228_n4798) );
  AND2X2 AND2X2_1369 ( .A(u2__abc_44228_n4796), .B(u2__abc_44228_n4799_1), .Y(u2__abc_44228_n4800) );
  AND2X2 AND2X2_137 ( .A(_abc_64468_n1011), .B(_abc_64468_n1010), .Y(_auto_iopadmap_cc_313_execute_65414_172_) );
  AND2X2 AND2X2_1370 ( .A(u2__abc_44228_n4801), .B(u2_remHi_186_), .Y(u2__abc_44228_n4802) );
  AND2X2 AND2X2_1371 ( .A(u2__abc_44228_n4803), .B(sqrto_186_), .Y(u2__abc_44228_n4804) );
  AND2X2 AND2X2_1372 ( .A(u2__abc_44228_n4806), .B(u2__abc_44228_n4800), .Y(u2__abc_44228_n4807) );
  AND2X2 AND2X2_1373 ( .A(u2__abc_44228_n4793), .B(u2__abc_44228_n4807), .Y(u2__abc_44228_n4808) );
  AND2X2 AND2X2_1374 ( .A(u2__abc_44228_n4809_1), .B(u2_remHi_183_), .Y(u2__abc_44228_n4810) );
  AND2X2 AND2X2_1375 ( .A(u2__abc_44228_n4812), .B(sqrto_183_), .Y(u2__abc_44228_n4813) );
  AND2X2 AND2X2_1376 ( .A(u2__abc_44228_n4811), .B(u2__abc_44228_n4814), .Y(u2__abc_44228_n4815) );
  AND2X2 AND2X2_1377 ( .A(u2__abc_44228_n4816), .B(u2_remHi_182_), .Y(u2__abc_44228_n4817) );
  AND2X2 AND2X2_1378 ( .A(u2__abc_44228_n4818_1), .B(sqrto_182_), .Y(u2__abc_44228_n4819) );
  AND2X2 AND2X2_1379 ( .A(u2__abc_44228_n4821), .B(u2__abc_44228_n4815), .Y(u2__abc_44228_n4822) );
  AND2X2 AND2X2_138 ( .A(_abc_64468_n1014), .B(_abc_64468_n1013), .Y(_auto_iopadmap_cc_313_execute_65414_173_) );
  AND2X2 AND2X2_1380 ( .A(u2__abc_44228_n4823), .B(u2_remHi_185_), .Y(u2__abc_44228_n4824) );
  AND2X2 AND2X2_1381 ( .A(u2__abc_44228_n4826), .B(sqrto_185_), .Y(u2__abc_44228_n4827_1) );
  AND2X2 AND2X2_1382 ( .A(u2__abc_44228_n4825), .B(u2__abc_44228_n4828), .Y(u2__abc_44228_n4829) );
  AND2X2 AND2X2_1383 ( .A(u2__abc_44228_n4830), .B(u2_remHi_184_), .Y(u2__abc_44228_n4831) );
  AND2X2 AND2X2_1384 ( .A(u2__abc_44228_n4832), .B(sqrto_184_), .Y(u2__abc_44228_n4833) );
  AND2X2 AND2X2_1385 ( .A(u2__abc_44228_n4835), .B(u2__abc_44228_n4829), .Y(u2__abc_44228_n4836_1) );
  AND2X2 AND2X2_1386 ( .A(u2__abc_44228_n4822), .B(u2__abc_44228_n4836_1), .Y(u2__abc_44228_n4837) );
  AND2X2 AND2X2_1387 ( .A(u2__abc_44228_n4808), .B(u2__abc_44228_n4837), .Y(u2__abc_44228_n4838) );
  AND2X2 AND2X2_1388 ( .A(u2__abc_44228_n4839), .B(u2_remHi_181_), .Y(u2__abc_44228_n4840) );
  AND2X2 AND2X2_1389 ( .A(u2__abc_44228_n4842), .B(sqrto_181_), .Y(u2__abc_44228_n4843) );
  AND2X2 AND2X2_139 ( .A(_abc_64468_n1017), .B(_abc_64468_n1016), .Y(_auto_iopadmap_cc_313_execute_65414_174_) );
  AND2X2 AND2X2_1390 ( .A(u2__abc_44228_n4841), .B(u2__abc_44228_n4844), .Y(u2__abc_44228_n4845) );
  AND2X2 AND2X2_1391 ( .A(u2__abc_44228_n4846_1), .B(u2_remHi_180_), .Y(u2__abc_44228_n4847) );
  AND2X2 AND2X2_1392 ( .A(u2__abc_44228_n4848), .B(sqrto_180_), .Y(u2__abc_44228_n4849) );
  AND2X2 AND2X2_1393 ( .A(u2__abc_44228_n4851), .B(u2__abc_44228_n4845), .Y(u2__abc_44228_n4852) );
  AND2X2 AND2X2_1394 ( .A(u2__abc_44228_n4853), .B(u2_remHi_179_), .Y(u2__abc_44228_n4854) );
  AND2X2 AND2X2_1395 ( .A(u2__abc_44228_n4856), .B(sqrto_179_), .Y(u2__abc_44228_n4857) );
  AND2X2 AND2X2_1396 ( .A(u2__abc_44228_n4855_1), .B(u2__abc_44228_n4858), .Y(u2__abc_44228_n4859) );
  AND2X2 AND2X2_1397 ( .A(u2__abc_44228_n4860), .B(u2_remHi_178_), .Y(u2__abc_44228_n4861) );
  AND2X2 AND2X2_1398 ( .A(u2__abc_44228_n4862), .B(sqrto_178_), .Y(u2__abc_44228_n4863) );
  AND2X2 AND2X2_1399 ( .A(u2__abc_44228_n4865), .B(u2__abc_44228_n4859), .Y(u2__abc_44228_n4866) );
  AND2X2 AND2X2_14 ( .A(_abc_64468_n753_bF_buf0), .B(sqrto_13_), .Y(_auto_iopadmap_cc_313_execute_65414_49_) );
  AND2X2 AND2X2_140 ( .A(_abc_64468_n1020), .B(_abc_64468_n1019), .Y(_auto_iopadmap_cc_313_execute_65414_175_) );
  AND2X2 AND2X2_1400 ( .A(u2__abc_44228_n4852), .B(u2__abc_44228_n4866), .Y(u2__abc_44228_n4867) );
  AND2X2 AND2X2_1401 ( .A(u2__abc_44228_n4868), .B(u2_remHi_177_), .Y(u2__abc_44228_n4869) );
  AND2X2 AND2X2_1402 ( .A(u2__abc_44228_n4871), .B(sqrto_177_), .Y(u2__abc_44228_n4872) );
  AND2X2 AND2X2_1403 ( .A(u2__abc_44228_n4870), .B(u2__abc_44228_n4873_1), .Y(u2__abc_44228_n4874) );
  AND2X2 AND2X2_1404 ( .A(u2__abc_44228_n4875), .B(u2_remHi_176_), .Y(u2__abc_44228_n4876) );
  AND2X2 AND2X2_1405 ( .A(u2__abc_44228_n4877), .B(sqrto_176_), .Y(u2__abc_44228_n4878) );
  AND2X2 AND2X2_1406 ( .A(u2__abc_44228_n4880), .B(u2__abc_44228_n4874), .Y(u2__abc_44228_n4881) );
  AND2X2 AND2X2_1407 ( .A(u2__abc_44228_n4882_1), .B(u2_remHi_175_), .Y(u2__abc_44228_n4883) );
  AND2X2 AND2X2_1408 ( .A(u2__abc_44228_n4885), .B(sqrto_175_), .Y(u2__abc_44228_n4886) );
  AND2X2 AND2X2_1409 ( .A(u2__abc_44228_n4884), .B(u2__abc_44228_n4887), .Y(u2__abc_44228_n4888) );
  AND2X2 AND2X2_141 ( .A(_abc_64468_n1023), .B(_abc_64468_n1022), .Y(_auto_iopadmap_cc_313_execute_65414_176_) );
  AND2X2 AND2X2_1410 ( .A(u2__abc_44228_n4889), .B(u2_remHi_174_), .Y(u2__abc_44228_n4890) );
  AND2X2 AND2X2_1411 ( .A(u2__abc_44228_n4891), .B(sqrto_174_), .Y(u2__abc_44228_n4892_1) );
  AND2X2 AND2X2_1412 ( .A(u2__abc_44228_n4894), .B(u2__abc_44228_n4888), .Y(u2__abc_44228_n4895) );
  AND2X2 AND2X2_1413 ( .A(u2__abc_44228_n4881), .B(u2__abc_44228_n4895), .Y(u2__abc_44228_n4896) );
  AND2X2 AND2X2_1414 ( .A(u2__abc_44228_n4867), .B(u2__abc_44228_n4896), .Y(u2__abc_44228_n4897) );
  AND2X2 AND2X2_1415 ( .A(u2__abc_44228_n4838), .B(u2__abc_44228_n4897), .Y(u2__abc_44228_n4898) );
  AND2X2 AND2X2_1416 ( .A(u2__abc_44228_n4899), .B(u2_remHi_173_), .Y(u2__abc_44228_n4900) );
  AND2X2 AND2X2_1417 ( .A(u2__abc_44228_n4902), .B(sqrto_173_), .Y(u2__abc_44228_n4903) );
  AND2X2 AND2X2_1418 ( .A(u2__abc_44228_n4901_1), .B(u2__abc_44228_n4904), .Y(u2__abc_44228_n4905) );
  AND2X2 AND2X2_1419 ( .A(u2__abc_44228_n4906), .B(u2_remHi_172_), .Y(u2__abc_44228_n4907) );
  AND2X2 AND2X2_142 ( .A(_abc_64468_n1026), .B(_abc_64468_n1025), .Y(_auto_iopadmap_cc_313_execute_65414_177_) );
  AND2X2 AND2X2_1420 ( .A(u2__abc_44228_n4908), .B(sqrto_172_), .Y(u2__abc_44228_n4909) );
  AND2X2 AND2X2_1421 ( .A(u2__abc_44228_n4911_1), .B(u2__abc_44228_n4905), .Y(u2__abc_44228_n4912) );
  AND2X2 AND2X2_1422 ( .A(u2__abc_44228_n4913), .B(u2_remHi_170_), .Y(u2__abc_44228_n4914) );
  AND2X2 AND2X2_1423 ( .A(u2__abc_44228_n4915), .B(sqrto_170_), .Y(u2__abc_44228_n4916) );
  AND2X2 AND2X2_1424 ( .A(u2__abc_44228_n4919), .B(u2_remHi_171_), .Y(u2__abc_44228_n4920) );
  AND2X2 AND2X2_1425 ( .A(u2__abc_44228_n4922), .B(sqrto_171_), .Y(u2__abc_44228_n4923) );
  AND2X2 AND2X2_1426 ( .A(u2__abc_44228_n4921_1), .B(u2__abc_44228_n4924), .Y(u2__abc_44228_n4925) );
  AND2X2 AND2X2_1427 ( .A(u2__abc_44228_n4918), .B(u2__abc_44228_n4925), .Y(u2__abc_44228_n4926) );
  AND2X2 AND2X2_1428 ( .A(u2__abc_44228_n4912), .B(u2__abc_44228_n4926), .Y(u2__abc_44228_n4927) );
  AND2X2 AND2X2_1429 ( .A(u2__abc_44228_n4928), .B(u2_remHi_169_), .Y(u2__abc_44228_n4929) );
  AND2X2 AND2X2_143 ( .A(_abc_64468_n1029), .B(_abc_64468_n1028), .Y(_auto_iopadmap_cc_313_execute_65414_178_) );
  AND2X2 AND2X2_1430 ( .A(u2__abc_44228_n4931), .B(sqrto_169_), .Y(u2__abc_44228_n4932) );
  AND2X2 AND2X2_1431 ( .A(u2__abc_44228_n4930_1), .B(u2__abc_44228_n4933), .Y(u2__abc_44228_n4934) );
  AND2X2 AND2X2_1432 ( .A(u2__abc_44228_n4935), .B(u2_remHi_168_), .Y(u2__abc_44228_n4936) );
  AND2X2 AND2X2_1433 ( .A(u2__abc_44228_n4937), .B(sqrto_168_), .Y(u2__abc_44228_n4938) );
  AND2X2 AND2X2_1434 ( .A(u2__abc_44228_n4940), .B(u2__abc_44228_n4934), .Y(u2__abc_44228_n4941) );
  AND2X2 AND2X2_1435 ( .A(u2__abc_44228_n4942), .B(u2_remHi_166_), .Y(u2__abc_44228_n4943) );
  AND2X2 AND2X2_1436 ( .A(u2__abc_44228_n4944), .B(sqrto_166_), .Y(u2__abc_44228_n4945) );
  AND2X2 AND2X2_1437 ( .A(u2__abc_44228_n4948_1), .B(u2_remHi_167_), .Y(u2__abc_44228_n4949) );
  AND2X2 AND2X2_1438 ( .A(u2__abc_44228_n4951), .B(sqrto_167_), .Y(u2__abc_44228_n4952) );
  AND2X2 AND2X2_1439 ( .A(u2__abc_44228_n4950), .B(u2__abc_44228_n4953), .Y(u2__abc_44228_n4954) );
  AND2X2 AND2X2_144 ( .A(_abc_64468_n1032), .B(_abc_64468_n1031), .Y(_auto_iopadmap_cc_313_execute_65414_179_) );
  AND2X2 AND2X2_1440 ( .A(u2__abc_44228_n4947), .B(u2__abc_44228_n4954), .Y(u2__abc_44228_n4955) );
  AND2X2 AND2X2_1441 ( .A(u2__abc_44228_n4941), .B(u2__abc_44228_n4955), .Y(u2__abc_44228_n4956) );
  AND2X2 AND2X2_1442 ( .A(u2__abc_44228_n4927), .B(u2__abc_44228_n4956), .Y(u2__abc_44228_n4957_1) );
  AND2X2 AND2X2_1443 ( .A(u2__abc_44228_n4958), .B(u2_remHi_165_), .Y(u2__abc_44228_n4959) );
  AND2X2 AND2X2_1444 ( .A(u2__abc_44228_n4961), .B(sqrto_165_), .Y(u2__abc_44228_n4962) );
  AND2X2 AND2X2_1445 ( .A(u2__abc_44228_n4960), .B(u2__abc_44228_n4963), .Y(u2__abc_44228_n4964) );
  AND2X2 AND2X2_1446 ( .A(u2__abc_44228_n4965), .B(u2_remHi_164_), .Y(u2__abc_44228_n4966) );
  AND2X2 AND2X2_1447 ( .A(u2__abc_44228_n4967_1), .B(sqrto_164_), .Y(u2__abc_44228_n4968) );
  AND2X2 AND2X2_1448 ( .A(u2__abc_44228_n4970), .B(u2__abc_44228_n4964), .Y(u2__abc_44228_n4971) );
  AND2X2 AND2X2_1449 ( .A(u2__abc_44228_n4972), .B(u2_remHi_162_), .Y(u2__abc_44228_n4973) );
  AND2X2 AND2X2_145 ( .A(_abc_64468_n1035), .B(_abc_64468_n1034), .Y(_auto_iopadmap_cc_313_execute_65414_180_) );
  AND2X2 AND2X2_1450 ( .A(u2__abc_44228_n4974), .B(sqrto_162_), .Y(u2__abc_44228_n4975) );
  AND2X2 AND2X2_1451 ( .A(u2__abc_44228_n4978), .B(u2_remHi_163_), .Y(u2__abc_44228_n4979) );
  AND2X2 AND2X2_1452 ( .A(u2__abc_44228_n4981), .B(sqrto_163_), .Y(u2__abc_44228_n4982) );
  AND2X2 AND2X2_1453 ( .A(u2__abc_44228_n4980), .B(u2__abc_44228_n4983), .Y(u2__abc_44228_n4984) );
  AND2X2 AND2X2_1454 ( .A(u2__abc_44228_n4977), .B(u2__abc_44228_n4984), .Y(u2__abc_44228_n4985) );
  AND2X2 AND2X2_1455 ( .A(u2__abc_44228_n4971), .B(u2__abc_44228_n4985), .Y(u2__abc_44228_n4986_1) );
  AND2X2 AND2X2_1456 ( .A(u2__abc_44228_n4987), .B(u2_remHi_161_), .Y(u2__abc_44228_n4988) );
  AND2X2 AND2X2_1457 ( .A(u2__abc_44228_n4990), .B(sqrto_161_), .Y(u2__abc_44228_n4991) );
  AND2X2 AND2X2_1458 ( .A(u2__abc_44228_n4989), .B(u2__abc_44228_n4992), .Y(u2__abc_44228_n4993) );
  AND2X2 AND2X2_1459 ( .A(u2__abc_44228_n4994), .B(u2_remHi_160_), .Y(u2__abc_44228_n4995) );
  AND2X2 AND2X2_146 ( .A(_abc_64468_n1038), .B(_abc_64468_n1037), .Y(_auto_iopadmap_cc_313_execute_65414_181_) );
  AND2X2 AND2X2_1460 ( .A(u2__abc_44228_n4996_1), .B(sqrto_160_), .Y(u2__abc_44228_n4997) );
  AND2X2 AND2X2_1461 ( .A(u2__abc_44228_n4999), .B(u2__abc_44228_n4993), .Y(u2__abc_44228_n5000) );
  AND2X2 AND2X2_1462 ( .A(u2__abc_44228_n5001), .B(u2_remHi_158_), .Y(u2__abc_44228_n5002) );
  AND2X2 AND2X2_1463 ( .A(u2__abc_44228_n5003), .B(sqrto_158_), .Y(u2__abc_44228_n5004) );
  AND2X2 AND2X2_1464 ( .A(u2__abc_44228_n5007), .B(u2_remHi_159_), .Y(u2__abc_44228_n5008) );
  AND2X2 AND2X2_1465 ( .A(u2__abc_44228_n5010), .B(sqrto_159_), .Y(u2__abc_44228_n5011) );
  AND2X2 AND2X2_1466 ( .A(u2__abc_44228_n5009), .B(u2__abc_44228_n5012), .Y(u2__abc_44228_n5013) );
  AND2X2 AND2X2_1467 ( .A(u2__abc_44228_n5006), .B(u2__abc_44228_n5013), .Y(u2__abc_44228_n5014_1) );
  AND2X2 AND2X2_1468 ( .A(u2__abc_44228_n5000), .B(u2__abc_44228_n5014_1), .Y(u2__abc_44228_n5015) );
  AND2X2 AND2X2_1469 ( .A(u2__abc_44228_n4986_1), .B(u2__abc_44228_n5015), .Y(u2__abc_44228_n5016) );
  AND2X2 AND2X2_147 ( .A(_abc_64468_n1041), .B(_abc_64468_n1040), .Y(_auto_iopadmap_cc_313_execute_65414_182_) );
  AND2X2 AND2X2_1470 ( .A(u2__abc_44228_n4957_1), .B(u2__abc_44228_n5016), .Y(u2__abc_44228_n5017) );
  AND2X2 AND2X2_1471 ( .A(u2__abc_44228_n4898), .B(u2__abc_44228_n5017), .Y(u2__abc_44228_n5018) );
  AND2X2 AND2X2_1472 ( .A(u2__abc_44228_n5019), .B(u2_remHi_157_), .Y(u2__abc_44228_n5020) );
  AND2X2 AND2X2_1473 ( .A(u2__abc_44228_n5022), .B(sqrto_157_), .Y(u2__abc_44228_n5023_1) );
  AND2X2 AND2X2_1474 ( .A(u2__abc_44228_n5021), .B(u2__abc_44228_n5024), .Y(u2__abc_44228_n5025) );
  AND2X2 AND2X2_1475 ( .A(u2__abc_44228_n5026), .B(u2_remHi_156_), .Y(u2__abc_44228_n5027) );
  AND2X2 AND2X2_1476 ( .A(u2__abc_44228_n5028), .B(sqrto_156_), .Y(u2__abc_44228_n5029) );
  AND2X2 AND2X2_1477 ( .A(u2__abc_44228_n5031), .B(u2__abc_44228_n5025), .Y(u2__abc_44228_n5032_1) );
  AND2X2 AND2X2_1478 ( .A(u2__abc_44228_n5033), .B(u2_remHi_155_), .Y(u2__abc_44228_n5034) );
  AND2X2 AND2X2_1479 ( .A(u2__abc_44228_n5036), .B(sqrto_155_), .Y(u2__abc_44228_n5037) );
  AND2X2 AND2X2_148 ( .A(_abc_64468_n1044), .B(_abc_64468_n1043), .Y(_auto_iopadmap_cc_313_execute_65414_183_) );
  AND2X2 AND2X2_1480 ( .A(u2__abc_44228_n5035), .B(u2__abc_44228_n5038), .Y(u2__abc_44228_n5039) );
  AND2X2 AND2X2_1481 ( .A(u2__abc_44228_n5040), .B(u2_remHi_154_), .Y(u2__abc_44228_n5041) );
  AND2X2 AND2X2_1482 ( .A(u2__abc_44228_n5042_1), .B(sqrto_154_), .Y(u2__abc_44228_n5043) );
  AND2X2 AND2X2_1483 ( .A(u2__abc_44228_n5045), .B(u2__abc_44228_n5039), .Y(u2__abc_44228_n5046) );
  AND2X2 AND2X2_1484 ( .A(u2__abc_44228_n5032_1), .B(u2__abc_44228_n5046), .Y(u2__abc_44228_n5047) );
  AND2X2 AND2X2_1485 ( .A(u2__abc_44228_n5048), .B(u2_remHi_153_), .Y(u2__abc_44228_n5049) );
  AND2X2 AND2X2_1486 ( .A(u2__abc_44228_n5051_1), .B(sqrto_153_), .Y(u2__abc_44228_n5052) );
  AND2X2 AND2X2_1487 ( .A(u2__abc_44228_n5050), .B(u2__abc_44228_n5053), .Y(u2__abc_44228_n5054) );
  AND2X2 AND2X2_1488 ( .A(u2__abc_44228_n5055), .B(u2_remHi_152_), .Y(u2__abc_44228_n5056) );
  AND2X2 AND2X2_1489 ( .A(u2__abc_44228_n5057), .B(sqrto_152_), .Y(u2__abc_44228_n5058) );
  AND2X2 AND2X2_149 ( .A(_abc_64468_n1047), .B(_abc_64468_n1046), .Y(_auto_iopadmap_cc_313_execute_65414_184_) );
  AND2X2 AND2X2_1490 ( .A(u2__abc_44228_n5060), .B(u2__abc_44228_n5054), .Y(u2__abc_44228_n5061_1) );
  AND2X2 AND2X2_1491 ( .A(u2__abc_44228_n5062), .B(u2_remHi_150_), .Y(u2__abc_44228_n5063) );
  AND2X2 AND2X2_1492 ( .A(u2__abc_44228_n5064), .B(sqrto_150_), .Y(u2__abc_44228_n5065) );
  AND2X2 AND2X2_1493 ( .A(u2__abc_44228_n5068), .B(u2_remHi_151_), .Y(u2__abc_44228_n5069) );
  AND2X2 AND2X2_1494 ( .A(u2__abc_44228_n5071_1), .B(sqrto_151_), .Y(u2__abc_44228_n5072) );
  AND2X2 AND2X2_1495 ( .A(u2__abc_44228_n5070), .B(u2__abc_44228_n5073), .Y(u2__abc_44228_n5074) );
  AND2X2 AND2X2_1496 ( .A(u2__abc_44228_n5067), .B(u2__abc_44228_n5074), .Y(u2__abc_44228_n5075) );
  AND2X2 AND2X2_1497 ( .A(u2__abc_44228_n5061_1), .B(u2__abc_44228_n5075), .Y(u2__abc_44228_n5076) );
  AND2X2 AND2X2_1498 ( .A(u2__abc_44228_n5047), .B(u2__abc_44228_n5076), .Y(u2__abc_44228_n5077) );
  AND2X2 AND2X2_1499 ( .A(u2__abc_44228_n5078), .B(u2_remHi_149_), .Y(u2__abc_44228_n5079) );
  AND2X2 AND2X2_15 ( .A(_abc_64468_n753_bF_buf13), .B(sqrto_14_), .Y(_auto_iopadmap_cc_313_execute_65414_50_) );
  AND2X2 AND2X2_150 ( .A(_abc_64468_n1050), .B(_abc_64468_n1049), .Y(_auto_iopadmap_cc_313_execute_65414_185_) );
  AND2X2 AND2X2_1500 ( .A(u2__abc_44228_n5081), .B(sqrto_149_), .Y(u2__abc_44228_n5082) );
  AND2X2 AND2X2_1501 ( .A(u2__abc_44228_n5080_1), .B(u2__abc_44228_n5083), .Y(u2__abc_44228_n5084) );
  AND2X2 AND2X2_1502 ( .A(u2__abc_44228_n5085), .B(u2_remHi_148_), .Y(u2__abc_44228_n5086) );
  AND2X2 AND2X2_1503 ( .A(u2__abc_44228_n5087), .B(sqrto_148_), .Y(u2__abc_44228_n5088) );
  AND2X2 AND2X2_1504 ( .A(u2__abc_44228_n5090), .B(u2__abc_44228_n5084), .Y(u2__abc_44228_n5091) );
  AND2X2 AND2X2_1505 ( .A(u2__abc_44228_n5092), .B(u2_remHi_146_), .Y(u2__abc_44228_n5093) );
  AND2X2 AND2X2_1506 ( .A(u2__abc_44228_n5094), .B(sqrto_146_), .Y(u2__abc_44228_n5095) );
  AND2X2 AND2X2_1507 ( .A(u2__abc_44228_n5098), .B(u2_remHi_147_), .Y(u2__abc_44228_n5099_1) );
  AND2X2 AND2X2_1508 ( .A(u2__abc_44228_n5101), .B(sqrto_147_), .Y(u2__abc_44228_n5102) );
  AND2X2 AND2X2_1509 ( .A(u2__abc_44228_n5100), .B(u2__abc_44228_n5103), .Y(u2__abc_44228_n5104) );
  AND2X2 AND2X2_151 ( .A(_abc_64468_n1053), .B(_abc_64468_n1052), .Y(_auto_iopadmap_cc_313_execute_65414_186_) );
  AND2X2 AND2X2_1510 ( .A(u2__abc_44228_n5097), .B(u2__abc_44228_n5104), .Y(u2__abc_44228_n5105) );
  AND2X2 AND2X2_1511 ( .A(u2__abc_44228_n5091), .B(u2__abc_44228_n5105), .Y(u2__abc_44228_n5106) );
  AND2X2 AND2X2_1512 ( .A(u2__abc_44228_n5107), .B(u2_remHi_145_), .Y(u2__abc_44228_n5108) );
  AND2X2 AND2X2_1513 ( .A(u2__abc_44228_n5110), .B(sqrto_145_), .Y(u2__abc_44228_n5111) );
  AND2X2 AND2X2_1514 ( .A(u2__abc_44228_n5109_1), .B(u2__abc_44228_n5112), .Y(u2__abc_44228_n5113) );
  AND2X2 AND2X2_1515 ( .A(u2__abc_44228_n5114), .B(u2_remHi_144_), .Y(u2__abc_44228_n5115) );
  AND2X2 AND2X2_1516 ( .A(u2__abc_44228_n5116), .B(sqrto_144_), .Y(u2__abc_44228_n5117) );
  AND2X2 AND2X2_1517 ( .A(u2__abc_44228_n5119), .B(u2__abc_44228_n5113), .Y(u2__abc_44228_n5120) );
  AND2X2 AND2X2_1518 ( .A(u2__abc_44228_n5121), .B(u2_remHi_143_), .Y(u2__abc_44228_n5122) );
  AND2X2 AND2X2_1519 ( .A(u2__abc_44228_n5124), .B(sqrto_143_), .Y(u2__abc_44228_n5125) );
  AND2X2 AND2X2_152 ( .A(_abc_64468_n1056), .B(_abc_64468_n1055), .Y(_auto_iopadmap_cc_313_execute_65414_187_) );
  AND2X2 AND2X2_1520 ( .A(u2__abc_44228_n5123), .B(u2__abc_44228_n5126), .Y(u2__abc_44228_n5127_1) );
  AND2X2 AND2X2_1521 ( .A(u2__abc_44228_n5128), .B(u2_remHi_142_), .Y(u2__abc_44228_n5129) );
  AND2X2 AND2X2_1522 ( .A(u2__abc_44228_n5130), .B(sqrto_142_), .Y(u2__abc_44228_n5131) );
  AND2X2 AND2X2_1523 ( .A(u2__abc_44228_n5133), .B(u2__abc_44228_n5127_1), .Y(u2__abc_44228_n5134) );
  AND2X2 AND2X2_1524 ( .A(u2__abc_44228_n5120), .B(u2__abc_44228_n5134), .Y(u2__abc_44228_n5135) );
  AND2X2 AND2X2_1525 ( .A(u2__abc_44228_n5106), .B(u2__abc_44228_n5135), .Y(u2__abc_44228_n5136_1) );
  AND2X2 AND2X2_1526 ( .A(u2__abc_44228_n5077), .B(u2__abc_44228_n5136_1), .Y(u2__abc_44228_n5137) );
  AND2X2 AND2X2_1527 ( .A(u2__abc_44228_n5138), .B(u2_remHi_141_), .Y(u2__abc_44228_n5139) );
  AND2X2 AND2X2_1528 ( .A(u2__abc_44228_n5141), .B(sqrto_141_), .Y(u2__abc_44228_n5142) );
  AND2X2 AND2X2_1529 ( .A(u2__abc_44228_n5140), .B(u2__abc_44228_n5143), .Y(u2__abc_44228_n5144) );
  AND2X2 AND2X2_153 ( .A(_abc_64468_n1059), .B(_abc_64468_n1058), .Y(_auto_iopadmap_cc_313_execute_65414_188_) );
  AND2X2 AND2X2_1530 ( .A(u2__abc_44228_n5145), .B(u2_remHi_140_), .Y(u2__abc_44228_n5146_1) );
  AND2X2 AND2X2_1531 ( .A(u2__abc_44228_n5147), .B(sqrto_140_), .Y(u2__abc_44228_n5148) );
  AND2X2 AND2X2_1532 ( .A(u2__abc_44228_n5150), .B(u2__abc_44228_n5144), .Y(u2__abc_44228_n5151) );
  AND2X2 AND2X2_1533 ( .A(u2__abc_44228_n5152), .B(u2_remHi_139_), .Y(u2__abc_44228_n5153) );
  AND2X2 AND2X2_1534 ( .A(u2__abc_44228_n5155_1), .B(sqrto_139_), .Y(u2__abc_44228_n5156) );
  AND2X2 AND2X2_1535 ( .A(u2__abc_44228_n5154), .B(u2__abc_44228_n5157), .Y(u2__abc_44228_n5158) );
  AND2X2 AND2X2_1536 ( .A(u2__abc_44228_n5159), .B(u2_remHi_138_), .Y(u2__abc_44228_n5160) );
  AND2X2 AND2X2_1537 ( .A(u2__abc_44228_n5161), .B(sqrto_138_), .Y(u2__abc_44228_n5162) );
  AND2X2 AND2X2_1538 ( .A(u2__abc_44228_n5164_1), .B(u2__abc_44228_n5158), .Y(u2__abc_44228_n5165) );
  AND2X2 AND2X2_1539 ( .A(u2__abc_44228_n5151), .B(u2__abc_44228_n5165), .Y(u2__abc_44228_n5166) );
  AND2X2 AND2X2_154 ( .A(_abc_64468_n1062), .B(_abc_64468_n1061), .Y(_auto_iopadmap_cc_313_execute_65414_189_) );
  AND2X2 AND2X2_1540 ( .A(u2__abc_44228_n5167), .B(u2_remHi_135_), .Y(u2__abc_44228_n5168) );
  AND2X2 AND2X2_1541 ( .A(u2__abc_44228_n5170), .B(sqrto_135_), .Y(u2__abc_44228_n5171) );
  AND2X2 AND2X2_1542 ( .A(u2__abc_44228_n5169), .B(u2__abc_44228_n5172), .Y(u2__abc_44228_n5173_1) );
  AND2X2 AND2X2_1543 ( .A(u2__abc_44228_n5174), .B(u2_remHi_134_), .Y(u2__abc_44228_n5175) );
  AND2X2 AND2X2_1544 ( .A(u2__abc_44228_n5176), .B(sqrto_134_), .Y(u2__abc_44228_n5177) );
  AND2X2 AND2X2_1545 ( .A(u2__abc_44228_n5179), .B(u2__abc_44228_n5173_1), .Y(u2__abc_44228_n5180) );
  AND2X2 AND2X2_1546 ( .A(u2__abc_44228_n5181), .B(u2_remHi_137_), .Y(u2__abc_44228_n5182_1) );
  AND2X2 AND2X2_1547 ( .A(u2__abc_44228_n5184), .B(sqrto_137_), .Y(u2__abc_44228_n5185) );
  AND2X2 AND2X2_1548 ( .A(u2__abc_44228_n5183), .B(u2__abc_44228_n5186), .Y(u2__abc_44228_n5187) );
  AND2X2 AND2X2_1549 ( .A(u2__abc_44228_n5188), .B(u2_remHi_136_), .Y(u2__abc_44228_n5189) );
  AND2X2 AND2X2_155 ( .A(_abc_64468_n1065), .B(_abc_64468_n1064), .Y(_auto_iopadmap_cc_313_execute_65414_190_) );
  AND2X2 AND2X2_1550 ( .A(u2__abc_44228_n5190), .B(sqrto_136_), .Y(u2__abc_44228_n5191) );
  AND2X2 AND2X2_1551 ( .A(u2__abc_44228_n5193), .B(u2__abc_44228_n5187), .Y(u2__abc_44228_n5194) );
  AND2X2 AND2X2_1552 ( .A(u2__abc_44228_n5180), .B(u2__abc_44228_n5194), .Y(u2__abc_44228_n5195) );
  AND2X2 AND2X2_1553 ( .A(u2__abc_44228_n5166), .B(u2__abc_44228_n5195), .Y(u2__abc_44228_n5196) );
  AND2X2 AND2X2_1554 ( .A(u2__abc_44228_n5197), .B(u2_remHi_133_), .Y(u2__abc_44228_n5198) );
  AND2X2 AND2X2_1555 ( .A(u2__abc_44228_n5200), .B(sqrto_133_), .Y(u2__abc_44228_n5201_1) );
  AND2X2 AND2X2_1556 ( .A(u2__abc_44228_n5199), .B(u2__abc_44228_n5202), .Y(u2__abc_44228_n5203) );
  AND2X2 AND2X2_1557 ( .A(u2__abc_44228_n5204), .B(u2_remHi_132_), .Y(u2__abc_44228_n5205) );
  AND2X2 AND2X2_1558 ( .A(u2__abc_44228_n5206), .B(sqrto_132_), .Y(u2__abc_44228_n5207) );
  AND2X2 AND2X2_1559 ( .A(u2__abc_44228_n5209), .B(u2__abc_44228_n5203), .Y(u2__abc_44228_n5210) );
  AND2X2 AND2X2_156 ( .A(_abc_64468_n1068), .B(_abc_64468_n1067), .Y(_auto_iopadmap_cc_313_execute_65414_191_) );
  AND2X2 AND2X2_1560 ( .A(u2__abc_44228_n5211_1), .B(u2_remHi_131_), .Y(u2__abc_44228_n5212) );
  AND2X2 AND2X2_1561 ( .A(u2__abc_44228_n5214), .B(sqrto_131_), .Y(u2__abc_44228_n5215) );
  AND2X2 AND2X2_1562 ( .A(u2__abc_44228_n5213), .B(u2__abc_44228_n5216), .Y(u2__abc_44228_n5217) );
  AND2X2 AND2X2_1563 ( .A(u2__abc_44228_n5218), .B(u2_remHi_130_), .Y(u2__abc_44228_n5219) );
  AND2X2 AND2X2_1564 ( .A(u2__abc_44228_n5220), .B(sqrto_130_), .Y(u2__abc_44228_n5221_1) );
  AND2X2 AND2X2_1565 ( .A(u2__abc_44228_n5223), .B(u2__abc_44228_n5217), .Y(u2__abc_44228_n5224) );
  AND2X2 AND2X2_1566 ( .A(u2__abc_44228_n5210), .B(u2__abc_44228_n5224), .Y(u2__abc_44228_n5225) );
  AND2X2 AND2X2_1567 ( .A(u2__abc_44228_n5227), .B(u2__abc_44228_n5229), .Y(u2__abc_44228_n5230_1) );
  AND2X2 AND2X2_1568 ( .A(u2__abc_44228_n5232), .B(u2__abc_44228_n5234), .Y(u2__abc_44228_n5235) );
  AND2X2 AND2X2_1569 ( .A(u2__abc_44228_n5230_1), .B(u2__abc_44228_n5235), .Y(u2__abc_44228_n5236) );
  AND2X2 AND2X2_157 ( .A(_abc_64468_n1071), .B(_abc_64468_n1070), .Y(_auto_iopadmap_cc_313_execute_65414_192_) );
  AND2X2 AND2X2_1570 ( .A(u2__abc_44228_n5237), .B(u2_remHi_127_), .Y(u2__abc_44228_n5238) );
  AND2X2 AND2X2_1571 ( .A(u2__abc_44228_n5240), .B(sqrto_127_), .Y(u2__abc_44228_n5241) );
  AND2X2 AND2X2_1572 ( .A(u2__abc_44228_n5239_1), .B(u2__abc_44228_n5242), .Y(u2__abc_44228_n5243) );
  AND2X2 AND2X2_1573 ( .A(u2__abc_44228_n5244), .B(u2_remHi_126_), .Y(u2__abc_44228_n5245) );
  AND2X2 AND2X2_1574 ( .A(u2__abc_44228_n5246), .B(sqrto_126_), .Y(u2__abc_44228_n5247) );
  AND2X2 AND2X2_1575 ( .A(u2__abc_44228_n5249), .B(u2__abc_44228_n5243), .Y(u2__abc_44228_n5250_1) );
  AND2X2 AND2X2_1576 ( .A(u2__abc_44228_n5250_1), .B(u2__abc_44228_n5236), .Y(u2__abc_44228_n5251) );
  AND2X2 AND2X2_1577 ( .A(u2__abc_44228_n5225), .B(u2__abc_44228_n5251), .Y(u2__abc_44228_n5252) );
  AND2X2 AND2X2_1578 ( .A(u2__abc_44228_n5196), .B(u2__abc_44228_n5252), .Y(u2__abc_44228_n5253) );
  AND2X2 AND2X2_1579 ( .A(u2__abc_44228_n5137), .B(u2__abc_44228_n5253), .Y(u2__abc_44228_n5254) );
  AND2X2 AND2X2_158 ( .A(_abc_64468_n1074), .B(_abc_64468_n1073), .Y(_auto_iopadmap_cc_313_execute_65414_193_) );
  AND2X2 AND2X2_1580 ( .A(u2__abc_44228_n5018), .B(u2__abc_44228_n5254), .Y(u2__abc_44228_n5255) );
  AND2X2 AND2X2_1581 ( .A(u2__abc_44228_n4779_1), .B(u2__abc_44228_n5255), .Y(u2__abc_44228_n5256) );
  AND2X2 AND2X2_1582 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5256), .Y(u2__abc_44228_n5257) );
  AND2X2 AND2X2_1583 ( .A(u2__abc_44228_n5258), .B(u2__abc_44228_n5242), .Y(u2__abc_44228_n5259) );
  AND2X2 AND2X2_1584 ( .A(u2__abc_44228_n5259), .B(u2__abc_44228_n5236), .Y(u2__abc_44228_n5260_1) );
  AND2X2 AND2X2_1585 ( .A(u2__abc_44228_n5262), .B(u2__abc_44228_n5229), .Y(u2__abc_44228_n5263) );
  AND2X2 AND2X2_1586 ( .A(u2__abc_44228_n5265), .B(u2__abc_44228_n5225), .Y(u2__abc_44228_n5266) );
  AND2X2 AND2X2_1587 ( .A(u2__abc_44228_n5267), .B(u2__abc_44228_n5216), .Y(u2__abc_44228_n5268) );
  AND2X2 AND2X2_1588 ( .A(u2__abc_44228_n5210), .B(u2__abc_44228_n5268), .Y(u2__abc_44228_n5269_1) );
  AND2X2 AND2X2_1589 ( .A(u2__abc_44228_n5202), .B(u2__abc_44228_n5205), .Y(u2__abc_44228_n5270) );
  AND2X2 AND2X2_159 ( .A(_abc_64468_n1077), .B(_abc_64468_n1076), .Y(_auto_iopadmap_cc_313_execute_65414_194_) );
  AND2X2 AND2X2_1590 ( .A(u2__abc_44228_n5273), .B(u2__abc_44228_n5196), .Y(u2__abc_44228_n5274) );
  AND2X2 AND2X2_1591 ( .A(u2__abc_44228_n5275), .B(u2__abc_44228_n5172), .Y(u2__abc_44228_n5276) );
  AND2X2 AND2X2_1592 ( .A(u2__abc_44228_n5194), .B(u2__abc_44228_n5276), .Y(u2__abc_44228_n5277) );
  AND2X2 AND2X2_1593 ( .A(u2__abc_44228_n5278_1), .B(u2__abc_44228_n5186), .Y(u2__abc_44228_n5279) );
  AND2X2 AND2X2_1594 ( .A(u2__abc_44228_n5280), .B(u2__abc_44228_n5166), .Y(u2__abc_44228_n5281) );
  AND2X2 AND2X2_1595 ( .A(u2__abc_44228_n5154), .B(u2__abc_44228_n5282), .Y(u2__abc_44228_n5283) );
  AND2X2 AND2X2_1596 ( .A(u2__abc_44228_n5284), .B(u2__abc_44228_n5157), .Y(u2__abc_44228_n5285) );
  AND2X2 AND2X2_1597 ( .A(u2__abc_44228_n5285), .B(u2__abc_44228_n5151), .Y(u2__abc_44228_n5286) );
  AND2X2 AND2X2_1598 ( .A(u2__abc_44228_n5287_1), .B(u2__abc_44228_n5143), .Y(u2__abc_44228_n5288) );
  AND2X2 AND2X2_1599 ( .A(u2__abc_44228_n5291), .B(u2__abc_44228_n5137), .Y(u2__abc_44228_n5292) );
  AND2X2 AND2X2_16 ( .A(_abc_64468_n753_bF_buf12), .B(sqrto_15_), .Y(_auto_iopadmap_cc_313_execute_65414_51_) );
  AND2X2 AND2X2_160 ( .A(_abc_64468_n1080), .B(_abc_64468_n1079), .Y(_auto_iopadmap_cc_313_execute_65414_195_) );
  AND2X2 AND2X2_1600 ( .A(u2__abc_44228_n5293), .B(u2__abc_44228_n5126), .Y(u2__abc_44228_n5294) );
  AND2X2 AND2X2_1601 ( .A(u2__abc_44228_n5120), .B(u2__abc_44228_n5294), .Y(u2__abc_44228_n5295) );
  AND2X2 AND2X2_1602 ( .A(u2__abc_44228_n5109_1), .B(u2__abc_44228_n5296), .Y(u2__abc_44228_n5297_1) );
  AND2X2 AND2X2_1603 ( .A(u2__abc_44228_n5298), .B(u2__abc_44228_n5112), .Y(u2__abc_44228_n5299) );
  AND2X2 AND2X2_1604 ( .A(u2__abc_44228_n5300), .B(u2__abc_44228_n5106), .Y(u2__abc_44228_n5301) );
  AND2X2 AND2X2_1605 ( .A(u2__abc_44228_n5302), .B(u2__abc_44228_n5100), .Y(u2__abc_44228_n5303) );
  AND2X2 AND2X2_1606 ( .A(u2__abc_44228_n5304), .B(u2__abc_44228_n5103), .Y(u2__abc_44228_n5305) );
  AND2X2 AND2X2_1607 ( .A(u2__abc_44228_n5305), .B(u2__abc_44228_n5091), .Y(u2__abc_44228_n5306_1) );
  AND2X2 AND2X2_1608 ( .A(u2__abc_44228_n5083), .B(u2__abc_44228_n5086), .Y(u2__abc_44228_n5307) );
  AND2X2 AND2X2_1609 ( .A(u2__abc_44228_n5310), .B(u2__abc_44228_n5077), .Y(u2__abc_44228_n5311) );
  AND2X2 AND2X2_161 ( .A(_abc_64468_n1083), .B(_abc_64468_n1082), .Y(_auto_iopadmap_cc_313_execute_65414_196_) );
  AND2X2 AND2X2_1610 ( .A(u2__abc_44228_n5312), .B(u2__abc_44228_n5053), .Y(u2__abc_44228_n5313) );
  AND2X2 AND2X2_1611 ( .A(u2__abc_44228_n5314), .B(u2__abc_44228_n5070), .Y(u2__abc_44228_n5315_1) );
  AND2X2 AND2X2_1612 ( .A(u2__abc_44228_n5316), .B(u2__abc_44228_n5073), .Y(u2__abc_44228_n5317) );
  AND2X2 AND2X2_1613 ( .A(u2__abc_44228_n5317), .B(u2__abc_44228_n5061_1), .Y(u2__abc_44228_n5318) );
  AND2X2 AND2X2_1614 ( .A(u2__abc_44228_n5319), .B(u2__abc_44228_n5047), .Y(u2__abc_44228_n5320) );
  AND2X2 AND2X2_1615 ( .A(u2__abc_44228_n5024), .B(u2__abc_44228_n5027), .Y(u2__abc_44228_n5321) );
  AND2X2 AND2X2_1616 ( .A(u2__abc_44228_n5324_1), .B(u2__abc_44228_n5035), .Y(u2__abc_44228_n5325) );
  AND2X2 AND2X2_1617 ( .A(u2__abc_44228_n5326), .B(u2__abc_44228_n5032_1), .Y(u2__abc_44228_n5327) );
  AND2X2 AND2X2_1618 ( .A(u2__abc_44228_n5331), .B(u2__abc_44228_n5018), .Y(u2__abc_44228_n5332) );
  AND2X2 AND2X2_1619 ( .A(u2__abc_44228_n5333_1), .B(u2__abc_44228_n5012), .Y(u2__abc_44228_n5334) );
  AND2X2 AND2X2_162 ( .A(_abc_64468_n1086), .B(_abc_64468_n1085), .Y(_auto_iopadmap_cc_313_execute_65414_197_) );
  AND2X2 AND2X2_1620 ( .A(u2__abc_44228_n5000), .B(u2__abc_44228_n5334), .Y(u2__abc_44228_n5335) );
  AND2X2 AND2X2_1621 ( .A(u2__abc_44228_n4992), .B(u2__abc_44228_n4995), .Y(u2__abc_44228_n5336) );
  AND2X2 AND2X2_1622 ( .A(u2__abc_44228_n5338), .B(u2__abc_44228_n4986_1), .Y(u2__abc_44228_n5339) );
  AND2X2 AND2X2_1623 ( .A(u2__abc_44228_n5340), .B(u2__abc_44228_n4980), .Y(u2__abc_44228_n5341) );
  AND2X2 AND2X2_1624 ( .A(u2__abc_44228_n5342), .B(u2__abc_44228_n4983), .Y(u2__abc_44228_n5343_1) );
  AND2X2 AND2X2_1625 ( .A(u2__abc_44228_n5343_1), .B(u2__abc_44228_n4971), .Y(u2__abc_44228_n5344) );
  AND2X2 AND2X2_1626 ( .A(u2__abc_44228_n4963), .B(u2__abc_44228_n4966), .Y(u2__abc_44228_n5345) );
  AND2X2 AND2X2_1627 ( .A(u2__abc_44228_n5348), .B(u2__abc_44228_n4957_1), .Y(u2__abc_44228_n5349) );
  AND2X2 AND2X2_1628 ( .A(u2__abc_44228_n5350), .B(u2__abc_44228_n4933), .Y(u2__abc_44228_n5351) );
  AND2X2 AND2X2_1629 ( .A(u2__abc_44228_n5352_1), .B(u2__abc_44228_n4950), .Y(u2__abc_44228_n5353) );
  AND2X2 AND2X2_163 ( .A(_abc_64468_n1089), .B(_abc_64468_n1088), .Y(_auto_iopadmap_cc_313_execute_65414_198_) );
  AND2X2 AND2X2_1630 ( .A(u2__abc_44228_n5354), .B(u2__abc_44228_n4953), .Y(u2__abc_44228_n5355) );
  AND2X2 AND2X2_1631 ( .A(u2__abc_44228_n5355), .B(u2__abc_44228_n4941), .Y(u2__abc_44228_n5356) );
  AND2X2 AND2X2_1632 ( .A(u2__abc_44228_n5357), .B(u2__abc_44228_n4927), .Y(u2__abc_44228_n5358) );
  AND2X2 AND2X2_1633 ( .A(u2__abc_44228_n5359), .B(u2__abc_44228_n4921_1), .Y(u2__abc_44228_n5360) );
  AND2X2 AND2X2_1634 ( .A(u2__abc_44228_n5361), .B(u2__abc_44228_n4924), .Y(u2__abc_44228_n5362_1) );
  AND2X2 AND2X2_1635 ( .A(u2__abc_44228_n5362_1), .B(u2__abc_44228_n4912), .Y(u2__abc_44228_n5363) );
  AND2X2 AND2X2_1636 ( .A(u2__abc_44228_n4904), .B(u2__abc_44228_n4907), .Y(u2__abc_44228_n5364) );
  AND2X2 AND2X2_1637 ( .A(u2__abc_44228_n5368), .B(u2__abc_44228_n4898), .Y(u2__abc_44228_n5369) );
  AND2X2 AND2X2_1638 ( .A(u2__abc_44228_n5371), .B(u2__abc_44228_n4884), .Y(u2__abc_44228_n5372_1) );
  AND2X2 AND2X2_1639 ( .A(u2__abc_44228_n5373), .B(u2__abc_44228_n4881), .Y(u2__abc_44228_n5374) );
  AND2X2 AND2X2_164 ( .A(_abc_64468_n1092), .B(_abc_64468_n1091), .Y(_auto_iopadmap_cc_313_execute_65414_199_) );
  AND2X2 AND2X2_1640 ( .A(u2__abc_44228_n4873_1), .B(u2__abc_44228_n4876), .Y(u2__abc_44228_n5375) );
  AND2X2 AND2X2_1641 ( .A(u2__abc_44228_n5377), .B(u2__abc_44228_n4867), .Y(u2__abc_44228_n5378) );
  AND2X2 AND2X2_1642 ( .A(u2__abc_44228_n5380), .B(u2__abc_44228_n4855_1), .Y(u2__abc_44228_n5381_1) );
  AND2X2 AND2X2_1643 ( .A(u2__abc_44228_n5382), .B(u2__abc_44228_n4852), .Y(u2__abc_44228_n5383) );
  AND2X2 AND2X2_1644 ( .A(u2__abc_44228_n4844), .B(u2__abc_44228_n4847), .Y(u2__abc_44228_n5384) );
  AND2X2 AND2X2_1645 ( .A(u2__abc_44228_n5387), .B(u2__abc_44228_n4838), .Y(u2__abc_44228_n5388) );
  AND2X2 AND2X2_1646 ( .A(u2__abc_44228_n5390_1), .B(u2__abc_44228_n4796), .Y(u2__abc_44228_n5391) );
  AND2X2 AND2X2_1647 ( .A(u2__abc_44228_n5392), .B(u2__abc_44228_n4793), .Y(u2__abc_44228_n5393) );
  AND2X2 AND2X2_1648 ( .A(u2__abc_44228_n4785), .B(u2__abc_44228_n4788_1), .Y(u2__abc_44228_n5394) );
  AND2X2 AND2X2_1649 ( .A(u2__abc_44228_n5398), .B(u2__abc_44228_n4811), .Y(u2__abc_44228_n5399) );
  AND2X2 AND2X2_165 ( .A(_abc_64468_n1095), .B(_abc_64468_n1094), .Y(_auto_iopadmap_cc_313_execute_65414_200_) );
  AND2X2 AND2X2_1650 ( .A(u2__abc_44228_n5400_1), .B(u2__abc_44228_n4836_1), .Y(u2__abc_44228_n5401) );
  AND2X2 AND2X2_1651 ( .A(u2__abc_44228_n4825), .B(u2__abc_44228_n5402), .Y(u2__abc_44228_n5403) );
  AND2X2 AND2X2_1652 ( .A(u2__abc_44228_n5404), .B(u2__abc_44228_n4828), .Y(u2__abc_44228_n5405) );
  AND2X2 AND2X2_1653 ( .A(u2__abc_44228_n5406), .B(u2__abc_44228_n4808), .Y(u2__abc_44228_n5407) );
  AND2X2 AND2X2_1654 ( .A(u2__abc_44228_n5411), .B(u2__abc_44228_n4779_1), .Y(u2__abc_44228_n5412) );
  AND2X2 AND2X2_1655 ( .A(u2__abc_44228_n5413), .B(u2__abc_44228_n4772), .Y(u2__abc_44228_n5414) );
  AND2X2 AND2X2_1656 ( .A(u2__abc_44228_n4760_1), .B(u2__abc_44228_n5414), .Y(u2__abc_44228_n5415) );
  AND2X2 AND2X2_1657 ( .A(u2__abc_44228_n4752), .B(u2__abc_44228_n4755), .Y(u2__abc_44228_n5416) );
  AND2X2 AND2X2_1658 ( .A(u2__abc_44228_n5418), .B(u2__abc_44228_n4746), .Y(u2__abc_44228_n5419_1) );
  AND2X2 AND2X2_1659 ( .A(u2__abc_44228_n5421), .B(u2__abc_44228_n4734), .Y(u2__abc_44228_n5422) );
  AND2X2 AND2X2_166 ( .A(_abc_64468_n1098), .B(_abc_64468_n1097), .Y(_auto_iopadmap_cc_313_execute_65414_201_) );
  AND2X2 AND2X2_1660 ( .A(u2__abc_44228_n5423), .B(u2__abc_44228_n4731_1), .Y(u2__abc_44228_n5424) );
  AND2X2 AND2X2_1661 ( .A(u2__abc_44228_n4723), .B(u2__abc_44228_n4726), .Y(u2__abc_44228_n5425) );
  AND2X2 AND2X2_1662 ( .A(u2__abc_44228_n5428_1), .B(u2__abc_44228_n4717), .Y(u2__abc_44228_n5429) );
  AND2X2 AND2X2_1663 ( .A(u2__abc_44228_n5430), .B(u2__abc_44228_n4710), .Y(u2__abc_44228_n5431) );
  AND2X2 AND2X2_1664 ( .A(u2__abc_44228_n5432), .B(u2__abc_44228_n4713_1), .Y(u2__abc_44228_n5433) );
  AND2X2 AND2X2_1665 ( .A(u2__abc_44228_n5433), .B(u2__abc_44228_n4701), .Y(u2__abc_44228_n5434) );
  AND2X2 AND2X2_1666 ( .A(u2__abc_44228_n4693), .B(u2__abc_44228_n4696), .Y(u2__abc_44228_n5435) );
  AND2X2 AND2X2_1667 ( .A(u2__abc_44228_n5437_1), .B(u2__abc_44228_n4687), .Y(u2__abc_44228_n5438) );
  AND2X2 AND2X2_1668 ( .A(u2__abc_44228_n5440), .B(u2__abc_44228_n4675), .Y(u2__abc_44228_n5441) );
  AND2X2 AND2X2_1669 ( .A(u2__abc_44228_n5442), .B(u2__abc_44228_n4672), .Y(u2__abc_44228_n5443) );
  AND2X2 AND2X2_167 ( .A(_abc_64468_n1101), .B(_abc_64468_n1100), .Y(_auto_iopadmap_cc_313_execute_65414_202_) );
  AND2X2 AND2X2_1670 ( .A(u2__abc_44228_n4664), .B(u2__abc_44228_n4667), .Y(u2__abc_44228_n5444) );
  AND2X2 AND2X2_1671 ( .A(u2__abc_44228_n5448), .B(u2__abc_44228_n4658), .Y(u2__abc_44228_n5449) );
  AND2X2 AND2X2_1672 ( .A(u2__abc_44228_n5451), .B(u2__abc_44228_n4644), .Y(u2__abc_44228_n5452) );
  AND2X2 AND2X2_1673 ( .A(u2__abc_44228_n5453), .B(u2__abc_44228_n4641), .Y(u2__abc_44228_n5454) );
  AND2X2 AND2X2_1674 ( .A(u2__abc_44228_n4633), .B(u2__abc_44228_n4636), .Y(u2__abc_44228_n5455) );
  AND2X2 AND2X2_1675 ( .A(u2__abc_44228_n5457), .B(u2__abc_44228_n4627), .Y(u2__abc_44228_n5458) );
  AND2X2 AND2X2_1676 ( .A(u2__abc_44228_n5459), .B(u2__abc_44228_n4621), .Y(u2__abc_44228_n5460) );
  AND2X2 AND2X2_1677 ( .A(u2__abc_44228_n5461), .B(u2__abc_44228_n4624), .Y(u2__abc_44228_n5462) );
  AND2X2 AND2X2_1678 ( .A(u2__abc_44228_n5462), .B(u2__abc_44228_n4612), .Y(u2__abc_44228_n5463) );
  AND2X2 AND2X2_1679 ( .A(u2__abc_44228_n4604), .B(u2__abc_44228_n4607), .Y(u2__abc_44228_n5464) );
  AND2X2 AND2X2_168 ( .A(_abc_64468_n1104), .B(_abc_64468_n1103), .Y(_auto_iopadmap_cc_313_execute_65414_203_) );
  AND2X2 AND2X2_1680 ( .A(u2__abc_44228_n5467), .B(u2__abc_44228_n4598), .Y(u2__abc_44228_n5468) );
  AND2X2 AND2X2_1681 ( .A(u2__abc_44228_n5469), .B(u2__abc_44228_n4591_1), .Y(u2__abc_44228_n5470) );
  AND2X2 AND2X2_1682 ( .A(u2__abc_44228_n5471), .B(u2__abc_44228_n4594), .Y(u2__abc_44228_n5472) );
  AND2X2 AND2X2_1683 ( .A(u2__abc_44228_n5472), .B(u2__abc_44228_n4582), .Y(u2__abc_44228_n5473) );
  AND2X2 AND2X2_1684 ( .A(u2__abc_44228_n4574), .B(u2__abc_44228_n4577), .Y(u2__abc_44228_n5474_1) );
  AND2X2 AND2X2_1685 ( .A(u2__abc_44228_n5476), .B(u2__abc_44228_n4568), .Y(u2__abc_44228_n5477) );
  AND2X2 AND2X2_1686 ( .A(u2__abc_44228_n4545_1), .B(u2__abc_44228_n4548), .Y(u2__abc_44228_n5478) );
  AND2X2 AND2X2_1687 ( .A(u2__abc_44228_n5480), .B(u2__abc_44228_n4562), .Y(u2__abc_44228_n5481) );
  AND2X2 AND2X2_1688 ( .A(u2__abc_44228_n5482), .B(u2__abc_44228_n4565), .Y(u2__abc_44228_n5483_1) );
  AND2X2 AND2X2_1689 ( .A(u2__abc_44228_n5483_1), .B(u2__abc_44228_n4553), .Y(u2__abc_44228_n5484) );
  AND2X2 AND2X2_169 ( .A(_abc_64468_n1107), .B(_abc_64468_n1106), .Y(_auto_iopadmap_cc_313_execute_65414_204_) );
  AND2X2 AND2X2_1690 ( .A(u2__abc_44228_n5488), .B(u2__abc_44228_n4539), .Y(u2__abc_44228_n5489) );
  AND2X2 AND2X2_1691 ( .A(u2__abc_44228_n5491), .B(u2__abc_44228_n4530), .Y(u2__abc_44228_n5492) );
  AND2X2 AND2X2_1692 ( .A(u2__abc_44228_n5493_1), .B(u2__abc_44228_n4521), .Y(u2__abc_44228_n5494) );
  AND2X2 AND2X2_1693 ( .A(u2__abc_44228_n4513), .B(u2__abc_44228_n4516), .Y(u2__abc_44228_n5495) );
  AND2X2 AND2X2_1694 ( .A(u2__abc_44228_n5497), .B(u2__abc_44228_n4507), .Y(u2__abc_44228_n5498) );
  AND2X2 AND2X2_1695 ( .A(u2__abc_44228_n5499), .B(u2__abc_44228_n4501), .Y(u2__abc_44228_n5500) );
  AND2X2 AND2X2_1696 ( .A(u2__abc_44228_n5501), .B(u2__abc_44228_n4504), .Y(u2__abc_44228_n5502_1) );
  AND2X2 AND2X2_1697 ( .A(u2__abc_44228_n5502_1), .B(u2__abc_44228_n4492), .Y(u2__abc_44228_n5503) );
  AND2X2 AND2X2_1698 ( .A(u2__abc_44228_n4484), .B(u2__abc_44228_n4487), .Y(u2__abc_44228_n5504) );
  AND2X2 AND2X2_1699 ( .A(u2__abc_44228_n5507), .B(u2__abc_44228_n4478), .Y(u2__abc_44228_n5508) );
  AND2X2 AND2X2_17 ( .A(_abc_64468_n753_bF_buf11), .B(sqrto_16_), .Y(_auto_iopadmap_cc_313_execute_65414_52_) );
  AND2X2 AND2X2_170 ( .A(_abc_64468_n1110), .B(_abc_64468_n1109), .Y(_auto_iopadmap_cc_313_execute_65414_205_) );
  AND2X2 AND2X2_1700 ( .A(u2__abc_44228_n5510), .B(u2__abc_44228_n4451_1), .Y(u2__abc_44228_n5511) );
  AND2X2 AND2X2_1701 ( .A(u2__abc_44228_n5512_1), .B(u2__abc_44228_n4476), .Y(u2__abc_44228_n5513) );
  AND2X2 AND2X2_1702 ( .A(u2__abc_44228_n4465), .B(u2__abc_44228_n5514), .Y(u2__abc_44228_n5515) );
  AND2X2 AND2X2_1703 ( .A(u2__abc_44228_n5516), .B(u2__abc_44228_n4468), .Y(u2__abc_44228_n5517) );
  AND2X2 AND2X2_1704 ( .A(u2__abc_44228_n5518), .B(u2__abc_44228_n4448), .Y(u2__abc_44228_n5519) );
  AND2X2 AND2X2_1705 ( .A(u2__abc_44228_n5520), .B(u2__abc_44228_n4442_1), .Y(u2__abc_44228_n5521) );
  AND2X2 AND2X2_1706 ( .A(u2__abc_44228_n5522_1), .B(u2__abc_44228_n4445), .Y(u2__abc_44228_n5523) );
  AND2X2 AND2X2_1707 ( .A(u2__abc_44228_n5523), .B(u2__abc_44228_n4433), .Y(u2__abc_44228_n5524) );
  AND2X2 AND2X2_1708 ( .A(u2__abc_44228_n4425), .B(u2__abc_44228_n4428), .Y(u2__abc_44228_n5525) );
  AND2X2 AND2X2_1709 ( .A(u2__abc_44228_n5529), .B(u2__abc_44228_n4419), .Y(u2__abc_44228_n5530) );
  AND2X2 AND2X2_171 ( .A(_abc_64468_n1113), .B(_abc_64468_n1112), .Y(_auto_iopadmap_cc_313_execute_65414_206_) );
  AND2X2 AND2X2_1710 ( .A(u2__abc_44228_n5531_1), .B(u2__abc_44228_n4352), .Y(u2__abc_44228_n5532) );
  AND2X2 AND2X2_1711 ( .A(u2__abc_44228_n5533), .B(u2__abc_44228_n4355), .Y(u2__abc_44228_n5534) );
  AND2X2 AND2X2_1712 ( .A(u2__abc_44228_n5534), .B(u2__abc_44228_n4343), .Y(u2__abc_44228_n5535) );
  AND2X2 AND2X2_1713 ( .A(u2__abc_44228_n4335), .B(u2__abc_44228_n4338_1), .Y(u2__abc_44228_n5536) );
  AND2X2 AND2X2_1714 ( .A(u2__abc_44228_n5538), .B(u2__abc_44228_n4329_1), .Y(u2__abc_44228_n5539) );
  AND2X2 AND2X2_1715 ( .A(u2__abc_44228_n5540_1), .B(u2__abc_44228_n4306), .Y(u2__abc_44228_n5541) );
  AND2X2 AND2X2_1716 ( .A(u2__abc_44228_n5542), .B(u2__abc_44228_n4323), .Y(u2__abc_44228_n5543) );
  AND2X2 AND2X2_1717 ( .A(u2__abc_44228_n5544), .B(u2__abc_44228_n4326), .Y(u2__abc_44228_n5545) );
  AND2X2 AND2X2_1718 ( .A(u2__abc_44228_n5545), .B(u2__abc_44228_n4314), .Y(u2__abc_44228_n5546) );
  AND2X2 AND2X2_1719 ( .A(u2__abc_44228_n5549_1), .B(u2__abc_44228_n4411), .Y(u2__abc_44228_n5550) );
  AND2X2 AND2X2_172 ( .A(_abc_64468_n1116), .B(_abc_64468_n1115), .Y(_auto_iopadmap_cc_313_execute_65414_207_) );
  AND2X2 AND2X2_1720 ( .A(u2__abc_44228_n5551), .B(u2__abc_44228_n4414_1), .Y(u2__abc_44228_n5552) );
  AND2X2 AND2X2_1721 ( .A(u2__abc_44228_n5552), .B(u2__abc_44228_n4402), .Y(u2__abc_44228_n5553) );
  AND2X2 AND2X2_1722 ( .A(u2__abc_44228_n4394), .B(u2__abc_44228_n4397), .Y(u2__abc_44228_n5554) );
  AND2X2 AND2X2_1723 ( .A(u2__abc_44228_n5556), .B(u2__abc_44228_n4388), .Y(u2__abc_44228_n5557) );
  AND2X2 AND2X2_1724 ( .A(u2__abc_44228_n5558_1), .B(u2__abc_44228_n4382), .Y(u2__abc_44228_n5559) );
  AND2X2 AND2X2_1725 ( .A(u2__abc_44228_n5560), .B(u2__abc_44228_n4385), .Y(u2__abc_44228_n5561) );
  AND2X2 AND2X2_1726 ( .A(u2__abc_44228_n5561), .B(u2__abc_44228_n4373), .Y(u2__abc_44228_n5562) );
  AND2X2 AND2X2_1727 ( .A(u2__abc_44228_n4365), .B(u2__abc_44228_n4368_1), .Y(u2__abc_44228_n5563) );
  AND2X2 AND2X2_1728 ( .A(u2__abc_44228_n5566), .B(u2__abc_44228_n4359_1), .Y(u2__abc_44228_n5567) );
  AND2X2 AND2X2_1729 ( .A(u2__abc_44228_n5573), .B(u2_remHi_381_), .Y(u2__abc_44228_n5574) );
  AND2X2 AND2X2_173 ( .A(_abc_64468_n1119), .B(_abc_64468_n1118), .Y(_auto_iopadmap_cc_313_execute_65414_208_) );
  AND2X2 AND2X2_1730 ( .A(u2__abc_44228_n5576), .B(u2_o_381_), .Y(u2__abc_44228_n5577_1) );
  AND2X2 AND2X2_1731 ( .A(u2__abc_44228_n5575), .B(u2__abc_44228_n5578), .Y(u2__abc_44228_n5579) );
  AND2X2 AND2X2_1732 ( .A(u2__abc_44228_n5580), .B(u2_remHi_380_), .Y(u2__abc_44228_n5581) );
  AND2X2 AND2X2_1733 ( .A(u2__abc_44228_n5582), .B(u2_o_380_), .Y(u2__abc_44228_n5583) );
  AND2X2 AND2X2_1734 ( .A(u2__abc_44228_n5585), .B(u2__abc_44228_n5579), .Y(u2__abc_44228_n5586) );
  AND2X2 AND2X2_1735 ( .A(u2__abc_44228_n5587_1), .B(u2_remHi_379_), .Y(u2__abc_44228_n5588) );
  AND2X2 AND2X2_1736 ( .A(u2__abc_44228_n5590), .B(u2_o_379_), .Y(u2__abc_44228_n5591) );
  AND2X2 AND2X2_1737 ( .A(u2__abc_44228_n5589), .B(u2__abc_44228_n5592), .Y(u2__abc_44228_n5593) );
  AND2X2 AND2X2_1738 ( .A(u2__abc_44228_n5594), .B(u2_remHi_378_), .Y(u2__abc_44228_n5595) );
  AND2X2 AND2X2_1739 ( .A(u2__abc_44228_n5596), .B(u2_o_378_), .Y(u2__abc_44228_n5597_1) );
  AND2X2 AND2X2_174 ( .A(_abc_64468_n1122), .B(_abc_64468_n1121), .Y(_auto_iopadmap_cc_313_execute_65414_209_) );
  AND2X2 AND2X2_1740 ( .A(u2__abc_44228_n5599), .B(u2__abc_44228_n5593), .Y(u2__abc_44228_n5600) );
  AND2X2 AND2X2_1741 ( .A(u2__abc_44228_n5586), .B(u2__abc_44228_n5600), .Y(u2__abc_44228_n5601) );
  AND2X2 AND2X2_1742 ( .A(u2__abc_44228_n5602), .B(u2_remHi_375_), .Y(u2__abc_44228_n5603) );
  AND2X2 AND2X2_1743 ( .A(u2__abc_44228_n5605), .B(u2_o_375_), .Y(u2__abc_44228_n5606_1) );
  AND2X2 AND2X2_1744 ( .A(u2__abc_44228_n5604), .B(u2__abc_44228_n5607), .Y(u2__abc_44228_n5608) );
  AND2X2 AND2X2_1745 ( .A(u2__abc_44228_n5609), .B(u2_remHi_374_), .Y(u2__abc_44228_n5610) );
  AND2X2 AND2X2_1746 ( .A(u2__abc_44228_n5611), .B(u2_o_374_), .Y(u2__abc_44228_n5612) );
  AND2X2 AND2X2_1747 ( .A(u2__abc_44228_n5614), .B(u2__abc_44228_n5608), .Y(u2__abc_44228_n5615_1) );
  AND2X2 AND2X2_1748 ( .A(u2__abc_44228_n5616), .B(u2_remHi_377_), .Y(u2__abc_44228_n5617) );
  AND2X2 AND2X2_1749 ( .A(u2__abc_44228_n5619), .B(u2_o_377_), .Y(u2__abc_44228_n5620) );
  AND2X2 AND2X2_175 ( .A(_abc_64468_n1125), .B(_abc_64468_n1124), .Y(_auto_iopadmap_cc_313_execute_65414_210_) );
  AND2X2 AND2X2_1750 ( .A(u2__abc_44228_n5618), .B(u2__abc_44228_n5621), .Y(u2__abc_44228_n5622) );
  AND2X2 AND2X2_1751 ( .A(u2__abc_44228_n5623), .B(u2_remHi_376_), .Y(u2__abc_44228_n5624_1) );
  AND2X2 AND2X2_1752 ( .A(u2__abc_44228_n5625), .B(u2_o_376_), .Y(u2__abc_44228_n5626) );
  AND2X2 AND2X2_1753 ( .A(u2__abc_44228_n5628), .B(u2__abc_44228_n5622), .Y(u2__abc_44228_n5629) );
  AND2X2 AND2X2_1754 ( .A(u2__abc_44228_n5615_1), .B(u2__abc_44228_n5629), .Y(u2__abc_44228_n5630) );
  AND2X2 AND2X2_1755 ( .A(u2__abc_44228_n5601), .B(u2__abc_44228_n5630), .Y(u2__abc_44228_n5631) );
  AND2X2 AND2X2_1756 ( .A(u2__abc_44228_n5632), .B(u2_remHi_373_), .Y(u2__abc_44228_n5633_1) );
  AND2X2 AND2X2_1757 ( .A(u2__abc_44228_n5635), .B(u2_o_373_), .Y(u2__abc_44228_n5636) );
  AND2X2 AND2X2_1758 ( .A(u2__abc_44228_n5634), .B(u2__abc_44228_n5637), .Y(u2__abc_44228_n5638) );
  AND2X2 AND2X2_1759 ( .A(u2__abc_44228_n5639), .B(u2_remHi_372_), .Y(u2__abc_44228_n5640) );
  AND2X2 AND2X2_176 ( .A(_abc_64468_n1128), .B(_abc_64468_n1127), .Y(_auto_iopadmap_cc_313_execute_65414_211_) );
  AND2X2 AND2X2_1760 ( .A(u2__abc_44228_n5641), .B(u2_o_372_), .Y(u2__abc_44228_n5642) );
  AND2X2 AND2X2_1761 ( .A(u2__abc_44228_n5644), .B(u2__abc_44228_n5638), .Y(u2__abc_44228_n5645) );
  AND2X2 AND2X2_1762 ( .A(u2__abc_44228_n5646), .B(u2_remHi_370_), .Y(u2__abc_44228_n5647) );
  AND2X2 AND2X2_1763 ( .A(u2__abc_44228_n5648), .B(u2_o_370_), .Y(u2__abc_44228_n5649) );
  AND2X2 AND2X2_1764 ( .A(u2__abc_44228_n5652_1), .B(u2_remHi_371_), .Y(u2__abc_44228_n5653) );
  AND2X2 AND2X2_1765 ( .A(u2__abc_44228_n5655), .B(u2_o_371_), .Y(u2__abc_44228_n5656) );
  AND2X2 AND2X2_1766 ( .A(u2__abc_44228_n5654), .B(u2__abc_44228_n5657), .Y(u2__abc_44228_n5658) );
  AND2X2 AND2X2_1767 ( .A(u2__abc_44228_n5651), .B(u2__abc_44228_n5658), .Y(u2__abc_44228_n5659) );
  AND2X2 AND2X2_1768 ( .A(u2__abc_44228_n5645), .B(u2__abc_44228_n5659), .Y(u2__abc_44228_n5660) );
  AND2X2 AND2X2_1769 ( .A(u2__abc_44228_n5661), .B(u2_remHi_367_), .Y(u2__abc_44228_n5662_1) );
  AND2X2 AND2X2_177 ( .A(_abc_64468_n1131), .B(_abc_64468_n1130), .Y(_auto_iopadmap_cc_313_execute_65414_212_) );
  AND2X2 AND2X2_1770 ( .A(u2__abc_44228_n5664), .B(u2_o_367_), .Y(u2__abc_44228_n5665) );
  AND2X2 AND2X2_1771 ( .A(u2__abc_44228_n5663), .B(u2__abc_44228_n5666), .Y(u2__abc_44228_n5667) );
  AND2X2 AND2X2_1772 ( .A(u2__abc_44228_n5668), .B(u2_remHi_366_), .Y(u2__abc_44228_n5669) );
  AND2X2 AND2X2_1773 ( .A(u2__abc_44228_n5670), .B(u2_o_366_), .Y(u2__abc_44228_n5671) );
  AND2X2 AND2X2_1774 ( .A(u2__abc_44228_n5673), .B(u2__abc_44228_n5667), .Y(u2__abc_44228_n5674) );
  AND2X2 AND2X2_1775 ( .A(u2__abc_44228_n5675), .B(u2_remHi_369_), .Y(u2__abc_44228_n5676) );
  AND2X2 AND2X2_1776 ( .A(u2__abc_44228_n5678), .B(u2_o_369_), .Y(u2__abc_44228_n5679) );
  AND2X2 AND2X2_1777 ( .A(u2__abc_44228_n5677), .B(u2__abc_44228_n5680), .Y(u2__abc_44228_n5681_1) );
  AND2X2 AND2X2_1778 ( .A(u2__abc_44228_n5682), .B(u2_remHi_368_), .Y(u2__abc_44228_n5683) );
  AND2X2 AND2X2_1779 ( .A(u2__abc_44228_n5684), .B(u2_o_368_), .Y(u2__abc_44228_n5685) );
  AND2X2 AND2X2_178 ( .A(_abc_64468_n1134), .B(_abc_64468_n1133), .Y(_auto_iopadmap_cc_313_execute_65414_213_) );
  AND2X2 AND2X2_1780 ( .A(u2__abc_44228_n5687), .B(u2__abc_44228_n5681_1), .Y(u2__abc_44228_n5688) );
  AND2X2 AND2X2_1781 ( .A(u2__abc_44228_n5674), .B(u2__abc_44228_n5688), .Y(u2__abc_44228_n5689) );
  AND2X2 AND2X2_1782 ( .A(u2__abc_44228_n5660), .B(u2__abc_44228_n5689), .Y(u2__abc_44228_n5690_1) );
  AND2X2 AND2X2_1783 ( .A(u2__abc_44228_n5631), .B(u2__abc_44228_n5690_1), .Y(u2__abc_44228_n5691) );
  AND2X2 AND2X2_1784 ( .A(u2__abc_44228_n5692), .B(u2_remHi_365_), .Y(u2__abc_44228_n5693) );
  AND2X2 AND2X2_1785 ( .A(u2__abc_44228_n5695), .B(u2_o_365_), .Y(u2__abc_44228_n5696) );
  AND2X2 AND2X2_1786 ( .A(u2__abc_44228_n5694), .B(u2__abc_44228_n5697), .Y(u2__abc_44228_n5698) );
  AND2X2 AND2X2_1787 ( .A(u2__abc_44228_n5699), .B(u2_remHi_364_), .Y(u2__abc_44228_n5700_1) );
  AND2X2 AND2X2_1788 ( .A(u2__abc_44228_n5701), .B(u2_o_364_), .Y(u2__abc_44228_n5702) );
  AND2X2 AND2X2_1789 ( .A(u2__abc_44228_n5704), .B(u2__abc_44228_n5698), .Y(u2__abc_44228_n5705) );
  AND2X2 AND2X2_179 ( .A(_abc_64468_n1137), .B(_abc_64468_n1136), .Y(_auto_iopadmap_cc_313_execute_65414_214_) );
  AND2X2 AND2X2_1790 ( .A(u2__abc_44228_n5706), .B(u2_remHi_363_), .Y(u2__abc_44228_n5707) );
  AND2X2 AND2X2_1791 ( .A(u2__abc_44228_n5709), .B(u2_o_363_), .Y(u2__abc_44228_n5710_1) );
  AND2X2 AND2X2_1792 ( .A(u2__abc_44228_n5708), .B(u2__abc_44228_n5711), .Y(u2__abc_44228_n5712) );
  AND2X2 AND2X2_1793 ( .A(u2__abc_44228_n5713), .B(u2_remHi_362_), .Y(u2__abc_44228_n5714) );
  AND2X2 AND2X2_1794 ( .A(u2__abc_44228_n5715), .B(u2_o_362_), .Y(u2__abc_44228_n5716) );
  AND2X2 AND2X2_1795 ( .A(u2__abc_44228_n5718), .B(u2__abc_44228_n5712), .Y(u2__abc_44228_n5719_1) );
  AND2X2 AND2X2_1796 ( .A(u2__abc_44228_n5705), .B(u2__abc_44228_n5719_1), .Y(u2__abc_44228_n5720) );
  AND2X2 AND2X2_1797 ( .A(u2__abc_44228_n5721), .B(u2_remHi_359_), .Y(u2__abc_44228_n5722) );
  AND2X2 AND2X2_1798 ( .A(u2__abc_44228_n5724), .B(u2_o_359_), .Y(u2__abc_44228_n5725) );
  AND2X2 AND2X2_1799 ( .A(u2__abc_44228_n5723), .B(u2__abc_44228_n5726), .Y(u2__abc_44228_n5727) );
  AND2X2 AND2X2_18 ( .A(_abc_64468_n753_bF_buf10), .B(sqrto_17_), .Y(_auto_iopadmap_cc_313_execute_65414_53_) );
  AND2X2 AND2X2_180 ( .A(_abc_64468_n1140), .B(_abc_64468_n1139), .Y(_auto_iopadmap_cc_313_execute_65414_215_) );
  AND2X2 AND2X2_1800 ( .A(u2__abc_44228_n5728_1), .B(u2_remHi_358_), .Y(u2__abc_44228_n5729) );
  AND2X2 AND2X2_1801 ( .A(u2__abc_44228_n5730), .B(u2_o_358_), .Y(u2__abc_44228_n5731) );
  AND2X2 AND2X2_1802 ( .A(u2__abc_44228_n5733), .B(u2__abc_44228_n5727), .Y(u2__abc_44228_n5734) );
  AND2X2 AND2X2_1803 ( .A(u2__abc_44228_n5735), .B(u2_remHi_361_), .Y(u2__abc_44228_n5736) );
  AND2X2 AND2X2_1804 ( .A(u2__abc_44228_n5738), .B(u2_o_361_), .Y(u2__abc_44228_n5739) );
  AND2X2 AND2X2_1805 ( .A(u2__abc_44228_n5737_1), .B(u2__abc_44228_n5740), .Y(u2__abc_44228_n5741) );
  AND2X2 AND2X2_1806 ( .A(u2__abc_44228_n5742), .B(u2_remHi_360_), .Y(u2__abc_44228_n5743) );
  AND2X2 AND2X2_1807 ( .A(u2__abc_44228_n5744), .B(u2_o_360_), .Y(u2__abc_44228_n5745) );
  AND2X2 AND2X2_1808 ( .A(u2__abc_44228_n5747_1), .B(u2__abc_44228_n5741), .Y(u2__abc_44228_n5748) );
  AND2X2 AND2X2_1809 ( .A(u2__abc_44228_n5734), .B(u2__abc_44228_n5748), .Y(u2__abc_44228_n5749) );
  AND2X2 AND2X2_181 ( .A(_abc_64468_n1143), .B(_abc_64468_n1142), .Y(_auto_iopadmap_cc_313_execute_65414_216_) );
  AND2X2 AND2X2_1810 ( .A(u2__abc_44228_n5720), .B(u2__abc_44228_n5749), .Y(u2__abc_44228_n5750) );
  AND2X2 AND2X2_1811 ( .A(u2__abc_44228_n5751), .B(u2_remHi_357_), .Y(u2__abc_44228_n5752) );
  AND2X2 AND2X2_1812 ( .A(u2__abc_44228_n5754), .B(u2_o_357_), .Y(u2__abc_44228_n5755) );
  AND2X2 AND2X2_1813 ( .A(u2__abc_44228_n5753), .B(u2__abc_44228_n5756_1), .Y(u2__abc_44228_n5757) );
  AND2X2 AND2X2_1814 ( .A(u2__abc_44228_n5758), .B(u2_remHi_356_), .Y(u2__abc_44228_n5759) );
  AND2X2 AND2X2_1815 ( .A(u2__abc_44228_n5760), .B(u2_o_356_), .Y(u2__abc_44228_n5761) );
  AND2X2 AND2X2_1816 ( .A(u2__abc_44228_n5763), .B(u2__abc_44228_n5757), .Y(u2__abc_44228_n5764) );
  AND2X2 AND2X2_1817 ( .A(u2__abc_44228_n5765_1), .B(u2_remHi_354_), .Y(u2__abc_44228_n5766) );
  AND2X2 AND2X2_1818 ( .A(u2__abc_44228_n5767), .B(u2_o_354_), .Y(u2__abc_44228_n5768) );
  AND2X2 AND2X2_1819 ( .A(u2__abc_44228_n5771), .B(u2_remHi_355_), .Y(u2__abc_44228_n5772) );
  AND2X2 AND2X2_182 ( .A(_abc_64468_n1146), .B(_abc_64468_n1145), .Y(_auto_iopadmap_cc_313_execute_65414_217_) );
  AND2X2 AND2X2_1820 ( .A(u2__abc_44228_n5774_1), .B(u2_o_355_), .Y(u2__abc_44228_n5775) );
  AND2X2 AND2X2_1821 ( .A(u2__abc_44228_n5773), .B(u2__abc_44228_n5776), .Y(u2__abc_44228_n5777) );
  AND2X2 AND2X2_1822 ( .A(u2__abc_44228_n5770), .B(u2__abc_44228_n5777), .Y(u2__abc_44228_n5778) );
  AND2X2 AND2X2_1823 ( .A(u2__abc_44228_n5764), .B(u2__abc_44228_n5778), .Y(u2__abc_44228_n5779) );
  AND2X2 AND2X2_1824 ( .A(u2__abc_44228_n5780), .B(u2_remHi_353_), .Y(u2__abc_44228_n5781) );
  AND2X2 AND2X2_1825 ( .A(u2__abc_44228_n5783_1), .B(u2_o_353_), .Y(u2__abc_44228_n5784) );
  AND2X2 AND2X2_1826 ( .A(u2__abc_44228_n5782), .B(u2__abc_44228_n5785), .Y(u2__abc_44228_n5786) );
  AND2X2 AND2X2_1827 ( .A(u2__abc_44228_n5787), .B(u2_remHi_352_), .Y(u2__abc_44228_n5788) );
  AND2X2 AND2X2_1828 ( .A(u2__abc_44228_n5789), .B(u2_o_352_), .Y(u2__abc_44228_n5790) );
  AND2X2 AND2X2_1829 ( .A(u2__abc_44228_n5792), .B(u2__abc_44228_n5786), .Y(u2__abc_44228_n5793_1) );
  AND2X2 AND2X2_183 ( .A(_abc_64468_n1149), .B(_abc_64468_n1148), .Y(_auto_iopadmap_cc_313_execute_65414_218_) );
  AND2X2 AND2X2_1830 ( .A(u2__abc_44228_n5794), .B(u2_remHi_351_), .Y(u2__abc_44228_n5795) );
  AND2X2 AND2X2_1831 ( .A(u2__abc_44228_n5797), .B(u2_o_351_), .Y(u2__abc_44228_n5798) );
  AND2X2 AND2X2_1832 ( .A(u2__abc_44228_n5796), .B(u2__abc_44228_n5799), .Y(u2__abc_44228_n5800) );
  AND2X2 AND2X2_1833 ( .A(u2__abc_44228_n5801), .B(u2_remHi_350_), .Y(u2__abc_44228_n5802_1) );
  AND2X2 AND2X2_1834 ( .A(u2__abc_44228_n5803), .B(u2_o_350_), .Y(u2__abc_44228_n5804) );
  AND2X2 AND2X2_1835 ( .A(u2__abc_44228_n5806), .B(u2__abc_44228_n5800), .Y(u2__abc_44228_n5807) );
  AND2X2 AND2X2_1836 ( .A(u2__abc_44228_n5793_1), .B(u2__abc_44228_n5807), .Y(u2__abc_44228_n5808) );
  AND2X2 AND2X2_1837 ( .A(u2__abc_44228_n5779), .B(u2__abc_44228_n5808), .Y(u2__abc_44228_n5809) );
  AND2X2 AND2X2_1838 ( .A(u2__abc_44228_n5750), .B(u2__abc_44228_n5809), .Y(u2__abc_44228_n5810) );
  AND2X2 AND2X2_1839 ( .A(u2__abc_44228_n5691), .B(u2__abc_44228_n5810), .Y(u2__abc_44228_n5811) );
  AND2X2 AND2X2_184 ( .A(_abc_64468_n1152), .B(_abc_64468_n1151), .Y(_auto_iopadmap_cc_313_execute_65414_219_) );
  AND2X2 AND2X2_1840 ( .A(u2__abc_44228_n5812_1), .B(u2_remHi_349_), .Y(u2__abc_44228_n5813) );
  AND2X2 AND2X2_1841 ( .A(u2__abc_44228_n5815), .B(u2_o_349_), .Y(u2__abc_44228_n5816) );
  AND2X2 AND2X2_1842 ( .A(u2__abc_44228_n5814), .B(u2__abc_44228_n5817), .Y(u2__abc_44228_n5818) );
  AND2X2 AND2X2_1843 ( .A(u2__abc_44228_n5819), .B(u2_remHi_348_), .Y(u2__abc_44228_n5820) );
  AND2X2 AND2X2_1844 ( .A(u2__abc_44228_n5821), .B(u2_o_348_), .Y(u2__abc_44228_n5822_1) );
  AND2X2 AND2X2_1845 ( .A(u2__abc_44228_n5824), .B(u2__abc_44228_n5818), .Y(u2__abc_44228_n5825) );
  AND2X2 AND2X2_1846 ( .A(u2__abc_44228_n5826), .B(u2_remHi_346_), .Y(u2__abc_44228_n5827) );
  AND2X2 AND2X2_1847 ( .A(u2__abc_44228_n5828), .B(u2_o_346_), .Y(u2__abc_44228_n5829) );
  AND2X2 AND2X2_1848 ( .A(u2__abc_44228_n5832), .B(u2_remHi_347_), .Y(u2__abc_44228_n5833) );
  AND2X2 AND2X2_1849 ( .A(u2__abc_44228_n5835), .B(u2_o_347_), .Y(u2__abc_44228_n5836) );
  AND2X2 AND2X2_185 ( .A(_abc_64468_n1155), .B(_abc_64468_n1154), .Y(_auto_iopadmap_cc_313_execute_65414_220_) );
  AND2X2 AND2X2_1850 ( .A(u2__abc_44228_n5834), .B(u2__abc_44228_n5837), .Y(u2__abc_44228_n5838_1) );
  AND2X2 AND2X2_1851 ( .A(u2__abc_44228_n5831), .B(u2__abc_44228_n5838_1), .Y(u2__abc_44228_n5839) );
  AND2X2 AND2X2_1852 ( .A(u2__abc_44228_n5825), .B(u2__abc_44228_n5839), .Y(u2__abc_44228_n5840) );
  AND2X2 AND2X2_1853 ( .A(u2__abc_44228_n5841), .B(u2_remHi_343_), .Y(u2__abc_44228_n5842) );
  AND2X2 AND2X2_1854 ( .A(u2__abc_44228_n5844), .B(u2_o_343_), .Y(u2__abc_44228_n5845_1) );
  AND2X2 AND2X2_1855 ( .A(u2__abc_44228_n5843), .B(u2__abc_44228_n5846), .Y(u2__abc_44228_n5847) );
  AND2X2 AND2X2_1856 ( .A(u2__abc_44228_n5848), .B(u2_remHi_342_), .Y(u2__abc_44228_n5849) );
  AND2X2 AND2X2_1857 ( .A(u2__abc_44228_n5850), .B(u2_o_342_), .Y(u2__abc_44228_n5851) );
  AND2X2 AND2X2_1858 ( .A(u2__abc_44228_n5853), .B(u2__abc_44228_n5847), .Y(u2__abc_44228_n5854_1) );
  AND2X2 AND2X2_1859 ( .A(u2__abc_44228_n5855), .B(u2_remHi_345_), .Y(u2__abc_44228_n5856) );
  AND2X2 AND2X2_186 ( .A(_abc_64468_n1158), .B(_abc_64468_n1157), .Y(_auto_iopadmap_cc_313_execute_65414_221_) );
  AND2X2 AND2X2_1860 ( .A(u2__abc_44228_n5858), .B(u2_o_345_), .Y(u2__abc_44228_n5859) );
  AND2X2 AND2X2_1861 ( .A(u2__abc_44228_n5857), .B(u2__abc_44228_n5860), .Y(u2__abc_44228_n5861) );
  AND2X2 AND2X2_1862 ( .A(u2__abc_44228_n5862), .B(u2_remHi_344_), .Y(u2__abc_44228_n5863_1) );
  AND2X2 AND2X2_1863 ( .A(u2__abc_44228_n5864), .B(u2_o_344_), .Y(u2__abc_44228_n5865) );
  AND2X2 AND2X2_1864 ( .A(u2__abc_44228_n5867), .B(u2__abc_44228_n5861), .Y(u2__abc_44228_n5868) );
  AND2X2 AND2X2_1865 ( .A(u2__abc_44228_n5854_1), .B(u2__abc_44228_n5868), .Y(u2__abc_44228_n5869) );
  AND2X2 AND2X2_1866 ( .A(u2__abc_44228_n5840), .B(u2__abc_44228_n5869), .Y(u2__abc_44228_n5870) );
  AND2X2 AND2X2_1867 ( .A(u2__abc_44228_n5871), .B(u2_remHi_341_), .Y(u2__abc_44228_n5872) );
  AND2X2 AND2X2_1868 ( .A(u2__abc_44228_n5874), .B(u2_o_341_), .Y(u2__abc_44228_n5875) );
  AND2X2 AND2X2_1869 ( .A(u2__abc_44228_n5873_1), .B(u2__abc_44228_n5876), .Y(u2__abc_44228_n5877) );
  AND2X2 AND2X2_187 ( .A(_abc_64468_n1161), .B(_abc_64468_n1160), .Y(_auto_iopadmap_cc_313_execute_65414_222_) );
  AND2X2 AND2X2_1870 ( .A(u2__abc_44228_n5878), .B(u2_remHi_340_), .Y(u2__abc_44228_n5879) );
  AND2X2 AND2X2_1871 ( .A(u2__abc_44228_n5880), .B(u2_o_340_), .Y(u2__abc_44228_n5881) );
  AND2X2 AND2X2_1872 ( .A(u2__abc_44228_n5883_1), .B(u2__abc_44228_n5877), .Y(u2__abc_44228_n5884) );
  AND2X2 AND2X2_1873 ( .A(u2__abc_44228_n5885), .B(u2_remHi_338_), .Y(u2__abc_44228_n5886) );
  AND2X2 AND2X2_1874 ( .A(u2__abc_44228_n5887), .B(u2_o_338_), .Y(u2__abc_44228_n5888) );
  AND2X2 AND2X2_1875 ( .A(u2__abc_44228_n5891), .B(u2_remHi_339_), .Y(u2__abc_44228_n5892_1) );
  AND2X2 AND2X2_1876 ( .A(u2__abc_44228_n5894), .B(u2_o_339_), .Y(u2__abc_44228_n5895) );
  AND2X2 AND2X2_1877 ( .A(u2__abc_44228_n5893), .B(u2__abc_44228_n5896), .Y(u2__abc_44228_n5897) );
  AND2X2 AND2X2_1878 ( .A(u2__abc_44228_n5890), .B(u2__abc_44228_n5897), .Y(u2__abc_44228_n5898) );
  AND2X2 AND2X2_1879 ( .A(u2__abc_44228_n5884), .B(u2__abc_44228_n5898), .Y(u2__abc_44228_n5899) );
  AND2X2 AND2X2_188 ( .A(_abc_64468_n1164), .B(_abc_64468_n1163), .Y(_auto_iopadmap_cc_313_execute_65414_223_) );
  AND2X2 AND2X2_1880 ( .A(u2__abc_44228_n5900), .B(u2_remHi_337_), .Y(u2__abc_44228_n5901_1) );
  AND2X2 AND2X2_1881 ( .A(u2__abc_44228_n5903), .B(u2_o_337_), .Y(u2__abc_44228_n5904) );
  AND2X2 AND2X2_1882 ( .A(u2__abc_44228_n5902), .B(u2__abc_44228_n5905), .Y(u2__abc_44228_n5906) );
  AND2X2 AND2X2_1883 ( .A(u2__abc_44228_n5907), .B(u2_remHi_336_), .Y(u2__abc_44228_n5908) );
  AND2X2 AND2X2_1884 ( .A(u2__abc_44228_n5909), .B(u2_o_336_), .Y(u2__abc_44228_n5910) );
  AND2X2 AND2X2_1885 ( .A(u2__abc_44228_n5912), .B(u2__abc_44228_n5906), .Y(u2__abc_44228_n5913) );
  AND2X2 AND2X2_1886 ( .A(u2__abc_44228_n5914), .B(u2_remHi_335_), .Y(u2__abc_44228_n5915) );
  AND2X2 AND2X2_1887 ( .A(u2__abc_44228_n5917), .B(u2_o_335_), .Y(u2__abc_44228_n5918) );
  AND2X2 AND2X2_1888 ( .A(u2__abc_44228_n5916), .B(u2__abc_44228_n5919), .Y(u2__abc_44228_n5920_1) );
  AND2X2 AND2X2_1889 ( .A(u2__abc_44228_n5921), .B(u2_remHi_334_), .Y(u2__abc_44228_n5922) );
  AND2X2 AND2X2_189 ( .A(_abc_64468_n753_bF_buf7), .B(sqrto_189_), .Y(_auto_iopadmap_cc_313_execute_65414_225_) );
  AND2X2 AND2X2_1890 ( .A(u2__abc_44228_n5923), .B(u2_o_334_), .Y(u2__abc_44228_n5924) );
  AND2X2 AND2X2_1891 ( .A(u2__abc_44228_n5926), .B(u2__abc_44228_n5920_1), .Y(u2__abc_44228_n5927) );
  AND2X2 AND2X2_1892 ( .A(u2__abc_44228_n5913), .B(u2__abc_44228_n5927), .Y(u2__abc_44228_n5928) );
  AND2X2 AND2X2_1893 ( .A(u2__abc_44228_n5899), .B(u2__abc_44228_n5928), .Y(u2__abc_44228_n5929) );
  AND2X2 AND2X2_1894 ( .A(u2__abc_44228_n5870), .B(u2__abc_44228_n5929), .Y(u2__abc_44228_n5930_1) );
  AND2X2 AND2X2_1895 ( .A(u2__abc_44228_n5931), .B(u2_remHi_333_), .Y(u2__abc_44228_n5932) );
  AND2X2 AND2X2_1896 ( .A(u2__abc_44228_n5934), .B(u2_o_333_), .Y(u2__abc_44228_n5935) );
  AND2X2 AND2X2_1897 ( .A(u2__abc_44228_n5933), .B(u2__abc_44228_n5936), .Y(u2__abc_44228_n5937) );
  AND2X2 AND2X2_1898 ( .A(u2__abc_44228_n5938_1), .B(u2_remHi_332_), .Y(u2__abc_44228_n5939) );
  AND2X2 AND2X2_1899 ( .A(u2__abc_44228_n5940), .B(u2_o_332_), .Y(u2__abc_44228_n5941) );
  AND2X2 AND2X2_19 ( .A(_abc_64468_n753_bF_buf9), .B(sqrto_18_), .Y(_auto_iopadmap_cc_313_execute_65414_54_) );
  AND2X2 AND2X2_190 ( .A(a_112_bF_buf9), .B(\a[0] ), .Y(fracta1_0_) );
  AND2X2 AND2X2_1900 ( .A(u2__abc_44228_n5943), .B(u2__abc_44228_n5937), .Y(u2__abc_44228_n5944) );
  AND2X2 AND2X2_1901 ( .A(u2__abc_44228_n5945), .B(u2_remHi_331_), .Y(u2__abc_44228_n5946) );
  AND2X2 AND2X2_1902 ( .A(u2__abc_44228_n5948_1), .B(u2_o_331_), .Y(u2__abc_44228_n5949) );
  AND2X2 AND2X2_1903 ( .A(u2__abc_44228_n5947), .B(u2__abc_44228_n5950), .Y(u2__abc_44228_n5951) );
  AND2X2 AND2X2_1904 ( .A(u2__abc_44228_n5952), .B(u2_remHi_330_), .Y(u2__abc_44228_n5953) );
  AND2X2 AND2X2_1905 ( .A(u2__abc_44228_n5954), .B(u2_o_330_), .Y(u2__abc_44228_n5955) );
  AND2X2 AND2X2_1906 ( .A(u2__abc_44228_n5957_1), .B(u2__abc_44228_n5951), .Y(u2__abc_44228_n5958) );
  AND2X2 AND2X2_1907 ( .A(u2__abc_44228_n5944), .B(u2__abc_44228_n5958), .Y(u2__abc_44228_n5959) );
  AND2X2 AND2X2_1908 ( .A(u2__abc_44228_n5960), .B(u2_remHi_329_), .Y(u2__abc_44228_n5961) );
  AND2X2 AND2X2_1909 ( .A(u2__abc_44228_n5963), .B(u2_o_329_), .Y(u2__abc_44228_n5964) );
  AND2X2 AND2X2_191 ( .A(_abc_64468_n1171), .B(_abc_64468_n1169), .Y(fracta1_1_) );
  AND2X2 AND2X2_1910 ( .A(u2__abc_44228_n5962), .B(u2__abc_44228_n5965), .Y(u2__abc_44228_n5966_1) );
  AND2X2 AND2X2_1911 ( .A(u2__abc_44228_n5967), .B(u2_remHi_328_), .Y(u2__abc_44228_n5968) );
  AND2X2 AND2X2_1912 ( .A(u2__abc_44228_n5969), .B(u2_o_328_), .Y(u2__abc_44228_n5970) );
  AND2X2 AND2X2_1913 ( .A(u2__abc_44228_n5972), .B(u2__abc_44228_n5966_1), .Y(u2__abc_44228_n5973) );
  AND2X2 AND2X2_1914 ( .A(u2__abc_44228_n5974), .B(u2_remHi_327_), .Y(u2__abc_44228_n5975_1) );
  AND2X2 AND2X2_1915 ( .A(u2__abc_44228_n5977), .B(u2_o_327_), .Y(u2__abc_44228_n5978) );
  AND2X2 AND2X2_1916 ( .A(u2__abc_44228_n5976), .B(u2__abc_44228_n5979), .Y(u2__abc_44228_n5980) );
  AND2X2 AND2X2_1917 ( .A(u2__abc_44228_n5981), .B(u2_remHi_326_), .Y(u2__abc_44228_n5982) );
  AND2X2 AND2X2_1918 ( .A(u2__abc_44228_n5983), .B(u2_o_326_), .Y(u2__abc_44228_n5984) );
  AND2X2 AND2X2_1919 ( .A(u2__abc_44228_n5986), .B(u2__abc_44228_n5980), .Y(u2__abc_44228_n5987) );
  AND2X2 AND2X2_192 ( .A(_abc_64468_n1174), .B(_abc_64468_n1173), .Y(fracta1_2_) );
  AND2X2 AND2X2_1920 ( .A(u2__abc_44228_n5973), .B(u2__abc_44228_n5987), .Y(u2__abc_44228_n5988) );
  AND2X2 AND2X2_1921 ( .A(u2__abc_44228_n5959), .B(u2__abc_44228_n5988), .Y(u2__abc_44228_n5989) );
  AND2X2 AND2X2_1922 ( .A(u2__abc_44228_n5990), .B(u2_remHi_325_), .Y(u2__abc_44228_n5991) );
  AND2X2 AND2X2_1923 ( .A(u2__abc_44228_n5993), .B(u2_o_325_), .Y(u2__abc_44228_n5994_1) );
  AND2X2 AND2X2_1924 ( .A(u2__abc_44228_n5992), .B(u2__abc_44228_n5995), .Y(u2__abc_44228_n5996) );
  AND2X2 AND2X2_1925 ( .A(u2__abc_44228_n5997), .B(u2_remHi_324_), .Y(u2__abc_44228_n5998) );
  AND2X2 AND2X2_1926 ( .A(u2__abc_44228_n5999), .B(u2_o_324_), .Y(u2__abc_44228_n6000) );
  AND2X2 AND2X2_1927 ( .A(u2__abc_44228_n6002), .B(u2__abc_44228_n5996), .Y(u2__abc_44228_n6003_1) );
  AND2X2 AND2X2_1928 ( .A(u2__abc_44228_n6004), .B(u2_remHi_322_), .Y(u2__abc_44228_n6005) );
  AND2X2 AND2X2_1929 ( .A(u2__abc_44228_n6006), .B(u2_o_322_), .Y(u2__abc_44228_n6007) );
  AND2X2 AND2X2_193 ( .A(_abc_64468_n1177), .B(_abc_64468_n1176), .Y(fracta1_3_) );
  AND2X2 AND2X2_1930 ( .A(u2__abc_44228_n6010), .B(u2_remHi_323_), .Y(u2__abc_44228_n6011) );
  AND2X2 AND2X2_1931 ( .A(u2__abc_44228_n6013), .B(u2_o_323_), .Y(u2__abc_44228_n6014) );
  AND2X2 AND2X2_1932 ( .A(u2__abc_44228_n6012_1), .B(u2__abc_44228_n6015), .Y(u2__abc_44228_n6016) );
  AND2X2 AND2X2_1933 ( .A(u2__abc_44228_n6009), .B(u2__abc_44228_n6016), .Y(u2__abc_44228_n6017) );
  AND2X2 AND2X2_1934 ( .A(u2__abc_44228_n6003_1), .B(u2__abc_44228_n6017), .Y(u2__abc_44228_n6018) );
  AND2X2 AND2X2_1935 ( .A(u2__abc_44228_n6019), .B(u2_remHi_321_), .Y(u2__abc_44228_n6020) );
  AND2X2 AND2X2_1936 ( .A(u2__abc_44228_n6022_1), .B(u2_o_321_), .Y(u2__abc_44228_n6023) );
  AND2X2 AND2X2_1937 ( .A(u2__abc_44228_n6021), .B(u2__abc_44228_n6024), .Y(u2__abc_44228_n6025) );
  AND2X2 AND2X2_1938 ( .A(u2__abc_44228_n6026), .B(u2_remHi_320_), .Y(u2__abc_44228_n6027) );
  AND2X2 AND2X2_1939 ( .A(u2__abc_44228_n6028), .B(u2_o_320_), .Y(u2__abc_44228_n6029) );
  AND2X2 AND2X2_194 ( .A(_abc_64468_n1180), .B(_abc_64468_n1179), .Y(fracta1_4_) );
  AND2X2 AND2X2_1940 ( .A(u2__abc_44228_n6031_1), .B(u2__abc_44228_n6025), .Y(u2__abc_44228_n6032) );
  AND2X2 AND2X2_1941 ( .A(u2__abc_44228_n6033), .B(u2_remHi_318_), .Y(u2__abc_44228_n6034) );
  AND2X2 AND2X2_1942 ( .A(u2__abc_44228_n6035), .B(u2_o_318_), .Y(u2__abc_44228_n6036) );
  AND2X2 AND2X2_1943 ( .A(u2__abc_44228_n6039), .B(u2_remHi_319_), .Y(u2__abc_44228_n6040_1) );
  AND2X2 AND2X2_1944 ( .A(u2__abc_44228_n6042), .B(u2_o_319_), .Y(u2__abc_44228_n6043) );
  AND2X2 AND2X2_1945 ( .A(u2__abc_44228_n6041), .B(u2__abc_44228_n6044), .Y(u2__abc_44228_n6045) );
  AND2X2 AND2X2_1946 ( .A(u2__abc_44228_n6038), .B(u2__abc_44228_n6045), .Y(u2__abc_44228_n6046) );
  AND2X2 AND2X2_1947 ( .A(u2__abc_44228_n6032), .B(u2__abc_44228_n6046), .Y(u2__abc_44228_n6047) );
  AND2X2 AND2X2_1948 ( .A(u2__abc_44228_n6018), .B(u2__abc_44228_n6047), .Y(u2__abc_44228_n6048) );
  AND2X2 AND2X2_1949 ( .A(u2__abc_44228_n5989), .B(u2__abc_44228_n6048), .Y(u2__abc_44228_n6049_1) );
  AND2X2 AND2X2_195 ( .A(_abc_64468_n1183), .B(_abc_64468_n1182), .Y(fracta1_5_) );
  AND2X2 AND2X2_1950 ( .A(u2__abc_44228_n5930_1), .B(u2__abc_44228_n6049_1), .Y(u2__abc_44228_n6050) );
  AND2X2 AND2X2_1951 ( .A(u2__abc_44228_n5811), .B(u2__abc_44228_n6050), .Y(u2__abc_44228_n6051) );
  AND2X2 AND2X2_1952 ( .A(u2__abc_44228_n6052), .B(u2_remHi_317_), .Y(u2__abc_44228_n6053) );
  AND2X2 AND2X2_1953 ( .A(u2__abc_44228_n6055), .B(u2_o_317_), .Y(u2__abc_44228_n6056) );
  AND2X2 AND2X2_1954 ( .A(u2__abc_44228_n6054), .B(u2__abc_44228_n6057), .Y(u2__abc_44228_n6058) );
  AND2X2 AND2X2_1955 ( .A(u2__abc_44228_n6059_1), .B(u2_remHi_316_), .Y(u2__abc_44228_n6060) );
  AND2X2 AND2X2_1956 ( .A(u2__abc_44228_n6061), .B(u2_o_316_), .Y(u2__abc_44228_n6062) );
  AND2X2 AND2X2_1957 ( .A(u2__abc_44228_n6064), .B(u2__abc_44228_n6058), .Y(u2__abc_44228_n6065) );
  AND2X2 AND2X2_1958 ( .A(u2__abc_44228_n6066), .B(u2_remHi_315_), .Y(u2__abc_44228_n6067) );
  AND2X2 AND2X2_1959 ( .A(u2__abc_44228_n6069), .B(u2_o_315_), .Y(u2__abc_44228_n6070) );
  AND2X2 AND2X2_196 ( .A(_abc_64468_n1186), .B(_abc_64468_n1185), .Y(fracta1_6_) );
  AND2X2 AND2X2_1960 ( .A(u2__abc_44228_n6068_1), .B(u2__abc_44228_n6071), .Y(u2__abc_44228_n6072) );
  AND2X2 AND2X2_1961 ( .A(u2__abc_44228_n6073), .B(u2_remHi_314_), .Y(u2__abc_44228_n6074) );
  AND2X2 AND2X2_1962 ( .A(u2__abc_44228_n6075), .B(u2_o_314_), .Y(u2__abc_44228_n6076) );
  AND2X2 AND2X2_1963 ( .A(u2__abc_44228_n6078_1), .B(u2__abc_44228_n6072), .Y(u2__abc_44228_n6079) );
  AND2X2 AND2X2_1964 ( .A(u2__abc_44228_n6065), .B(u2__abc_44228_n6079), .Y(u2__abc_44228_n6080) );
  AND2X2 AND2X2_1965 ( .A(u2__abc_44228_n6081), .B(u2_remHi_313_), .Y(u2__abc_44228_n6082) );
  AND2X2 AND2X2_1966 ( .A(u2__abc_44228_n6084), .B(u2_o_313_), .Y(u2__abc_44228_n6085) );
  AND2X2 AND2X2_1967 ( .A(u2__abc_44228_n6083), .B(u2__abc_44228_n6086_1), .Y(u2__abc_44228_n6087) );
  AND2X2 AND2X2_1968 ( .A(u2__abc_44228_n6088), .B(u2_remHi_312_), .Y(u2__abc_44228_n6089) );
  AND2X2 AND2X2_1969 ( .A(u2__abc_44228_n6090), .B(u2_o_312_), .Y(u2__abc_44228_n6091) );
  AND2X2 AND2X2_197 ( .A(_abc_64468_n1189), .B(_abc_64468_n1188), .Y(fracta1_7_) );
  AND2X2 AND2X2_1970 ( .A(u2__abc_44228_n6093), .B(u2__abc_44228_n6087), .Y(u2__abc_44228_n6094) );
  AND2X2 AND2X2_1971 ( .A(u2__abc_44228_n6095), .B(u2_remHi_311_), .Y(u2__abc_44228_n6096_1) );
  AND2X2 AND2X2_1972 ( .A(u2__abc_44228_n6098), .B(u2_o_311_), .Y(u2__abc_44228_n6099) );
  AND2X2 AND2X2_1973 ( .A(u2__abc_44228_n6097), .B(u2__abc_44228_n6100), .Y(u2__abc_44228_n6101) );
  AND2X2 AND2X2_1974 ( .A(u2__abc_44228_n6102), .B(u2_remHi_310_), .Y(u2__abc_44228_n6103) );
  AND2X2 AND2X2_1975 ( .A(u2__abc_44228_n6104_1), .B(u2_o_310_), .Y(u2__abc_44228_n6105) );
  AND2X2 AND2X2_1976 ( .A(u2__abc_44228_n6107), .B(u2__abc_44228_n6101), .Y(u2__abc_44228_n6108) );
  AND2X2 AND2X2_1977 ( .A(u2__abc_44228_n6094), .B(u2__abc_44228_n6108), .Y(u2__abc_44228_n6109) );
  AND2X2 AND2X2_1978 ( .A(u2__abc_44228_n6080), .B(u2__abc_44228_n6109), .Y(u2__abc_44228_n6110) );
  AND2X2 AND2X2_1979 ( .A(u2__abc_44228_n6111), .B(u2_remHi_309_), .Y(u2__abc_44228_n6112) );
  AND2X2 AND2X2_198 ( .A(_abc_64468_n1192), .B(_abc_64468_n1191), .Y(fracta1_8_) );
  AND2X2 AND2X2_1980 ( .A(u2__abc_44228_n6114), .B(u2_o_309_), .Y(u2__abc_44228_n6115) );
  AND2X2 AND2X2_1981 ( .A(u2__abc_44228_n6113_1), .B(u2__abc_44228_n6116), .Y(u2__abc_44228_n6117) );
  AND2X2 AND2X2_1982 ( .A(u2__abc_44228_n6118), .B(u2_remHi_308_), .Y(u2__abc_44228_n6119) );
  AND2X2 AND2X2_1983 ( .A(u2__abc_44228_n6120), .B(u2_o_308_), .Y(u2__abc_44228_n6121) );
  AND2X2 AND2X2_1984 ( .A(u2__abc_44228_n6123), .B(u2__abc_44228_n6117), .Y(u2__abc_44228_n6124) );
  AND2X2 AND2X2_1985 ( .A(u2__abc_44228_n6125), .B(u2_remHi_306_), .Y(u2__abc_44228_n6126) );
  AND2X2 AND2X2_1986 ( .A(u2__abc_44228_n6127), .B(u2_o_306_), .Y(u2__abc_44228_n6128) );
  AND2X2 AND2X2_1987 ( .A(u2__abc_44228_n6131), .B(u2_remHi_307_), .Y(u2__abc_44228_n6132_1) );
  AND2X2 AND2X2_1988 ( .A(u2__abc_44228_n6134), .B(u2_o_307_), .Y(u2__abc_44228_n6135) );
  AND2X2 AND2X2_1989 ( .A(u2__abc_44228_n6133), .B(u2__abc_44228_n6136), .Y(u2__abc_44228_n6137) );
  AND2X2 AND2X2_199 ( .A(_abc_64468_n1195), .B(_abc_64468_n1194), .Y(fracta1_9_) );
  AND2X2 AND2X2_1990 ( .A(u2__abc_44228_n6130), .B(u2__abc_44228_n6137), .Y(u2__abc_44228_n6138) );
  AND2X2 AND2X2_1991 ( .A(u2__abc_44228_n6124), .B(u2__abc_44228_n6138), .Y(u2__abc_44228_n6139) );
  AND2X2 AND2X2_1992 ( .A(u2__abc_44228_n6140), .B(u2_remHi_305_), .Y(u2__abc_44228_n6141_1) );
  AND2X2 AND2X2_1993 ( .A(u2__abc_44228_n6143), .B(u2_o_305_), .Y(u2__abc_44228_n6144) );
  AND2X2 AND2X2_1994 ( .A(u2__abc_44228_n6142), .B(u2__abc_44228_n6145), .Y(u2__abc_44228_n6146) );
  AND2X2 AND2X2_1995 ( .A(u2__abc_44228_n6147), .B(u2_remHi_304_), .Y(u2__abc_44228_n6148) );
  AND2X2 AND2X2_1996 ( .A(u2__abc_44228_n6149), .B(u2_o_304_), .Y(u2__abc_44228_n6150) );
  AND2X2 AND2X2_1997 ( .A(u2__abc_44228_n6152), .B(u2__abc_44228_n6146), .Y(u2__abc_44228_n6153) );
  AND2X2 AND2X2_1998 ( .A(u2__abc_44228_n6154), .B(u2_remHi_302_), .Y(u2__abc_44228_n6155) );
  AND2X2 AND2X2_1999 ( .A(u2__abc_44228_n6156), .B(u2_o_302_), .Y(u2__abc_44228_n6157) );
  AND2X2 AND2X2_2 ( .A(_abc_64468_n753_bF_buf12), .B(sqrto_1_), .Y(_auto_iopadmap_cc_313_execute_65414_37_) );
  AND2X2 AND2X2_20 ( .A(_abc_64468_n753_bF_buf8), .B(sqrto_19_), .Y(_auto_iopadmap_cc_313_execute_65414_55_) );
  AND2X2 AND2X2_200 ( .A(_abc_64468_n1198), .B(_abc_64468_n1197), .Y(fracta1_10_) );
  AND2X2 AND2X2_2000 ( .A(u2__abc_44228_n6160), .B(u2_remHi_303_), .Y(u2__abc_44228_n6161) );
  AND2X2 AND2X2_2001 ( .A(u2__abc_44228_n6163), .B(u2_o_303_), .Y(u2__abc_44228_n6164) );
  AND2X2 AND2X2_2002 ( .A(u2__abc_44228_n6162), .B(u2__abc_44228_n6165), .Y(u2__abc_44228_n6166) );
  AND2X2 AND2X2_2003 ( .A(u2__abc_44228_n6159_1), .B(u2__abc_44228_n6166), .Y(u2__abc_44228_n6167) );
  AND2X2 AND2X2_2004 ( .A(u2__abc_44228_n6153), .B(u2__abc_44228_n6167), .Y(u2__abc_44228_n6168) );
  AND2X2 AND2X2_2005 ( .A(u2__abc_44228_n6139), .B(u2__abc_44228_n6168), .Y(u2__abc_44228_n6169_1) );
  AND2X2 AND2X2_2006 ( .A(u2__abc_44228_n6110), .B(u2__abc_44228_n6169_1), .Y(u2__abc_44228_n6170) );
  AND2X2 AND2X2_2007 ( .A(u2__abc_44228_n6171), .B(u2_remHi_301_), .Y(u2__abc_44228_n6172) );
  AND2X2 AND2X2_2008 ( .A(u2__abc_44228_n6174), .B(u2_o_301_), .Y(u2__abc_44228_n6175) );
  AND2X2 AND2X2_2009 ( .A(u2__abc_44228_n6173), .B(u2__abc_44228_n6176), .Y(u2__abc_44228_n6177) );
  AND2X2 AND2X2_201 ( .A(_abc_64468_n1201), .B(_abc_64468_n1200), .Y(fracta1_11_) );
  AND2X2 AND2X2_2010 ( .A(u2__abc_44228_n6178_1), .B(u2_remHi_300_), .Y(u2__abc_44228_n6179) );
  AND2X2 AND2X2_2011 ( .A(u2__abc_44228_n6180), .B(u2_o_300_), .Y(u2__abc_44228_n6181) );
  AND2X2 AND2X2_2012 ( .A(u2__abc_44228_n6183), .B(u2__abc_44228_n6177), .Y(u2__abc_44228_n6184) );
  AND2X2 AND2X2_2013 ( .A(u2__abc_44228_n6185), .B(u2_remHi_299_), .Y(u2__abc_44228_n6186) );
  AND2X2 AND2X2_2014 ( .A(u2__abc_44228_n6188), .B(u2_o_299_), .Y(u2__abc_44228_n6189) );
  AND2X2 AND2X2_2015 ( .A(u2__abc_44228_n6187_1), .B(u2__abc_44228_n6190), .Y(u2__abc_44228_n6191) );
  AND2X2 AND2X2_2016 ( .A(u2__abc_44228_n6192), .B(u2_remHi_298_), .Y(u2__abc_44228_n6193) );
  AND2X2 AND2X2_2017 ( .A(u2__abc_44228_n6194), .B(u2_o_298_), .Y(u2__abc_44228_n6195) );
  AND2X2 AND2X2_2018 ( .A(u2__abc_44228_n6197), .B(u2__abc_44228_n6191), .Y(u2__abc_44228_n6198) );
  AND2X2 AND2X2_2019 ( .A(u2__abc_44228_n6184), .B(u2__abc_44228_n6198), .Y(u2__abc_44228_n6199) );
  AND2X2 AND2X2_202 ( .A(_abc_64468_n1204), .B(_abc_64468_n1203), .Y(fracta1_12_) );
  AND2X2 AND2X2_2020 ( .A(u2__abc_44228_n6200), .B(u2_remHi_295_), .Y(u2__abc_44228_n6201) );
  AND2X2 AND2X2_2021 ( .A(u2__abc_44228_n6203), .B(u2_o_295_), .Y(u2__abc_44228_n6204) );
  AND2X2 AND2X2_2022 ( .A(u2__abc_44228_n6202), .B(u2__abc_44228_n6205), .Y(u2__abc_44228_n6206_1) );
  AND2X2 AND2X2_2023 ( .A(u2__abc_44228_n6207), .B(u2_remHi_294_), .Y(u2__abc_44228_n6208) );
  AND2X2 AND2X2_2024 ( .A(u2__abc_44228_n6209), .B(u2_o_294_), .Y(u2__abc_44228_n6210) );
  AND2X2 AND2X2_2025 ( .A(u2__abc_44228_n6212), .B(u2__abc_44228_n6206_1), .Y(u2__abc_44228_n6213) );
  AND2X2 AND2X2_2026 ( .A(u2__abc_44228_n6214_1), .B(u2_remHi_297_), .Y(u2__abc_44228_n6215) );
  AND2X2 AND2X2_2027 ( .A(u2__abc_44228_n6217), .B(u2_o_297_), .Y(u2__abc_44228_n6218) );
  AND2X2 AND2X2_2028 ( .A(u2__abc_44228_n6216), .B(u2__abc_44228_n6219), .Y(u2__abc_44228_n6220) );
  AND2X2 AND2X2_2029 ( .A(u2__abc_44228_n6221), .B(u2_remHi_296_), .Y(u2__abc_44228_n6222) );
  AND2X2 AND2X2_203 ( .A(_abc_64468_n1207), .B(_abc_64468_n1206), .Y(fracta1_13_) );
  AND2X2 AND2X2_2030 ( .A(u2__abc_44228_n6223), .B(u2_o_296_), .Y(u2__abc_44228_n6224_1) );
  AND2X2 AND2X2_2031 ( .A(u2__abc_44228_n6226), .B(u2__abc_44228_n6220), .Y(u2__abc_44228_n6227) );
  AND2X2 AND2X2_2032 ( .A(u2__abc_44228_n6213), .B(u2__abc_44228_n6227), .Y(u2__abc_44228_n6228) );
  AND2X2 AND2X2_2033 ( .A(u2__abc_44228_n6199), .B(u2__abc_44228_n6228), .Y(u2__abc_44228_n6229) );
  AND2X2 AND2X2_2034 ( .A(u2__abc_44228_n6230), .B(u2_remHi_293_), .Y(u2__abc_44228_n6231) );
  AND2X2 AND2X2_2035 ( .A(u2__abc_44228_n6233), .B(u2_o_293_), .Y(u2__abc_44228_n6234) );
  AND2X2 AND2X2_2036 ( .A(u2__abc_44228_n6232_1), .B(u2__abc_44228_n6235), .Y(u2__abc_44228_n6236) );
  AND2X2 AND2X2_2037 ( .A(u2__abc_44228_n6237), .B(u2_remHi_292_), .Y(u2__abc_44228_n6238) );
  AND2X2 AND2X2_2038 ( .A(u2__abc_44228_n6239), .B(u2_o_292_), .Y(u2__abc_44228_n6240) );
  AND2X2 AND2X2_2039 ( .A(u2__abc_44228_n6242_1), .B(u2__abc_44228_n6236), .Y(u2__abc_44228_n6243) );
  AND2X2 AND2X2_204 ( .A(_abc_64468_n1210), .B(_abc_64468_n1209), .Y(fracta1_14_) );
  AND2X2 AND2X2_2040 ( .A(u2__abc_44228_n6244), .B(u2_remHi_291_), .Y(u2__abc_44228_n6245) );
  AND2X2 AND2X2_2041 ( .A(u2__abc_44228_n6247), .B(u2_o_291_), .Y(u2__abc_44228_n6248) );
  AND2X2 AND2X2_2042 ( .A(u2__abc_44228_n6246), .B(u2__abc_44228_n6249), .Y(u2__abc_44228_n6250) );
  AND2X2 AND2X2_2043 ( .A(u2__abc_44228_n6251_1), .B(u2_remHi_290_), .Y(u2__abc_44228_n6252) );
  AND2X2 AND2X2_2044 ( .A(u2__abc_44228_n6253), .B(u2_o_290_), .Y(u2__abc_44228_n6254) );
  AND2X2 AND2X2_2045 ( .A(u2__abc_44228_n6256), .B(u2__abc_44228_n6250), .Y(u2__abc_44228_n6257) );
  AND2X2 AND2X2_2046 ( .A(u2__abc_44228_n6243), .B(u2__abc_44228_n6257), .Y(u2__abc_44228_n6258) );
  AND2X2 AND2X2_2047 ( .A(u2__abc_44228_n6259), .B(u2_remHi_289_), .Y(u2__abc_44228_n6260_1) );
  AND2X2 AND2X2_2048 ( .A(u2__abc_44228_n6262), .B(u2_o_289_), .Y(u2__abc_44228_n6263) );
  AND2X2 AND2X2_2049 ( .A(u2__abc_44228_n6261), .B(u2__abc_44228_n6264), .Y(u2__abc_44228_n6265) );
  AND2X2 AND2X2_205 ( .A(_abc_64468_n1213), .B(_abc_64468_n1212), .Y(fracta1_15_) );
  AND2X2 AND2X2_2050 ( .A(u2__abc_44228_n6266), .B(u2_remHi_288_), .Y(u2__abc_44228_n6267) );
  AND2X2 AND2X2_2051 ( .A(u2__abc_44228_n6268), .B(u2_o_288_), .Y(u2__abc_44228_n6269_1) );
  AND2X2 AND2X2_2052 ( .A(u2__abc_44228_n6271), .B(u2__abc_44228_n6265), .Y(u2__abc_44228_n6272) );
  AND2X2 AND2X2_2053 ( .A(u2__abc_44228_n6273), .B(u2_remHi_287_), .Y(u2__abc_44228_n6274) );
  AND2X2 AND2X2_2054 ( .A(u2__abc_44228_n6276), .B(u2_o_287_), .Y(u2__abc_44228_n6277) );
  AND2X2 AND2X2_2055 ( .A(u2__abc_44228_n6275), .B(u2__abc_44228_n6278), .Y(u2__abc_44228_n6279_1) );
  AND2X2 AND2X2_2056 ( .A(u2__abc_44228_n6280), .B(u2_remHi_286_), .Y(u2__abc_44228_n6281) );
  AND2X2 AND2X2_2057 ( .A(u2__abc_44228_n6282), .B(u2_o_286_), .Y(u2__abc_44228_n6283) );
  AND2X2 AND2X2_2058 ( .A(u2__abc_44228_n6285), .B(u2__abc_44228_n6279_1), .Y(u2__abc_44228_n6286) );
  AND2X2 AND2X2_2059 ( .A(u2__abc_44228_n6272), .B(u2__abc_44228_n6286), .Y(u2__abc_44228_n6287_1) );
  AND2X2 AND2X2_206 ( .A(_abc_64468_n1216), .B(_abc_64468_n1215), .Y(fracta1_16_) );
  AND2X2 AND2X2_2060 ( .A(u2__abc_44228_n6258), .B(u2__abc_44228_n6287_1), .Y(u2__abc_44228_n6288) );
  AND2X2 AND2X2_2061 ( .A(u2__abc_44228_n6229), .B(u2__abc_44228_n6288), .Y(u2__abc_44228_n6289) );
  AND2X2 AND2X2_2062 ( .A(u2__abc_44228_n6170), .B(u2__abc_44228_n6289), .Y(u2__abc_44228_n6290) );
  AND2X2 AND2X2_2063 ( .A(u2__abc_44228_n6291), .B(u2_remHi_285_), .Y(u2__abc_44228_n6292) );
  AND2X2 AND2X2_2064 ( .A(u2__abc_44228_n6294), .B(u2_o_285_), .Y(u2__abc_44228_n6295) );
  AND2X2 AND2X2_2065 ( .A(u2__abc_44228_n6293), .B(u2__abc_44228_n6296_1), .Y(u2__abc_44228_n6297) );
  AND2X2 AND2X2_2066 ( .A(u2__abc_44228_n6298), .B(u2_remHi_284_), .Y(u2__abc_44228_n6299) );
  AND2X2 AND2X2_2067 ( .A(u2__abc_44228_n6300), .B(u2_o_284_), .Y(u2__abc_44228_n6301) );
  AND2X2 AND2X2_2068 ( .A(u2__abc_44228_n6303), .B(u2__abc_44228_n6297), .Y(u2__abc_44228_n6304) );
  AND2X2 AND2X2_2069 ( .A(u2__abc_44228_n6305_1), .B(u2_remHi_283_), .Y(u2__abc_44228_n6306) );
  AND2X2 AND2X2_207 ( .A(_abc_64468_n1219), .B(_abc_64468_n1218), .Y(fracta1_17_) );
  AND2X2 AND2X2_2070 ( .A(u2__abc_44228_n6308), .B(u2_o_283_), .Y(u2__abc_44228_n6309) );
  AND2X2 AND2X2_2071 ( .A(u2__abc_44228_n6307), .B(u2__abc_44228_n6310), .Y(u2__abc_44228_n6311) );
  AND2X2 AND2X2_2072 ( .A(u2__abc_44228_n6312), .B(u2_remHi_282_), .Y(u2__abc_44228_n6313) );
  AND2X2 AND2X2_2073 ( .A(u2__abc_44228_n6314), .B(u2_o_282_), .Y(u2__abc_44228_n6315_1) );
  AND2X2 AND2X2_2074 ( .A(u2__abc_44228_n6317), .B(u2__abc_44228_n6311), .Y(u2__abc_44228_n6318) );
  AND2X2 AND2X2_2075 ( .A(u2__abc_44228_n6304), .B(u2__abc_44228_n6318), .Y(u2__abc_44228_n6319) );
  AND2X2 AND2X2_2076 ( .A(u2__abc_44228_n6320), .B(u2_remHi_279_), .Y(u2__abc_44228_n6321) );
  AND2X2 AND2X2_2077 ( .A(u2__abc_44228_n6323), .B(u2_o_279_), .Y(u2__abc_44228_n6324_1) );
  AND2X2 AND2X2_2078 ( .A(u2__abc_44228_n6322), .B(u2__abc_44228_n6325), .Y(u2__abc_44228_n6326) );
  AND2X2 AND2X2_2079 ( .A(u2__abc_44228_n6327), .B(u2_remHi_278_), .Y(u2__abc_44228_n6328) );
  AND2X2 AND2X2_208 ( .A(_abc_64468_n1222), .B(_abc_64468_n1221), .Y(fracta1_18_) );
  AND2X2 AND2X2_2080 ( .A(u2__abc_44228_n6329), .B(u2_o_278_), .Y(u2__abc_44228_n6330) );
  AND2X2 AND2X2_2081 ( .A(u2__abc_44228_n6332), .B(u2__abc_44228_n6326), .Y(u2__abc_44228_n6333_1) );
  AND2X2 AND2X2_2082 ( .A(u2__abc_44228_n6334), .B(u2_remHi_281_), .Y(u2__abc_44228_n6335) );
  AND2X2 AND2X2_2083 ( .A(u2__abc_44228_n6337), .B(u2_o_281_), .Y(u2__abc_44228_n6338) );
  AND2X2 AND2X2_2084 ( .A(u2__abc_44228_n6336), .B(u2__abc_44228_n6339), .Y(u2__abc_44228_n6340) );
  AND2X2 AND2X2_2085 ( .A(u2__abc_44228_n6341), .B(u2_remHi_280_), .Y(u2__abc_44228_n6342_1) );
  AND2X2 AND2X2_2086 ( .A(u2__abc_44228_n6343), .B(u2_o_280_), .Y(u2__abc_44228_n6344) );
  AND2X2 AND2X2_2087 ( .A(u2__abc_44228_n6346), .B(u2__abc_44228_n6340), .Y(u2__abc_44228_n6347) );
  AND2X2 AND2X2_2088 ( .A(u2__abc_44228_n6333_1), .B(u2__abc_44228_n6347), .Y(u2__abc_44228_n6348) );
  AND2X2 AND2X2_2089 ( .A(u2__abc_44228_n6319), .B(u2__abc_44228_n6348), .Y(u2__abc_44228_n6349) );
  AND2X2 AND2X2_209 ( .A(_abc_64468_n1225), .B(_abc_64468_n1224), .Y(fracta1_19_) );
  AND2X2 AND2X2_2090 ( .A(u2__abc_44228_n6350), .B(u2_remHi_277_), .Y(u2__abc_44228_n6351) );
  AND2X2 AND2X2_2091 ( .A(u2__abc_44228_n6353), .B(u2_o_277_), .Y(u2__abc_44228_n6354) );
  AND2X2 AND2X2_2092 ( .A(u2__abc_44228_n6352_1), .B(u2__abc_44228_n6355), .Y(u2__abc_44228_n6356) );
  AND2X2 AND2X2_2093 ( .A(u2__abc_44228_n6357), .B(u2_remHi_276_), .Y(u2__abc_44228_n6358) );
  AND2X2 AND2X2_2094 ( .A(u2__abc_44228_n6359), .B(u2_o_276_), .Y(u2__abc_44228_n6360) );
  AND2X2 AND2X2_2095 ( .A(u2__abc_44228_n6362), .B(u2__abc_44228_n6356), .Y(u2__abc_44228_n6363) );
  AND2X2 AND2X2_2096 ( .A(u2__abc_44228_n6364), .B(u2_remHi_275_), .Y(u2__abc_44228_n6365) );
  AND2X2 AND2X2_2097 ( .A(u2__abc_44228_n6367), .B(u2_o_275_), .Y(u2__abc_44228_n6368) );
  AND2X2 AND2X2_2098 ( .A(u2__abc_44228_n6366), .B(u2__abc_44228_n6369), .Y(u2__abc_44228_n6370) );
  AND2X2 AND2X2_2099 ( .A(u2__abc_44228_n6371_1), .B(u2_remHi_274_), .Y(u2__abc_44228_n6372) );
  AND2X2 AND2X2_21 ( .A(_abc_64468_n753_bF_buf7), .B(sqrto_20_), .Y(_auto_iopadmap_cc_313_execute_65414_56_) );
  AND2X2 AND2X2_210 ( .A(_abc_64468_n1228), .B(_abc_64468_n1227), .Y(fracta1_20_) );
  AND2X2 AND2X2_2100 ( .A(u2__abc_44228_n6373), .B(u2_o_274_), .Y(u2__abc_44228_n6374) );
  AND2X2 AND2X2_2101 ( .A(u2__abc_44228_n6376), .B(u2__abc_44228_n6370), .Y(u2__abc_44228_n6377) );
  AND2X2 AND2X2_2102 ( .A(u2__abc_44228_n6363), .B(u2__abc_44228_n6377), .Y(u2__abc_44228_n6378) );
  AND2X2 AND2X2_2103 ( .A(u2__abc_44228_n6379_1), .B(u2_remHi_273_), .Y(u2__abc_44228_n6380) );
  AND2X2 AND2X2_2104 ( .A(u2__abc_44228_n6382), .B(u2_o_273_), .Y(u2__abc_44228_n6383) );
  AND2X2 AND2X2_2105 ( .A(u2__abc_44228_n6381), .B(u2__abc_44228_n6384), .Y(u2__abc_44228_n6385) );
  AND2X2 AND2X2_2106 ( .A(u2__abc_44228_n6386), .B(u2_remHi_272_), .Y(u2__abc_44228_n6387) );
  AND2X2 AND2X2_2107 ( .A(u2__abc_44228_n6388), .B(u2_o_272_), .Y(u2__abc_44228_n6389_1) );
  AND2X2 AND2X2_2108 ( .A(u2__abc_44228_n6391), .B(u2__abc_44228_n6385), .Y(u2__abc_44228_n6392) );
  AND2X2 AND2X2_2109 ( .A(u2__abc_44228_n6393), .B(u2_remHi_270_), .Y(u2__abc_44228_n6394) );
  AND2X2 AND2X2_211 ( .A(_abc_64468_n1231), .B(_abc_64468_n1230), .Y(fracta1_21_) );
  AND2X2 AND2X2_2110 ( .A(u2__abc_44228_n6395), .B(u2_o_270_), .Y(u2__abc_44228_n6396) );
  AND2X2 AND2X2_2111 ( .A(u2__abc_44228_n6399), .B(u2_remHi_271_), .Y(u2__abc_44228_n6400) );
  AND2X2 AND2X2_2112 ( .A(u2__abc_44228_n6402), .B(u2_o_271_), .Y(u2__abc_44228_n6403) );
  AND2X2 AND2X2_2113 ( .A(u2__abc_44228_n6401), .B(u2__abc_44228_n6404), .Y(u2__abc_44228_n6405) );
  AND2X2 AND2X2_2114 ( .A(u2__abc_44228_n6398), .B(u2__abc_44228_n6405), .Y(u2__abc_44228_n6406_1) );
  AND2X2 AND2X2_2115 ( .A(u2__abc_44228_n6392), .B(u2__abc_44228_n6406_1), .Y(u2__abc_44228_n6407) );
  AND2X2 AND2X2_2116 ( .A(u2__abc_44228_n6378), .B(u2__abc_44228_n6407), .Y(u2__abc_44228_n6408) );
  AND2X2 AND2X2_2117 ( .A(u2__abc_44228_n6349), .B(u2__abc_44228_n6408), .Y(u2__abc_44228_n6409) );
  AND2X2 AND2X2_2118 ( .A(u2__abc_44228_n6410), .B(u2_remHi_269_), .Y(u2__abc_44228_n6411) );
  AND2X2 AND2X2_2119 ( .A(u2__abc_44228_n6413), .B(u2_o_269_), .Y(u2__abc_44228_n6414) );
  AND2X2 AND2X2_212 ( .A(_abc_64468_n1234), .B(_abc_64468_n1233), .Y(fracta1_22_) );
  AND2X2 AND2X2_2120 ( .A(u2__abc_44228_n6412), .B(u2__abc_44228_n6415_1), .Y(u2__abc_44228_n6416) );
  AND2X2 AND2X2_2121 ( .A(u2__abc_44228_n6417), .B(u2_remHi_268_), .Y(u2__abc_44228_n6418) );
  AND2X2 AND2X2_2122 ( .A(u2__abc_44228_n6419), .B(u2_o_268_), .Y(u2__abc_44228_n6420) );
  AND2X2 AND2X2_2123 ( .A(u2__abc_44228_n6422), .B(u2__abc_44228_n6416), .Y(u2__abc_44228_n6423) );
  AND2X2 AND2X2_2124 ( .A(u2__abc_44228_n6424), .B(u2_remHi_267_), .Y(u2__abc_44228_n6425_1) );
  AND2X2 AND2X2_2125 ( .A(u2__abc_44228_n6427), .B(u2_o_267_), .Y(u2__abc_44228_n6428) );
  AND2X2 AND2X2_2126 ( .A(u2__abc_44228_n6426), .B(u2__abc_44228_n6429), .Y(u2__abc_44228_n6430) );
  AND2X2 AND2X2_2127 ( .A(u2__abc_44228_n6431), .B(u2_remHi_266_), .Y(u2__abc_44228_n6432) );
  AND2X2 AND2X2_2128 ( .A(u2__abc_44228_n6433), .B(u2_o_266_), .Y(u2__abc_44228_n6434) );
  AND2X2 AND2X2_2129 ( .A(u2__abc_44228_n6436), .B(u2__abc_44228_n6430), .Y(u2__abc_44228_n6437) );
  AND2X2 AND2X2_213 ( .A(_abc_64468_n1237), .B(_abc_64468_n1236), .Y(fracta1_23_) );
  AND2X2 AND2X2_2130 ( .A(u2__abc_44228_n6423), .B(u2__abc_44228_n6437), .Y(u2__abc_44228_n6438) );
  AND2X2 AND2X2_2131 ( .A(u2__abc_44228_n6439), .B(u2_remHi_265_), .Y(u2__abc_44228_n6440) );
  AND2X2 AND2X2_2132 ( .A(u2__abc_44228_n6442), .B(u2_o_265_), .Y(u2__abc_44228_n6443) );
  AND2X2 AND2X2_2133 ( .A(u2__abc_44228_n6441), .B(u2__abc_44228_n6444), .Y(u2__abc_44228_n6445_1) );
  AND2X2 AND2X2_2134 ( .A(u2__abc_44228_n6446), .B(u2_remHi_264_), .Y(u2__abc_44228_n6447) );
  AND2X2 AND2X2_2135 ( .A(u2__abc_44228_n6448), .B(u2_o_264_), .Y(u2__abc_44228_n6449) );
  AND2X2 AND2X2_2136 ( .A(u2__abc_44228_n6451), .B(u2__abc_44228_n6445_1), .Y(u2__abc_44228_n6452) );
  AND2X2 AND2X2_2137 ( .A(u2__abc_44228_n6453_1), .B(u2_remHi_263_), .Y(u2__abc_44228_n6454) );
  AND2X2 AND2X2_2138 ( .A(u2__abc_44228_n6456), .B(u2_o_263_), .Y(u2__abc_44228_n6457) );
  AND2X2 AND2X2_2139 ( .A(u2__abc_44228_n6455), .B(u2__abc_44228_n6458), .Y(u2__abc_44228_n6459) );
  AND2X2 AND2X2_214 ( .A(_abc_64468_n1240), .B(_abc_64468_n1239), .Y(fracta1_24_) );
  AND2X2 AND2X2_2140 ( .A(u2__abc_44228_n6460), .B(u2_remHi_262_), .Y(u2__abc_44228_n6461) );
  AND2X2 AND2X2_2141 ( .A(u2__abc_44228_n6462), .B(u2_o_262_), .Y(u2__abc_44228_n6463_1) );
  AND2X2 AND2X2_2142 ( .A(u2__abc_44228_n6465), .B(u2__abc_44228_n6459), .Y(u2__abc_44228_n6466) );
  AND2X2 AND2X2_2143 ( .A(u2__abc_44228_n6452), .B(u2__abc_44228_n6466), .Y(u2__abc_44228_n6467) );
  AND2X2 AND2X2_2144 ( .A(u2__abc_44228_n6438), .B(u2__abc_44228_n6467), .Y(u2__abc_44228_n6468) );
  AND2X2 AND2X2_2145 ( .A(u2__abc_44228_n6469), .B(u2_remHi_261_), .Y(u2__abc_44228_n6470) );
  AND2X2 AND2X2_2146 ( .A(u2__abc_44228_n6472), .B(u2_o_261_), .Y(u2__abc_44228_n6473) );
  AND2X2 AND2X2_2147 ( .A(u2__abc_44228_n6471_1), .B(u2__abc_44228_n6474), .Y(u2__abc_44228_n6475) );
  AND2X2 AND2X2_2148 ( .A(u2__abc_44228_n6476), .B(u2_remHi_260_), .Y(u2__abc_44228_n6477) );
  AND2X2 AND2X2_2149 ( .A(u2__abc_44228_n6478), .B(u2_o_260_), .Y(u2__abc_44228_n6479) );
  AND2X2 AND2X2_215 ( .A(_abc_64468_n1243), .B(_abc_64468_n1242), .Y(fracta1_25_) );
  AND2X2 AND2X2_2150 ( .A(u2__abc_44228_n6481), .B(u2__abc_44228_n6475), .Y(u2__abc_44228_n6482) );
  AND2X2 AND2X2_2151 ( .A(u2__abc_44228_n6483), .B(u2_remHi_259_), .Y(u2__abc_44228_n6484) );
  AND2X2 AND2X2_2152 ( .A(u2__abc_44228_n6486), .B(u2_o_259_), .Y(u2__abc_44228_n6487) );
  AND2X2 AND2X2_2153 ( .A(u2__abc_44228_n6485), .B(u2__abc_44228_n6488), .Y(u2__abc_44228_n6489_1) );
  AND2X2 AND2X2_2154 ( .A(u2__abc_44228_n6490), .B(u2_remHi_258_), .Y(u2__abc_44228_n6491) );
  AND2X2 AND2X2_2155 ( .A(u2__abc_44228_n6492), .B(u2_o_258_), .Y(u2__abc_44228_n6493) );
  AND2X2 AND2X2_2156 ( .A(u2__abc_44228_n6495), .B(u2__abc_44228_n6489_1), .Y(u2__abc_44228_n6496) );
  AND2X2 AND2X2_2157 ( .A(u2__abc_44228_n6482), .B(u2__abc_44228_n6496), .Y(u2__abc_44228_n6497) );
  AND2X2 AND2X2_2158 ( .A(u2__abc_44228_n6498), .B(u2_remHi_257_), .Y(u2__abc_44228_n6499_1) );
  AND2X2 AND2X2_2159 ( .A(u2__abc_44228_n6501), .B(u2_o_257_), .Y(u2__abc_44228_n6502) );
  AND2X2 AND2X2_216 ( .A(_abc_64468_n1246), .B(_abc_64468_n1245), .Y(fracta1_26_) );
  AND2X2 AND2X2_2160 ( .A(u2__abc_44228_n6500), .B(u2__abc_44228_n6503), .Y(u2__abc_44228_n6504) );
  AND2X2 AND2X2_2161 ( .A(u2__abc_44228_n6505), .B(u2_remHi_256_), .Y(u2__abc_44228_n6506) );
  AND2X2 AND2X2_2162 ( .A(u2__abc_44228_n6507_1), .B(u2_o_256_), .Y(u2__abc_44228_n6508) );
  AND2X2 AND2X2_2163 ( .A(u2__abc_44228_n6510), .B(u2__abc_44228_n6504), .Y(u2__abc_44228_n6511) );
  AND2X2 AND2X2_2164 ( .A(u2__abc_44228_n6512), .B(u2_remHi_255_), .Y(u2__abc_44228_n6513) );
  AND2X2 AND2X2_2165 ( .A(u2__abc_44228_n6515), .B(u2_o_255_), .Y(u2__abc_44228_n6516) );
  AND2X2 AND2X2_2166 ( .A(u2__abc_44228_n6514), .B(u2__abc_44228_n6517_1), .Y(u2__abc_44228_n6518) );
  AND2X2 AND2X2_2167 ( .A(u2__abc_44228_n6519), .B(u2_remHi_254_), .Y(u2__abc_44228_n6520) );
  AND2X2 AND2X2_2168 ( .A(u2__abc_44228_n6521), .B(u2_o_254_), .Y(u2__abc_44228_n6522) );
  AND2X2 AND2X2_2169 ( .A(u2__abc_44228_n6524), .B(u2__abc_44228_n6518), .Y(u2__abc_44228_n6525_1) );
  AND2X2 AND2X2_217 ( .A(_abc_64468_n1249), .B(_abc_64468_n1248), .Y(fracta1_27_) );
  AND2X2 AND2X2_2170 ( .A(u2__abc_44228_n6511), .B(u2__abc_44228_n6525_1), .Y(u2__abc_44228_n6526) );
  AND2X2 AND2X2_2171 ( .A(u2__abc_44228_n6497), .B(u2__abc_44228_n6526), .Y(u2__abc_44228_n6527) );
  AND2X2 AND2X2_2172 ( .A(u2__abc_44228_n6468), .B(u2__abc_44228_n6527), .Y(u2__abc_44228_n6528) );
  AND2X2 AND2X2_2173 ( .A(u2__abc_44228_n6409), .B(u2__abc_44228_n6528), .Y(u2__abc_44228_n6529) );
  AND2X2 AND2X2_2174 ( .A(u2__abc_44228_n6290), .B(u2__abc_44228_n6529), .Y(u2__abc_44228_n6530) );
  AND2X2 AND2X2_2175 ( .A(u2__abc_44228_n6051), .B(u2__abc_44228_n6530), .Y(u2__abc_44228_n6531) );
  AND2X2 AND2X2_2176 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6531), .Y(u2__abc_44228_n6532) );
  AND2X2 AND2X2_2177 ( .A(u2__abc_44228_n6534), .B(u2__abc_44228_n6514), .Y(u2__abc_44228_n6535_1) );
  AND2X2 AND2X2_2178 ( .A(u2__abc_44228_n6536), .B(u2__abc_44228_n6511), .Y(u2__abc_44228_n6537) );
  AND2X2 AND2X2_2179 ( .A(u2__abc_44228_n6503), .B(u2__abc_44228_n6506), .Y(u2__abc_44228_n6538) );
  AND2X2 AND2X2_218 ( .A(_abc_64468_n1252), .B(_abc_64468_n1251), .Y(fracta1_28_) );
  AND2X2 AND2X2_2180 ( .A(u2__abc_44228_n6540), .B(u2__abc_44228_n6497), .Y(u2__abc_44228_n6541) );
  AND2X2 AND2X2_2181 ( .A(u2__abc_44228_n6543_1), .B(u2__abc_44228_n6485), .Y(u2__abc_44228_n6544) );
  AND2X2 AND2X2_2182 ( .A(u2__abc_44228_n6545), .B(u2__abc_44228_n6482), .Y(u2__abc_44228_n6546) );
  AND2X2 AND2X2_2183 ( .A(u2__abc_44228_n6474), .B(u2__abc_44228_n6477), .Y(u2__abc_44228_n6547) );
  AND2X2 AND2X2_2184 ( .A(u2__abc_44228_n6550), .B(u2__abc_44228_n6468), .Y(u2__abc_44228_n6551) );
  AND2X2 AND2X2_2185 ( .A(u2__abc_44228_n6552_1), .B(u2__abc_44228_n6444), .Y(u2__abc_44228_n6553) );
  AND2X2 AND2X2_2186 ( .A(u2__abc_44228_n6455), .B(u2__abc_44228_n6554), .Y(u2__abc_44228_n6555) );
  AND2X2 AND2X2_2187 ( .A(u2__abc_44228_n6556), .B(u2__abc_44228_n6458), .Y(u2__abc_44228_n6557) );
  AND2X2 AND2X2_2188 ( .A(u2__abc_44228_n6557), .B(u2__abc_44228_n6452), .Y(u2__abc_44228_n6558) );
  AND2X2 AND2X2_2189 ( .A(u2__abc_44228_n6559), .B(u2__abc_44228_n6438), .Y(u2__abc_44228_n6560) );
  AND2X2 AND2X2_219 ( .A(_abc_64468_n1255), .B(_abc_64468_n1254), .Y(fracta1_29_) );
  AND2X2 AND2X2_2190 ( .A(u2__abc_44228_n6562), .B(u2__abc_44228_n6426), .Y(u2__abc_44228_n6563) );
  AND2X2 AND2X2_2191 ( .A(u2__abc_44228_n6564), .B(u2__abc_44228_n6423), .Y(u2__abc_44228_n6565) );
  AND2X2 AND2X2_2192 ( .A(u2__abc_44228_n6415_1), .B(u2__abc_44228_n6418), .Y(u2__abc_44228_n6566) );
  AND2X2 AND2X2_2193 ( .A(u2__abc_44228_n6570), .B(u2__abc_44228_n6409), .Y(u2__abc_44228_n6571_1) );
  AND2X2 AND2X2_2194 ( .A(u2__abc_44228_n6572), .B(u2__abc_44228_n6401), .Y(u2__abc_44228_n6573) );
  AND2X2 AND2X2_2195 ( .A(u2__abc_44228_n6574), .B(u2__abc_44228_n6404), .Y(u2__abc_44228_n6575) );
  AND2X2 AND2X2_2196 ( .A(u2__abc_44228_n6575), .B(u2__abc_44228_n6392), .Y(u2__abc_44228_n6576) );
  AND2X2 AND2X2_2197 ( .A(u2__abc_44228_n6384), .B(u2__abc_44228_n6387), .Y(u2__abc_44228_n6577) );
  AND2X2 AND2X2_2198 ( .A(u2__abc_44228_n6579_1), .B(u2__abc_44228_n6378), .Y(u2__abc_44228_n6580) );
  AND2X2 AND2X2_2199 ( .A(u2__abc_44228_n6582), .B(u2__abc_44228_n6366), .Y(u2__abc_44228_n6583) );
  AND2X2 AND2X2_22 ( .A(_abc_64468_n753_bF_buf6), .B(sqrto_21_), .Y(_auto_iopadmap_cc_313_execute_65414_57_) );
  AND2X2 AND2X2_220 ( .A(_abc_64468_n1258), .B(_abc_64468_n1257), .Y(fracta1_30_) );
  AND2X2 AND2X2_2200 ( .A(u2__abc_44228_n6584), .B(u2__abc_44228_n6363), .Y(u2__abc_44228_n6585) );
  AND2X2 AND2X2_2201 ( .A(u2__abc_44228_n6355), .B(u2__abc_44228_n6358), .Y(u2__abc_44228_n6586) );
  AND2X2 AND2X2_2202 ( .A(u2__abc_44228_n6589), .B(u2__abc_44228_n6349), .Y(u2__abc_44228_n6590) );
  AND2X2 AND2X2_2203 ( .A(u2__abc_44228_n6592), .B(u2__abc_44228_n6322), .Y(u2__abc_44228_n6593) );
  AND2X2 AND2X2_2204 ( .A(u2__abc_44228_n6594), .B(u2__abc_44228_n6347), .Y(u2__abc_44228_n6595) );
  AND2X2 AND2X2_2205 ( .A(u2__abc_44228_n6336), .B(u2__abc_44228_n6596), .Y(u2__abc_44228_n6597_1) );
  AND2X2 AND2X2_2206 ( .A(u2__abc_44228_n6598), .B(u2__abc_44228_n6339), .Y(u2__abc_44228_n6599) );
  AND2X2 AND2X2_2207 ( .A(u2__abc_44228_n6600), .B(u2__abc_44228_n6319), .Y(u2__abc_44228_n6601) );
  AND2X2 AND2X2_2208 ( .A(u2__abc_44228_n6296_1), .B(u2__abc_44228_n6299), .Y(u2__abc_44228_n6602) );
  AND2X2 AND2X2_2209 ( .A(u2__abc_44228_n6307), .B(u2__abc_44228_n6604), .Y(u2__abc_44228_n6605) );
  AND2X2 AND2X2_221 ( .A(_abc_64468_n1261), .B(_abc_64468_n1260), .Y(fracta1_31_) );
  AND2X2 AND2X2_2210 ( .A(u2__abc_44228_n6606), .B(u2__abc_44228_n6310), .Y(u2__abc_44228_n6607_1) );
  AND2X2 AND2X2_2211 ( .A(u2__abc_44228_n6607_1), .B(u2__abc_44228_n6304), .Y(u2__abc_44228_n6608) );
  AND2X2 AND2X2_2212 ( .A(u2__abc_44228_n6612), .B(u2__abc_44228_n6290), .Y(u2__abc_44228_n6613) );
  AND2X2 AND2X2_2213 ( .A(u2__abc_44228_n6615), .B(u2__abc_44228_n6275), .Y(u2__abc_44228_n6616_1) );
  AND2X2 AND2X2_2214 ( .A(u2__abc_44228_n6617), .B(u2__abc_44228_n6272), .Y(u2__abc_44228_n6618) );
  AND2X2 AND2X2_2215 ( .A(u2__abc_44228_n6264), .B(u2__abc_44228_n6267), .Y(u2__abc_44228_n6619) );
  AND2X2 AND2X2_2216 ( .A(u2__abc_44228_n6621), .B(u2__abc_44228_n6258), .Y(u2__abc_44228_n6622) );
  AND2X2 AND2X2_2217 ( .A(u2__abc_44228_n6624), .B(u2__abc_44228_n6246), .Y(u2__abc_44228_n6625_1) );
  AND2X2 AND2X2_2218 ( .A(u2__abc_44228_n6626), .B(u2__abc_44228_n6243), .Y(u2__abc_44228_n6627) );
  AND2X2 AND2X2_2219 ( .A(u2__abc_44228_n6235), .B(u2__abc_44228_n6238), .Y(u2__abc_44228_n6628) );
  AND2X2 AND2X2_222 ( .A(_abc_64468_n1264), .B(_abc_64468_n1263), .Y(fracta1_32_) );
  AND2X2 AND2X2_2220 ( .A(u2__abc_44228_n6631), .B(u2__abc_44228_n6229), .Y(u2__abc_44228_n6632) );
  AND2X2 AND2X2_2221 ( .A(u2__abc_44228_n6634_1), .B(u2__abc_44228_n6202), .Y(u2__abc_44228_n6635) );
  AND2X2 AND2X2_2222 ( .A(u2__abc_44228_n6636), .B(u2__abc_44228_n6227), .Y(u2__abc_44228_n6637) );
  AND2X2 AND2X2_2223 ( .A(u2__abc_44228_n6216), .B(u2__abc_44228_n6638), .Y(u2__abc_44228_n6639) );
  AND2X2 AND2X2_2224 ( .A(u2__abc_44228_n6640), .B(u2__abc_44228_n6219), .Y(u2__abc_44228_n6641) );
  AND2X2 AND2X2_2225 ( .A(u2__abc_44228_n6642), .B(u2__abc_44228_n6199), .Y(u2__abc_44228_n6643) );
  AND2X2 AND2X2_2226 ( .A(u2__abc_44228_n6187_1), .B(u2__abc_44228_n6644_1), .Y(u2__abc_44228_n6645) );
  AND2X2 AND2X2_2227 ( .A(u2__abc_44228_n6646), .B(u2__abc_44228_n6190), .Y(u2__abc_44228_n6647) );
  AND2X2 AND2X2_2228 ( .A(u2__abc_44228_n6647), .B(u2__abc_44228_n6184), .Y(u2__abc_44228_n6648) );
  AND2X2 AND2X2_2229 ( .A(u2__abc_44228_n6176), .B(u2__abc_44228_n6179), .Y(u2__abc_44228_n6649) );
  AND2X2 AND2X2_223 ( .A(_abc_64468_n1267), .B(_abc_64468_n1266), .Y(fracta1_33_) );
  AND2X2 AND2X2_2230 ( .A(u2__abc_44228_n6653_1), .B(u2__abc_44228_n6170), .Y(u2__abc_44228_n6654) );
  AND2X2 AND2X2_2231 ( .A(u2__abc_44228_n6656), .B(u2__abc_44228_n6162), .Y(u2__abc_44228_n6657) );
  AND2X2 AND2X2_2232 ( .A(u2__abc_44228_n6658), .B(u2__abc_44228_n6153), .Y(u2__abc_44228_n6659) );
  AND2X2 AND2X2_2233 ( .A(u2__abc_44228_n6145), .B(u2__abc_44228_n6148), .Y(u2__abc_44228_n6660) );
  AND2X2 AND2X2_2234 ( .A(u2__abc_44228_n6662), .B(u2__abc_44228_n6139), .Y(u2__abc_44228_n6663_1) );
  AND2X2 AND2X2_2235 ( .A(u2__abc_44228_n6665), .B(u2__abc_44228_n6133), .Y(u2__abc_44228_n6666) );
  AND2X2 AND2X2_2236 ( .A(u2__abc_44228_n6667), .B(u2__abc_44228_n6124), .Y(u2__abc_44228_n6668) );
  AND2X2 AND2X2_2237 ( .A(u2__abc_44228_n6116), .B(u2__abc_44228_n6119), .Y(u2__abc_44228_n6669) );
  AND2X2 AND2X2_2238 ( .A(u2__abc_44228_n6672), .B(u2__abc_44228_n6110), .Y(u2__abc_44228_n6673) );
  AND2X2 AND2X2_2239 ( .A(u2__abc_44228_n6675), .B(u2__abc_44228_n6097), .Y(u2__abc_44228_n6676) );
  AND2X2 AND2X2_224 ( .A(_abc_64468_n1270), .B(_abc_64468_n1269), .Y(fracta1_34_) );
  AND2X2 AND2X2_2240 ( .A(u2__abc_44228_n6677), .B(u2__abc_44228_n6094), .Y(u2__abc_44228_n6678) );
  AND2X2 AND2X2_2241 ( .A(u2__abc_44228_n6083), .B(u2__abc_44228_n6679), .Y(u2__abc_44228_n6680) );
  AND2X2 AND2X2_2242 ( .A(u2__abc_44228_n6681_1), .B(u2__abc_44228_n6086_1), .Y(u2__abc_44228_n6682) );
  AND2X2 AND2X2_2243 ( .A(u2__abc_44228_n6683), .B(u2__abc_44228_n6080), .Y(u2__abc_44228_n6684) );
  AND2X2 AND2X2_2244 ( .A(u2__abc_44228_n6057), .B(u2__abc_44228_n6060), .Y(u2__abc_44228_n6685) );
  AND2X2 AND2X2_2245 ( .A(u2__abc_44228_n6688), .B(u2__abc_44228_n6068_1), .Y(u2__abc_44228_n6689_1) );
  AND2X2 AND2X2_2246 ( .A(u2__abc_44228_n6690), .B(u2__abc_44228_n6065), .Y(u2__abc_44228_n6691) );
  AND2X2 AND2X2_2247 ( .A(u2__abc_44228_n6696), .B(u2__abc_44228_n6051), .Y(u2__abc_44228_n6697) );
  AND2X2 AND2X2_2248 ( .A(u2__abc_44228_n6698_1), .B(u2__abc_44228_n6041), .Y(u2__abc_44228_n6699) );
  AND2X2 AND2X2_2249 ( .A(u2__abc_44228_n6700), .B(u2__abc_44228_n6044), .Y(u2__abc_44228_n6701) );
  AND2X2 AND2X2_225 ( .A(_abc_64468_n1273), .B(_abc_64468_n1272), .Y(fracta1_35_) );
  AND2X2 AND2X2_2250 ( .A(u2__abc_44228_n6701), .B(u2__abc_44228_n6032), .Y(u2__abc_44228_n6702) );
  AND2X2 AND2X2_2251 ( .A(u2__abc_44228_n6024), .B(u2__abc_44228_n6027), .Y(u2__abc_44228_n6703) );
  AND2X2 AND2X2_2252 ( .A(u2__abc_44228_n6705), .B(u2__abc_44228_n6018), .Y(u2__abc_44228_n6706) );
  AND2X2 AND2X2_2253 ( .A(u2__abc_44228_n6707_1), .B(u2__abc_44228_n6012_1), .Y(u2__abc_44228_n6708) );
  AND2X2 AND2X2_2254 ( .A(u2__abc_44228_n6709), .B(u2__abc_44228_n6015), .Y(u2__abc_44228_n6710) );
  AND2X2 AND2X2_2255 ( .A(u2__abc_44228_n6710), .B(u2__abc_44228_n6003_1), .Y(u2__abc_44228_n6711) );
  AND2X2 AND2X2_2256 ( .A(u2__abc_44228_n5995), .B(u2__abc_44228_n5998), .Y(u2__abc_44228_n6712) );
  AND2X2 AND2X2_2257 ( .A(u2__abc_44228_n6715), .B(u2__abc_44228_n5989), .Y(u2__abc_44228_n6716) );
  AND2X2 AND2X2_2258 ( .A(u2__abc_44228_n6717_1), .B(u2__abc_44228_n5965), .Y(u2__abc_44228_n6718) );
  AND2X2 AND2X2_2259 ( .A(u2__abc_44228_n5976), .B(u2__abc_44228_n6719), .Y(u2__abc_44228_n6720) );
  AND2X2 AND2X2_226 ( .A(_abc_64468_n1276), .B(_abc_64468_n1275), .Y(fracta1_36_) );
  AND2X2 AND2X2_2260 ( .A(u2__abc_44228_n6721), .B(u2__abc_44228_n5979), .Y(u2__abc_44228_n6722) );
  AND2X2 AND2X2_2261 ( .A(u2__abc_44228_n6722), .B(u2__abc_44228_n5973), .Y(u2__abc_44228_n6723) );
  AND2X2 AND2X2_2262 ( .A(u2__abc_44228_n6724), .B(u2__abc_44228_n5959), .Y(u2__abc_44228_n6725_1) );
  AND2X2 AND2X2_2263 ( .A(u2__abc_44228_n5947), .B(u2__abc_44228_n6726), .Y(u2__abc_44228_n6727) );
  AND2X2 AND2X2_2264 ( .A(u2__abc_44228_n6728), .B(u2__abc_44228_n5950), .Y(u2__abc_44228_n6729) );
  AND2X2 AND2X2_2265 ( .A(u2__abc_44228_n6729), .B(u2__abc_44228_n5944), .Y(u2__abc_44228_n6730) );
  AND2X2 AND2X2_2266 ( .A(u2__abc_44228_n5936), .B(u2__abc_44228_n5939), .Y(u2__abc_44228_n6731) );
  AND2X2 AND2X2_2267 ( .A(u2__abc_44228_n6735_1), .B(u2__abc_44228_n5930_1), .Y(u2__abc_44228_n6736) );
  AND2X2 AND2X2_2268 ( .A(u2__abc_44228_n6738), .B(u2__abc_44228_n5916), .Y(u2__abc_44228_n6739) );
  AND2X2 AND2X2_2269 ( .A(u2__abc_44228_n6740), .B(u2__abc_44228_n5913), .Y(u2__abc_44228_n6741) );
  AND2X2 AND2X2_227 ( .A(_abc_64468_n1279), .B(_abc_64468_n1278), .Y(fracta1_37_) );
  AND2X2 AND2X2_2270 ( .A(u2__abc_44228_n5905), .B(u2__abc_44228_n5908), .Y(u2__abc_44228_n6742) );
  AND2X2 AND2X2_2271 ( .A(u2__abc_44228_n6744), .B(u2__abc_44228_n5899), .Y(u2__abc_44228_n6745) );
  AND2X2 AND2X2_2272 ( .A(u2__abc_44228_n6746), .B(u2__abc_44228_n5893), .Y(u2__abc_44228_n6747) );
  AND2X2 AND2X2_2273 ( .A(u2__abc_44228_n6748), .B(u2__abc_44228_n5896), .Y(u2__abc_44228_n6749) );
  AND2X2 AND2X2_2274 ( .A(u2__abc_44228_n6749), .B(u2__abc_44228_n5884), .Y(u2__abc_44228_n6750) );
  AND2X2 AND2X2_2275 ( .A(u2__abc_44228_n5876), .B(u2__abc_44228_n5879), .Y(u2__abc_44228_n6751) );
  AND2X2 AND2X2_2276 ( .A(u2__abc_44228_n6754), .B(u2__abc_44228_n5870), .Y(u2__abc_44228_n6755) );
  AND2X2 AND2X2_2277 ( .A(u2__abc_44228_n6757), .B(u2__abc_44228_n5843), .Y(u2__abc_44228_n6758) );
  AND2X2 AND2X2_2278 ( .A(u2__abc_44228_n6759), .B(u2__abc_44228_n5868), .Y(u2__abc_44228_n6760) );
  AND2X2 AND2X2_2279 ( .A(u2__abc_44228_n5857), .B(u2__abc_44228_n6761_1), .Y(u2__abc_44228_n6762) );
  AND2X2 AND2X2_228 ( .A(_abc_64468_n1282), .B(_abc_64468_n1281), .Y(fracta1_38_) );
  AND2X2 AND2X2_2280 ( .A(u2__abc_44228_n6763), .B(u2__abc_44228_n5860), .Y(u2__abc_44228_n6764) );
  AND2X2 AND2X2_2281 ( .A(u2__abc_44228_n6765), .B(u2__abc_44228_n5840), .Y(u2__abc_44228_n6766) );
  AND2X2 AND2X2_2282 ( .A(u2__abc_44228_n5817), .B(u2__abc_44228_n5820), .Y(u2__abc_44228_n6767) );
  AND2X2 AND2X2_2283 ( .A(u2__abc_44228_n6769), .B(u2__abc_44228_n5834), .Y(u2__abc_44228_n6770_1) );
  AND2X2 AND2X2_2284 ( .A(u2__abc_44228_n6771), .B(u2__abc_44228_n5837), .Y(u2__abc_44228_n6772) );
  AND2X2 AND2X2_2285 ( .A(u2__abc_44228_n6772), .B(u2__abc_44228_n5825), .Y(u2__abc_44228_n6773) );
  AND2X2 AND2X2_2286 ( .A(u2__abc_44228_n6777), .B(u2__abc_44228_n5811), .Y(u2__abc_44228_n6778) );
  AND2X2 AND2X2_2287 ( .A(u2__abc_44228_n6780), .B(u2__abc_44228_n5796), .Y(u2__abc_44228_n6781) );
  AND2X2 AND2X2_2288 ( .A(u2__abc_44228_n6782), .B(u2__abc_44228_n5793_1), .Y(u2__abc_44228_n6783) );
  AND2X2 AND2X2_2289 ( .A(u2__abc_44228_n5785), .B(u2__abc_44228_n5788), .Y(u2__abc_44228_n6784) );
  AND2X2 AND2X2_229 ( .A(_abc_64468_n1285), .B(_abc_64468_n1284), .Y(fracta1_39_) );
  AND2X2 AND2X2_2290 ( .A(u2__abc_44228_n6786), .B(u2__abc_44228_n5779), .Y(u2__abc_44228_n6787) );
  AND2X2 AND2X2_2291 ( .A(u2__abc_44228_n6788), .B(u2__abc_44228_n5773), .Y(u2__abc_44228_n6789_1) );
  AND2X2 AND2X2_2292 ( .A(u2__abc_44228_n6790), .B(u2__abc_44228_n5776), .Y(u2__abc_44228_n6791) );
  AND2X2 AND2X2_2293 ( .A(u2__abc_44228_n6791), .B(u2__abc_44228_n5764), .Y(u2__abc_44228_n6792) );
  AND2X2 AND2X2_2294 ( .A(u2__abc_44228_n5756_1), .B(u2__abc_44228_n5759), .Y(u2__abc_44228_n6793) );
  AND2X2 AND2X2_2295 ( .A(u2__abc_44228_n6796), .B(u2__abc_44228_n5750), .Y(u2__abc_44228_n6797_1) );
  AND2X2 AND2X2_2296 ( .A(u2__abc_44228_n6799), .B(u2__abc_44228_n5723), .Y(u2__abc_44228_n6800) );
  AND2X2 AND2X2_2297 ( .A(u2__abc_44228_n6801), .B(u2__abc_44228_n5748), .Y(u2__abc_44228_n6802) );
  AND2X2 AND2X2_2298 ( .A(u2__abc_44228_n5737_1), .B(u2__abc_44228_n6803), .Y(u2__abc_44228_n6804) );
  AND2X2 AND2X2_2299 ( .A(u2__abc_44228_n6805), .B(u2__abc_44228_n5740), .Y(u2__abc_44228_n6806) );
  AND2X2 AND2X2_23 ( .A(_abc_64468_n753_bF_buf5), .B(sqrto_22_), .Y(_auto_iopadmap_cc_313_execute_65414_58_) );
  AND2X2 AND2X2_230 ( .A(_abc_64468_n1288), .B(_abc_64468_n1287), .Y(fracta1_40_) );
  AND2X2 AND2X2_2300 ( .A(u2__abc_44228_n6807_1), .B(u2__abc_44228_n5720), .Y(u2__abc_44228_n6808) );
  AND2X2 AND2X2_2301 ( .A(u2__abc_44228_n5697), .B(u2__abc_44228_n5700_1), .Y(u2__abc_44228_n6809) );
  AND2X2 AND2X2_2302 ( .A(u2__abc_44228_n6812), .B(u2__abc_44228_n5708), .Y(u2__abc_44228_n6813) );
  AND2X2 AND2X2_2303 ( .A(u2__abc_44228_n6814), .B(u2__abc_44228_n5705), .Y(u2__abc_44228_n6815_1) );
  AND2X2 AND2X2_2304 ( .A(u2__abc_44228_n6818), .B(u2__abc_44228_n5691), .Y(u2__abc_44228_n6819) );
  AND2X2 AND2X2_2305 ( .A(u2__abc_44228_n6821), .B(u2__abc_44228_n5663), .Y(u2__abc_44228_n6822) );
  AND2X2 AND2X2_2306 ( .A(u2__abc_44228_n6823), .B(u2__abc_44228_n5688), .Y(u2__abc_44228_n6824) );
  AND2X2 AND2X2_2307 ( .A(u2__abc_44228_n5677), .B(u2__abc_44228_n6825_1), .Y(u2__abc_44228_n6826) );
  AND2X2 AND2X2_2308 ( .A(u2__abc_44228_n6827), .B(u2__abc_44228_n5680), .Y(u2__abc_44228_n6828) );
  AND2X2 AND2X2_2309 ( .A(u2__abc_44228_n6829), .B(u2__abc_44228_n5660), .Y(u2__abc_44228_n6830) );
  AND2X2 AND2X2_231 ( .A(_abc_64468_n1291), .B(_abc_64468_n1290), .Y(fracta1_41_) );
  AND2X2 AND2X2_2310 ( .A(u2__abc_44228_n6831), .B(u2__abc_44228_n5654), .Y(u2__abc_44228_n6832) );
  AND2X2 AND2X2_2311 ( .A(u2__abc_44228_n6833_1), .B(u2__abc_44228_n5657), .Y(u2__abc_44228_n6834) );
  AND2X2 AND2X2_2312 ( .A(u2__abc_44228_n6834), .B(u2__abc_44228_n5645), .Y(u2__abc_44228_n6835) );
  AND2X2 AND2X2_2313 ( .A(u2__abc_44228_n5637), .B(u2__abc_44228_n5640), .Y(u2__abc_44228_n6836) );
  AND2X2 AND2X2_2314 ( .A(u2__abc_44228_n6839), .B(u2__abc_44228_n5631), .Y(u2__abc_44228_n6840) );
  AND2X2 AND2X2_2315 ( .A(u2__abc_44228_n6842_1), .B(u2__abc_44228_n5604), .Y(u2__abc_44228_n6843) );
  AND2X2 AND2X2_2316 ( .A(u2__abc_44228_n6844), .B(u2__abc_44228_n5629), .Y(u2__abc_44228_n6845) );
  AND2X2 AND2X2_2317 ( .A(u2__abc_44228_n5618), .B(u2__abc_44228_n6846), .Y(u2__abc_44228_n6847) );
  AND2X2 AND2X2_2318 ( .A(u2__abc_44228_n6848), .B(u2__abc_44228_n5621), .Y(u2__abc_44228_n6849) );
  AND2X2 AND2X2_2319 ( .A(u2__abc_44228_n6850), .B(u2__abc_44228_n5601), .Y(u2__abc_44228_n6851_1) );
  AND2X2 AND2X2_232 ( .A(_abc_64468_n1294), .B(_abc_64468_n1293), .Y(fracta1_42_) );
  AND2X2 AND2X2_2320 ( .A(u2__abc_44228_n5578), .B(u2__abc_44228_n5581), .Y(u2__abc_44228_n6852) );
  AND2X2 AND2X2_2321 ( .A(u2__abc_44228_n5589), .B(u2__abc_44228_n6854), .Y(u2__abc_44228_n6855) );
  AND2X2 AND2X2_2322 ( .A(u2__abc_44228_n6856), .B(u2__abc_44228_n5592), .Y(u2__abc_44228_n6857) );
  AND2X2 AND2X2_2323 ( .A(u2__abc_44228_n6857), .B(u2__abc_44228_n5586), .Y(u2__abc_44228_n6858) );
  AND2X2 AND2X2_2324 ( .A(u2__abc_44228_n6866), .B(u2_remHi_445_), .Y(u2__abc_44228_n6867) );
  AND2X2 AND2X2_2325 ( .A(u2__abc_44228_n6869_1), .B(u2_o_445_), .Y(u2__abc_44228_n6870) );
  AND2X2 AND2X2_2326 ( .A(u2__abc_44228_n6868), .B(u2__abc_44228_n6871), .Y(u2__abc_44228_n6872) );
  AND2X2 AND2X2_2327 ( .A(u2__abc_44228_n6873), .B(u2_remHi_444_), .Y(u2__abc_44228_n6874) );
  AND2X2 AND2X2_2328 ( .A(u2__abc_44228_n6875), .B(u2_o_444_), .Y(u2__abc_44228_n6876) );
  AND2X2 AND2X2_2329 ( .A(u2__abc_44228_n6878_1), .B(u2__abc_44228_n6872), .Y(u2__abc_44228_n6879) );
  AND2X2 AND2X2_233 ( .A(_abc_64468_n1297), .B(_abc_64468_n1296), .Y(fracta1_43_) );
  AND2X2 AND2X2_2330 ( .A(u2__abc_44228_n6880), .B(u2_remHi_443_), .Y(u2__abc_44228_n6881) );
  AND2X2 AND2X2_2331 ( .A(u2__abc_44228_n6883), .B(u2_o_443_), .Y(u2__abc_44228_n6884) );
  AND2X2 AND2X2_2332 ( .A(u2__abc_44228_n6882), .B(u2__abc_44228_n6885), .Y(u2__abc_44228_n6886) );
  AND2X2 AND2X2_2333 ( .A(u2__abc_44228_n6887_1), .B(u2_remHi_442_), .Y(u2__abc_44228_n6888) );
  AND2X2 AND2X2_2334 ( .A(u2__abc_44228_n6889), .B(u2_o_442_), .Y(u2__abc_44228_n6890) );
  AND2X2 AND2X2_2335 ( .A(u2__abc_44228_n6892), .B(u2__abc_44228_n6886), .Y(u2__abc_44228_n6893) );
  AND2X2 AND2X2_2336 ( .A(u2__abc_44228_n6879), .B(u2__abc_44228_n6893), .Y(u2__abc_44228_n6894) );
  AND2X2 AND2X2_2337 ( .A(u2__abc_44228_n6895), .B(u2_remHi_441_), .Y(u2__abc_44228_n6896) );
  AND2X2 AND2X2_2338 ( .A(u2__abc_44228_n6898), .B(u2_o_441_), .Y(u2__abc_44228_n6899) );
  AND2X2 AND2X2_2339 ( .A(u2__abc_44228_n6897_1), .B(u2__abc_44228_n6900), .Y(u2__abc_44228_n6901) );
  AND2X2 AND2X2_234 ( .A(_abc_64468_n1300), .B(_abc_64468_n1299), .Y(fracta1_44_) );
  AND2X2 AND2X2_2340 ( .A(u2__abc_44228_n6902), .B(u2_remHi_440_), .Y(u2__abc_44228_n6903) );
  AND2X2 AND2X2_2341 ( .A(u2__abc_44228_n6904), .B(u2_o_440_), .Y(u2__abc_44228_n6905) );
  AND2X2 AND2X2_2342 ( .A(u2__abc_44228_n6907), .B(u2__abc_44228_n6901), .Y(u2__abc_44228_n6908) );
  AND2X2 AND2X2_2343 ( .A(u2__abc_44228_n6909), .B(u2_remHi_439_), .Y(u2__abc_44228_n6910) );
  AND2X2 AND2X2_2344 ( .A(u2__abc_44228_n6912), .B(u2_o_439_), .Y(u2__abc_44228_n6913) );
  AND2X2 AND2X2_2345 ( .A(u2__abc_44228_n6911), .B(u2__abc_44228_n6914), .Y(u2__abc_44228_n6915_1) );
  AND2X2 AND2X2_2346 ( .A(u2__abc_44228_n6916), .B(u2_remHi_438_), .Y(u2__abc_44228_n6917) );
  AND2X2 AND2X2_2347 ( .A(u2__abc_44228_n6918), .B(u2_o_438_), .Y(u2__abc_44228_n6919) );
  AND2X2 AND2X2_2348 ( .A(u2__abc_44228_n6921), .B(u2__abc_44228_n6915_1), .Y(u2__abc_44228_n6922) );
  AND2X2 AND2X2_2349 ( .A(u2__abc_44228_n6908), .B(u2__abc_44228_n6922), .Y(u2__abc_44228_n6923) );
  AND2X2 AND2X2_235 ( .A(_abc_64468_n1303), .B(_abc_64468_n1302), .Y(fracta1_45_) );
  AND2X2 AND2X2_2350 ( .A(u2__abc_44228_n6894), .B(u2__abc_44228_n6923), .Y(u2__abc_44228_n6924_1) );
  AND2X2 AND2X2_2351 ( .A(u2__abc_44228_n6925), .B(u2_remHi_437_), .Y(u2__abc_44228_n6926) );
  AND2X2 AND2X2_2352 ( .A(u2__abc_44228_n6928), .B(u2_o_437_), .Y(u2__abc_44228_n6929) );
  AND2X2 AND2X2_2353 ( .A(u2__abc_44228_n6927), .B(u2__abc_44228_n6930), .Y(u2__abc_44228_n6931) );
  AND2X2 AND2X2_2354 ( .A(u2__abc_44228_n6932), .B(u2_remHi_436_), .Y(u2__abc_44228_n6933) );
  AND2X2 AND2X2_2355 ( .A(u2__abc_44228_n6934_1), .B(u2_o_436_), .Y(u2__abc_44228_n6935) );
  AND2X2 AND2X2_2356 ( .A(u2__abc_44228_n6937), .B(u2__abc_44228_n6931), .Y(u2__abc_44228_n6938) );
  AND2X2 AND2X2_2357 ( .A(u2__abc_44228_n6939), .B(u2_remHi_434_), .Y(u2__abc_44228_n6940) );
  AND2X2 AND2X2_2358 ( .A(u2__abc_44228_n6941), .B(u2_o_434_), .Y(u2__abc_44228_n6942) );
  AND2X2 AND2X2_2359 ( .A(u2__abc_44228_n6945), .B(u2_remHi_435_), .Y(u2__abc_44228_n6946) );
  AND2X2 AND2X2_236 ( .A(_abc_64468_n1306), .B(_abc_64468_n1305), .Y(fracta1_46_) );
  AND2X2 AND2X2_2360 ( .A(u2__abc_44228_n6948), .B(u2_o_435_), .Y(u2__abc_44228_n6949) );
  AND2X2 AND2X2_2361 ( .A(u2__abc_44228_n6947), .B(u2__abc_44228_n6950), .Y(u2__abc_44228_n6951) );
  AND2X2 AND2X2_2362 ( .A(u2__abc_44228_n6944), .B(u2__abc_44228_n6951), .Y(u2__abc_44228_n6952) );
  AND2X2 AND2X2_2363 ( .A(u2__abc_44228_n6938), .B(u2__abc_44228_n6952), .Y(u2__abc_44228_n6953_1) );
  AND2X2 AND2X2_2364 ( .A(u2__abc_44228_n6954), .B(u2_remHi_431_), .Y(u2__abc_44228_n6955) );
  AND2X2 AND2X2_2365 ( .A(u2__abc_44228_n6957), .B(u2_o_431_), .Y(u2__abc_44228_n6958) );
  AND2X2 AND2X2_2366 ( .A(u2__abc_44228_n6956), .B(u2__abc_44228_n6959), .Y(u2__abc_44228_n6960) );
  AND2X2 AND2X2_2367 ( .A(u2__abc_44228_n6961_1), .B(u2_remHi_430_), .Y(u2__abc_44228_n6962) );
  AND2X2 AND2X2_2368 ( .A(u2__abc_44228_n6963), .B(u2_o_430_), .Y(u2__abc_44228_n6964) );
  AND2X2 AND2X2_2369 ( .A(u2__abc_44228_n6966), .B(u2__abc_44228_n6960), .Y(u2__abc_44228_n6967) );
  AND2X2 AND2X2_237 ( .A(_abc_64468_n1309), .B(_abc_64468_n1308), .Y(fracta1_47_) );
  AND2X2 AND2X2_2370 ( .A(u2__abc_44228_n6968), .B(u2_remHi_433_), .Y(u2__abc_44228_n6969) );
  AND2X2 AND2X2_2371 ( .A(u2__abc_44228_n6971_1), .B(u2_o_433_), .Y(u2__abc_44228_n6972) );
  AND2X2 AND2X2_2372 ( .A(u2__abc_44228_n6970), .B(u2__abc_44228_n6973), .Y(u2__abc_44228_n6974) );
  AND2X2 AND2X2_2373 ( .A(u2__abc_44228_n6975), .B(u2_remHi_432_), .Y(u2__abc_44228_n6976) );
  AND2X2 AND2X2_2374 ( .A(u2__abc_44228_n6977), .B(u2_o_432_), .Y(u2__abc_44228_n6978) );
  AND2X2 AND2X2_2375 ( .A(u2__abc_44228_n6980), .B(u2__abc_44228_n6974), .Y(u2__abc_44228_n6981) );
  AND2X2 AND2X2_2376 ( .A(u2__abc_44228_n6967), .B(u2__abc_44228_n6981), .Y(u2__abc_44228_n6982) );
  AND2X2 AND2X2_2377 ( .A(u2__abc_44228_n6953_1), .B(u2__abc_44228_n6982), .Y(u2__abc_44228_n6983) );
  AND2X2 AND2X2_2378 ( .A(u2__abc_44228_n6924_1), .B(u2__abc_44228_n6983), .Y(u2__abc_44228_n6984) );
  AND2X2 AND2X2_2379 ( .A(u2__abc_44228_n6985), .B(u2_remHi_429_), .Y(u2__abc_44228_n6986) );
  AND2X2 AND2X2_238 ( .A(_abc_64468_n1312), .B(_abc_64468_n1311), .Y(fracta1_48_) );
  AND2X2 AND2X2_2380 ( .A(u2__abc_44228_n6988_1), .B(u2_o_429_), .Y(u2__abc_44228_n6989) );
  AND2X2 AND2X2_2381 ( .A(u2__abc_44228_n6987), .B(u2__abc_44228_n6990), .Y(u2__abc_44228_n6991) );
  AND2X2 AND2X2_2382 ( .A(u2__abc_44228_n6992), .B(u2_remHi_428_), .Y(u2__abc_44228_n6993) );
  AND2X2 AND2X2_2383 ( .A(u2__abc_44228_n6994), .B(u2_o_428_), .Y(u2__abc_44228_n6995) );
  AND2X2 AND2X2_2384 ( .A(u2__abc_44228_n6997_1), .B(u2__abc_44228_n6991), .Y(u2__abc_44228_n6998) );
  AND2X2 AND2X2_2385 ( .A(u2__abc_44228_n6999), .B(u2_remHi_427_), .Y(u2__abc_44228_n7000) );
  AND2X2 AND2X2_2386 ( .A(u2__abc_44228_n7002), .B(u2_o_427_), .Y(u2__abc_44228_n7003) );
  AND2X2 AND2X2_2387 ( .A(u2__abc_44228_n7001), .B(u2__abc_44228_n7004), .Y(u2__abc_44228_n7005) );
  AND2X2 AND2X2_2388 ( .A(u2__abc_44228_n7006), .B(u2_remHi_426_), .Y(u2__abc_44228_n7007_1) );
  AND2X2 AND2X2_2389 ( .A(u2__abc_44228_n7008), .B(u2_o_426_), .Y(u2__abc_44228_n7009) );
  AND2X2 AND2X2_239 ( .A(_abc_64468_n1315), .B(_abc_64468_n1314), .Y(fracta1_49_) );
  AND2X2 AND2X2_2390 ( .A(u2__abc_44228_n7011), .B(u2__abc_44228_n7005), .Y(u2__abc_44228_n7012) );
  AND2X2 AND2X2_2391 ( .A(u2__abc_44228_n6998), .B(u2__abc_44228_n7012), .Y(u2__abc_44228_n7013) );
  AND2X2 AND2X2_2392 ( .A(u2__abc_44228_n7014_1), .B(u2_remHi_425_), .Y(u2__abc_44228_n7015) );
  AND2X2 AND2X2_2393 ( .A(u2__abc_44228_n7017), .B(u2_o_425_), .Y(u2__abc_44228_n7018) );
  AND2X2 AND2X2_2394 ( .A(u2__abc_44228_n7016), .B(u2__abc_44228_n7019), .Y(u2__abc_44228_n7020) );
  AND2X2 AND2X2_2395 ( .A(u2__abc_44228_n7021), .B(u2_remHi_424_), .Y(u2__abc_44228_n7022_1) );
  AND2X2 AND2X2_2396 ( .A(u2__abc_44228_n7023), .B(u2_o_424_), .Y(u2__abc_44228_n7024) );
  AND2X2 AND2X2_2397 ( .A(u2__abc_44228_n7026), .B(u2__abc_44228_n7020), .Y(u2__abc_44228_n7027) );
  AND2X2 AND2X2_2398 ( .A(u2__abc_44228_n7028), .B(u2_remHi_423_), .Y(u2__abc_44228_n7029) );
  AND2X2 AND2X2_2399 ( .A(u2__abc_44228_n7031), .B(u2_o_423_), .Y(u2__abc_44228_n7032_1) );
  AND2X2 AND2X2_24 ( .A(_abc_64468_n753_bF_buf4), .B(sqrto_23_), .Y(_auto_iopadmap_cc_313_execute_65414_59_) );
  AND2X2 AND2X2_240 ( .A(_abc_64468_n1318), .B(_abc_64468_n1317), .Y(fracta1_50_) );
  AND2X2 AND2X2_2400 ( .A(u2__abc_44228_n7030), .B(u2__abc_44228_n7033), .Y(u2__abc_44228_n7034) );
  AND2X2 AND2X2_2401 ( .A(u2__abc_44228_n7035), .B(u2_remHi_422_), .Y(u2__abc_44228_n7036) );
  AND2X2 AND2X2_2402 ( .A(u2__abc_44228_n7037), .B(u2_o_422_), .Y(u2__abc_44228_n7038) );
  AND2X2 AND2X2_2403 ( .A(u2__abc_44228_n7040), .B(u2__abc_44228_n7034), .Y(u2__abc_44228_n7041) );
  AND2X2 AND2X2_2404 ( .A(u2__abc_44228_n7027), .B(u2__abc_44228_n7041), .Y(u2__abc_44228_n7042_1) );
  AND2X2 AND2X2_2405 ( .A(u2__abc_44228_n7013), .B(u2__abc_44228_n7042_1), .Y(u2__abc_44228_n7043) );
  AND2X2 AND2X2_2406 ( .A(u2__abc_44228_n7044), .B(u2_remHi_421_), .Y(u2__abc_44228_n7045) );
  AND2X2 AND2X2_2407 ( .A(u2__abc_44228_n7047), .B(u2_o_421_), .Y(u2__abc_44228_n7048) );
  AND2X2 AND2X2_2408 ( .A(u2__abc_44228_n7046), .B(u2__abc_44228_n7049), .Y(u2__abc_44228_n7050_1) );
  AND2X2 AND2X2_2409 ( .A(u2__abc_44228_n7051), .B(u2_remHi_420_), .Y(u2__abc_44228_n7052) );
  AND2X2 AND2X2_241 ( .A(_abc_64468_n1321), .B(_abc_64468_n1320), .Y(fracta1_51_) );
  AND2X2 AND2X2_2410 ( .A(u2__abc_44228_n7053), .B(u2_o_420_), .Y(u2__abc_44228_n7054) );
  AND2X2 AND2X2_2411 ( .A(u2__abc_44228_n7056), .B(u2__abc_44228_n7050_1), .Y(u2__abc_44228_n7057) );
  AND2X2 AND2X2_2412 ( .A(u2__abc_44228_n7058), .B(u2_remHi_419_), .Y(u2__abc_44228_n7059_1) );
  AND2X2 AND2X2_2413 ( .A(u2__abc_44228_n7061), .B(u2_o_419_), .Y(u2__abc_44228_n7062) );
  AND2X2 AND2X2_2414 ( .A(u2__abc_44228_n7060), .B(u2__abc_44228_n7063), .Y(u2__abc_44228_n7064) );
  AND2X2 AND2X2_2415 ( .A(u2__abc_44228_n7065), .B(u2_remHi_418_), .Y(u2__abc_44228_n7066) );
  AND2X2 AND2X2_2416 ( .A(u2__abc_44228_n7067), .B(u2_o_418_), .Y(u2__abc_44228_n7068_1) );
  AND2X2 AND2X2_2417 ( .A(u2__abc_44228_n7070), .B(u2__abc_44228_n7064), .Y(u2__abc_44228_n7071) );
  AND2X2 AND2X2_2418 ( .A(u2__abc_44228_n7057), .B(u2__abc_44228_n7071), .Y(u2__abc_44228_n7072) );
  AND2X2 AND2X2_2419 ( .A(u2__abc_44228_n7073), .B(u2_remHi_417_), .Y(u2__abc_44228_n7074) );
  AND2X2 AND2X2_242 ( .A(_abc_64468_n1324), .B(_abc_64468_n1323), .Y(fracta1_52_) );
  AND2X2 AND2X2_2420 ( .A(u2__abc_44228_n7076), .B(u2_o_417_), .Y(u2__abc_44228_n7077) );
  AND2X2 AND2X2_2421 ( .A(u2__abc_44228_n7075), .B(u2__abc_44228_n7078_1), .Y(u2__abc_44228_n7079) );
  AND2X2 AND2X2_2422 ( .A(u2__abc_44228_n7080), .B(u2_remHi_416_), .Y(u2__abc_44228_n7081) );
  AND2X2 AND2X2_2423 ( .A(u2__abc_44228_n7082), .B(u2_o_416_), .Y(u2__abc_44228_n7083) );
  AND2X2 AND2X2_2424 ( .A(u2__abc_44228_n7085), .B(u2__abc_44228_n7079), .Y(u2__abc_44228_n7086) );
  AND2X2 AND2X2_2425 ( .A(u2__abc_44228_n7087), .B(u2_remHi_414_), .Y(u2__abc_44228_n7088_1) );
  AND2X2 AND2X2_2426 ( .A(u2__abc_44228_n7089), .B(u2_o_414_), .Y(u2__abc_44228_n7090) );
  AND2X2 AND2X2_2427 ( .A(u2__abc_44228_n7093), .B(u2_remHi_415_), .Y(u2__abc_44228_n7094) );
  AND2X2 AND2X2_2428 ( .A(u2__abc_44228_n7096), .B(u2_o_415_), .Y(u2__abc_44228_n7097) );
  AND2X2 AND2X2_2429 ( .A(u2__abc_44228_n7095), .B(u2__abc_44228_n7098_1), .Y(u2__abc_44228_n7099) );
  AND2X2 AND2X2_243 ( .A(_abc_64468_n1327), .B(_abc_64468_n1326), .Y(fracta1_53_) );
  AND2X2 AND2X2_2430 ( .A(u2__abc_44228_n7092), .B(u2__abc_44228_n7099), .Y(u2__abc_44228_n7100) );
  AND2X2 AND2X2_2431 ( .A(u2__abc_44228_n7086), .B(u2__abc_44228_n7100), .Y(u2__abc_44228_n7101) );
  AND2X2 AND2X2_2432 ( .A(u2__abc_44228_n7072), .B(u2__abc_44228_n7101), .Y(u2__abc_44228_n7102) );
  AND2X2 AND2X2_2433 ( .A(u2__abc_44228_n7043), .B(u2__abc_44228_n7102), .Y(u2__abc_44228_n7103) );
  AND2X2 AND2X2_2434 ( .A(u2__abc_44228_n6984), .B(u2__abc_44228_n7103), .Y(u2__abc_44228_n7104) );
  AND2X2 AND2X2_2435 ( .A(u2__abc_44228_n7105), .B(u2_remHi_413_), .Y(u2__abc_44228_n7106_1) );
  AND2X2 AND2X2_2436 ( .A(u2__abc_44228_n7108), .B(u2_o_413_), .Y(u2__abc_44228_n7109) );
  AND2X2 AND2X2_2437 ( .A(u2__abc_44228_n7107), .B(u2__abc_44228_n7110), .Y(u2__abc_44228_n7111) );
  AND2X2 AND2X2_2438 ( .A(u2__abc_44228_n7112), .B(u2_remHi_412_), .Y(u2__abc_44228_n7113) );
  AND2X2 AND2X2_2439 ( .A(u2__abc_44228_n7114), .B(u2_o_412_), .Y(u2__abc_44228_n7115) );
  AND2X2 AND2X2_244 ( .A(_abc_64468_n1330), .B(_abc_64468_n1329), .Y(fracta1_54_) );
  AND2X2 AND2X2_2440 ( .A(u2__abc_44228_n7117), .B(u2__abc_44228_n7111), .Y(u2__abc_44228_n7118) );
  AND2X2 AND2X2_2441 ( .A(u2__abc_44228_n7119), .B(u2_remHi_411_), .Y(u2__abc_44228_n7120) );
  AND2X2 AND2X2_2442 ( .A(u2__abc_44228_n7122), .B(u2_o_411_), .Y(u2__abc_44228_n7123) );
  AND2X2 AND2X2_2443 ( .A(u2__abc_44228_n7121), .B(u2__abc_44228_n7124), .Y(u2__abc_44228_n7125_1) );
  AND2X2 AND2X2_2444 ( .A(u2__abc_44228_n7126), .B(u2_remHi_410_), .Y(u2__abc_44228_n7127) );
  AND2X2 AND2X2_2445 ( .A(u2__abc_44228_n7128), .B(u2_o_410_), .Y(u2__abc_44228_n7129) );
  AND2X2 AND2X2_2446 ( .A(u2__abc_44228_n7131), .B(u2__abc_44228_n7125_1), .Y(u2__abc_44228_n7132) );
  AND2X2 AND2X2_2447 ( .A(u2__abc_44228_n7118), .B(u2__abc_44228_n7132), .Y(u2__abc_44228_n7133) );
  AND2X2 AND2X2_2448 ( .A(u2__abc_44228_n7134_1), .B(u2_remHi_409_), .Y(u2__abc_44228_n7135) );
  AND2X2 AND2X2_2449 ( .A(u2__abc_44228_n7137), .B(u2_o_409_), .Y(u2__abc_44228_n7138) );
  AND2X2 AND2X2_245 ( .A(_abc_64468_n1333), .B(_abc_64468_n1332), .Y(fracta1_55_) );
  AND2X2 AND2X2_2450 ( .A(u2__abc_44228_n7136), .B(u2__abc_44228_n7139), .Y(u2__abc_44228_n7140) );
  AND2X2 AND2X2_2451 ( .A(u2__abc_44228_n7141), .B(u2_remHi_408_), .Y(u2__abc_44228_n7142) );
  AND2X2 AND2X2_2452 ( .A(u2__abc_44228_n7143_1), .B(u2_o_408_), .Y(u2__abc_44228_n7144) );
  AND2X2 AND2X2_2453 ( .A(u2__abc_44228_n7146), .B(u2__abc_44228_n7140), .Y(u2__abc_44228_n7147) );
  AND2X2 AND2X2_2454 ( .A(u2__abc_44228_n7148), .B(u2_remHi_407_), .Y(u2__abc_44228_n7149) );
  AND2X2 AND2X2_2455 ( .A(u2__abc_44228_n7151), .B(u2_o_407_), .Y(u2__abc_44228_n7152) );
  AND2X2 AND2X2_2456 ( .A(u2__abc_44228_n7150), .B(u2__abc_44228_n7153_1), .Y(u2__abc_44228_n7154) );
  AND2X2 AND2X2_2457 ( .A(u2__abc_44228_n7155), .B(u2_remHi_406_), .Y(u2__abc_44228_n7156) );
  AND2X2 AND2X2_2458 ( .A(u2__abc_44228_n7157), .B(u2_o_406_), .Y(u2__abc_44228_n7158) );
  AND2X2 AND2X2_2459 ( .A(u2__abc_44228_n7160), .B(u2__abc_44228_n7154), .Y(u2__abc_44228_n7161_1) );
  AND2X2 AND2X2_246 ( .A(_abc_64468_n1336), .B(_abc_64468_n1335), .Y(fracta1_56_) );
  AND2X2 AND2X2_2460 ( .A(u2__abc_44228_n7147), .B(u2__abc_44228_n7161_1), .Y(u2__abc_44228_n7162) );
  AND2X2 AND2X2_2461 ( .A(u2__abc_44228_n7133), .B(u2__abc_44228_n7162), .Y(u2__abc_44228_n7163) );
  AND2X2 AND2X2_2462 ( .A(u2__abc_44228_n7164), .B(u2_remHi_405_), .Y(u2__abc_44228_n7165) );
  AND2X2 AND2X2_2463 ( .A(u2__abc_44228_n7167), .B(u2_o_405_), .Y(u2__abc_44228_n7168) );
  AND2X2 AND2X2_2464 ( .A(u2__abc_44228_n7166), .B(u2__abc_44228_n7169), .Y(u2__abc_44228_n7170_1) );
  AND2X2 AND2X2_2465 ( .A(u2__abc_44228_n7171), .B(u2_remHi_404_), .Y(u2__abc_44228_n7172) );
  AND2X2 AND2X2_2466 ( .A(u2__abc_44228_n7173), .B(u2_o_404_), .Y(u2__abc_44228_n7174) );
  AND2X2 AND2X2_2467 ( .A(u2__abc_44228_n7176), .B(u2__abc_44228_n7170_1), .Y(u2__abc_44228_n7177) );
  AND2X2 AND2X2_2468 ( .A(u2__abc_44228_n7178), .B(u2_remHi_403_), .Y(u2__abc_44228_n7179_1) );
  AND2X2 AND2X2_2469 ( .A(u2__abc_44228_n7181), .B(u2_o_403_), .Y(u2__abc_44228_n7182) );
  AND2X2 AND2X2_247 ( .A(_abc_64468_n1339), .B(_abc_64468_n1338), .Y(fracta1_57_) );
  AND2X2 AND2X2_2470 ( .A(u2__abc_44228_n7180), .B(u2__abc_44228_n7183), .Y(u2__abc_44228_n7184) );
  AND2X2 AND2X2_2471 ( .A(u2__abc_44228_n7185), .B(u2_remHi_402_), .Y(u2__abc_44228_n7186) );
  AND2X2 AND2X2_2472 ( .A(u2__abc_44228_n7187), .B(u2_o_402_), .Y(u2__abc_44228_n7188) );
  AND2X2 AND2X2_2473 ( .A(u2__abc_44228_n7190), .B(u2__abc_44228_n7184), .Y(u2__abc_44228_n7191) );
  AND2X2 AND2X2_2474 ( .A(u2__abc_44228_n7177), .B(u2__abc_44228_n7191), .Y(u2__abc_44228_n7192) );
  AND2X2 AND2X2_2475 ( .A(u2__abc_44228_n7193), .B(u2_remHi_401_), .Y(u2__abc_44228_n7194) );
  AND2X2 AND2X2_2476 ( .A(u2__abc_44228_n7196), .B(u2_o_401_), .Y(u2__abc_44228_n7197_1) );
  AND2X2 AND2X2_2477 ( .A(u2__abc_44228_n7195), .B(u2__abc_44228_n7198), .Y(u2__abc_44228_n7199) );
  AND2X2 AND2X2_2478 ( .A(u2__abc_44228_n7200), .B(u2_remHi_400_), .Y(u2__abc_44228_n7201) );
  AND2X2 AND2X2_2479 ( .A(u2__abc_44228_n7202), .B(u2_o_400_), .Y(u2__abc_44228_n7203) );
  AND2X2 AND2X2_248 ( .A(_abc_64468_n1342), .B(_abc_64468_n1341), .Y(fracta1_58_) );
  AND2X2 AND2X2_2480 ( .A(u2__abc_44228_n7205), .B(u2__abc_44228_n7199), .Y(u2__abc_44228_n7206_1) );
  AND2X2 AND2X2_2481 ( .A(u2__abc_44228_n7207), .B(u2_remHi_398_), .Y(u2__abc_44228_n7208) );
  AND2X2 AND2X2_2482 ( .A(u2__abc_44228_n7209), .B(u2_o_398_), .Y(u2__abc_44228_n7210) );
  AND2X2 AND2X2_2483 ( .A(u2__abc_44228_n7213), .B(u2_remHi_399_), .Y(u2__abc_44228_n7214) );
  AND2X2 AND2X2_2484 ( .A(u2__abc_44228_n7216), .B(u2_o_399_), .Y(u2__abc_44228_n7217) );
  AND2X2 AND2X2_2485 ( .A(u2__abc_44228_n7215_1), .B(u2__abc_44228_n7218), .Y(u2__abc_44228_n7219) );
  AND2X2 AND2X2_2486 ( .A(u2__abc_44228_n7212), .B(u2__abc_44228_n7219), .Y(u2__abc_44228_n7220) );
  AND2X2 AND2X2_2487 ( .A(u2__abc_44228_n7206_1), .B(u2__abc_44228_n7220), .Y(u2__abc_44228_n7221) );
  AND2X2 AND2X2_2488 ( .A(u2__abc_44228_n7192), .B(u2__abc_44228_n7221), .Y(u2__abc_44228_n7222) );
  AND2X2 AND2X2_2489 ( .A(u2__abc_44228_n7163), .B(u2__abc_44228_n7222), .Y(u2__abc_44228_n7223) );
  AND2X2 AND2X2_249 ( .A(_abc_64468_n1345), .B(_abc_64468_n1344), .Y(fracta1_59_) );
  AND2X2 AND2X2_2490 ( .A(u2__abc_44228_n7224), .B(u2_remHi_397_), .Y(u2__abc_44228_n7225_1) );
  AND2X2 AND2X2_2491 ( .A(u2__abc_44228_n7227), .B(u2_o_397_), .Y(u2__abc_44228_n7228) );
  AND2X2 AND2X2_2492 ( .A(u2__abc_44228_n7226), .B(u2__abc_44228_n7229), .Y(u2__abc_44228_n7230) );
  AND2X2 AND2X2_2493 ( .A(u2__abc_44228_n7231), .B(u2_remHi_396_), .Y(u2__abc_44228_n7232) );
  AND2X2 AND2X2_2494 ( .A(u2__abc_44228_n7233), .B(u2_o_396_), .Y(u2__abc_44228_n7234_1) );
  AND2X2 AND2X2_2495 ( .A(u2__abc_44228_n7236), .B(u2__abc_44228_n7230), .Y(u2__abc_44228_n7237) );
  AND2X2 AND2X2_2496 ( .A(u2__abc_44228_n7238), .B(u2_remHi_394_), .Y(u2__abc_44228_n7239) );
  AND2X2 AND2X2_2497 ( .A(u2__abc_44228_n7240), .B(u2_o_394_), .Y(u2__abc_44228_n7241) );
  AND2X2 AND2X2_2498 ( .A(u2__abc_44228_n7244_1), .B(u2_remHi_395_), .Y(u2__abc_44228_n7245) );
  AND2X2 AND2X2_2499 ( .A(u2__abc_44228_n7247), .B(u2_o_395_), .Y(u2__abc_44228_n7248) );
  AND2X2 AND2X2_25 ( .A(_abc_64468_n753_bF_buf3), .B(sqrto_24_), .Y(_auto_iopadmap_cc_313_execute_65414_60_) );
  AND2X2 AND2X2_250 ( .A(_abc_64468_n1348), .B(_abc_64468_n1347), .Y(fracta1_60_) );
  AND2X2 AND2X2_2500 ( .A(u2__abc_44228_n7246), .B(u2__abc_44228_n7249), .Y(u2__abc_44228_n7250) );
  AND2X2 AND2X2_2501 ( .A(u2__abc_44228_n7243), .B(u2__abc_44228_n7250), .Y(u2__abc_44228_n7251) );
  AND2X2 AND2X2_2502 ( .A(u2__abc_44228_n7237), .B(u2__abc_44228_n7251), .Y(u2__abc_44228_n7252_1) );
  AND2X2 AND2X2_2503 ( .A(u2__abc_44228_n7253), .B(u2_remHi_393_), .Y(u2__abc_44228_n7254) );
  AND2X2 AND2X2_2504 ( .A(u2__abc_44228_n7256), .B(u2_o_393_), .Y(u2__abc_44228_n7257) );
  AND2X2 AND2X2_2505 ( .A(u2__abc_44228_n7255), .B(u2__abc_44228_n7258), .Y(u2__abc_44228_n7259) );
  AND2X2 AND2X2_2506 ( .A(u2__abc_44228_n7260), .B(u2_remHi_392_), .Y(u2__abc_44228_n7261) );
  AND2X2 AND2X2_2507 ( .A(u2__abc_44228_n7262_1), .B(u2_o_392_), .Y(u2__abc_44228_n7263) );
  AND2X2 AND2X2_2508 ( .A(u2__abc_44228_n7265), .B(u2__abc_44228_n7259), .Y(u2__abc_44228_n7266) );
  AND2X2 AND2X2_2509 ( .A(u2__abc_44228_n7267), .B(u2_remHi_390_), .Y(u2__abc_44228_n7268) );
  AND2X2 AND2X2_251 ( .A(_abc_64468_n1351), .B(_abc_64468_n1350), .Y(fracta1_61_) );
  AND2X2 AND2X2_2510 ( .A(u2__abc_44228_n7269), .B(u2_o_390_), .Y(u2__abc_44228_n7270) );
  AND2X2 AND2X2_2511 ( .A(u2__abc_44228_n7273), .B(u2_remHi_391_), .Y(u2__abc_44228_n7274) );
  AND2X2 AND2X2_2512 ( .A(u2__abc_44228_n7276), .B(u2_o_391_), .Y(u2__abc_44228_n7277) );
  AND2X2 AND2X2_2513 ( .A(u2__abc_44228_n7275), .B(u2__abc_44228_n7278), .Y(u2__abc_44228_n7279) );
  AND2X2 AND2X2_2514 ( .A(u2__abc_44228_n7272), .B(u2__abc_44228_n7279), .Y(u2__abc_44228_n7280_1) );
  AND2X2 AND2X2_2515 ( .A(u2__abc_44228_n7266), .B(u2__abc_44228_n7280_1), .Y(u2__abc_44228_n7281) );
  AND2X2 AND2X2_2516 ( .A(u2__abc_44228_n7252_1), .B(u2__abc_44228_n7281), .Y(u2__abc_44228_n7282) );
  AND2X2 AND2X2_2517 ( .A(u2__abc_44228_n7283), .B(u2_remHi_389_), .Y(u2__abc_44228_n7284) );
  AND2X2 AND2X2_2518 ( .A(u2__abc_44228_n7286), .B(u2_o_389_), .Y(u2__abc_44228_n7287) );
  AND2X2 AND2X2_2519 ( .A(u2__abc_44228_n7285), .B(u2__abc_44228_n7288), .Y(u2__abc_44228_n7289_1) );
  AND2X2 AND2X2_252 ( .A(_abc_64468_n1354), .B(_abc_64468_n1353), .Y(fracta1_62_) );
  AND2X2 AND2X2_2520 ( .A(u2__abc_44228_n7290), .B(u2_remHi_388_), .Y(u2__abc_44228_n7291) );
  AND2X2 AND2X2_2521 ( .A(u2__abc_44228_n7292), .B(u2_o_388_), .Y(u2__abc_44228_n7293) );
  AND2X2 AND2X2_2522 ( .A(u2__abc_44228_n7295), .B(u2__abc_44228_n7289_1), .Y(u2__abc_44228_n7296) );
  AND2X2 AND2X2_2523 ( .A(u2__abc_44228_n7297), .B(u2_remHi_386_), .Y(u2__abc_44228_n7298) );
  AND2X2 AND2X2_2524 ( .A(u2__abc_44228_n7299_1), .B(u2_o_386_), .Y(u2__abc_44228_n7300) );
  AND2X2 AND2X2_2525 ( .A(u2__abc_44228_n7303), .B(u2_remHi_387_), .Y(u2__abc_44228_n7304) );
  AND2X2 AND2X2_2526 ( .A(u2__abc_44228_n7306), .B(u2_o_387_), .Y(u2__abc_44228_n7307) );
  AND2X2 AND2X2_2527 ( .A(u2__abc_44228_n7305), .B(u2__abc_44228_n7308), .Y(u2__abc_44228_n7309_1) );
  AND2X2 AND2X2_2528 ( .A(u2__abc_44228_n7302), .B(u2__abc_44228_n7309_1), .Y(u2__abc_44228_n7310) );
  AND2X2 AND2X2_2529 ( .A(u2__abc_44228_n7296), .B(u2__abc_44228_n7310), .Y(u2__abc_44228_n7311) );
  AND2X2 AND2X2_253 ( .A(_abc_64468_n1357), .B(_abc_64468_n1356), .Y(fracta1_63_) );
  AND2X2 AND2X2_2530 ( .A(u2__abc_44228_n7312), .B(u2_remHi_385_), .Y(u2__abc_44228_n7313) );
  AND2X2 AND2X2_2531 ( .A(u2__abc_44228_n7315), .B(u2_o_385_), .Y(u2__abc_44228_n7316) );
  AND2X2 AND2X2_2532 ( .A(u2__abc_44228_n7314), .B(u2__abc_44228_n7317), .Y(u2__abc_44228_n7318) );
  AND2X2 AND2X2_2533 ( .A(u2__abc_44228_n7319_1), .B(u2_remHi_384_), .Y(u2__abc_44228_n7320) );
  AND2X2 AND2X2_2534 ( .A(u2__abc_44228_n7321), .B(u2_o_384_), .Y(u2__abc_44228_n7322) );
  AND2X2 AND2X2_2535 ( .A(u2__abc_44228_n7324), .B(u2__abc_44228_n7318), .Y(u2__abc_44228_n7325) );
  AND2X2 AND2X2_2536 ( .A(u2__abc_44228_n7326), .B(u2_remHi_383_), .Y(u2__abc_44228_n7327_1) );
  AND2X2 AND2X2_2537 ( .A(u2__abc_44228_n7329), .B(u2_o_383_), .Y(u2__abc_44228_n7330) );
  AND2X2 AND2X2_2538 ( .A(u2__abc_44228_n7328), .B(u2__abc_44228_n7331), .Y(u2__abc_44228_n7332) );
  AND2X2 AND2X2_2539 ( .A(u2__abc_44228_n7333), .B(u2_remHi_382_), .Y(u2__abc_44228_n7334) );
  AND2X2 AND2X2_254 ( .A(_abc_64468_n1360), .B(_abc_64468_n1359), .Y(fracta1_64_) );
  AND2X2 AND2X2_2540 ( .A(u2__abc_44228_n7335), .B(u2_o_382_), .Y(u2__abc_44228_n7336) );
  AND2X2 AND2X2_2541 ( .A(u2__abc_44228_n7338), .B(u2__abc_44228_n7332), .Y(u2__abc_44228_n7339) );
  AND2X2 AND2X2_2542 ( .A(u2__abc_44228_n7325), .B(u2__abc_44228_n7339), .Y(u2__abc_44228_n7340) );
  AND2X2 AND2X2_2543 ( .A(u2__abc_44228_n7311), .B(u2__abc_44228_n7340), .Y(u2__abc_44228_n7341) );
  AND2X2 AND2X2_2544 ( .A(u2__abc_44228_n7282), .B(u2__abc_44228_n7341), .Y(u2__abc_44228_n7342) );
  AND2X2 AND2X2_2545 ( .A(u2__abc_44228_n7223), .B(u2__abc_44228_n7342), .Y(u2__abc_44228_n7343) );
  AND2X2 AND2X2_2546 ( .A(u2__abc_44228_n7104), .B(u2__abc_44228_n7343), .Y(u2__abc_44228_n7344) );
  AND2X2 AND2X2_2547 ( .A(u2__abc_44228_n6865), .B(u2__abc_44228_n7344), .Y(u2__abc_44228_n7345) );
  AND2X2 AND2X2_2548 ( .A(u2__abc_44228_n7347), .B(u2__abc_44228_n7328), .Y(u2__abc_44228_n7348) );
  AND2X2 AND2X2_2549 ( .A(u2__abc_44228_n7349), .B(u2__abc_44228_n7325), .Y(u2__abc_44228_n7350) );
  AND2X2 AND2X2_255 ( .A(_abc_64468_n1363), .B(_abc_64468_n1362), .Y(fracta1_65_) );
  AND2X2 AND2X2_2550 ( .A(u2__abc_44228_n7317), .B(u2__abc_44228_n7320), .Y(u2__abc_44228_n7351) );
  AND2X2 AND2X2_2551 ( .A(u2__abc_44228_n7353), .B(u2__abc_44228_n7311), .Y(u2__abc_44228_n7354) );
  AND2X2 AND2X2_2552 ( .A(u2__abc_44228_n7355_1), .B(u2__abc_44228_n7305), .Y(u2__abc_44228_n7356) );
  AND2X2 AND2X2_2553 ( .A(u2__abc_44228_n7357), .B(u2__abc_44228_n7308), .Y(u2__abc_44228_n7358) );
  AND2X2 AND2X2_2554 ( .A(u2__abc_44228_n7358), .B(u2__abc_44228_n7296), .Y(u2__abc_44228_n7359) );
  AND2X2 AND2X2_2555 ( .A(u2__abc_44228_n7288), .B(u2__abc_44228_n7291), .Y(u2__abc_44228_n7360) );
  AND2X2 AND2X2_2556 ( .A(u2__abc_44228_n7363), .B(u2__abc_44228_n7282), .Y(u2__abc_44228_n7364_1) );
  AND2X2 AND2X2_2557 ( .A(u2__abc_44228_n7365), .B(u2__abc_44228_n7275), .Y(u2__abc_44228_n7366) );
  AND2X2 AND2X2_2558 ( .A(u2__abc_44228_n7367), .B(u2__abc_44228_n7278), .Y(u2__abc_44228_n7368) );
  AND2X2 AND2X2_2559 ( .A(u2__abc_44228_n7368), .B(u2__abc_44228_n7266), .Y(u2__abc_44228_n7369) );
  AND2X2 AND2X2_256 ( .A(_abc_64468_n1366), .B(_abc_64468_n1365), .Y(fracta1_66_) );
  AND2X2 AND2X2_2560 ( .A(u2__abc_44228_n7258), .B(u2__abc_44228_n7261), .Y(u2__abc_44228_n7370) );
  AND2X2 AND2X2_2561 ( .A(u2__abc_44228_n7372), .B(u2__abc_44228_n7252_1), .Y(u2__abc_44228_n7373) );
  AND2X2 AND2X2_2562 ( .A(u2__abc_44228_n7229), .B(u2__abc_44228_n7232), .Y(u2__abc_44228_n7374_1) );
  AND2X2 AND2X2_2563 ( .A(u2__abc_44228_n7376), .B(u2__abc_44228_n7246), .Y(u2__abc_44228_n7377) );
  AND2X2 AND2X2_2564 ( .A(u2__abc_44228_n7378), .B(u2__abc_44228_n7249), .Y(u2__abc_44228_n7379) );
  AND2X2 AND2X2_2565 ( .A(u2__abc_44228_n7379), .B(u2__abc_44228_n7237), .Y(u2__abc_44228_n7380) );
  AND2X2 AND2X2_2566 ( .A(u2__abc_44228_n7383), .B(u2__abc_44228_n7223), .Y(u2__abc_44228_n7384) );
  AND2X2 AND2X2_2567 ( .A(u2__abc_44228_n7385), .B(u2__abc_44228_n7215_1), .Y(u2__abc_44228_n7386) );
  AND2X2 AND2X2_2568 ( .A(u2__abc_44228_n7387), .B(u2__abc_44228_n7218), .Y(u2__abc_44228_n7388) );
  AND2X2 AND2X2_2569 ( .A(u2__abc_44228_n7388), .B(u2__abc_44228_n7206_1), .Y(u2__abc_44228_n7389) );
  AND2X2 AND2X2_257 ( .A(_abc_64468_n1369), .B(_abc_64468_n1368), .Y(fracta1_67_) );
  AND2X2 AND2X2_2570 ( .A(u2__abc_44228_n7198), .B(u2__abc_44228_n7201), .Y(u2__abc_44228_n7390) );
  AND2X2 AND2X2_2571 ( .A(u2__abc_44228_n7392_1), .B(u2__abc_44228_n7192), .Y(u2__abc_44228_n7393) );
  AND2X2 AND2X2_2572 ( .A(u2__abc_44228_n7395), .B(u2__abc_44228_n7180), .Y(u2__abc_44228_n7396) );
  AND2X2 AND2X2_2573 ( .A(u2__abc_44228_n7397), .B(u2__abc_44228_n7177), .Y(u2__abc_44228_n7398) );
  AND2X2 AND2X2_2574 ( .A(u2__abc_44228_n7169), .B(u2__abc_44228_n7172), .Y(u2__abc_44228_n7399) );
  AND2X2 AND2X2_2575 ( .A(u2__abc_44228_n7402), .B(u2__abc_44228_n7163), .Y(u2__abc_44228_n7403) );
  AND2X2 AND2X2_2576 ( .A(u2__abc_44228_n7404), .B(u2__abc_44228_n7139), .Y(u2__abc_44228_n7405) );
  AND2X2 AND2X2_2577 ( .A(u2__abc_44228_n7150), .B(u2__abc_44228_n7406), .Y(u2__abc_44228_n7407) );
  AND2X2 AND2X2_2578 ( .A(u2__abc_44228_n7408), .B(u2__abc_44228_n7153_1), .Y(u2__abc_44228_n7409) );
  AND2X2 AND2X2_2579 ( .A(u2__abc_44228_n7409), .B(u2__abc_44228_n7147), .Y(u2__abc_44228_n7410_1) );
  AND2X2 AND2X2_258 ( .A(_abc_64468_n1372), .B(_abc_64468_n1371), .Y(fracta1_68_) );
  AND2X2 AND2X2_2580 ( .A(u2__abc_44228_n7411), .B(u2__abc_44228_n7133), .Y(u2__abc_44228_n7412) );
  AND2X2 AND2X2_2581 ( .A(u2__abc_44228_n7121), .B(u2__abc_44228_n7413), .Y(u2__abc_44228_n7414) );
  AND2X2 AND2X2_2582 ( .A(u2__abc_44228_n7415), .B(u2__abc_44228_n7124), .Y(u2__abc_44228_n7416) );
  AND2X2 AND2X2_2583 ( .A(u2__abc_44228_n7416), .B(u2__abc_44228_n7118), .Y(u2__abc_44228_n7417) );
  AND2X2 AND2X2_2584 ( .A(u2__abc_44228_n7110), .B(u2__abc_44228_n7113), .Y(u2__abc_44228_n7418) );
  AND2X2 AND2X2_2585 ( .A(u2__abc_44228_n7423), .B(u2__abc_44228_n7104), .Y(u2__abc_44228_n7424) );
  AND2X2 AND2X2_2586 ( .A(u2__abc_44228_n7425), .B(u2__abc_44228_n7095), .Y(u2__abc_44228_n7426) );
  AND2X2 AND2X2_2587 ( .A(u2__abc_44228_n7427), .B(u2__abc_44228_n7098_1), .Y(u2__abc_44228_n7428_1) );
  AND2X2 AND2X2_2588 ( .A(u2__abc_44228_n7428_1), .B(u2__abc_44228_n7086), .Y(u2__abc_44228_n7429) );
  AND2X2 AND2X2_2589 ( .A(u2__abc_44228_n7078_1), .B(u2__abc_44228_n7081), .Y(u2__abc_44228_n7430) );
  AND2X2 AND2X2_259 ( .A(_abc_64468_n1375), .B(_abc_64468_n1374), .Y(fracta1_69_) );
  AND2X2 AND2X2_2590 ( .A(u2__abc_44228_n7432), .B(u2__abc_44228_n7072), .Y(u2__abc_44228_n7433) );
  AND2X2 AND2X2_2591 ( .A(u2__abc_44228_n7435), .B(u2__abc_44228_n7060), .Y(u2__abc_44228_n7436) );
  AND2X2 AND2X2_2592 ( .A(u2__abc_44228_n7437_1), .B(u2__abc_44228_n7057), .Y(u2__abc_44228_n7438) );
  AND2X2 AND2X2_2593 ( .A(u2__abc_44228_n7049), .B(u2__abc_44228_n7052), .Y(u2__abc_44228_n7439) );
  AND2X2 AND2X2_2594 ( .A(u2__abc_44228_n7442), .B(u2__abc_44228_n7043), .Y(u2__abc_44228_n7443) );
  AND2X2 AND2X2_2595 ( .A(u2__abc_44228_n7445), .B(u2__abc_44228_n7030), .Y(u2__abc_44228_n7446) );
  AND2X2 AND2X2_2596 ( .A(u2__abc_44228_n7447_1), .B(u2__abc_44228_n7027), .Y(u2__abc_44228_n7448) );
  AND2X2 AND2X2_2597 ( .A(u2__abc_44228_n7016), .B(u2__abc_44228_n7449), .Y(u2__abc_44228_n7450) );
  AND2X2 AND2X2_2598 ( .A(u2__abc_44228_n7451), .B(u2__abc_44228_n7019), .Y(u2__abc_44228_n7452) );
  AND2X2 AND2X2_2599 ( .A(u2__abc_44228_n7453), .B(u2__abc_44228_n7013), .Y(u2__abc_44228_n7454) );
  AND2X2 AND2X2_26 ( .A(_abc_64468_n753_bF_buf2), .B(sqrto_25_), .Y(_auto_iopadmap_cc_313_execute_65414_61_) );
  AND2X2 AND2X2_260 ( .A(_abc_64468_n1378), .B(_abc_64468_n1377), .Y(fracta1_70_) );
  AND2X2 AND2X2_2600 ( .A(u2__abc_44228_n6990), .B(u2__abc_44228_n6993), .Y(u2__abc_44228_n7455_1) );
  AND2X2 AND2X2_2601 ( .A(u2__abc_44228_n7001), .B(u2__abc_44228_n7457), .Y(u2__abc_44228_n7458) );
  AND2X2 AND2X2_2602 ( .A(u2__abc_44228_n7459), .B(u2__abc_44228_n7004), .Y(u2__abc_44228_n7460) );
  AND2X2 AND2X2_2603 ( .A(u2__abc_44228_n7460), .B(u2__abc_44228_n6998), .Y(u2__abc_44228_n7461) );
  AND2X2 AND2X2_2604 ( .A(u2__abc_44228_n7464_1), .B(u2__abc_44228_n6984), .Y(u2__abc_44228_n7465) );
  AND2X2 AND2X2_2605 ( .A(u2__abc_44228_n7467), .B(u2__abc_44228_n6956), .Y(u2__abc_44228_n7468) );
  AND2X2 AND2X2_2606 ( .A(u2__abc_44228_n7469), .B(u2__abc_44228_n6981), .Y(u2__abc_44228_n7470) );
  AND2X2 AND2X2_2607 ( .A(u2__abc_44228_n6970), .B(u2__abc_44228_n7471), .Y(u2__abc_44228_n7472) );
  AND2X2 AND2X2_2608 ( .A(u2__abc_44228_n7473_1), .B(u2__abc_44228_n6973), .Y(u2__abc_44228_n7474) );
  AND2X2 AND2X2_2609 ( .A(u2__abc_44228_n7475), .B(u2__abc_44228_n6953_1), .Y(u2__abc_44228_n7476) );
  AND2X2 AND2X2_261 ( .A(_abc_64468_n1381), .B(_abc_64468_n1380), .Y(fracta1_71_) );
  AND2X2 AND2X2_2610 ( .A(u2__abc_44228_n7477), .B(u2__abc_44228_n6947), .Y(u2__abc_44228_n7478) );
  AND2X2 AND2X2_2611 ( .A(u2__abc_44228_n7479), .B(u2__abc_44228_n6950), .Y(u2__abc_44228_n7480) );
  AND2X2 AND2X2_2612 ( .A(u2__abc_44228_n7480), .B(u2__abc_44228_n6938), .Y(u2__abc_44228_n7481) );
  AND2X2 AND2X2_2613 ( .A(u2__abc_44228_n6930), .B(u2__abc_44228_n6933), .Y(u2__abc_44228_n7482) );
  AND2X2 AND2X2_2614 ( .A(u2__abc_44228_n7485), .B(u2__abc_44228_n6924_1), .Y(u2__abc_44228_n7486) );
  AND2X2 AND2X2_2615 ( .A(u2__abc_44228_n7487), .B(u2__abc_44228_n6900), .Y(u2__abc_44228_n7488) );
  AND2X2 AND2X2_2616 ( .A(u2__abc_44228_n6911), .B(u2__abc_44228_n7489), .Y(u2__abc_44228_n7490) );
  AND2X2 AND2X2_2617 ( .A(u2__abc_44228_n7491), .B(u2__abc_44228_n6914), .Y(u2__abc_44228_n7492) );
  AND2X2 AND2X2_2618 ( .A(u2__abc_44228_n7492), .B(u2__abc_44228_n6908), .Y(u2__abc_44228_n7493_1) );
  AND2X2 AND2X2_2619 ( .A(u2__abc_44228_n7494), .B(u2__abc_44228_n6894), .Y(u2__abc_44228_n7495) );
  AND2X2 AND2X2_262 ( .A(_abc_64468_n1384), .B(_abc_64468_n1383), .Y(fracta1_72_) );
  AND2X2 AND2X2_2620 ( .A(u2__abc_44228_n7497), .B(u2__abc_44228_n6882), .Y(u2__abc_44228_n7498) );
  AND2X2 AND2X2_2621 ( .A(u2__abc_44228_n7499), .B(u2__abc_44228_n6879), .Y(u2__abc_44228_n7500) );
  AND2X2 AND2X2_2622 ( .A(u2__abc_44228_n6871), .B(u2__abc_44228_n6874), .Y(u2__abc_44228_n7501) );
  AND2X2 AND2X2_2623 ( .A(u2__abc_44228_n7509), .B(u2_remHi_449_), .Y(u2__abc_44228_n7510) );
  AND2X2 AND2X2_2624 ( .A(u2__abc_44228_n7512), .B(u2_o_449_), .Y(u2__abc_44228_n7513) );
  AND2X2 AND2X2_2625 ( .A(u2__abc_44228_n7511_1), .B(u2__abc_44228_n7514), .Y(u2__abc_44228_n7515) );
  AND2X2 AND2X2_2626 ( .A(u2__abc_44228_n7516), .B(u2_remHi_448_), .Y(u2__abc_44228_n7517) );
  AND2X2 AND2X2_2627 ( .A(u2__abc_44228_n7518), .B(u2_o_448_), .Y(u2__abc_44228_n7519) );
  AND2X2 AND2X2_2628 ( .A(u2__abc_44228_n7521_1), .B(u2__abc_44228_n7515), .Y(u2__abc_44228_n7522) );
  AND2X2 AND2X2_2629 ( .A(u2__abc_44228_n7523), .B(u2_remHi_446_), .Y(u2__abc_44228_n7524) );
  AND2X2 AND2X2_263 ( .A(_abc_64468_n1387), .B(_abc_64468_n1386), .Y(fracta1_73_) );
  AND2X2 AND2X2_2630 ( .A(u2__abc_44228_n7525), .B(u2_o_446_), .Y(u2__abc_44228_n7526) );
  AND2X2 AND2X2_2631 ( .A(u2__abc_44228_n7529), .B(u2_remHi_447_), .Y(u2__abc_44228_n7530_1) );
  AND2X2 AND2X2_2632 ( .A(u2__abc_44228_n7532), .B(u2_o_447_), .Y(u2__abc_44228_n7533) );
  AND2X2 AND2X2_2633 ( .A(u2__abc_44228_n7531), .B(u2__abc_44228_n7534), .Y(u2__abc_44228_n7535) );
  AND2X2 AND2X2_2634 ( .A(u2__abc_44228_n7528), .B(u2__abc_44228_n7535), .Y(u2__abc_44228_n7536) );
  AND2X2 AND2X2_2635 ( .A(u2__abc_44228_n7522), .B(u2__abc_44228_n7536), .Y(u2__abc_44228_n7537) );
  AND2X2 AND2X2_2636 ( .A(u2__abc_44228_n7508), .B(u2__abc_44228_n7537), .Y(u2__abc_44228_n7538) );
  AND2X2 AND2X2_2637 ( .A(u2__abc_44228_n7539), .B(u2__abc_44228_n7531), .Y(u2__abc_44228_n7540_1) );
  AND2X2 AND2X2_2638 ( .A(u2__abc_44228_n7542), .B(u2__abc_44228_n7522), .Y(u2__abc_44228_n7543) );
  AND2X2 AND2X2_2639 ( .A(u2__abc_44228_n7514), .B(u2__abc_44228_n7517), .Y(u2__abc_44228_n7544) );
  AND2X2 AND2X2_264 ( .A(_abc_64468_n1390), .B(_abc_64468_n1389), .Y(fracta1_74_) );
  AND2X2 AND2X2_2640 ( .A(u2__abc_44228_n7548_1_bF_buf57), .B(u2_remHiShift_0_), .Y(u2__abc_44228_n7549) );
  AND2X2 AND2X2_2641 ( .A(u2__abc_44228_n7547_bF_buf56), .B(u2__abc_44228_n7550), .Y(u2__abc_44228_n7551) );
  AND2X2 AND2X2_2642 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n7554), .Y(u2__abc_44228_n7555) );
  AND2X2 AND2X2_2643 ( .A(u2__abc_44228_n7556), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n7557) );
  AND2X2 AND2X2_2644 ( .A(u2__abc_44228_n7553), .B(u2__abc_44228_n7557), .Y(u2__abc_44228_n7558_1) );
  AND2X2 AND2X2_2645 ( .A(u2__abc_44228_n7559), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_remHi_0__FF_INPUT) );
  AND2X2 AND2X2_2646 ( .A(u2__abc_44228_n3062_bF_buf91), .B(u2_remHi_1_), .Y(u2__abc_44228_n7561) );
  AND2X2 AND2X2_2647 ( .A(u2__abc_44228_n7562), .B(u2__abc_44228_n7563), .Y(u2__abc_44228_n7564) );
  AND2X2 AND2X2_2648 ( .A(u2__abc_44228_n7547_bF_buf55), .B(u2__abc_44228_n7564), .Y(u2__abc_44228_n7565) );
  AND2X2 AND2X2_2649 ( .A(u2__abc_44228_n7548_1_bF_buf56), .B(u2_remHiShift_1_), .Y(u2__abc_44228_n7566) );
  AND2X2 AND2X2_265 ( .A(_abc_64468_n1393), .B(_abc_64468_n1392), .Y(fracta1_75_) );
  AND2X2 AND2X2_2650 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n3072), .Y(u2__abc_44228_n7569) );
  AND2X2 AND2X2_2651 ( .A(u2__abc_44228_n7570), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n7571) );
  AND2X2 AND2X2_2652 ( .A(u2__abc_44228_n7568), .B(u2__abc_44228_n7571), .Y(u2__abc_44228_n7572) );
  AND2X2 AND2X2_2653 ( .A(u2__abc_44228_n7573), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_remHi_1__FF_INPUT) );
  AND2X2 AND2X2_2654 ( .A(u2__abc_44228_n3062_bF_buf90), .B(u2_remHi_2_), .Y(u2__abc_44228_n7575) );
  AND2X2 AND2X2_2655 ( .A(u2__abc_44228_n3071), .B(u2__abc_44228_n3081), .Y(u2__abc_44228_n7576_1) );
  AND2X2 AND2X2_2656 ( .A(u2__abc_44228_n7577), .B(u2__abc_44228_n7578), .Y(u2__abc_44228_n7579) );
  AND2X2 AND2X2_2657 ( .A(u2__abc_44228_n7547_bF_buf54), .B(u2__abc_44228_n7579), .Y(u2__abc_44228_n7580) );
  AND2X2 AND2X2_2658 ( .A(u2__abc_44228_n7548_1_bF_buf55), .B(u2_remHi_0_), .Y(u2__abc_44228_n7581) );
  AND2X2 AND2X2_2659 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n7584), .Y(u2__abc_44228_n7585) );
  AND2X2 AND2X2_266 ( .A(_abc_64468_n1396), .B(_abc_64468_n1395), .Y(fracta1_76_) );
  AND2X2 AND2X2_2660 ( .A(u2__abc_44228_n7586_1), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n7587) );
  AND2X2 AND2X2_2661 ( .A(u2__abc_44228_n7583), .B(u2__abc_44228_n7587), .Y(u2__abc_44228_n7588) );
  AND2X2 AND2X2_2662 ( .A(u2__abc_44228_n7589), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_remHi_2__FF_INPUT) );
  AND2X2 AND2X2_2663 ( .A(u2__abc_44228_n3062_bF_buf89), .B(u2_remHi_3_), .Y(u2__abc_44228_n7591) );
  AND2X2 AND2X2_2664 ( .A(u2__abc_44228_n7577), .B(u2__abc_44228_n3079), .Y(u2__abc_44228_n7592) );
  AND2X2 AND2X2_2665 ( .A(u2__abc_44228_n7594), .B(u2__abc_44228_n7596), .Y(u2__abc_44228_n7597_1) );
  AND2X2 AND2X2_2666 ( .A(u2__abc_44228_n7547_bF_buf53), .B(u2__abc_44228_n7597_1), .Y(u2__abc_44228_n7598) );
  AND2X2 AND2X2_2667 ( .A(u2__abc_44228_n7548_1_bF_buf54), .B(u2_remHi_1_), .Y(u2__abc_44228_n7599) );
  AND2X2 AND2X2_2668 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n7602), .Y(u2__abc_44228_n7603) );
  AND2X2 AND2X2_2669 ( .A(u2__abc_44228_n7604), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n7605_1) );
  AND2X2 AND2X2_267 ( .A(_abc_64468_n1399), .B(_abc_64468_n1398), .Y(fracta1_77_) );
  AND2X2 AND2X2_2670 ( .A(u2__abc_44228_n7601), .B(u2__abc_44228_n7605_1), .Y(u2__abc_44228_n7606) );
  AND2X2 AND2X2_2671 ( .A(u2__abc_44228_n7607), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_remHi_3__FF_INPUT) );
  AND2X2 AND2X2_2672 ( .A(u2__abc_44228_n3062_bF_buf88), .B(u2_remHi_4_), .Y(u2__abc_44228_n7609) );
  AND2X2 AND2X2_2673 ( .A(u2__abc_44228_n3087), .B(u2__abc_44228_n3108), .Y(u2__abc_44228_n7611) );
  AND2X2 AND2X2_2674 ( .A(u2__abc_44228_n7612), .B(u2__abc_44228_n7610), .Y(u2__abc_44228_n7613) );
  AND2X2 AND2X2_2675 ( .A(u2__abc_44228_n7547_bF_buf52), .B(u2__abc_44228_n7613), .Y(u2__abc_44228_n7614) );
  AND2X2 AND2X2_2676 ( .A(u2__abc_44228_n7548_1_bF_buf53), .B(u2_remHi_2_), .Y(u2__abc_44228_n7615_1) );
  AND2X2 AND2X2_2677 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n3093), .Y(u2__abc_44228_n7618) );
  AND2X2 AND2X2_2678 ( .A(u2__abc_44228_n7619), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n7620) );
  AND2X2 AND2X2_2679 ( .A(u2__abc_44228_n7617), .B(u2__abc_44228_n7620), .Y(u2__abc_44228_n7621) );
  AND2X2 AND2X2_268 ( .A(_abc_64468_n1402), .B(_abc_64468_n1401), .Y(fracta1_78_) );
  AND2X2 AND2X2_2680 ( .A(u2__abc_44228_n7622_1), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_remHi_4__FF_INPUT) );
  AND2X2 AND2X2_2681 ( .A(u2__abc_44228_n3062_bF_buf87), .B(u2_remHi_5_), .Y(u2__abc_44228_n7624) );
  AND2X2 AND2X2_2682 ( .A(u2__abc_44228_n7612), .B(u2__abc_44228_n3106), .Y(u2__abc_44228_n7626) );
  AND2X2 AND2X2_2683 ( .A(u2__abc_44228_n7629_1), .B(u2__abc_44228_n7627), .Y(u2__abc_44228_n7630_1) );
  AND2X2 AND2X2_2684 ( .A(u2__abc_44228_n7547_bF_buf51), .B(u2__abc_44228_n7630_1), .Y(u2__abc_44228_n7631) );
  AND2X2 AND2X2_2685 ( .A(u2__abc_44228_n7548_1_bF_buf52), .B(u2_remHi_3_), .Y(u2__abc_44228_n7632) );
  AND2X2 AND2X2_2686 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n3088), .Y(u2__abc_44228_n7635) );
  AND2X2 AND2X2_2687 ( .A(u2__abc_44228_n7636_1), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n7637_1) );
  AND2X2 AND2X2_2688 ( .A(u2__abc_44228_n7634), .B(u2__abc_44228_n7637_1), .Y(u2__abc_44228_n7638) );
  AND2X2 AND2X2_2689 ( .A(u2__abc_44228_n7639), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_remHi_5__FF_INPUT) );
  AND2X2 AND2X2_269 ( .A(_abc_64468_n1405), .B(_abc_64468_n1404), .Y(fracta1_79_) );
  AND2X2 AND2X2_2690 ( .A(u2__abc_44228_n3062_bF_buf86), .B(u2_remHi_6_), .Y(u2__abc_44228_n7641) );
  AND2X2 AND2X2_2691 ( .A(u2__abc_44228_n3087), .B(u2__abc_44228_n3109), .Y(u2__abc_44228_n7642) );
  AND2X2 AND2X2_2692 ( .A(u2__abc_44228_n7643_1), .B(u2__abc_44228_n3097), .Y(u2__abc_44228_n7644_1) );
  AND2X2 AND2X2_2693 ( .A(u2__abc_44228_n7645), .B(u2__abc_44228_n7646), .Y(u2__abc_44228_n7647) );
  AND2X2 AND2X2_2694 ( .A(u2__abc_44228_n7547_bF_buf50), .B(u2__abc_44228_n7647), .Y(u2__abc_44228_n7648) );
  AND2X2 AND2X2_2695 ( .A(u2__abc_44228_n7548_1_bF_buf51), .B(u2_remHi_4_), .Y(u2__abc_44228_n7649) );
  AND2X2 AND2X2_2696 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n3163), .Y(u2__abc_44228_n7652) );
  AND2X2 AND2X2_2697 ( .A(u2__abc_44228_n7653), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n7654) );
  AND2X2 AND2X2_2698 ( .A(u2__abc_44228_n7651_1), .B(u2__abc_44228_n7654), .Y(u2__abc_44228_n7655) );
  AND2X2 AND2X2_2699 ( .A(u2__abc_44228_n7656), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_remHi_6__FF_INPUT) );
  AND2X2 AND2X2_27 ( .A(_abc_64468_n753_bF_buf1), .B(sqrto_26_), .Y(_auto_iopadmap_cc_313_execute_65414_62_) );
  AND2X2 AND2X2_270 ( .A(_abc_64468_n1408), .B(_abc_64468_n1407), .Y(fracta1_80_) );
  AND2X2 AND2X2_2700 ( .A(u2__abc_44228_n3062_bF_buf85), .B(u2_remHi_7_), .Y(u2__abc_44228_n7658_1) );
  AND2X2 AND2X2_2701 ( .A(u2__abc_44228_n7645), .B(u2__abc_44228_n3094), .Y(u2__abc_44228_n7659) );
  AND2X2 AND2X2_2702 ( .A(u2__abc_44228_n7661), .B(u2__abc_44228_n7663), .Y(u2__abc_44228_n7664_1) );
  AND2X2 AND2X2_2703 ( .A(u2__abc_44228_n7547_bF_buf49), .B(u2__abc_44228_n7664_1), .Y(u2__abc_44228_n7665_1) );
  AND2X2 AND2X2_2704 ( .A(u2__abc_44228_n7548_1_bF_buf50), .B(u2_remHi_5_), .Y(u2__abc_44228_n7666) );
  AND2X2 AND2X2_2705 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n3170), .Y(u2__abc_44228_n7669) );
  AND2X2 AND2X2_2706 ( .A(u2__abc_44228_n7670), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n7671_1) );
  AND2X2 AND2X2_2707 ( .A(u2__abc_44228_n7668), .B(u2__abc_44228_n7671_1), .Y(u2__abc_44228_n7672_1) );
  AND2X2 AND2X2_2708 ( .A(u2__abc_44228_n7673), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_remHi_7__FF_INPUT) );
  AND2X2 AND2X2_2709 ( .A(u2__abc_44228_n3062_bF_buf84), .B(u2_remHi_8_), .Y(u2__abc_44228_n7675) );
  AND2X2 AND2X2_271 ( .A(_abc_64468_n1411), .B(_abc_64468_n1410), .Y(fracta1_81_) );
  AND2X2 AND2X2_2710 ( .A(u2__abc_44228_n3120), .B(u2__abc_44228_n3166), .Y(u2__abc_44228_n7676) );
  AND2X2 AND2X2_2711 ( .A(u2__abc_44228_n7677), .B(u2__abc_44228_n7678_1), .Y(u2__abc_44228_n7679_1) );
  AND2X2 AND2X2_2712 ( .A(u2__abc_44228_n7547_bF_buf48), .B(u2__abc_44228_n7679_1), .Y(u2__abc_44228_n7680) );
  AND2X2 AND2X2_2713 ( .A(u2__abc_44228_n7548_1_bF_buf49), .B(u2_remHi_6_), .Y(u2__abc_44228_n7681) );
  AND2X2 AND2X2_2714 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n3155), .Y(u2__abc_44228_n7684) );
  AND2X2 AND2X2_2715 ( .A(u2__abc_44228_n7685_1), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n7686_1) );
  AND2X2 AND2X2_2716 ( .A(u2__abc_44228_n7683), .B(u2__abc_44228_n7686_1), .Y(u2__abc_44228_n7687) );
  AND2X2 AND2X2_2717 ( .A(u2__abc_44228_n7688), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_remHi_8__FF_INPUT) );
  AND2X2 AND2X2_2718 ( .A(u2__abc_44228_n3062_bF_buf83), .B(u2_remHi_9_), .Y(u2__abc_44228_n7690) );
  AND2X2 AND2X2_2719 ( .A(u2__abc_44228_n7692_1), .B(u2__abc_44228_n7691), .Y(u2__abc_44228_n7693_1) );
  AND2X2 AND2X2_272 ( .A(_abc_64468_n1414), .B(_abc_64468_n1413), .Y(fracta1_82_) );
  AND2X2 AND2X2_2720 ( .A(u2__abc_44228_n7694), .B(u2__abc_44228_n3173), .Y(u2__abc_44228_n7695) );
  AND2X2 AND2X2_2721 ( .A(u2__abc_44228_n7547_bF_buf47), .B(u2__abc_44228_n7696), .Y(u2__abc_44228_n7697) );
  AND2X2 AND2X2_2722 ( .A(u2__abc_44228_n7548_1_bF_buf48), .B(u2_remHi_7_), .Y(u2__abc_44228_n7698) );
  AND2X2 AND2X2_2723 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n3150), .Y(u2__abc_44228_n7701) );
  AND2X2 AND2X2_2724 ( .A(u2__abc_44228_n7702), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n7703) );
  AND2X2 AND2X2_2725 ( .A(u2__abc_44228_n7700_1), .B(u2__abc_44228_n7703), .Y(u2__abc_44228_n7704) );
  AND2X2 AND2X2_2726 ( .A(u2__abc_44228_n7705), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_remHi_9__FF_INPUT) );
  AND2X2 AND2X2_2727 ( .A(u2__abc_44228_n3062_bF_buf82), .B(u2_remHi_10_), .Y(u2__abc_44228_n7707_1) );
  AND2X2 AND2X2_2728 ( .A(u2__abc_44228_n3120), .B(u2__abc_44228_n3174), .Y(u2__abc_44228_n7708) );
  AND2X2 AND2X2_2729 ( .A(u2__abc_44228_n7709), .B(u2__abc_44228_n3159), .Y(u2__abc_44228_n7711) );
  AND2X2 AND2X2_273 ( .A(_abc_64468_n1417), .B(_abc_64468_n1416), .Y(fracta1_83_) );
  AND2X2 AND2X2_2730 ( .A(u2__abc_44228_n7712), .B(u2__abc_44228_n7710), .Y(u2__abc_44228_n7713_1) );
  AND2X2 AND2X2_2731 ( .A(u2__abc_44228_n7547_bF_buf46), .B(u2__abc_44228_n7713_1), .Y(u2__abc_44228_n7714_1) );
  AND2X2 AND2X2_2732 ( .A(u2__abc_44228_n7548_1_bF_buf47), .B(u2_remHi_8_), .Y(u2__abc_44228_n7715) );
  AND2X2 AND2X2_2733 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n3144), .Y(u2__abc_44228_n7718) );
  AND2X2 AND2X2_2734 ( .A(u2__abc_44228_n7719), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n7720_1) );
  AND2X2 AND2X2_2735 ( .A(u2__abc_44228_n7717), .B(u2__abc_44228_n7720_1), .Y(u2__abc_44228_n7721_1) );
  AND2X2 AND2X2_2736 ( .A(u2__abc_44228_n7722), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_remHi_10__FF_INPUT) );
  AND2X2 AND2X2_2737 ( .A(u2__abc_44228_n3062_bF_buf81), .B(u2_remHi_11_), .Y(u2__abc_44228_n7724) );
  AND2X2 AND2X2_2738 ( .A(u2__abc_44228_n7712), .B(u2__abc_44228_n3156), .Y(u2__abc_44228_n7725) );
  AND2X2 AND2X2_2739 ( .A(u2__abc_44228_n7727_1), .B(u2__abc_44228_n7729), .Y(u2__abc_44228_n7730) );
  AND2X2 AND2X2_274 ( .A(_abc_64468_n1420), .B(_abc_64468_n1419), .Y(fracta1_84_) );
  AND2X2 AND2X2_2740 ( .A(u2__abc_44228_n7547_bF_buf45), .B(u2__abc_44228_n7730), .Y(u2__abc_44228_n7731) );
  AND2X2 AND2X2_2741 ( .A(u2__abc_44228_n7548_1_bF_buf46), .B(u2_remHi_9_), .Y(u2__abc_44228_n7732) );
  AND2X2 AND2X2_2742 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n3138), .Y(u2__abc_44228_n7735_1) );
  AND2X2 AND2X2_2743 ( .A(u2__abc_44228_n7736), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n7737) );
  AND2X2 AND2X2_2744 ( .A(u2__abc_44228_n7734_1), .B(u2__abc_44228_n7737), .Y(u2__abc_44228_n7738) );
  AND2X2 AND2X2_2745 ( .A(u2__abc_44228_n7739), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_remHi_11__FF_INPUT) );
  AND2X2 AND2X2_2746 ( .A(u2__abc_44228_n3062_bF_buf80), .B(u2_remHi_12_), .Y(u2__abc_44228_n7741_1) );
  AND2X2 AND2X2_2747 ( .A(u2__abc_44228_n3120), .B(u2__abc_44228_n3175), .Y(u2__abc_44228_n7742_1) );
  AND2X2 AND2X2_2748 ( .A(u2__abc_44228_n7743), .B(u2__abc_44228_n3147), .Y(u2__abc_44228_n7744) );
  AND2X2 AND2X2_2749 ( .A(u2__abc_44228_n7745), .B(u2__abc_44228_n7746), .Y(u2__abc_44228_n7747) );
  AND2X2 AND2X2_275 ( .A(_abc_64468_n1423), .B(_abc_64468_n1422), .Y(fracta1_85_) );
  AND2X2 AND2X2_2750 ( .A(u2__abc_44228_n7547_bF_buf44), .B(u2__abc_44228_n7747), .Y(u2__abc_44228_n7748_1) );
  AND2X2 AND2X2_2751 ( .A(u2__abc_44228_n7548_1_bF_buf45), .B(u2_remHi_10_), .Y(u2__abc_44228_n7749_1) );
  AND2X2 AND2X2_2752 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n3130), .Y(u2__abc_44228_n7752) );
  AND2X2 AND2X2_2753 ( .A(u2__abc_44228_n7753), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n7754) );
  AND2X2 AND2X2_2754 ( .A(u2__abc_44228_n7751), .B(u2__abc_44228_n7754), .Y(u2__abc_44228_n7755_1) );
  AND2X2 AND2X2_2755 ( .A(u2__abc_44228_n7756_1), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_remHi_12__FF_INPUT) );
  AND2X2 AND2X2_2756 ( .A(u2__abc_44228_n3062_bF_buf79), .B(u2_remHi_13_), .Y(u2__abc_44228_n7758) );
  AND2X2 AND2X2_2757 ( .A(u2__abc_44228_n7763_1), .B(u2__abc_44228_n7760), .Y(u2__abc_44228_n7764) );
  AND2X2 AND2X2_2758 ( .A(u2__abc_44228_n7547_bF_buf43), .B(u2__abc_44228_n7764), .Y(u2__abc_44228_n7765) );
  AND2X2 AND2X2_2759 ( .A(u2__abc_44228_n7548_1_bF_buf44), .B(u2_remHi_11_), .Y(u2__abc_44228_n7766) );
  AND2X2 AND2X2_276 ( .A(_abc_64468_n1426), .B(_abc_64468_n1425), .Y(fracta1_86_) );
  AND2X2 AND2X2_2760 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n3124), .Y(u2__abc_44228_n7769_1) );
  AND2X2 AND2X2_2761 ( .A(u2__abc_44228_n7770_1), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n7771) );
  AND2X2 AND2X2_2762 ( .A(u2__abc_44228_n7768), .B(u2__abc_44228_n7771), .Y(u2__abc_44228_n7772) );
  AND2X2 AND2X2_2763 ( .A(u2__abc_44228_n7773), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_remHi_13__FF_INPUT) );
  AND2X2 AND2X2_2764 ( .A(u2__abc_44228_n3062_bF_buf78), .B(u2_remHi_14_), .Y(u2__abc_44228_n7775) );
  AND2X2 AND2X2_2765 ( .A(u2__abc_44228_n7743), .B(u2__abc_44228_n3148), .Y(u2__abc_44228_n7776_1) );
  AND2X2 AND2X2_2766 ( .A(u2__abc_44228_n7777_1), .B(u2__abc_44228_n3133), .Y(u2__abc_44228_n7779) );
  AND2X2 AND2X2_2767 ( .A(u2__abc_44228_n7780), .B(u2__abc_44228_n7778), .Y(u2__abc_44228_n7781) );
  AND2X2 AND2X2_2768 ( .A(u2__abc_44228_n7547_bF_buf42), .B(u2__abc_44228_n7781), .Y(u2__abc_44228_n7782) );
  AND2X2 AND2X2_2769 ( .A(u2__abc_44228_n7548_1_bF_buf43), .B(u2_remHi_12_), .Y(u2__abc_44228_n7783_1) );
  AND2X2 AND2X2_277 ( .A(_abc_64468_n1429), .B(_abc_64468_n1428), .Y(fracta1_87_) );
  AND2X2 AND2X2_2770 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n3303), .Y(u2__abc_44228_n7786) );
  AND2X2 AND2X2_2771 ( .A(u2__abc_44228_n7787), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n7788) );
  AND2X2 AND2X2_2772 ( .A(u2__abc_44228_n7785), .B(u2__abc_44228_n7788), .Y(u2__abc_44228_n7789) );
  AND2X2 AND2X2_2773 ( .A(u2__abc_44228_n7790_1), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_remHi_14__FF_INPUT) );
  AND2X2 AND2X2_2774 ( .A(u2__abc_44228_n3062_bF_buf77), .B(u2_remHi_15_), .Y(u2__abc_44228_n7792) );
  AND2X2 AND2X2_2775 ( .A(u2__abc_44228_n7796), .B(u2__abc_44228_n7797_1), .Y(u2__abc_44228_n7798_1) );
  AND2X2 AND2X2_2776 ( .A(u2__abc_44228_n7547_bF_buf41), .B(u2__abc_44228_n7798_1), .Y(u2__abc_44228_n7799) );
  AND2X2 AND2X2_2777 ( .A(u2__abc_44228_n7548_1_bF_buf42), .B(u2_remHi_13_), .Y(u2__abc_44228_n7800) );
  AND2X2 AND2X2_2778 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n3297), .Y(u2__abc_44228_n7803) );
  AND2X2 AND2X2_2779 ( .A(u2__abc_44228_n7804_1), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n7805_1) );
  AND2X2 AND2X2_278 ( .A(_abc_64468_n1432), .B(_abc_64468_n1431), .Y(fracta1_88_) );
  AND2X2 AND2X2_2780 ( .A(u2__abc_44228_n7802), .B(u2__abc_44228_n7805_1), .Y(u2__abc_44228_n7806) );
  AND2X2 AND2X2_2781 ( .A(u2__abc_44228_n7807), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_remHi_15__FF_INPUT) );
  AND2X2 AND2X2_2782 ( .A(u2__abc_44228_n3062_bF_buf76), .B(u2_remHi_16_), .Y(u2__abc_44228_n7809) );
  AND2X2 AND2X2_2783 ( .A(u2__abc_44228_n3194), .B(u2__abc_44228_n3306), .Y(u2__abc_44228_n7811_1) );
  AND2X2 AND2X2_2784 ( .A(u2__abc_44228_n7812_1), .B(u2__abc_44228_n7810), .Y(u2__abc_44228_n7813) );
  AND2X2 AND2X2_2785 ( .A(u2__abc_44228_n7547_bF_buf40), .B(u2__abc_44228_n7813), .Y(u2__abc_44228_n7814) );
  AND2X2 AND2X2_2786 ( .A(u2__abc_44228_n7548_1_bF_buf41), .B(u2_remHi_14_), .Y(u2__abc_44228_n7815) );
  AND2X2 AND2X2_2787 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n3288), .Y(u2__abc_44228_n7818_1) );
  AND2X2 AND2X2_2788 ( .A(u2__abc_44228_n7819_1), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n7820) );
  AND2X2 AND2X2_2789 ( .A(u2__abc_44228_n7817), .B(u2__abc_44228_n7820), .Y(u2__abc_44228_n7821) );
  AND2X2 AND2X2_279 ( .A(_abc_64468_n1435), .B(_abc_64468_n1434), .Y(fracta1_89_) );
  AND2X2 AND2X2_2790 ( .A(u2__abc_44228_n7822), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_remHi_16__FF_INPUT) );
  AND2X2 AND2X2_2791 ( .A(u2__abc_44228_n3062_bF_buf75), .B(u2_remHi_17_), .Y(u2__abc_44228_n7824) );
  AND2X2 AND2X2_2792 ( .A(u2__abc_44228_n7829), .B(u2__abc_44228_n7826_1), .Y(u2__abc_44228_n7830) );
  AND2X2 AND2X2_2793 ( .A(u2__abc_44228_n7547_bF_buf39), .B(u2__abc_44228_n7830), .Y(u2__abc_44228_n7831) );
  AND2X2 AND2X2_2794 ( .A(u2__abc_44228_n7548_1_bF_buf40), .B(u2_remHi_15_), .Y(u2__abc_44228_n7832_1) );
  AND2X2 AND2X2_2795 ( .A(u2__abc_44228_n2983_bF_buf104), .B(u2__abc_44228_n3283), .Y(u2__abc_44228_n7835) );
  AND2X2 AND2X2_2796 ( .A(u2__abc_44228_n7836), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n7837) );
  AND2X2 AND2X2_2797 ( .A(u2__abc_44228_n7834), .B(u2__abc_44228_n7837), .Y(u2__abc_44228_n7838) );
  AND2X2 AND2X2_2798 ( .A(u2__abc_44228_n7839_1), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_remHi_17__FF_INPUT) );
  AND2X2 AND2X2_2799 ( .A(u2__abc_44228_n3062_bF_buf74), .B(u2_remHi_18_), .Y(u2__abc_44228_n7841) );
  AND2X2 AND2X2_28 ( .A(_abc_64468_n753_bF_buf0), .B(sqrto_27_), .Y(_auto_iopadmap_cc_313_execute_65414_63_) );
  AND2X2 AND2X2_280 ( .A(_abc_64468_n1438), .B(_abc_64468_n1437), .Y(fracta1_90_) );
  AND2X2 AND2X2_2800 ( .A(u2__abc_44228_n3194), .B(u2__abc_44228_n3307), .Y(u2__abc_44228_n7842) );
  AND2X2 AND2X2_2801 ( .A(u2__abc_44228_n7843), .B(u2__abc_44228_n3292), .Y(u2__abc_44228_n7845_1) );
  AND2X2 AND2X2_2802 ( .A(u2__abc_44228_n7846), .B(u2__abc_44228_n7844), .Y(u2__abc_44228_n7847) );
  AND2X2 AND2X2_2803 ( .A(u2__abc_44228_n7547_bF_buf38), .B(u2__abc_44228_n7847), .Y(u2__abc_44228_n7848) );
  AND2X2 AND2X2_2804 ( .A(u2__abc_44228_n7548_1_bF_buf39), .B(u2_remHi_16_), .Y(u2__abc_44228_n7849) );
  AND2X2 AND2X2_2805 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n3270), .Y(u2__abc_44228_n7852) );
  AND2X2 AND2X2_2806 ( .A(u2__abc_44228_n7853), .B(u2__abc_44228_n2972_bF_buf87), .Y(u2__abc_44228_n7854) );
  AND2X2 AND2X2_2807 ( .A(u2__abc_44228_n7851_1), .B(u2__abc_44228_n7854), .Y(u2__abc_44228_n7855) );
  AND2X2 AND2X2_2808 ( .A(u2__abc_44228_n7856_1), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_remHi_18__FF_INPUT) );
  AND2X2 AND2X2_2809 ( .A(u2__abc_44228_n3062_bF_buf73), .B(u2_remHi_19_), .Y(u2__abc_44228_n7858) );
  AND2X2 AND2X2_281 ( .A(_abc_64468_n1441), .B(_abc_64468_n1440), .Y(fracta1_91_) );
  AND2X2 AND2X2_2810 ( .A(u2__abc_44228_n7846), .B(u2__abc_44228_n3289), .Y(u2__abc_44228_n7859) );
  AND2X2 AND2X2_2811 ( .A(u2__abc_44228_n7861_1), .B(u2__abc_44228_n7863), .Y(u2__abc_44228_n7864) );
  AND2X2 AND2X2_2812 ( .A(u2__abc_44228_n7547_bF_buf37), .B(u2__abc_44228_n7864), .Y(u2__abc_44228_n7865) );
  AND2X2 AND2X2_2813 ( .A(u2__abc_44228_n7548_1_bF_buf38), .B(u2_remHi_17_), .Y(u2__abc_44228_n7866) );
  AND2X2 AND2X2_2814 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n3277), .Y(u2__abc_44228_n7869) );
  AND2X2 AND2X2_2815 ( .A(u2__abc_44228_n7870), .B(u2__abc_44228_n2972_bF_buf86), .Y(u2__abc_44228_n7871) );
  AND2X2 AND2X2_2816 ( .A(u2__abc_44228_n7868), .B(u2__abc_44228_n7871), .Y(u2__abc_44228_n7872_1) );
  AND2X2 AND2X2_2817 ( .A(u2__abc_44228_n7873_1), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_remHi_19__FF_INPUT) );
  AND2X2 AND2X2_2818 ( .A(u2__abc_44228_n3062_bF_buf72), .B(u2_remHi_20_), .Y(u2__abc_44228_n7875) );
  AND2X2 AND2X2_2819 ( .A(u2__abc_44228_n3194), .B(u2__abc_44228_n3308), .Y(u2__abc_44228_n7876) );
  AND2X2 AND2X2_282 ( .A(_abc_64468_n1444), .B(_abc_64468_n1443), .Y(fracta1_92_) );
  AND2X2 AND2X2_2820 ( .A(u2__abc_44228_n7877), .B(u2__abc_44228_n3273), .Y(u2__abc_44228_n7878_1) );
  AND2X2 AND2X2_2821 ( .A(u2__abc_44228_n7879), .B(u2__abc_44228_n7880), .Y(u2__abc_44228_n7881) );
  AND2X2 AND2X2_2822 ( .A(u2__abc_44228_n7547_bF_buf36), .B(u2__abc_44228_n7881), .Y(u2__abc_44228_n7882) );
  AND2X2 AND2X2_2823 ( .A(u2__abc_44228_n7548_1_bF_buf37), .B(u2_remHi_18_), .Y(u2__abc_44228_n7883_1) );
  AND2X2 AND2X2_2824 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n3263), .Y(u2__abc_44228_n7886) );
  AND2X2 AND2X2_2825 ( .A(u2__abc_44228_n7887), .B(u2__abc_44228_n2972_bF_buf85), .Y(u2__abc_44228_n7888) );
  AND2X2 AND2X2_2826 ( .A(u2__abc_44228_n7885), .B(u2__abc_44228_n7888), .Y(u2__abc_44228_n7889_1) );
  AND2X2 AND2X2_2827 ( .A(u2__abc_44228_n7890), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_remHi_20__FF_INPUT) );
  AND2X2 AND2X2_2828 ( .A(u2__abc_44228_n3062_bF_buf71), .B(u2_remHi_21_), .Y(u2__abc_44228_n7892) );
  AND2X2 AND2X2_2829 ( .A(u2__abc_44228_n7894_1), .B(u2__abc_44228_n7893), .Y(u2__abc_44228_n7895_1) );
  AND2X2 AND2X2_283 ( .A(_abc_64468_n1447), .B(_abc_64468_n1446), .Y(fracta1_93_) );
  AND2X2 AND2X2_2830 ( .A(u2__abc_44228_n7896), .B(u2__abc_44228_n3280), .Y(u2__abc_44228_n7897) );
  AND2X2 AND2X2_2831 ( .A(u2__abc_44228_n7547_bF_buf35), .B(u2__abc_44228_n7898), .Y(u2__abc_44228_n7899) );
  AND2X2 AND2X2_2832 ( .A(u2__abc_44228_n7548_1_bF_buf36), .B(u2_remHi_19_), .Y(u2__abc_44228_n7900_1) );
  AND2X2 AND2X2_2833 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n3257), .Y(u2__abc_44228_n7903) );
  AND2X2 AND2X2_2834 ( .A(u2__abc_44228_n7904), .B(u2__abc_44228_n2972_bF_buf84), .Y(u2__abc_44228_n7905_1) );
  AND2X2 AND2X2_2835 ( .A(u2__abc_44228_n7902), .B(u2__abc_44228_n7905_1), .Y(u2__abc_44228_n7906_1) );
  AND2X2 AND2X2_2836 ( .A(u2__abc_44228_n7907), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_remHi_21__FF_INPUT) );
  AND2X2 AND2X2_2837 ( .A(u2__abc_44228_n3062_bF_buf70), .B(u2_remHi_22_), .Y(u2__abc_44228_n7909) );
  AND2X2 AND2X2_2838 ( .A(u2__abc_44228_n7877), .B(u2__abc_44228_n3281), .Y(u2__abc_44228_n7910) );
  AND2X2 AND2X2_2839 ( .A(u2__abc_44228_n7911_1), .B(u2__abc_44228_n3266), .Y(u2__abc_44228_n7913) );
  AND2X2 AND2X2_284 ( .A(_abc_64468_n1450), .B(_abc_64468_n1449), .Y(fracta1_94_) );
  AND2X2 AND2X2_2840 ( .A(u2__abc_44228_n7914), .B(u2__abc_44228_n7912), .Y(u2__abc_44228_n7915) );
  AND2X2 AND2X2_2841 ( .A(u2__abc_44228_n7547_bF_buf34), .B(u2__abc_44228_n7915), .Y(u2__abc_44228_n7916_1) );
  AND2X2 AND2X2_2842 ( .A(u2__abc_44228_n7548_1_bF_buf35), .B(u2_remHi_20_), .Y(u2__abc_44228_n7917_1) );
  AND2X2 AND2X2_2843 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n3233), .Y(u2__abc_44228_n7920) );
  AND2X2 AND2X2_2844 ( .A(u2__abc_44228_n7921), .B(u2__abc_44228_n2972_bF_buf83), .Y(u2__abc_44228_n7922_1) );
  AND2X2 AND2X2_2845 ( .A(u2__abc_44228_n7919), .B(u2__abc_44228_n7922_1), .Y(u2__abc_44228_n7923) );
  AND2X2 AND2X2_2846 ( .A(u2__abc_44228_n7924), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_remHi_22__FF_INPUT) );
  AND2X2 AND2X2_2847 ( .A(u2__abc_44228_n3062_bF_buf69), .B(u2_remHi_23_), .Y(u2__abc_44228_n7926) );
  AND2X2 AND2X2_2848 ( .A(u2__abc_44228_n7928_1), .B(u2__abc_44228_n7927_1), .Y(u2__abc_44228_n7929) );
  AND2X2 AND2X2_2849 ( .A(u2__abc_44228_n7930), .B(u2__abc_44228_n3260), .Y(u2__abc_44228_n7931) );
  AND2X2 AND2X2_285 ( .A(_abc_64468_n1453), .B(_abc_64468_n1452), .Y(fracta1_95_) );
  AND2X2 AND2X2_2850 ( .A(u2__abc_44228_n7547_bF_buf33), .B(u2__abc_44228_n7932), .Y(u2__abc_44228_n7933_1) );
  AND2X2 AND2X2_2851 ( .A(u2__abc_44228_n7548_1_bF_buf34), .B(u2_remHi_21_), .Y(u2__abc_44228_n7934) );
  AND2X2 AND2X2_2852 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n3227), .Y(u2__abc_44228_n7937) );
  AND2X2 AND2X2_2853 ( .A(u2__abc_44228_n7938_1), .B(u2__abc_44228_n2972_bF_buf82), .Y(u2__abc_44228_n7939_1) );
  AND2X2 AND2X2_2854 ( .A(u2__abc_44228_n7936), .B(u2__abc_44228_n7939_1), .Y(u2__abc_44228_n7940) );
  AND2X2 AND2X2_2855 ( .A(u2__abc_44228_n7941), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_remHi_23__FF_INPUT) );
  AND2X2 AND2X2_2856 ( .A(u2__abc_44228_n3062_bF_buf68), .B(u2_remHi_24_), .Y(u2__abc_44228_n7943) );
  AND2X2 AND2X2_2857 ( .A(u2__abc_44228_n3194), .B(u2__abc_44228_n3309), .Y(u2__abc_44228_n7944_1) );
  AND2X2 AND2X2_2858 ( .A(u2__abc_44228_n7945), .B(u2__abc_44228_n3236), .Y(u2__abc_44228_n7947) );
  AND2X2 AND2X2_2859 ( .A(u2__abc_44228_n7948), .B(u2__abc_44228_n7946), .Y(u2__abc_44228_n7949_1) );
  AND2X2 AND2X2_286 ( .A(_abc_64468_n1456), .B(_abc_64468_n1455), .Y(fracta1_96_) );
  AND2X2 AND2X2_2860 ( .A(u2__abc_44228_n7547_bF_buf32), .B(u2__abc_44228_n7949_1), .Y(u2__abc_44228_n7950_1) );
  AND2X2 AND2X2_2861 ( .A(u2__abc_44228_n7548_1_bF_buf33), .B(u2_remHi_22_), .Y(u2__abc_44228_n7951) );
  AND2X2 AND2X2_2862 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n3247), .Y(u2__abc_44228_n7954) );
  AND2X2 AND2X2_2863 ( .A(u2__abc_44228_n7955_1), .B(u2__abc_44228_n2972_bF_buf81), .Y(u2__abc_44228_n7956) );
  AND2X2 AND2X2_2864 ( .A(u2__abc_44228_n7953), .B(u2__abc_44228_n7956), .Y(u2__abc_44228_n7957) );
  AND2X2 AND2X2_2865 ( .A(u2__abc_44228_n7958), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_remHi_24__FF_INPUT) );
  AND2X2 AND2X2_2866 ( .A(u2__abc_44228_n3062_bF_buf67), .B(u2_remHi_25_), .Y(u2__abc_44228_n7960_1) );
  AND2X2 AND2X2_2867 ( .A(u2__abc_44228_n7964), .B(u2__abc_44228_n7965), .Y(u2__abc_44228_n7966_1) );
  AND2X2 AND2X2_2868 ( .A(u2__abc_44228_n7547_bF_buf31), .B(u2__abc_44228_n7966_1), .Y(u2__abc_44228_n7967) );
  AND2X2 AND2X2_2869 ( .A(u2__abc_44228_n7548_1_bF_buf32), .B(u2_remHi_23_), .Y(u2__abc_44228_n7968) );
  AND2X2 AND2X2_287 ( .A(_abc_64468_n1459), .B(_abc_64468_n1458), .Y(fracta1_97_) );
  AND2X2 AND2X2_2870 ( .A(u2__abc_44228_n2983_bF_buf88), .B(u2__abc_44228_n3241), .Y(u2__abc_44228_n7971_1) );
  AND2X2 AND2X2_2871 ( .A(u2__abc_44228_n7972_1), .B(u2__abc_44228_n2972_bF_buf80), .Y(u2__abc_44228_n7973) );
  AND2X2 AND2X2_2872 ( .A(u2__abc_44228_n7970), .B(u2__abc_44228_n7973), .Y(u2__abc_44228_n7974) );
  AND2X2 AND2X2_2873 ( .A(u2__abc_44228_n7975), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_remHi_25__FF_INPUT) );
  AND2X2 AND2X2_2874 ( .A(u2__abc_44228_n3062_bF_buf66), .B(u2_remHi_26_), .Y(u2__abc_44228_n7977_1) );
  AND2X2 AND2X2_2875 ( .A(u2__abc_44228_n7945), .B(u2__abc_44228_n3237), .Y(u2__abc_44228_n7978) );
  AND2X2 AND2X2_2876 ( .A(u2__abc_44228_n7979), .B(u2__abc_44228_n3250), .Y(u2__abc_44228_n7981) );
  AND2X2 AND2X2_2877 ( .A(u2__abc_44228_n7982_1), .B(u2__abc_44228_n7980), .Y(u2__abc_44228_n7983_1) );
  AND2X2 AND2X2_2878 ( .A(u2__abc_44228_n7547_bF_buf30), .B(u2__abc_44228_n7983_1), .Y(u2__abc_44228_n7984) );
  AND2X2 AND2X2_2879 ( .A(u2__abc_44228_n7548_1_bF_buf31), .B(u2_remHi_24_), .Y(u2__abc_44228_n7985) );
  AND2X2 AND2X2_288 ( .A(_abc_64468_n1462), .B(_abc_64468_n1461), .Y(fracta1_98_) );
  AND2X2 AND2X2_2880 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n3211), .Y(u2__abc_44228_n7988_1) );
  AND2X2 AND2X2_2881 ( .A(u2__abc_44228_n7989), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n7990) );
  AND2X2 AND2X2_2882 ( .A(u2__abc_44228_n7987), .B(u2__abc_44228_n7990), .Y(u2__abc_44228_n7991) );
  AND2X2 AND2X2_2883 ( .A(u2__abc_44228_n7992), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_remHi_26__FF_INPUT) );
  AND2X2 AND2X2_2884 ( .A(u2__abc_44228_n3062_bF_buf65), .B(u2_remHi_27_), .Y(u2__abc_44228_n7994_1) );
  AND2X2 AND2X2_2885 ( .A(u2__abc_44228_n7982_1), .B(u2__abc_44228_n3332), .Y(u2__abc_44228_n7995) );
  AND2X2 AND2X2_2886 ( .A(u2__abc_44228_n7997), .B(u2__abc_44228_n7999_1), .Y(u2__abc_44228_n8000) );
  AND2X2 AND2X2_2887 ( .A(u2__abc_44228_n7547_bF_buf29), .B(u2__abc_44228_n8000), .Y(u2__abc_44228_n8001) );
  AND2X2 AND2X2_2888 ( .A(u2__abc_44228_n7548_1_bF_buf30), .B(u2_remHi_25_), .Y(u2__abc_44228_n8002) );
  AND2X2 AND2X2_2889 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n3218), .Y(u2__abc_44228_n8005_1) );
  AND2X2 AND2X2_289 ( .A(_abc_64468_n1465), .B(_abc_64468_n1464), .Y(fracta1_99_) );
  AND2X2 AND2X2_2890 ( .A(u2__abc_44228_n8006), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n8007) );
  AND2X2 AND2X2_2891 ( .A(u2__abc_44228_n8004_1), .B(u2__abc_44228_n8007), .Y(u2__abc_44228_n8008) );
  AND2X2 AND2X2_2892 ( .A(u2__abc_44228_n8009), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_remHi_27__FF_INPUT) );
  AND2X2 AND2X2_2893 ( .A(u2__abc_44228_n3062_bF_buf64), .B(u2_remHi_28_), .Y(u2__abc_44228_n8011) );
  AND2X2 AND2X2_2894 ( .A(u2__abc_44228_n7548_1_bF_buf29), .B(u2_remHi_26_), .Y(u2__abc_44228_n8012) );
  AND2X2 AND2X2_2895 ( .A(u2__abc_44228_n7982_1), .B(u2__abc_44228_n3333), .Y(u2__abc_44228_n8013) );
  AND2X2 AND2X2_2896 ( .A(u2__abc_44228_n8015_1), .B(u2__abc_44228_n3214), .Y(u2__abc_44228_n8016_1) );
  AND2X2 AND2X2_2897 ( .A(u2__abc_44228_n8017), .B(u2__abc_44228_n8018), .Y(u2__abc_44228_n8019) );
  AND2X2 AND2X2_2898 ( .A(u2__abc_44228_n7547_bF_buf28), .B(u2__abc_44228_n8019), .Y(u2__abc_44228_n8020) );
  AND2X2 AND2X2_2899 ( .A(u2__abc_44228_n2983_bF_buf82), .B(u2__abc_44228_n3204), .Y(u2__abc_44228_n8023) );
  AND2X2 AND2X2_29 ( .A(_abc_64468_n753_bF_buf13), .B(sqrto_28_), .Y(_auto_iopadmap_cc_313_execute_65414_64_) );
  AND2X2 AND2X2_290 ( .A(_abc_64468_n1468), .B(_abc_64468_n1467), .Y(fracta1_100_) );
  AND2X2 AND2X2_2900 ( .A(u2__abc_44228_n8024), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n8025) );
  AND2X2 AND2X2_2901 ( .A(u2__abc_44228_n8022), .B(u2__abc_44228_n8025), .Y(u2__abc_44228_n8026_1) );
  AND2X2 AND2X2_2902 ( .A(u2__abc_44228_n8027_1), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_remHi_28__FF_INPUT) );
  AND2X2 AND2X2_2903 ( .A(u2__abc_44228_n3062_bF_buf63), .B(u2_remHi_29_), .Y(u2__abc_44228_n8029) );
  AND2X2 AND2X2_2904 ( .A(u2__abc_44228_n8017), .B(u2__abc_44228_n3338), .Y(u2__abc_44228_n8032_1) );
  AND2X2 AND2X2_2905 ( .A(u2__abc_44228_n8033), .B(u2__abc_44228_n8031), .Y(u2__abc_44228_n8034) );
  AND2X2 AND2X2_2906 ( .A(u2__abc_44228_n8032_1), .B(u2__abc_44228_n3221), .Y(u2__abc_44228_n8035) );
  AND2X2 AND2X2_2907 ( .A(u2__abc_44228_n8037_1), .B(u2__abc_44228_n8030), .Y(u2__abc_44228_n8038_1) );
  AND2X2 AND2X2_2908 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n3198), .Y(u2__abc_44228_n8040) );
  AND2X2 AND2X2_2909 ( .A(u2__abc_44228_n8041), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n8042) );
  AND2X2 AND2X2_291 ( .A(_abc_64468_n1471), .B(_abc_64468_n1470), .Y(fracta1_101_) );
  AND2X2 AND2X2_2910 ( .A(u2__abc_44228_n8039), .B(u2__abc_44228_n8042), .Y(u2__abc_44228_n8043_1) );
  AND2X2 AND2X2_2911 ( .A(u2__abc_44228_n8044), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_remHi_29__FF_INPUT) );
  AND2X2 AND2X2_2912 ( .A(u2__abc_44228_n3062_bF_buf62), .B(u2_remHi_30_), .Y(u2__abc_44228_n8046) );
  AND2X2 AND2X2_2913 ( .A(u2__abc_44228_n8017), .B(u2__abc_44228_n3339), .Y(u2__abc_44228_n8047) );
  AND2X2 AND2X2_2914 ( .A(u2__abc_44228_n8049_1), .B(u2__abc_44228_n3207), .Y(u2__abc_44228_n8051) );
  AND2X2 AND2X2_2915 ( .A(u2__abc_44228_n8052), .B(u2__abc_44228_n8050), .Y(u2__abc_44228_n8053) );
  AND2X2 AND2X2_2916 ( .A(u2__abc_44228_n8054_1), .B(u2__abc_44228_n8055), .Y(u2__abc_44228_n8056) );
  AND2X2 AND2X2_2917 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n3569), .Y(u2__abc_44228_n8058) );
  AND2X2 AND2X2_2918 ( .A(u2__abc_44228_n8059_1), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n8060_1) );
  AND2X2 AND2X2_2919 ( .A(u2__abc_44228_n8057), .B(u2__abc_44228_n8060_1), .Y(u2__abc_44228_n8061) );
  AND2X2 AND2X2_292 ( .A(_abc_64468_n1474), .B(_abc_64468_n1473), .Y(fracta1_102_) );
  AND2X2 AND2X2_2920 ( .A(u2__abc_44228_n8062), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_remHi_30__FF_INPUT) );
  AND2X2 AND2X2_2921 ( .A(u2__abc_44228_n3062_bF_buf61), .B(u2_remHi_31_), .Y(u2__abc_44228_n8064) );
  AND2X2 AND2X2_2922 ( .A(u2__abc_44228_n8068), .B(u2__abc_44228_n8069), .Y(u2__abc_44228_n8070_1) );
  AND2X2 AND2X2_2923 ( .A(u2__abc_44228_n8070_1), .B(u2__abc_44228_n7547_bF_buf25), .Y(u2__abc_44228_n8071_1) );
  AND2X2 AND2X2_2924 ( .A(u2__abc_44228_n7548_1_bF_buf26), .B(u2_remHi_29_), .Y(u2__abc_44228_n8072) );
  AND2X2 AND2X2_2925 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n3576), .Y(u2__abc_44228_n8075) );
  AND2X2 AND2X2_2926 ( .A(u2__abc_44228_n8076_1), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n8077) );
  AND2X2 AND2X2_2927 ( .A(u2__abc_44228_n8074), .B(u2__abc_44228_n8077), .Y(u2__abc_44228_n8078) );
  AND2X2 AND2X2_2928 ( .A(u2__abc_44228_n8079), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_remHi_31__FF_INPUT) );
  AND2X2 AND2X2_2929 ( .A(u2__abc_44228_n3062_bF_buf60), .B(u2_remHi_32_), .Y(u2__abc_44228_n8081_1) );
  AND2X2 AND2X2_293 ( .A(_abc_64468_n1477), .B(_abc_64468_n1476), .Y(fracta1_103_) );
  AND2X2 AND2X2_2930 ( .A(u2__abc_44228_n3348), .B(u2__abc_44228_n3572), .Y(u2__abc_44228_n8082_1) );
  AND2X2 AND2X2_2931 ( .A(u2__abc_44228_n8083), .B(u2__abc_44228_n8084), .Y(u2__abc_44228_n8085) );
  AND2X2 AND2X2_2932 ( .A(u2__abc_44228_n7547_bF_buf24), .B(u2__abc_44228_n8085), .Y(u2__abc_44228_n8086) );
  AND2X2 AND2X2_2933 ( .A(u2__abc_44228_n7548_1_bF_buf25), .B(u2_remHi_30_), .Y(u2__abc_44228_n8087_1) );
  AND2X2 AND2X2_2934 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n3561), .Y(u2__abc_44228_n8090) );
  AND2X2 AND2X2_2935 ( .A(u2__abc_44228_n8091), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n8092_1) );
  AND2X2 AND2X2_2936 ( .A(u2__abc_44228_n8089), .B(u2__abc_44228_n8092_1), .Y(u2__abc_44228_n8093_1) );
  AND2X2 AND2X2_2937 ( .A(u2__abc_44228_n8094), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_remHi_32__FF_INPUT) );
  AND2X2 AND2X2_2938 ( .A(u2__abc_44228_n3062_bF_buf59), .B(u2_remHi_33_), .Y(u2__abc_44228_n8096) );
  AND2X2 AND2X2_2939 ( .A(u2__abc_44228_n8101), .B(u2__abc_44228_n8098_1), .Y(u2__abc_44228_n8102) );
  AND2X2 AND2X2_294 ( .A(_abc_64468_n1480), .B(_abc_64468_n1479), .Y(fracta1_104_) );
  AND2X2 AND2X2_2940 ( .A(u2__abc_44228_n7547_bF_buf23), .B(u2__abc_44228_n8102), .Y(u2__abc_44228_n8103_1) );
  AND2X2 AND2X2_2941 ( .A(u2__abc_44228_n7548_1_bF_buf24), .B(u2_remHi_31_), .Y(u2__abc_44228_n8104_1) );
  AND2X2 AND2X2_2942 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n3556), .Y(u2__abc_44228_n8107) );
  AND2X2 AND2X2_2943 ( .A(u2__abc_44228_n8108), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n8109_1) );
  AND2X2 AND2X2_2944 ( .A(u2__abc_44228_n8106), .B(u2__abc_44228_n8109_1), .Y(u2__abc_44228_n8110) );
  AND2X2 AND2X2_2945 ( .A(u2__abc_44228_n8111), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_remHi_33__FF_INPUT) );
  AND2X2 AND2X2_2946 ( .A(u2__abc_44228_n3062_bF_buf58), .B(u2_remHi_34_), .Y(u2__abc_44228_n8113) );
  AND2X2 AND2X2_2947 ( .A(u2__abc_44228_n3348), .B(u2__abc_44228_n3580_1), .Y(u2__abc_44228_n8114_1) );
  AND2X2 AND2X2_2948 ( .A(u2__abc_44228_n8115_1), .B(u2__abc_44228_n3565), .Y(u2__abc_44228_n8117) );
  AND2X2 AND2X2_2949 ( .A(u2__abc_44228_n8118), .B(u2__abc_44228_n8116), .Y(u2__abc_44228_n8119) );
  AND2X2 AND2X2_295 ( .A(_abc_64468_n1483), .B(_abc_64468_n1482), .Y(fracta1_105_) );
  AND2X2 AND2X2_2950 ( .A(u2__abc_44228_n7547_bF_buf22), .B(u2__abc_44228_n8119), .Y(u2__abc_44228_n8120_1) );
  AND2X2 AND2X2_2951 ( .A(u2__abc_44228_n7548_1_bF_buf23), .B(u2_remHi_32_), .Y(u2__abc_44228_n8121) );
  AND2X2 AND2X2_2952 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n3543), .Y(u2__abc_44228_n8124) );
  AND2X2 AND2X2_2953 ( .A(u2__abc_44228_n8125_1), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n8126_1) );
  AND2X2 AND2X2_2954 ( .A(u2__abc_44228_n8123), .B(u2__abc_44228_n8126_1), .Y(u2__abc_44228_n8127) );
  AND2X2 AND2X2_2955 ( .A(u2__abc_44228_n8128), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_remHi_34__FF_INPUT) );
  AND2X2 AND2X2_2956 ( .A(u2__abc_44228_n3062_bF_buf57), .B(u2_remHi_35_), .Y(u2__abc_44228_n8130) );
  AND2X2 AND2X2_2957 ( .A(u2__abc_44228_n7548_1_bF_buf22), .B(u2_remHi_33_), .Y(u2__abc_44228_n8131_1) );
  AND2X2 AND2X2_2958 ( .A(u2__abc_44228_n8118), .B(u2__abc_44228_n3562_1), .Y(u2__abc_44228_n8133) );
  AND2X2 AND2X2_2959 ( .A(u2__abc_44228_n8136_1), .B(u2__abc_44228_n8134), .Y(u2__abc_44228_n8137_1) );
  AND2X2 AND2X2_296 ( .A(_abc_64468_n1486), .B(_abc_64468_n1485), .Y(fracta1_106_) );
  AND2X2 AND2X2_2960 ( .A(u2__abc_44228_n7547_bF_buf21), .B(u2__abc_44228_n8137_1), .Y(u2__abc_44228_n8138) );
  AND2X2 AND2X2_2961 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n3550), .Y(u2__abc_44228_n8141) );
  AND2X2 AND2X2_2962 ( .A(u2__abc_44228_n8142_1), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n8143) );
  AND2X2 AND2X2_2963 ( .A(u2__abc_44228_n8140), .B(u2__abc_44228_n8143), .Y(u2__abc_44228_n8144) );
  AND2X2 AND2X2_2964 ( .A(u2__abc_44228_n8145), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_remHi_35__FF_INPUT) );
  AND2X2 AND2X2_2965 ( .A(u2__abc_44228_n3062_bF_buf56), .B(u2_remHi_36_), .Y(u2__abc_44228_n8147_1) );
  AND2X2 AND2X2_2966 ( .A(u2__abc_44228_n3348), .B(u2__abc_44228_n3581), .Y(u2__abc_44228_n8148_1) );
  AND2X2 AND2X2_2967 ( .A(u2__abc_44228_n8149), .B(u2__abc_44228_n3546), .Y(u2__abc_44228_n8150) );
  AND2X2 AND2X2_2968 ( .A(u2__abc_44228_n8151), .B(u2__abc_44228_n8152), .Y(u2__abc_44228_n8153_1) );
  AND2X2 AND2X2_2969 ( .A(u2__abc_44228_n7547_bF_buf20), .B(u2__abc_44228_n8153_1), .Y(u2__abc_44228_n8154) );
  AND2X2 AND2X2_297 ( .A(_abc_64468_n1489), .B(_abc_64468_n1488), .Y(fracta1_107_) );
  AND2X2 AND2X2_2970 ( .A(u2__abc_44228_n7548_1_bF_buf21), .B(u2_remHi_34_), .Y(u2__abc_44228_n8155) );
  AND2X2 AND2X2_2971 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n3536), .Y(u2__abc_44228_n8158_1) );
  AND2X2 AND2X2_2972 ( .A(u2__abc_44228_n8159_1), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n8160) );
  AND2X2 AND2X2_2973 ( .A(u2__abc_44228_n8157), .B(u2__abc_44228_n8160), .Y(u2__abc_44228_n8161) );
  AND2X2 AND2X2_2974 ( .A(u2__abc_44228_n8162), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_remHi_36__FF_INPUT) );
  AND2X2 AND2X2_2975 ( .A(u2__abc_44228_n3062_bF_buf55), .B(u2_remHi_37_), .Y(u2__abc_44228_n8164_1) );
  AND2X2 AND2X2_2976 ( .A(u2__abc_44228_n8151), .B(u2__abc_44228_n3595), .Y(u2__abc_44228_n8166) );
  AND2X2 AND2X2_2977 ( .A(u2__abc_44228_n8169_1), .B(u2__abc_44228_n8167), .Y(u2__abc_44228_n8170_1) );
  AND2X2 AND2X2_2978 ( .A(u2__abc_44228_n7547_bF_buf19), .B(u2__abc_44228_n8170_1), .Y(u2__abc_44228_n8171) );
  AND2X2 AND2X2_2979 ( .A(u2__abc_44228_n7548_1_bF_buf20), .B(u2_remHi_35_), .Y(u2__abc_44228_n8172) );
  AND2X2 AND2X2_298 ( .A(_abc_64468_n1492), .B(_abc_64468_n1491), .Y(fracta1_108_) );
  AND2X2 AND2X2_2980 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n3530), .Y(u2__abc_44228_n8175_1) );
  AND2X2 AND2X2_2981 ( .A(u2__abc_44228_n8176), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n8177) );
  AND2X2 AND2X2_2982 ( .A(u2__abc_44228_n8174), .B(u2__abc_44228_n8177), .Y(u2__abc_44228_n8178) );
  AND2X2 AND2X2_2983 ( .A(u2__abc_44228_n8179), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_remHi_37__FF_INPUT) );
  AND2X2 AND2X2_2984 ( .A(u2__abc_44228_n3062_bF_buf54), .B(u2_remHi_38_), .Y(u2__abc_44228_n8181_1) );
  AND2X2 AND2X2_2985 ( .A(u2__abc_44228_n7548_1_bF_buf19), .B(u2_remHi_36_), .Y(u2__abc_44228_n8182) );
  AND2X2 AND2X2_2986 ( .A(u2__abc_44228_n8151), .B(u2__abc_44228_n3596), .Y(u2__abc_44228_n8183) );
  AND2X2 AND2X2_2987 ( .A(u2__abc_44228_n8185), .B(u2__abc_44228_n3539), .Y(u2__abc_44228_n8187) );
  AND2X2 AND2X2_2988 ( .A(u2__abc_44228_n8188), .B(u2__abc_44228_n8186_1), .Y(u2__abc_44228_n8189) );
  AND2X2 AND2X2_2989 ( .A(u2__abc_44228_n7547_bF_buf18), .B(u2__abc_44228_n8189), .Y(u2__abc_44228_n8190) );
  AND2X2 AND2X2_299 ( .A(_abc_64468_n1495), .B(_abc_64468_n1494), .Y(fracta1_109_) );
  AND2X2 AND2X2_2990 ( .A(u2__abc_44228_n2983_bF_buf62), .B(u2__abc_44228_n3506), .Y(u2__abc_44228_n8193) );
  AND2X2 AND2X2_2991 ( .A(u2__abc_44228_n8194), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n8195) );
  AND2X2 AND2X2_2992 ( .A(u2__abc_44228_n8192_1), .B(u2__abc_44228_n8195), .Y(u2__abc_44228_n8196) );
  AND2X2 AND2X2_2993 ( .A(u2__abc_44228_n8197_1), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_remHi_38__FF_INPUT) );
  AND2X2 AND2X2_2994 ( .A(u2__abc_44228_n3062_bF_buf53), .B(u2_remHi_39_), .Y(u2__abc_44228_n8199) );
  AND2X2 AND2X2_2995 ( .A(u2__abc_44228_n8201), .B(u2__abc_44228_n8200), .Y(u2__abc_44228_n8202_1) );
  AND2X2 AND2X2_2996 ( .A(u2__abc_44228_n8203_1), .B(u2__abc_44228_n3533), .Y(u2__abc_44228_n8204) );
  AND2X2 AND2X2_2997 ( .A(u2__abc_44228_n7547_bF_buf17), .B(u2__abc_44228_n8205), .Y(u2__abc_44228_n8206) );
  AND2X2 AND2X2_2998 ( .A(u2__abc_44228_n2979), .B(u2_cnt_7_), .Y(u2__abc_44228_n8207) );
  AND2X2 AND2X2_2999 ( .A(u2__abc_44228_n2978), .B(u2__abc_44228_n3048), .Y(u2__abc_44228_n8208_1) );
  AND2X2 AND2X2_3 ( .A(_abc_64468_n753_bF_buf11), .B(sqrto_2_), .Y(_auto_iopadmap_cc_313_execute_65414_38_) );
  AND2X2 AND2X2_30 ( .A(_abc_64468_n753_bF_buf12), .B(sqrto_29_), .Y(_auto_iopadmap_cc_313_execute_65414_65_) );
  AND2X2 AND2X2_300 ( .A(_abc_64468_n1498), .B(_abc_64468_n1497), .Y(fracta1_110_) );
  AND2X2 AND2X2_3000 ( .A(u2__abc_44228_n8208_1), .B(u2__abc_44228_n8207), .Y(u2__abc_44228_n8209) );
  AND2X2 AND2X2_3001 ( .A(u2__abc_44228_n7548_1_bF_buf18), .B(u2_remHi_37_), .Y(u2__abc_44228_n8210) );
  AND2X2 AND2X2_3002 ( .A(u2__abc_44228_n2983_bF_buf61), .B(u2__abc_44228_n3500), .Y(u2__abc_44228_n8213_1) );
  AND2X2 AND2X2_3003 ( .A(u2__abc_44228_n8214_1), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n8215) );
  AND2X2 AND2X2_3004 ( .A(u2__abc_44228_n8212), .B(u2__abc_44228_n8215), .Y(u2__abc_44228_n8216) );
  AND2X2 AND2X2_3005 ( .A(u2__abc_44228_n8217), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_remHi_39__FF_INPUT) );
  AND2X2 AND2X2_3006 ( .A(u2__abc_44228_n3062_bF_buf52), .B(u2_remHi_40_), .Y(u2__abc_44228_n8219_1) );
  AND2X2 AND2X2_3007 ( .A(u2__abc_44228_n3348), .B(u2__abc_44228_n3582), .Y(u2__abc_44228_n8220) );
  AND2X2 AND2X2_3008 ( .A(u2__abc_44228_n8221), .B(u2__abc_44228_n3509), .Y(u2__abc_44228_n8223) );
  AND2X2 AND2X2_3009 ( .A(u2__abc_44228_n8224_1), .B(u2__abc_44228_n8222), .Y(u2__abc_44228_n8225_1) );
  AND2X2 AND2X2_301 ( .A(_abc_64468_n1501), .B(_abc_64468_n1500), .Y(fracta1_111_) );
  AND2X2 AND2X2_3010 ( .A(u2__abc_44228_n7547_bF_buf16), .B(u2__abc_44228_n8225_1), .Y(u2__abc_44228_n8226) );
  AND2X2 AND2X2_3011 ( .A(u2__abc_44228_n7548_1_bF_buf17), .B(u2_remHi_38_), .Y(u2__abc_44228_n8227) );
  AND2X2 AND2X2_3012 ( .A(u2__abc_44228_n2983_bF_buf59), .B(u2__abc_44228_n3520), .Y(u2__abc_44228_n8230_1) );
  AND2X2 AND2X2_3013 ( .A(u2__abc_44228_n8231), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n8232) );
  AND2X2 AND2X2_3014 ( .A(u2__abc_44228_n8229), .B(u2__abc_44228_n8232), .Y(u2__abc_44228_n8233) );
  AND2X2 AND2X2_3015 ( .A(u2__abc_44228_n8234), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_remHi_40__FF_INPUT) );
  AND2X2 AND2X2_3016 ( .A(u2__abc_44228_n3062_bF_buf51), .B(u2_remHi_41_), .Y(u2__abc_44228_n8236_1) );
  AND2X2 AND2X2_3017 ( .A(u2__abc_44228_n8240), .B(u2__abc_44228_n8241_1), .Y(u2__abc_44228_n8242) );
  AND2X2 AND2X2_3018 ( .A(u2__abc_44228_n7547_bF_buf15), .B(u2__abc_44228_n8242), .Y(u2__abc_44228_n8243) );
  AND2X2 AND2X2_3019 ( .A(u2__abc_44228_n7548_1_bF_buf16), .B(u2_remHi_39_), .Y(u2__abc_44228_n8244) );
  AND2X2 AND2X2_302 ( .A(_abc_64468_n1504), .B(_abc_64468_n1503), .Y(fracta1_112_) );
  AND2X2 AND2X2_3020 ( .A(u2__abc_44228_n2983_bF_buf57), .B(u2__abc_44228_n3514), .Y(u2__abc_44228_n8247_1) );
  AND2X2 AND2X2_3021 ( .A(u2__abc_44228_n8248), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n8249) );
  AND2X2 AND2X2_3022 ( .A(u2__abc_44228_n8246_1), .B(u2__abc_44228_n8249), .Y(u2__abc_44228_n8250) );
  AND2X2 AND2X2_3023 ( .A(u2__abc_44228_n8251), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_remHi_41__FF_INPUT) );
  AND2X2 AND2X2_3024 ( .A(u2__abc_44228_n3062_bF_buf50), .B(u2_remHi_42_), .Y(u2__abc_44228_n8253) );
  AND2X2 AND2X2_3025 ( .A(u2__abc_44228_n8221), .B(u2__abc_44228_n3510), .Y(u2__abc_44228_n8254) );
  AND2X2 AND2X2_3026 ( .A(u2__abc_44228_n8255), .B(u2__abc_44228_n3523_1), .Y(u2__abc_44228_n8257_1) );
  AND2X2 AND2X2_3027 ( .A(u2__abc_44228_n8258_1), .B(u2__abc_44228_n8256), .Y(u2__abc_44228_n8259) );
  AND2X2 AND2X2_3028 ( .A(u2__abc_44228_n7547_bF_buf14), .B(u2__abc_44228_n8259), .Y(u2__abc_44228_n8260) );
  AND2X2 AND2X2_3029 ( .A(u2__abc_44228_n7548_1_bF_buf15), .B(u2_remHi_40_), .Y(u2__abc_44228_n8261) );
  AND2X2 AND2X2_303 ( .A(_abc_64468_n1170_bF_buf7), .B(fracta_112_), .Y(fracta1_113_) );
  AND2X2 AND2X2_3030 ( .A(u2__abc_44228_n2983_bF_buf55), .B(u2__abc_44228_n3484_1), .Y(u2__abc_44228_n8264) );
  AND2X2 AND2X2_3031 ( .A(u2__abc_44228_n8265), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n8266) );
  AND2X2 AND2X2_3032 ( .A(u2__abc_44228_n8263_1), .B(u2__abc_44228_n8266), .Y(u2__abc_44228_n8267) );
  AND2X2 AND2X2_3033 ( .A(u2__abc_44228_n8268_1), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_remHi_42__FF_INPUT) );
  AND2X2 AND2X2_3034 ( .A(u2__abc_44228_n3062_bF_buf49), .B(u2_remHi_43_), .Y(u2__abc_44228_n8270) );
  AND2X2 AND2X2_3035 ( .A(u2__abc_44228_n8258_1), .B(u2__abc_44228_n3608_1), .Y(u2__abc_44228_n8272) );
  AND2X2 AND2X2_3036 ( .A(u2__abc_44228_n8273), .B(u2__abc_44228_n8271), .Y(u2__abc_44228_n8274_1) );
  AND2X2 AND2X2_3037 ( .A(u2__abc_44228_n8272), .B(u2__abc_44228_n3517), .Y(u2__abc_44228_n8275) );
  AND2X2 AND2X2_3038 ( .A(u2__abc_44228_n7547_bF_buf13), .B(u2__abc_44228_n8276), .Y(u2__abc_44228_n8277) );
  AND2X2 AND2X2_3039 ( .A(u2__abc_44228_n7548_1_bF_buf14), .B(u2_remHi_41_), .Y(u2__abc_44228_n8278) );
  AND2X2 AND2X2_304 ( .A(_abc_64468_n1170_bF_buf6), .B(_abc_64468_n1508), .Y(_abc_64468_n1509) );
  AND2X2 AND2X2_3040 ( .A(u2__abc_44228_n2983_bF_buf53), .B(u2__abc_44228_n3491), .Y(u2__abc_44228_n8281) );
  AND2X2 AND2X2_3041 ( .A(u2__abc_44228_n8282), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n8283) );
  AND2X2 AND2X2_3042 ( .A(u2__abc_44228_n8280_1), .B(u2__abc_44228_n8283), .Y(u2__abc_44228_n8284) );
  AND2X2 AND2X2_3043 ( .A(u2__abc_44228_n8285_1), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_remHi_43__FF_INPUT) );
  AND2X2 AND2X2_3044 ( .A(u2__abc_44228_n3062_bF_buf48), .B(u2_remHi_44_), .Y(u2__abc_44228_n8287) );
  AND2X2 AND2X2_3045 ( .A(u2__abc_44228_n8258_1), .B(u2__abc_44228_n3609), .Y(u2__abc_44228_n8288) );
  AND2X2 AND2X2_3046 ( .A(u2__abc_44228_n8290_1), .B(u2__abc_44228_n3487), .Y(u2__abc_44228_n8291_1) );
  AND2X2 AND2X2_3047 ( .A(u2__abc_44228_n8292), .B(u2__abc_44228_n8293), .Y(u2__abc_44228_n8294) );
  AND2X2 AND2X2_3048 ( .A(u2__abc_44228_n7547_bF_buf12), .B(u2__abc_44228_n8294), .Y(u2__abc_44228_n8295) );
  AND2X2 AND2X2_3049 ( .A(u2__abc_44228_n7548_1_bF_buf13), .B(u2_remHi_42_), .Y(u2__abc_44228_n8296_1) );
  AND2X2 AND2X2_305 ( .A(a_112_bF_buf4), .B(\a[113] ), .Y(_abc_64468_n1510) );
  AND2X2 AND2X2_3050 ( .A(u2__abc_44228_n2983_bF_buf51), .B(u2__abc_44228_n3477), .Y(u2__abc_44228_n8299) );
  AND2X2 AND2X2_3051 ( .A(u2__abc_44228_n8300), .B(u2__abc_44228_n2972_bF_buf61), .Y(u2__abc_44228_n8301_1) );
  AND2X2 AND2X2_3052 ( .A(u2__abc_44228_n8298), .B(u2__abc_44228_n8301_1), .Y(u2__abc_44228_n8302_1) );
  AND2X2 AND2X2_3053 ( .A(u2__abc_44228_n8303), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_remHi_44__FF_INPUT) );
  AND2X2 AND2X2_3054 ( .A(u2__abc_44228_n3062_bF_buf47), .B(u2_remHi_45_), .Y(u2__abc_44228_n8305) );
  AND2X2 AND2X2_3055 ( .A(u2__abc_44228_n8292), .B(u2__abc_44228_n3616), .Y(u2__abc_44228_n8307_1) );
  AND2X2 AND2X2_3056 ( .A(u2__abc_44228_n8310), .B(u2__abc_44228_n8308), .Y(u2__abc_44228_n8311) );
  AND2X2 AND2X2_3057 ( .A(u2__abc_44228_n8311), .B(u2__abc_44228_n7547_bF_buf11), .Y(u2__abc_44228_n8312_1) );
  AND2X2 AND2X2_3058 ( .A(u2__abc_44228_n7548_1_bF_buf12), .B(u2_remHi_43_), .Y(u2__abc_44228_n8313_1) );
  AND2X2 AND2X2_3059 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2__abc_44228_n3471), .Y(u2__abc_44228_n8316) );
  AND2X2 AND2X2_306 ( .A(_abc_64468_n1512), .B(_abc_64468_n1507), .Y(_auto_iopadmap_cc_313_execute_65414_226_) );
  AND2X2 AND2X2_3060 ( .A(u2__abc_44228_n8317), .B(u2__abc_44228_n2972_bF_buf60), .Y(u2__abc_44228_n8318_1) );
  AND2X2 AND2X2_3061 ( .A(u2__abc_44228_n8315), .B(u2__abc_44228_n8318_1), .Y(u2__abc_44228_n8319) );
  AND2X2 AND2X2_3062 ( .A(u2__abc_44228_n8320), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_remHi_45__FF_INPUT) );
  AND2X2 AND2X2_3063 ( .A(u2__abc_44228_n3062_bF_buf46), .B(u2_remHi_46_), .Y(u2__abc_44228_n8322) );
  AND2X2 AND2X2_3064 ( .A(u2__abc_44228_n8292), .B(u2__abc_44228_n3617_1), .Y(u2__abc_44228_n8323_1) );
  AND2X2 AND2X2_3065 ( .A(u2__abc_44228_n8325), .B(u2__abc_44228_n3480), .Y(u2__abc_44228_n8327) );
  AND2X2 AND2X2_3066 ( .A(u2__abc_44228_n8328), .B(u2__abc_44228_n8326), .Y(u2__abc_44228_n8329_1) );
  AND2X2 AND2X2_3067 ( .A(u2__abc_44228_n8330), .B(u2__abc_44228_n8331), .Y(u2__abc_44228_n8332) );
  AND2X2 AND2X2_3068 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n3460), .Y(u2__abc_44228_n8334_1) );
  AND2X2 AND2X2_3069 ( .A(u2__abc_44228_n8335_1), .B(u2__abc_44228_n2972_bF_buf59), .Y(u2__abc_44228_n8336) );
  AND2X2 AND2X2_307 ( .A(_abc_64468_n1515), .B(_abc_64468_n753_bF_buf5), .Y(_abc_64468_n1516) );
  AND2X2 AND2X2_3070 ( .A(u2__abc_44228_n8333), .B(u2__abc_44228_n8336), .Y(u2__abc_44228_n8337) );
  AND2X2 AND2X2_3071 ( .A(u2__abc_44228_n8338), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_remHi_46__FF_INPUT) );
  AND2X2 AND2X2_3072 ( .A(u2__abc_44228_n3062_bF_buf45), .B(u2_remHi_47_), .Y(u2__abc_44228_n8340_1) );
  AND2X2 AND2X2_3073 ( .A(u2__abc_44228_n8345_1), .B(u2__abc_44228_n7547_bF_buf9), .Y(u2__abc_44228_n8346_1) );
  AND2X2 AND2X2_3074 ( .A(u2__abc_44228_n8346_1), .B(u2__abc_44228_n8344), .Y(u2__abc_44228_n8347) );
  AND2X2 AND2X2_3075 ( .A(u2__abc_44228_n7548_1_bF_buf10), .B(u2_remHi_45_), .Y(u2__abc_44228_n8348) );
  AND2X2 AND2X2_3076 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n3454), .Y(u2__abc_44228_n8351_1) );
  AND2X2 AND2X2_3077 ( .A(u2__abc_44228_n8352), .B(u2__abc_44228_n2972_bF_buf58), .Y(u2__abc_44228_n8353) );
  AND2X2 AND2X2_3078 ( .A(u2__abc_44228_n8350), .B(u2__abc_44228_n8353), .Y(u2__abc_44228_n8354) );
  AND2X2 AND2X2_3079 ( .A(u2__abc_44228_n8355), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_remHi_47__FF_INPUT) );
  AND2X2 AND2X2_308 ( .A(_abc_64468_n1519), .B(_abc_64468_n753_bF_buf4), .Y(_abc_64468_n1520) );
  AND2X2 AND2X2_3080 ( .A(u2__abc_44228_n3062_bF_buf44), .B(u2_remHi_48_), .Y(u2__abc_44228_n8357_1) );
  AND2X2 AND2X2_3081 ( .A(u2__abc_44228_n3348), .B(u2__abc_44228_n3583), .Y(u2__abc_44228_n8358) );
  AND2X2 AND2X2_3082 ( .A(u2__abc_44228_n8359), .B(u2__abc_44228_n3463), .Y(u2__abc_44228_n8360) );
  AND2X2 AND2X2_3083 ( .A(u2__abc_44228_n8361), .B(u2__abc_44228_n8362_1), .Y(u2__abc_44228_n8363) );
  AND2X2 AND2X2_3084 ( .A(u2__abc_44228_n7547_bF_buf8), .B(u2__abc_44228_n8363), .Y(u2__abc_44228_n8364) );
  AND2X2 AND2X2_3085 ( .A(u2__abc_44228_n7548_1_bF_buf9), .B(u2_remHi_46_), .Y(u2__abc_44228_n8365) );
  AND2X2 AND2X2_3086 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n3446), .Y(u2__abc_44228_n8368_1) );
  AND2X2 AND2X2_3087 ( .A(u2__abc_44228_n8369), .B(u2__abc_44228_n2972_bF_buf57), .Y(u2__abc_44228_n8370) );
  AND2X2 AND2X2_3088 ( .A(u2__abc_44228_n8367_1), .B(u2__abc_44228_n8370), .Y(u2__abc_44228_n8371) );
  AND2X2 AND2X2_3089 ( .A(u2__abc_44228_n8372), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_remHi_48__FF_INPUT) );
  AND2X2 AND2X2_309 ( .A(_abc_64468_n1517), .B(_abc_64468_n1521), .Y(_auto_iopadmap_cc_313_execute_65414_227_) );
  AND2X2 AND2X2_3090 ( .A(u2__abc_44228_n3062_bF_buf43), .B(u2_remHi_49_), .Y(u2__abc_44228_n8374) );
  AND2X2 AND2X2_3091 ( .A(u2__abc_44228_n8378_1), .B(u2__abc_44228_n8379_1), .Y(u2__abc_44228_n8380) );
  AND2X2 AND2X2_3092 ( .A(u2__abc_44228_n7547_bF_buf7), .B(u2__abc_44228_n8380), .Y(u2__abc_44228_n8381) );
  AND2X2 AND2X2_3093 ( .A(u2__abc_44228_n7548_1_bF_buf8), .B(u2_remHi_47_), .Y(u2__abc_44228_n8382) );
  AND2X2 AND2X2_3094 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n3440), .Y(u2__abc_44228_n8385) );
  AND2X2 AND2X2_3095 ( .A(u2__abc_44228_n8386), .B(u2__abc_44228_n2972_bF_buf56), .Y(u2__abc_44228_n8387) );
  AND2X2 AND2X2_3096 ( .A(u2__abc_44228_n8384_1), .B(u2__abc_44228_n8387), .Y(u2__abc_44228_n8388) );
  AND2X2 AND2X2_3097 ( .A(u2__abc_44228_n8389_1), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_remHi_49__FF_INPUT) );
  AND2X2 AND2X2_3098 ( .A(u2__abc_44228_n3062_bF_buf42), .B(u2_remHi_50_), .Y(u2__abc_44228_n8391) );
  AND2X2 AND2X2_3099 ( .A(u2__abc_44228_n8359), .B(u2__abc_44228_n3464), .Y(u2__abc_44228_n8392) );
  AND2X2 AND2X2_31 ( .A(_abc_64468_n753_bF_buf11), .B(sqrto_30_), .Y(_auto_iopadmap_cc_313_execute_65414_66_) );
  AND2X2 AND2X2_310 ( .A(_abc_64468_n1514), .B(_abc_64468_n1523), .Y(_abc_64468_n1524) );
  AND2X2 AND2X2_3100 ( .A(u2__abc_44228_n8393), .B(u2__abc_44228_n3449_1), .Y(u2__abc_44228_n8395_1) );
  AND2X2 AND2X2_3101 ( .A(u2__abc_44228_n8396), .B(u2__abc_44228_n8394), .Y(u2__abc_44228_n8397) );
  AND2X2 AND2X2_3102 ( .A(u2__abc_44228_n7547_bF_buf6), .B(u2__abc_44228_n8397), .Y(u2__abc_44228_n8398) );
  AND2X2 AND2X2_3103 ( .A(u2__abc_44228_n7548_1_bF_buf7), .B(u2_remHi_48_), .Y(u2__abc_44228_n8399) );
  AND2X2 AND2X2_3104 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n3424), .Y(u2__abc_44228_n8402) );
  AND2X2 AND2X2_3105 ( .A(u2__abc_44228_n8403), .B(u2__abc_44228_n2972_bF_buf55), .Y(u2__abc_44228_n8404) );
  AND2X2 AND2X2_3106 ( .A(u2__abc_44228_n8401_1), .B(u2__abc_44228_n8404), .Y(u2__abc_44228_n8405) );
  AND2X2 AND2X2_3107 ( .A(u2__abc_44228_n8406_1), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_remHi_50__FF_INPUT) );
  AND2X2 AND2X2_3108 ( .A(u2__abc_44228_n3062_bF_buf41), .B(u2_remHi_51_), .Y(u2__abc_44228_n8408) );
  AND2X2 AND2X2_3109 ( .A(u2__abc_44228_n8410), .B(u2__abc_44228_n8409), .Y(u2__abc_44228_n8411_1) );
  AND2X2 AND2X2_311 ( .A(_abc_64468_n1510), .B(\a[114] ), .Y(_abc_64468_n1526) );
  AND2X2 AND2X2_3110 ( .A(u2__abc_44228_n8412_1), .B(u2__abc_44228_n3443), .Y(u2__abc_44228_n8413) );
  AND2X2 AND2X2_3111 ( .A(u2__abc_44228_n7547_bF_buf5), .B(u2__abc_44228_n8414), .Y(u2__abc_44228_n8415) );
  AND2X2 AND2X2_3112 ( .A(u2__abc_44228_n7548_1_bF_buf6), .B(u2_remHi_49_), .Y(u2__abc_44228_n8416) );
  AND2X2 AND2X2_3113 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n3431), .Y(u2__abc_44228_n8419) );
  AND2X2 AND2X2_3114 ( .A(u2__abc_44228_n8420), .B(u2__abc_44228_n2972_bF_buf54), .Y(u2__abc_44228_n8421) );
  AND2X2 AND2X2_3115 ( .A(u2__abc_44228_n8418), .B(u2__abc_44228_n8421), .Y(u2__abc_44228_n8422_1) );
  AND2X2 AND2X2_3116 ( .A(u2__abc_44228_n8423_1), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_remHi_51__FF_INPUT) );
  AND2X2 AND2X2_3117 ( .A(u2__abc_44228_n3062_bF_buf40), .B(u2_remHi_52_), .Y(u2__abc_44228_n8425) );
  AND2X2 AND2X2_3118 ( .A(u2__abc_44228_n8359), .B(u2__abc_44228_n3465), .Y(u2__abc_44228_n8426) );
  AND2X2 AND2X2_3119 ( .A(u2__abc_44228_n8427), .B(u2__abc_44228_n3427), .Y(u2__abc_44228_n8428_1) );
  AND2X2 AND2X2_312 ( .A(_abc_64468_n1526), .B(_abc_64468_n1525), .Y(_abc_64468_n1528) );
  AND2X2 AND2X2_3120 ( .A(u2__abc_44228_n8429), .B(u2__abc_44228_n8430), .Y(u2__abc_44228_n8431) );
  AND2X2 AND2X2_3121 ( .A(u2__abc_44228_n7547_bF_buf4), .B(u2__abc_44228_n8431), .Y(u2__abc_44228_n8432) );
  AND2X2 AND2X2_3122 ( .A(u2__abc_44228_n7548_1_bF_buf5), .B(u2_remHi_50_), .Y(u2__abc_44228_n8433_1) );
  AND2X2 AND2X2_3123 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n3417), .Y(u2__abc_44228_n8436) );
  AND2X2 AND2X2_3124 ( .A(u2__abc_44228_n8437), .B(u2__abc_44228_n2972_bF_buf53), .Y(u2__abc_44228_n8438) );
  AND2X2 AND2X2_3125 ( .A(u2__abc_44228_n8435), .B(u2__abc_44228_n8438), .Y(u2__abc_44228_n8439_1) );
  AND2X2 AND2X2_3126 ( .A(u2__abc_44228_n8440), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_remHi_52__FF_INPUT) );
  AND2X2 AND2X2_3127 ( .A(u2__abc_44228_n3062_bF_buf39), .B(u2_remHi_53_), .Y(u2__abc_44228_n8442) );
  AND2X2 AND2X2_3128 ( .A(u2__abc_44228_n8429), .B(u2__abc_44228_n3632), .Y(u2__abc_44228_n8443) );
  AND2X2 AND2X2_3129 ( .A(u2__abc_44228_n8443), .B(u2__abc_44228_n3434), .Y(u2__abc_44228_n8444_1) );
  AND2X2 AND2X2_313 ( .A(_abc_64468_n1529), .B(_abc_64468_n1527), .Y(_abc_64468_n1530) );
  AND2X2 AND2X2_3130 ( .A(u2__abc_44228_n8446), .B(u2__abc_44228_n8445_1), .Y(u2__abc_44228_n8447) );
  AND2X2 AND2X2_3131 ( .A(u2__abc_44228_n7547_bF_buf3), .B(u2__abc_44228_n8448), .Y(u2__abc_44228_n8449) );
  AND2X2 AND2X2_3132 ( .A(u2__abc_44228_n7548_1_bF_buf4), .B(u2_remHi_51_), .Y(u2__abc_44228_n8450_1) );
  AND2X2 AND2X2_3133 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n3411), .Y(u2__abc_44228_n8453) );
  AND2X2 AND2X2_3134 ( .A(u2__abc_44228_n8454), .B(u2__abc_44228_n2972_bF_buf52), .Y(u2__abc_44228_n8455_1) );
  AND2X2 AND2X2_3135 ( .A(u2__abc_44228_n8452), .B(u2__abc_44228_n8455_1), .Y(u2__abc_44228_n8456_1) );
  AND2X2 AND2X2_3136 ( .A(u2__abc_44228_n8457), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_remHi_53__FF_INPUT) );
  AND2X2 AND2X2_3137 ( .A(u2__abc_44228_n3062_bF_buf38), .B(u2_remHi_54_), .Y(u2__abc_44228_n8459) );
  AND2X2 AND2X2_3138 ( .A(u2__abc_44228_n8429), .B(u2__abc_44228_n3633), .Y(u2__abc_44228_n8460) );
  AND2X2 AND2X2_3139 ( .A(u2__abc_44228_n8462), .B(u2__abc_44228_n3420), .Y(u2__abc_44228_n8464) );
  AND2X2 AND2X2_314 ( .A(_abc_64468_n1530), .B(_abc_64468_n1524), .Y(_abc_64468_n1531) );
  AND2X2 AND2X2_3140 ( .A(u2__abc_44228_n8465), .B(u2__abc_44228_n8463), .Y(u2__abc_44228_n8466_1) );
  AND2X2 AND2X2_3141 ( .A(u2__abc_44228_n7547_bF_buf2), .B(u2__abc_44228_n8466_1), .Y(u2__abc_44228_n8467_1) );
  AND2X2 AND2X2_3142 ( .A(u2__abc_44228_n7548_1_bF_buf3), .B(u2_remHi_52_), .Y(u2__abc_44228_n8468) );
  AND2X2 AND2X2_3143 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n3401), .Y(u2__abc_44228_n8471) );
  AND2X2 AND2X2_3144 ( .A(u2__abc_44228_n8472_1), .B(u2__abc_44228_n2972_bF_buf51), .Y(u2__abc_44228_n8473) );
  AND2X2 AND2X2_3145 ( .A(u2__abc_44228_n8470), .B(u2__abc_44228_n8473), .Y(u2__abc_44228_n8474) );
  AND2X2 AND2X2_3146 ( .A(u2__abc_44228_n8475), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_remHi_54__FF_INPUT) );
  AND2X2 AND2X2_3147 ( .A(u2__abc_44228_n3062_bF_buf37), .B(u2_remHi_55_), .Y(u2__abc_44228_n8477_1) );
  AND2X2 AND2X2_3148 ( .A(u2__abc_44228_n8481), .B(u2__abc_44228_n8482), .Y(u2__abc_44228_n8483_1) );
  AND2X2 AND2X2_3149 ( .A(u2__abc_44228_n8483_1), .B(u2__abc_44228_n7547_bF_buf1), .Y(u2__abc_44228_n8484) );
  AND2X2 AND2X2_315 ( .A(_abc_64468_n1532), .B(\a[115] ), .Y(_abc_64468_n1533) );
  AND2X2 AND2X2_3150 ( .A(u2__abc_44228_n7548_1_bF_buf2), .B(u2_remHi_53_), .Y(u2__abc_44228_n8485) );
  AND2X2 AND2X2_3151 ( .A(u2__abc_44228_n2983_bF_buf31), .B(u2__abc_44228_n3395), .Y(u2__abc_44228_n8488_1) );
  AND2X2 AND2X2_3152 ( .A(u2__abc_44228_n8489_1), .B(u2__abc_44228_n2972_bF_buf50), .Y(u2__abc_44228_n8490) );
  AND2X2 AND2X2_3153 ( .A(u2__abc_44228_n8487), .B(u2__abc_44228_n8490), .Y(u2__abc_44228_n8491) );
  AND2X2 AND2X2_3154 ( .A(u2__abc_44228_n8492), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_remHi_55__FF_INPUT) );
  AND2X2 AND2X2_3155 ( .A(u2__abc_44228_n3062_bF_buf36), .B(u2_remHi_56_), .Y(u2__abc_44228_n8494_1) );
  AND2X2 AND2X2_3156 ( .A(u2__abc_44228_n8359), .B(u2__abc_44228_n3466), .Y(u2__abc_44228_n8495) );
  AND2X2 AND2X2_3157 ( .A(u2__abc_44228_n8496), .B(u2__abc_44228_n3404), .Y(u2__abc_44228_n8498) );
  AND2X2 AND2X2_3158 ( .A(u2__abc_44228_n8499_1), .B(u2__abc_44228_n8497), .Y(u2__abc_44228_n8500_1) );
  AND2X2 AND2X2_3159 ( .A(u2__abc_44228_n7547_bF_buf0), .B(u2__abc_44228_n8500_1), .Y(u2__abc_44228_n8501) );
  AND2X2 AND2X2_316 ( .A(_abc_64468_n1534), .B(_abc_64468_n753_bF_buf3), .Y(_abc_64468_n1535) );
  AND2X2 AND2X2_3160 ( .A(u2__abc_44228_n7548_1_bF_buf1), .B(u2_remHi_54_), .Y(u2__abc_44228_n8502) );
  AND2X2 AND2X2_3161 ( .A(u2__abc_44228_n2983_bF_buf29), .B(u2__abc_44228_n3387), .Y(u2__abc_44228_n8505_1) );
  AND2X2 AND2X2_3162 ( .A(u2__abc_44228_n8506), .B(u2__abc_44228_n2972_bF_buf49), .Y(u2__abc_44228_n8507) );
  AND2X2 AND2X2_3163 ( .A(u2__abc_44228_n8504), .B(u2__abc_44228_n8507), .Y(u2__abc_44228_n8508) );
  AND2X2 AND2X2_3164 ( .A(u2__abc_44228_n8509), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_remHi_56__FF_INPUT) );
  AND2X2 AND2X2_3165 ( .A(u2__abc_44228_n3062_bF_buf35), .B(u2_remHi_57_), .Y(u2__abc_44228_n8511_1) );
  AND2X2 AND2X2_3166 ( .A(u2__abc_44228_n7548_1_bF_buf0), .B(u2_remHi_55_), .Y(u2__abc_44228_n8512) );
  AND2X2 AND2X2_3167 ( .A(u2__abc_44228_n8499_1), .B(u2__abc_44228_n3642), .Y(u2__abc_44228_n8514) );
  AND2X2 AND2X2_3168 ( .A(u2__abc_44228_n8517), .B(u2__abc_44228_n8515), .Y(u2__abc_44228_n8518) );
  AND2X2 AND2X2_3169 ( .A(u2__abc_44228_n7547_bF_buf57), .B(u2__abc_44228_n8518), .Y(u2__abc_44228_n8519) );
  AND2X2 AND2X2_317 ( .A(aNan_bF_buf5), .B(\a[114] ), .Y(_abc_64468_n1536) );
  AND2X2 AND2X2_3170 ( .A(u2__abc_44228_n2983_bF_buf27), .B(u2__abc_44228_n3381), .Y(u2__abc_44228_n8522_1) );
  AND2X2 AND2X2_3171 ( .A(u2__abc_44228_n8523), .B(u2__abc_44228_n2972_bF_buf48), .Y(u2__abc_44228_n8524) );
  AND2X2 AND2X2_3172 ( .A(u2__abc_44228_n8521_1), .B(u2__abc_44228_n8524), .Y(u2__abc_44228_n8525) );
  AND2X2 AND2X2_3173 ( .A(u2__abc_44228_n8526), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_remHi_57__FF_INPUT) );
  AND2X2 AND2X2_3174 ( .A(u2__abc_44228_n3062_bF_buf34), .B(u2_remHi_58_), .Y(u2__abc_44228_n8528) );
  AND2X2 AND2X2_3175 ( .A(u2__abc_44228_n8496), .B(u2__abc_44228_n3405), .Y(u2__abc_44228_n8529) );
  AND2X2 AND2X2_3176 ( .A(u2__abc_44228_n8530), .B(u2__abc_44228_n3390), .Y(u2__abc_44228_n8532_1) );
  AND2X2 AND2X2_3177 ( .A(u2__abc_44228_n8533_1), .B(u2__abc_44228_n8531), .Y(u2__abc_44228_n8534) );
  AND2X2 AND2X2_3178 ( .A(u2__abc_44228_n8535), .B(u2__abc_44228_n8536), .Y(u2__abc_44228_n8537) );
  AND2X2 AND2X2_3179 ( .A(u2__abc_44228_n2983_bF_buf25), .B(u2__abc_44228_n3365), .Y(u2__abc_44228_n8539) );
  AND2X2 AND2X2_318 ( .A(_abc_64468_n1526), .B(\a[115] ), .Y(_abc_64468_n1539) );
  AND2X2 AND2X2_3180 ( .A(u2__abc_44228_n8540), .B(u2__abc_44228_n2972_bF_buf47), .Y(u2__abc_44228_n8541) );
  AND2X2 AND2X2_3181 ( .A(u2__abc_44228_n8538_1), .B(u2__abc_44228_n8541), .Y(u2__abc_44228_n8542) );
  AND2X2 AND2X2_3182 ( .A(u2__abc_44228_n8543_1), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_remHi_58__FF_INPUT) );
  AND2X2 AND2X2_3183 ( .A(u2__abc_44228_n3062_bF_buf33), .B(u2_remHi_59_), .Y(u2__abc_44228_n8545) );
  AND2X2 AND2X2_3184 ( .A(u2__abc_44228_n8533_1), .B(u2__abc_44228_n3647_1), .Y(u2__abc_44228_n8546) );
  AND2X2 AND2X2_3185 ( .A(u2__abc_44228_n8548), .B(u2__abc_44228_n8550), .Y(u2__abc_44228_n8551) );
  AND2X2 AND2X2_3186 ( .A(u2__abc_44228_n7547_bF_buf55), .B(u2__abc_44228_n8551), .Y(u2__abc_44228_n8552) );
  AND2X2 AND2X2_3187 ( .A(u2__abc_44228_n7548_1_bF_buf56), .B(u2_remHi_57_), .Y(u2__abc_44228_n8553) );
  AND2X2 AND2X2_3188 ( .A(u2__abc_44228_n2983_bF_buf23), .B(u2__abc_44228_n3372), .Y(u2__abc_44228_n8556) );
  AND2X2 AND2X2_3189 ( .A(u2__abc_44228_n8557), .B(u2__abc_44228_n2972_bF_buf46), .Y(u2__abc_44228_n8558) );
  AND2X2 AND2X2_319 ( .A(_abc_64468_n1539), .B(_abc_64468_n1538), .Y(_abc_64468_n1541) );
  AND2X2 AND2X2_3190 ( .A(u2__abc_44228_n8555_1), .B(u2__abc_44228_n8558), .Y(u2__abc_44228_n8559) );
  AND2X2 AND2X2_3191 ( .A(u2__abc_44228_n8560_1), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_remHi_59__FF_INPUT) );
  AND2X2 AND2X2_3192 ( .A(u2__abc_44228_n3062_bF_buf32), .B(u2_remHi_60_), .Y(u2__abc_44228_n8562) );
  AND2X2 AND2X2_3193 ( .A(u2__abc_44228_n8533_1), .B(u2__abc_44228_n3648), .Y(u2__abc_44228_n8563) );
  AND2X2 AND2X2_3194 ( .A(u2__abc_44228_n8565_1), .B(u2__abc_44228_n3368), .Y(u2__abc_44228_n8566_1) );
  AND2X2 AND2X2_3195 ( .A(u2__abc_44228_n8567), .B(u2__abc_44228_n8568), .Y(u2__abc_44228_n8569) );
  AND2X2 AND2X2_3196 ( .A(u2__abc_44228_n8570), .B(u2__abc_44228_n8571_1), .Y(u2__abc_44228_n8572) );
  AND2X2 AND2X2_3197 ( .A(u2__abc_44228_n2983_bF_buf21), .B(u2__abc_44228_n3358), .Y(u2__abc_44228_n8574) );
  AND2X2 AND2X2_3198 ( .A(u2__abc_44228_n8575), .B(u2__abc_44228_n2972_bF_buf45), .Y(u2__abc_44228_n8576_1) );
  AND2X2 AND2X2_3199 ( .A(u2__abc_44228_n8573), .B(u2__abc_44228_n8576_1), .Y(u2__abc_44228_n8577_1) );
  AND2X2 AND2X2_32 ( .A(_abc_64468_n753_bF_buf10), .B(sqrto_31_), .Y(_auto_iopadmap_cc_313_execute_65414_67_) );
  AND2X2 AND2X2_320 ( .A(_abc_64468_n1542), .B(_abc_64468_n1540), .Y(_abc_64468_n1543) );
  AND2X2 AND2X2_3200 ( .A(u2__abc_44228_n8578), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_remHi_60__FF_INPUT) );
  AND2X2 AND2X2_3201 ( .A(u2__abc_44228_n3062_bF_buf31), .B(u2_remHi_61_), .Y(u2__abc_44228_n8580) );
  AND2X2 AND2X2_3202 ( .A(u2__abc_44228_n8567), .B(u2__abc_44228_n3655), .Y(u2__abc_44228_n8581) );
  AND2X2 AND2X2_3203 ( .A(u2__abc_44228_n8585), .B(u2__abc_44228_n7547_bF_buf53), .Y(u2__abc_44228_n8586) );
  AND2X2 AND2X2_3204 ( .A(u2__abc_44228_n8586), .B(u2__abc_44228_n8583), .Y(u2__abc_44228_n8587_1) );
  AND2X2 AND2X2_3205 ( .A(u2__abc_44228_n7548_1_bF_buf54), .B(u2_remHi_59_), .Y(u2__abc_44228_n8588_1) );
  AND2X2 AND2X2_3206 ( .A(u2__abc_44228_n2983_bF_buf19), .B(u2__abc_44228_n3352), .Y(u2__abc_44228_n8591) );
  AND2X2 AND2X2_3207 ( .A(u2__abc_44228_n8592), .B(u2__abc_44228_n2972_bF_buf44), .Y(u2__abc_44228_n8593_1) );
  AND2X2 AND2X2_3208 ( .A(u2__abc_44228_n8590), .B(u2__abc_44228_n8593_1), .Y(u2__abc_44228_n8594) );
  AND2X2 AND2X2_3209 ( .A(u2__abc_44228_n8595), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_remHi_61__FF_INPUT) );
  AND2X2 AND2X2_321 ( .A(_abc_64468_n1531), .B(_abc_64468_n1543), .Y(_abc_64468_n1544) );
  AND2X2 AND2X2_3210 ( .A(u2__abc_44228_n3062_bF_buf30), .B(u2_remHi_62_), .Y(u2__abc_44228_n8597) );
  AND2X2 AND2X2_3211 ( .A(u2__abc_44228_n8567), .B(u2__abc_44228_n3656_1), .Y(u2__abc_44228_n8598_1) );
  AND2X2 AND2X2_3212 ( .A(u2__abc_44228_n8600), .B(u2__abc_44228_n3361), .Y(u2__abc_44228_n8602) );
  AND2X2 AND2X2_3213 ( .A(u2__abc_44228_n8603), .B(u2__abc_44228_n8601), .Y(u2__abc_44228_n8604_1) );
  AND2X2 AND2X2_3214 ( .A(u2__abc_44228_n8604_1), .B(u2__abc_44228_n7547_bF_buf52), .Y(u2__abc_44228_n8605) );
  AND2X2 AND2X2_3215 ( .A(u2__abc_44228_n7548_1_bF_buf53), .B(u2_remHi_60_), .Y(u2__abc_44228_n8606) );
  AND2X2 AND2X2_3216 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n4131), .Y(u2__abc_44228_n8609_1) );
  AND2X2 AND2X2_3217 ( .A(u2__abc_44228_n8610_1), .B(u2__abc_44228_n2972_bF_buf43), .Y(u2__abc_44228_n8611) );
  AND2X2 AND2X2_3218 ( .A(u2__abc_44228_n8608), .B(u2__abc_44228_n8611), .Y(u2__abc_44228_n8612) );
  AND2X2 AND2X2_3219 ( .A(u2__abc_44228_n8613), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_remHi_62__FF_INPUT) );
  AND2X2 AND2X2_322 ( .A(_abc_64468_n1545), .B(_abc_64468_n1546), .Y(_abc_64468_n1547) );
  AND2X2 AND2X2_3220 ( .A(u2__abc_44228_n3062_bF_buf29), .B(u2_remHi_63_), .Y(u2__abc_44228_n8615_1) );
  AND2X2 AND2X2_3221 ( .A(u2__abc_44228_n8620_1), .B(u2__abc_44228_n7547_bF_buf51), .Y(u2__abc_44228_n8621_1) );
  AND2X2 AND2X2_3222 ( .A(u2__abc_44228_n8621_1), .B(u2__abc_44228_n8619), .Y(u2__abc_44228_n8622) );
  AND2X2 AND2X2_3223 ( .A(u2__abc_44228_n7548_1_bF_buf52), .B(u2_remHi_61_), .Y(u2__abc_44228_n8623) );
  AND2X2 AND2X2_3224 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n4125), .Y(u2__abc_44228_n8626_1) );
  AND2X2 AND2X2_3225 ( .A(u2__abc_44228_n8627), .B(u2__abc_44228_n2972_bF_buf42), .Y(u2__abc_44228_n8628) );
  AND2X2 AND2X2_3226 ( .A(u2__abc_44228_n8625), .B(u2__abc_44228_n8628), .Y(u2__abc_44228_n8629) );
  AND2X2 AND2X2_3227 ( .A(u2__abc_44228_n8630), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_remHi_63__FF_INPUT) );
  AND2X2 AND2X2_3228 ( .A(u2__abc_44228_n3062_bF_buf28), .B(u2_remHi_64_), .Y(u2__abc_44228_n8632_1) );
  AND2X2 AND2X2_3229 ( .A(u2__abc_44228_n3664), .B(u2__abc_44228_n4134), .Y(u2__abc_44228_n8634) );
  AND2X2 AND2X2_323 ( .A(_abc_64468_n1549), .B(_abc_64468_n1550), .Y(_auto_iopadmap_cc_313_execute_65414_229_) );
  AND2X2 AND2X2_3230 ( .A(u2__abc_44228_n8635), .B(u2__abc_44228_n8633), .Y(u2__abc_44228_n8636) );
  AND2X2 AND2X2_3231 ( .A(u2__abc_44228_n7547_bF_buf50), .B(u2__abc_44228_n8636), .Y(u2__abc_44228_n8637_1) );
  AND2X2 AND2X2_3232 ( .A(u2__abc_44228_n7548_1_bF_buf51), .B(u2_remHi_62_), .Y(u2__abc_44228_n8638) );
  AND2X2 AND2X2_3233 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n4116), .Y(u2__abc_44228_n8641) );
  AND2X2 AND2X2_3234 ( .A(u2__abc_44228_n8642_1), .B(u2__abc_44228_n2972_bF_buf41), .Y(u2__abc_44228_n8643_1) );
  AND2X2 AND2X2_3235 ( .A(u2__abc_44228_n8640), .B(u2__abc_44228_n8643_1), .Y(u2__abc_44228_n8644) );
  AND2X2 AND2X2_3236 ( .A(u2__abc_44228_n8645), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_remHi_64__FF_INPUT) );
  AND2X2 AND2X2_3237 ( .A(u2__abc_44228_n3062_bF_buf27), .B(u2_remHi_65_), .Y(u2__abc_44228_n8647) );
  AND2X2 AND2X2_3238 ( .A(u2__abc_44228_n8651), .B(u2__abc_44228_n8652), .Y(u2__abc_44228_n8653_1) );
  AND2X2 AND2X2_3239 ( .A(u2__abc_44228_n7547_bF_buf49), .B(u2__abc_44228_n8653_1), .Y(u2__abc_44228_n8654_1) );
  AND2X2 AND2X2_324 ( .A(_abc_64468_n1539), .B(\a[116] ), .Y(_abc_64468_n1553) );
  AND2X2 AND2X2_3240 ( .A(u2__abc_44228_n7548_1_bF_buf50), .B(u2_remHi_63_), .Y(u2__abc_44228_n8655) );
  AND2X2 AND2X2_3241 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n4111), .Y(u2__abc_44228_n8658) );
  AND2X2 AND2X2_3242 ( .A(u2__abc_44228_n8659_1), .B(u2__abc_44228_n2972_bF_buf40), .Y(u2__abc_44228_n8660) );
  AND2X2 AND2X2_3243 ( .A(u2__abc_44228_n8657), .B(u2__abc_44228_n8660), .Y(u2__abc_44228_n8661) );
  AND2X2 AND2X2_3244 ( .A(u2__abc_44228_n8662), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_remHi_65__FF_INPUT) );
  AND2X2 AND2X2_3245 ( .A(u2__abc_44228_n3062_bF_buf26), .B(u2_remHi_66_), .Y(u2__abc_44228_n8664_1) );
  AND2X2 AND2X2_3246 ( .A(u2__abc_44228_n3664), .B(u2__abc_44228_n4135), .Y(u2__abc_44228_n8665_1) );
  AND2X2 AND2X2_3247 ( .A(u2__abc_44228_n8666), .B(u2__abc_44228_n4120), .Y(u2__abc_44228_n8668) );
  AND2X2 AND2X2_3248 ( .A(u2__abc_44228_n8669), .B(u2__abc_44228_n8667), .Y(u2__abc_44228_n8670_1) );
  AND2X2 AND2X2_3249 ( .A(u2__abc_44228_n7547_bF_buf48), .B(u2__abc_44228_n8670_1), .Y(u2__abc_44228_n8671) );
  AND2X2 AND2X2_325 ( .A(_abc_64468_n1553), .B(\a[117] ), .Y(_abc_64468_n1554) );
  AND2X2 AND2X2_3250 ( .A(u2__abc_44228_n7548_1_bF_buf49), .B(u2_remHi_64_), .Y(u2__abc_44228_n8672) );
  AND2X2 AND2X2_3251 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n4105), .Y(u2__abc_44228_n8675_1) );
  AND2X2 AND2X2_3252 ( .A(u2__abc_44228_n8676_1), .B(u2__abc_44228_n2972_bF_buf39), .Y(u2__abc_44228_n8677) );
  AND2X2 AND2X2_3253 ( .A(u2__abc_44228_n8674), .B(u2__abc_44228_n8677), .Y(u2__abc_44228_n8678) );
  AND2X2 AND2X2_3254 ( .A(u2__abc_44228_n8679), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_remHi_66__FF_INPUT) );
  AND2X2 AND2X2_3255 ( .A(u2__abc_44228_n3062_bF_buf25), .B(u2_remHi_67_), .Y(u2__abc_44228_n8681_1) );
  AND2X2 AND2X2_3256 ( .A(u2__abc_44228_n8669), .B(u2__abc_44228_n4117), .Y(u2__abc_44228_n8683) );
  AND2X2 AND2X2_3257 ( .A(u2__abc_44228_n8684), .B(u2__abc_44228_n8682), .Y(u2__abc_44228_n8685) );
  AND2X2 AND2X2_3258 ( .A(u2__abc_44228_n8683), .B(u2__abc_44228_n4115), .Y(u2__abc_44228_n8686_1) );
  AND2X2 AND2X2_3259 ( .A(u2__abc_44228_n7547_bF_buf47), .B(u2__abc_44228_n8687_1), .Y(u2__abc_44228_n8688) );
  AND2X2 AND2X2_326 ( .A(_abc_64468_n1556), .B(_abc_64468_n1555), .Y(_abc_64468_n1557) );
  AND2X2 AND2X2_3260 ( .A(u2__abc_44228_n7548_1_bF_buf48), .B(u2_remHi_65_), .Y(u2__abc_44228_n8689) );
  AND2X2 AND2X2_3261 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n4099), .Y(u2__abc_44228_n8692_1) );
  AND2X2 AND2X2_3262 ( .A(u2__abc_44228_n8693), .B(u2__abc_44228_n2972_bF_buf38), .Y(u2__abc_44228_n8694) );
  AND2X2 AND2X2_3263 ( .A(u2__abc_44228_n8691), .B(u2__abc_44228_n8694), .Y(u2__abc_44228_n8695) );
  AND2X2 AND2X2_3264 ( .A(u2__abc_44228_n8696), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_remHi_67__FF_INPUT) );
  AND2X2 AND2X2_3265 ( .A(u2__abc_44228_n3062_bF_buf24), .B(u2_remHi_68_), .Y(u2__abc_44228_n8698_1) );
  AND2X2 AND2X2_3266 ( .A(u2__abc_44228_n3664), .B(u2__abc_44228_n4136), .Y(u2__abc_44228_n8699) );
  AND2X2 AND2X2_3267 ( .A(u2__abc_44228_n8700), .B(u2__abc_44228_n4108), .Y(u2__abc_44228_n8701) );
  AND2X2 AND2X2_3268 ( .A(u2__abc_44228_n8702), .B(u2__abc_44228_n8703_1), .Y(u2__abc_44228_n8704) );
  AND2X2 AND2X2_3269 ( .A(u2__abc_44228_n7547_bF_buf46), .B(u2__abc_44228_n8704), .Y(u2__abc_44228_n8705) );
  AND2X2 AND2X2_327 ( .A(_abc_64468_n1559), .B(_abc_64468_n1552), .Y(_abc_64468_n1560) );
  AND2X2 AND2X2_3270 ( .A(u2__abc_44228_n7548_1_bF_buf47), .B(u2_remHi_66_), .Y(u2__abc_44228_n8706) );
  AND2X2 AND2X2_3271 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n4091), .Y(u2__abc_44228_n8709_1) );
  AND2X2 AND2X2_3272 ( .A(u2__abc_44228_n8710), .B(u2__abc_44228_n2972_bF_buf37), .Y(u2__abc_44228_n8711) );
  AND2X2 AND2X2_3273 ( .A(u2__abc_44228_n8708_1), .B(u2__abc_44228_n8711), .Y(u2__abc_44228_n8712) );
  AND2X2 AND2X2_3274 ( .A(u2__abc_44228_n8713), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_remHi_68__FF_INPUT) );
  AND2X2 AND2X2_3275 ( .A(u2__abc_44228_n3062_bF_buf23), .B(u2_remHi_69_), .Y(u2__abc_44228_n8715) );
  AND2X2 AND2X2_3276 ( .A(u2__abc_44228_n8717), .B(u2__abc_44228_n8716), .Y(u2__abc_44228_n8718) );
  AND2X2 AND2X2_3277 ( .A(u2__abc_44228_n8719_1), .B(u2__abc_44228_n4102), .Y(u2__abc_44228_n8720_1) );
  AND2X2 AND2X2_3278 ( .A(u2__abc_44228_n7547_bF_buf45), .B(u2__abc_44228_n8721), .Y(u2__abc_44228_n8722) );
  AND2X2 AND2X2_3279 ( .A(u2__abc_44228_n7548_1_bF_buf46), .B(u2_remHi_67_), .Y(u2__abc_44228_n8723) );
  AND2X2 AND2X2_328 ( .A(_abc_64468_n1558), .B(_abc_64468_n1544), .Y(_abc_64468_n1561) );
  AND2X2 AND2X2_3280 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n4085), .Y(u2__abc_44228_n8726) );
  AND2X2 AND2X2_3281 ( .A(u2__abc_44228_n8727), .B(u2__abc_44228_n2972_bF_buf36), .Y(u2__abc_44228_n8728) );
  AND2X2 AND2X2_3282 ( .A(u2__abc_44228_n8725_1), .B(u2__abc_44228_n8728), .Y(u2__abc_44228_n8729) );
  AND2X2 AND2X2_3283 ( .A(u2__abc_44228_n8730_1), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_remHi_69__FF_INPUT) );
  AND2X2 AND2X2_3284 ( .A(u2__abc_44228_n3062_bF_buf22), .B(u2_remHi_70_), .Y(u2__abc_44228_n8732) );
  AND2X2 AND2X2_3285 ( .A(u2__abc_44228_n7548_1_bF_buf45), .B(u2_remHi_68_), .Y(u2__abc_44228_n8733) );
  AND2X2 AND2X2_3286 ( .A(u2__abc_44228_n8700), .B(u2__abc_44228_n4109_1), .Y(u2__abc_44228_n8734) );
  AND2X2 AND2X2_3287 ( .A(u2__abc_44228_n8735), .B(u2__abc_44228_n4094), .Y(u2__abc_44228_n8737) );
  AND2X2 AND2X2_3288 ( .A(u2__abc_44228_n8738), .B(u2__abc_44228_n8736_1), .Y(u2__abc_44228_n8739) );
  AND2X2 AND2X2_3289 ( .A(u2__abc_44228_n7547_bF_buf44), .B(u2__abc_44228_n8739), .Y(u2__abc_44228_n8740) );
  AND2X2 AND2X2_329 ( .A(_abc_64468_n1563), .B(_abc_64468_n1564), .Y(_auto_iopadmap_cc_313_execute_65414_230_) );
  AND2X2 AND2X2_3290 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n4061_1), .Y(u2__abc_44228_n8743) );
  AND2X2 AND2X2_3291 ( .A(u2__abc_44228_n8744), .B(u2__abc_44228_n2972_bF_buf35), .Y(u2__abc_44228_n8745) );
  AND2X2 AND2X2_3292 ( .A(u2__abc_44228_n8742_1), .B(u2__abc_44228_n8745), .Y(u2__abc_44228_n8746) );
  AND2X2 AND2X2_3293 ( .A(u2__abc_44228_n8747_1), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_remHi_70__FF_INPUT) );
  AND2X2 AND2X2_3294 ( .A(u2__abc_44228_n3062_bF_buf21), .B(u2_remHi_71_), .Y(u2__abc_44228_n8749) );
  AND2X2 AND2X2_3295 ( .A(u2__abc_44228_n7548_1_bF_buf44), .B(u2_remHi_69_), .Y(u2__abc_44228_n8750) );
  AND2X2 AND2X2_3296 ( .A(u2__abc_44228_n8752_1), .B(u2__abc_44228_n8751), .Y(u2__abc_44228_n8753_1) );
  AND2X2 AND2X2_3297 ( .A(u2__abc_44228_n8754), .B(u2__abc_44228_n4088), .Y(u2__abc_44228_n8755) );
  AND2X2 AND2X2_3298 ( .A(u2__abc_44228_n7547_bF_buf43), .B(u2__abc_44228_n8756), .Y(u2__abc_44228_n8757) );
  AND2X2 AND2X2_3299 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n4055), .Y(u2__abc_44228_n8760) );
  AND2X2 AND2X2_33 ( .A(_abc_64468_n753_bF_buf9), .B(sqrto_32_), .Y(_auto_iopadmap_cc_313_execute_65414_68_) );
  AND2X2 AND2X2_330 ( .A(aNan_bF_buf2), .B(\a[117] ), .Y(_abc_64468_n1566) );
  AND2X2 AND2X2_3300 ( .A(u2__abc_44228_n8761), .B(u2__abc_44228_n2972_bF_buf34), .Y(u2__abc_44228_n8762) );
  AND2X2 AND2X2_3301 ( .A(u2__abc_44228_n8759), .B(u2__abc_44228_n8762), .Y(u2__abc_44228_n8763_1) );
  AND2X2 AND2X2_3302 ( .A(u2__abc_44228_n8764_1), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_remHi_71__FF_INPUT) );
  AND2X2 AND2X2_3303 ( .A(u2__abc_44228_n3062_bF_buf20), .B(u2_remHi_72_), .Y(u2__abc_44228_n8766) );
  AND2X2 AND2X2_3304 ( .A(u2__abc_44228_n3664), .B(u2__abc_44228_n4137), .Y(u2__abc_44228_n8767) );
  AND2X2 AND2X2_3305 ( .A(u2__abc_44228_n8768), .B(u2__abc_44228_n4064), .Y(u2__abc_44228_n8770) );
  AND2X2 AND2X2_3306 ( .A(u2__abc_44228_n8771), .B(u2__abc_44228_n8769_1), .Y(u2__abc_44228_n8772) );
  AND2X2 AND2X2_3307 ( .A(u2__abc_44228_n7547_bF_buf42), .B(u2__abc_44228_n8772), .Y(u2__abc_44228_n8773) );
  AND2X2 AND2X2_3308 ( .A(u2__abc_44228_n7548_1_bF_buf43), .B(u2_remHi_70_), .Y(u2__abc_44228_n8774_1) );
  AND2X2 AND2X2_3309 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n4075), .Y(u2__abc_44228_n8777) );
  AND2X2 AND2X2_331 ( .A(_abc_64468_n1554), .B(_abc_64468_n1568), .Y(_abc_64468_n1570) );
  AND2X2 AND2X2_3310 ( .A(u2__abc_44228_n8778), .B(u2__abc_44228_n2972_bF_buf33), .Y(u2__abc_44228_n8779) );
  AND2X2 AND2X2_3311 ( .A(u2__abc_44228_n8776), .B(u2__abc_44228_n8779), .Y(u2__abc_44228_n8780_1) );
  AND2X2 AND2X2_3312 ( .A(u2__abc_44228_n8781), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_remHi_72__FF_INPUT) );
  AND2X2 AND2X2_3313 ( .A(u2__abc_44228_n3062_bF_buf19), .B(u2_remHi_73_), .Y(u2__abc_44228_n8783) );
  AND2X2 AND2X2_3314 ( .A(u2__abc_44228_n8785_1), .B(u2__abc_44228_n8784), .Y(u2__abc_44228_n8786_1) );
  AND2X2 AND2X2_3315 ( .A(u2__abc_44228_n8787), .B(u2__abc_44228_n4058), .Y(u2__abc_44228_n8788) );
  AND2X2 AND2X2_3316 ( .A(u2__abc_44228_n7547_bF_buf41), .B(u2__abc_44228_n8789), .Y(u2__abc_44228_n8790) );
  AND2X2 AND2X2_3317 ( .A(u2__abc_44228_n7548_1_bF_buf42), .B(u2_remHi_71_), .Y(u2__abc_44228_n8791_1) );
  AND2X2 AND2X2_3318 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n4069), .Y(u2__abc_44228_n8794) );
  AND2X2 AND2X2_3319 ( .A(u2__abc_44228_n8795), .B(u2__abc_44228_n2972_bF_buf32), .Y(u2__abc_44228_n8796_1) );
  AND2X2 AND2X2_332 ( .A(_abc_64468_n1571), .B(_abc_64468_n1569), .Y(_abc_64468_n1572) );
  AND2X2 AND2X2_3320 ( .A(u2__abc_44228_n8793), .B(u2__abc_44228_n8796_1), .Y(u2__abc_44228_n8797_1) );
  AND2X2 AND2X2_3321 ( .A(u2__abc_44228_n8798), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_remHi_73__FF_INPUT) );
  AND2X2 AND2X2_3322 ( .A(u2__abc_44228_n3062_bF_buf18), .B(u2_remHi_74_), .Y(u2__abc_44228_n8800) );
  AND2X2 AND2X2_3323 ( .A(u2__abc_44228_n7548_1_bF_buf41), .B(u2_remHi_72_), .Y(u2__abc_44228_n8801) );
  AND2X2 AND2X2_3324 ( .A(u2__abc_44228_n8768), .B(u2__abc_44228_n4065), .Y(u2__abc_44228_n8802_1) );
  AND2X2 AND2X2_3325 ( .A(u2__abc_44228_n8803), .B(u2__abc_44228_n4078), .Y(u2__abc_44228_n8805) );
  AND2X2 AND2X2_3326 ( .A(u2__abc_44228_n8806), .B(u2__abc_44228_n8804), .Y(u2__abc_44228_n8807_1) );
  AND2X2 AND2X2_3327 ( .A(u2__abc_44228_n7547_bF_buf40), .B(u2__abc_44228_n8807_1), .Y(u2__abc_44228_n8808_1) );
  AND2X2 AND2X2_3328 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n4039), .Y(u2__abc_44228_n8811) );
  AND2X2 AND2X2_3329 ( .A(u2__abc_44228_n8812), .B(u2__abc_44228_n2972_bF_buf31), .Y(u2__abc_44228_n8813_1) );
  AND2X2 AND2X2_333 ( .A(_abc_64468_n1567), .B(_abc_64468_n1573), .Y(_abc_64468_n1574) );
  AND2X2 AND2X2_3330 ( .A(u2__abc_44228_n8810), .B(u2__abc_44228_n8813_1), .Y(u2__abc_44228_n8814) );
  AND2X2 AND2X2_3331 ( .A(u2__abc_44228_n8815), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_remHi_74__FF_INPUT) );
  AND2X2 AND2X2_3332 ( .A(u2__abc_44228_n3062_bF_buf17), .B(u2_remHi_75_), .Y(u2__abc_44228_n8817) );
  AND2X2 AND2X2_3333 ( .A(u2__abc_44228_n7548_1_bF_buf40), .B(u2_remHi_73_), .Y(u2__abc_44228_n8818_1) );
  AND2X2 AND2X2_3334 ( .A(u2__abc_44228_n8806), .B(u2__abc_44228_n4162), .Y(u2__abc_44228_n8820) );
  AND2X2 AND2X2_3335 ( .A(u2__abc_44228_n8821), .B(u2__abc_44228_n8819_1), .Y(u2__abc_44228_n8822) );
  AND2X2 AND2X2_3336 ( .A(u2__abc_44228_n8820), .B(u2__abc_44228_n4072), .Y(u2__abc_44228_n8823) );
  AND2X2 AND2X2_3337 ( .A(u2__abc_44228_n7547_bF_buf39), .B(u2__abc_44228_n8824_1), .Y(u2__abc_44228_n8825) );
  AND2X2 AND2X2_3338 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n4046), .Y(u2__abc_44228_n8828) );
  AND2X2 AND2X2_3339 ( .A(u2__abc_44228_n8829_1), .B(u2__abc_44228_n2972_bF_buf30), .Y(u2__abc_44228_n8830_1) );
  AND2X2 AND2X2_334 ( .A(_abc_64468_n1561), .B(_abc_64468_n1572), .Y(_abc_64468_n1575) );
  AND2X2 AND2X2_3340 ( .A(u2__abc_44228_n8827), .B(u2__abc_44228_n8830_1), .Y(u2__abc_44228_n8831) );
  AND2X2 AND2X2_3341 ( .A(u2__abc_44228_n8832), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_remHi_75__FF_INPUT) );
  AND2X2 AND2X2_3342 ( .A(u2__abc_44228_n3062_bF_buf16), .B(u2_remHi_76_), .Y(u2__abc_44228_n8834) );
  AND2X2 AND2X2_3343 ( .A(u2__abc_44228_n8806), .B(u2__abc_44228_n4163), .Y(u2__abc_44228_n8835_1) );
  AND2X2 AND2X2_3344 ( .A(u2__abc_44228_n8837), .B(u2__abc_44228_n4042), .Y(u2__abc_44228_n8838) );
  AND2X2 AND2X2_3345 ( .A(u2__abc_44228_n8839), .B(u2__abc_44228_n8840_1), .Y(u2__abc_44228_n8841_1) );
  AND2X2 AND2X2_3346 ( .A(u2__abc_44228_n8842), .B(u2__abc_44228_n8843), .Y(u2__abc_44228_n8844) );
  AND2X2 AND2X2_3347 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n4032), .Y(u2__abc_44228_n8846_1) );
  AND2X2 AND2X2_3348 ( .A(u2__abc_44228_n8847), .B(u2__abc_44228_n2972_bF_buf29), .Y(u2__abc_44228_n8848) );
  AND2X2 AND2X2_3349 ( .A(u2__abc_44228_n8845), .B(u2__abc_44228_n8848), .Y(u2__abc_44228_n8849) );
  AND2X2 AND2X2_335 ( .A(_abc_64468_n1576), .B(_abc_64468_n753_bF_buf0), .Y(_abc_64468_n1577) );
  AND2X2 AND2X2_3350 ( .A(u2__abc_44228_n8850), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_remHi_76__FF_INPUT) );
  AND2X2 AND2X2_3351 ( .A(u2__abc_44228_n3062_bF_buf15), .B(u2_remHi_77_), .Y(u2__abc_44228_n8852_1) );
  AND2X2 AND2X2_3352 ( .A(u2__abc_44228_n8839), .B(u2__abc_44228_n4169), .Y(u2__abc_44228_n8853) );
  AND2X2 AND2X2_3353 ( .A(u2__abc_44228_n8857_1), .B(u2__abc_44228_n7547_bF_buf37), .Y(u2__abc_44228_n8858) );
  AND2X2 AND2X2_3354 ( .A(u2__abc_44228_n8858), .B(u2__abc_44228_n8855), .Y(u2__abc_44228_n8859) );
  AND2X2 AND2X2_3355 ( .A(u2__abc_44228_n7548_1_bF_buf38), .B(u2_remHi_75_), .Y(u2__abc_44228_n8860) );
  AND2X2 AND2X2_3356 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n4026), .Y(u2__abc_44228_n8863_1) );
  AND2X2 AND2X2_3357 ( .A(u2__abc_44228_n8864), .B(u2__abc_44228_n2972_bF_buf28), .Y(u2__abc_44228_n8865) );
  AND2X2 AND2X2_3358 ( .A(u2__abc_44228_n8862_1), .B(u2__abc_44228_n8865), .Y(u2__abc_44228_n8866) );
  AND2X2 AND2X2_3359 ( .A(u2__abc_44228_n8867), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_remHi_77__FF_INPUT) );
  AND2X2 AND2X2_336 ( .A(_abc_64468_n1554), .B(\a[118] ), .Y(_abc_64468_n1581) );
  AND2X2 AND2X2_3360 ( .A(u2__abc_44228_n3062_bF_buf14), .B(u2_remHi_78_), .Y(u2__abc_44228_n8869) );
  AND2X2 AND2X2_3361 ( .A(u2__abc_44228_n8839), .B(u2__abc_44228_n4170), .Y(u2__abc_44228_n8870) );
  AND2X2 AND2X2_3362 ( .A(u2__abc_44228_n8872), .B(u2__abc_44228_n4035), .Y(u2__abc_44228_n8874_1) );
  AND2X2 AND2X2_3363 ( .A(u2__abc_44228_n8875), .B(u2__abc_44228_n8873_1), .Y(u2__abc_44228_n8876) );
  AND2X2 AND2X2_3364 ( .A(u2__abc_44228_n8876), .B(u2__abc_44228_n7547_bF_buf36), .Y(u2__abc_44228_n8877) );
  AND2X2 AND2X2_3365 ( .A(u2__abc_44228_n7548_1_bF_buf37), .B(u2_remHi_76_), .Y(u2__abc_44228_n8878) );
  AND2X2 AND2X2_3366 ( .A(u2__abc_44228_n2983_bF_buf129), .B(u2__abc_44228_n4008), .Y(u2__abc_44228_n8881) );
  AND2X2 AND2X2_3367 ( .A(u2__abc_44228_n8882), .B(u2__abc_44228_n2972_bF_buf27), .Y(u2__abc_44228_n8883) );
  AND2X2 AND2X2_3368 ( .A(u2__abc_44228_n8880), .B(u2__abc_44228_n8883), .Y(u2__abc_44228_n8884_1) );
  AND2X2 AND2X2_3369 ( .A(u2__abc_44228_n8885_1), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_remHi_78__FF_INPUT) );
  AND2X2 AND2X2_337 ( .A(_abc_64468_n1581), .B(_abc_64468_n1580), .Y(_abc_64468_n1583) );
  AND2X2 AND2X2_3370 ( .A(u2__abc_44228_n3062_bF_buf13), .B(u2_remHi_79_), .Y(u2__abc_44228_n8887) );
  AND2X2 AND2X2_3371 ( .A(u2__abc_44228_n8875), .B(u2__abc_44228_n8889), .Y(u2__abc_44228_n8890_1) );
  AND2X2 AND2X2_3372 ( .A(u2__abc_44228_n8893), .B(u2__abc_44228_n7547_bF_buf35), .Y(u2__abc_44228_n8894) );
  AND2X2 AND2X2_3373 ( .A(u2__abc_44228_n8894), .B(u2__abc_44228_n8891), .Y(u2__abc_44228_n8895_1) );
  AND2X2 AND2X2_3374 ( .A(u2__abc_44228_n7548_1_bF_buf36), .B(u2_remHi_77_), .Y(u2__abc_44228_n8896_1) );
  AND2X2 AND2X2_3375 ( .A(u2__abc_44228_n2983_bF_buf127), .B(u2__abc_44228_n4015_1), .Y(u2__abc_44228_n8899) );
  AND2X2 AND2X2_3376 ( .A(u2__abc_44228_n8900), .B(u2__abc_44228_n2972_bF_buf26), .Y(u2__abc_44228_n8901_1) );
  AND2X2 AND2X2_3377 ( .A(u2__abc_44228_n8898), .B(u2__abc_44228_n8901_1), .Y(u2__abc_44228_n8902) );
  AND2X2 AND2X2_3378 ( .A(u2__abc_44228_n8903), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_remHi_79__FF_INPUT) );
  AND2X2 AND2X2_3379 ( .A(u2__abc_44228_n3062_bF_buf12), .B(u2_remHi_80_), .Y(u2__abc_44228_n8905) );
  AND2X2 AND2X2_338 ( .A(_abc_64468_n1584), .B(_abc_64468_n1582), .Y(_abc_64468_n1585) );
  AND2X2 AND2X2_3380 ( .A(u2__abc_44228_n3664), .B(u2__abc_44228_n4138_1), .Y(u2__abc_44228_n8906_1) );
  AND2X2 AND2X2_3381 ( .A(u2__abc_44228_n8907_1), .B(u2__abc_44228_n4011), .Y(u2__abc_44228_n8908) );
  AND2X2 AND2X2_3382 ( .A(u2__abc_44228_n8909), .B(u2__abc_44228_n8910), .Y(u2__abc_44228_n8911) );
  AND2X2 AND2X2_3383 ( .A(u2__abc_44228_n7547_bF_buf34), .B(u2__abc_44228_n8911), .Y(u2__abc_44228_n8912_1) );
  AND2X2 AND2X2_3384 ( .A(u2__abc_44228_n7548_1_bF_buf35), .B(u2_remHi_78_), .Y(u2__abc_44228_n8913) );
  AND2X2 AND2X2_3385 ( .A(u2__abc_44228_n2983_bF_buf125), .B(u2__abc_44228_n4001), .Y(u2__abc_44228_n8916) );
  AND2X2 AND2X2_3386 ( .A(u2__abc_44228_n8917_1), .B(u2__abc_44228_n2972_bF_buf25), .Y(u2__abc_44228_n8918_1) );
  AND2X2 AND2X2_3387 ( .A(u2__abc_44228_n8915), .B(u2__abc_44228_n8918_1), .Y(u2__abc_44228_n8919) );
  AND2X2 AND2X2_3388 ( .A(u2__abc_44228_n8920), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_remHi_80__FF_INPUT) );
  AND2X2 AND2X2_3389 ( .A(u2__abc_44228_n3062_bF_buf11), .B(u2_remHi_81_), .Y(u2__abc_44228_n8922) );
  AND2X2 AND2X2_339 ( .A(_abc_64468_n1579), .B(_abc_64468_n1586), .Y(_abc_64468_n1587) );
  AND2X2 AND2X2_3390 ( .A(u2__abc_44228_n8909), .B(u2__abc_44228_n4179), .Y(u2__abc_44228_n8924) );
  AND2X2 AND2X2_3391 ( .A(u2__abc_44228_n8925), .B(u2__abc_44228_n8923_1), .Y(u2__abc_44228_n8926) );
  AND2X2 AND2X2_3392 ( .A(u2__abc_44228_n8924), .B(u2__abc_44228_n4018), .Y(u2__abc_44228_n8927) );
  AND2X2 AND2X2_3393 ( .A(u2__abc_44228_n7547_bF_buf33), .B(u2__abc_44228_n8928_1), .Y(u2__abc_44228_n8929_1) );
  AND2X2 AND2X2_3394 ( .A(u2__abc_44228_n7548_1_bF_buf34), .B(u2_remHi_79_), .Y(u2__abc_44228_n8930) );
  AND2X2 AND2X2_3395 ( .A(u2__abc_44228_n2983_bF_buf123), .B(u2__abc_44228_n3995_1), .Y(u2__abc_44228_n8933) );
  AND2X2 AND2X2_3396 ( .A(u2__abc_44228_n8934_1), .B(u2__abc_44228_n2972_bF_buf24), .Y(u2__abc_44228_n8935) );
  AND2X2 AND2X2_3397 ( .A(u2__abc_44228_n8932), .B(u2__abc_44228_n8935), .Y(u2__abc_44228_n8936) );
  AND2X2 AND2X2_3398 ( .A(u2__abc_44228_n8937), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_remHi_81__FF_INPUT) );
  AND2X2 AND2X2_3399 ( .A(u2__abc_44228_n3062_bF_buf10), .B(u2_remHi_82_), .Y(u2__abc_44228_n8939_1) );
  AND2X2 AND2X2_34 ( .A(_abc_64468_n753_bF_buf8), .B(sqrto_33_), .Y(_auto_iopadmap_cc_313_execute_65414_69_) );
  AND2X2 AND2X2_340 ( .A(_abc_64468_n1575), .B(_abc_64468_n1585), .Y(_abc_64468_n1588) );
  AND2X2 AND2X2_3400 ( .A(u2__abc_44228_n8909), .B(u2__abc_44228_n4180), .Y(u2__abc_44228_n8940_1) );
  AND2X2 AND2X2_3401 ( .A(u2__abc_44228_n8942), .B(u2__abc_44228_n4004), .Y(u2__abc_44228_n8944) );
  AND2X2 AND2X2_3402 ( .A(u2__abc_44228_n8945_1), .B(u2__abc_44228_n8943), .Y(u2__abc_44228_n8946) );
  AND2X2 AND2X2_3403 ( .A(u2__abc_44228_n7547_bF_buf32), .B(u2__abc_44228_n8946), .Y(u2__abc_44228_n8947) );
  AND2X2 AND2X2_3404 ( .A(u2__abc_44228_n7548_1_bF_buf33), .B(u2_remHi_80_), .Y(u2__abc_44228_n8948) );
  AND2X2 AND2X2_3405 ( .A(u2__abc_44228_n2983_bF_buf121), .B(u2__abc_44228_n3979), .Y(u2__abc_44228_n8951_1) );
  AND2X2 AND2X2_3406 ( .A(u2__abc_44228_n8952), .B(u2__abc_44228_n2972_bF_buf23), .Y(u2__abc_44228_n8953) );
  AND2X2 AND2X2_3407 ( .A(u2__abc_44228_n8950_1), .B(u2__abc_44228_n8953), .Y(u2__abc_44228_n8954) );
  AND2X2 AND2X2_3408 ( .A(u2__abc_44228_n8955), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_remHi_82__FF_INPUT) );
  AND2X2 AND2X2_3409 ( .A(u2__abc_44228_n3062_bF_buf9), .B(u2_remHi_83_), .Y(u2__abc_44228_n8957) );
  AND2X2 AND2X2_341 ( .A(_abc_64468_n1589), .B(_abc_64468_n753_bF_buf13), .Y(_abc_64468_n1590) );
  AND2X2 AND2X2_3410 ( .A(u2__abc_44228_n8962_1), .B(u2__abc_44228_n8959), .Y(u2__abc_44228_n8963) );
  AND2X2 AND2X2_3411 ( .A(u2__abc_44228_n8964), .B(u2__abc_44228_n8965), .Y(u2__abc_44228_n8966) );
  AND2X2 AND2X2_3412 ( .A(u2__abc_44228_n2983_bF_buf119), .B(u2__abc_44228_n3986_1), .Y(u2__abc_44228_n8968) );
  AND2X2 AND2X2_3413 ( .A(u2__abc_44228_n8969), .B(u2__abc_44228_n2972_bF_buf22), .Y(u2__abc_44228_n8970) );
  AND2X2 AND2X2_3414 ( .A(u2__abc_44228_n8967_1), .B(u2__abc_44228_n8970), .Y(u2__abc_44228_n8971) );
  AND2X2 AND2X2_3415 ( .A(u2__abc_44228_n8972_1), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_remHi_83__FF_INPUT) );
  AND2X2 AND2X2_3416 ( .A(u2__abc_44228_n3062_bF_buf8), .B(u2_remHi_84_), .Y(u2__abc_44228_n8974) );
  AND2X2 AND2X2_3417 ( .A(u2__abc_44228_n7548_1_bF_buf31), .B(u2_remHi_82_), .Y(u2__abc_44228_n8975) );
  AND2X2 AND2X2_3418 ( .A(u2__abc_44228_n8907_1), .B(u2__abc_44228_n4020), .Y(u2__abc_44228_n8976) );
  AND2X2 AND2X2_3419 ( .A(u2__abc_44228_n8977), .B(u2__abc_44228_n3982), .Y(u2__abc_44228_n8978_1) );
  AND2X2 AND2X2_342 ( .A(aNan_bF_buf1), .B(\a[118] ), .Y(_abc_64468_n1591) );
  AND2X2 AND2X2_3420 ( .A(u2__abc_44228_n8979), .B(u2__abc_44228_n8980), .Y(u2__abc_44228_n8981) );
  AND2X2 AND2X2_3421 ( .A(u2__abc_44228_n7547_bF_buf30), .B(u2__abc_44228_n8981), .Y(u2__abc_44228_n8982) );
  AND2X2 AND2X2_3422 ( .A(u2__abc_44228_n2983_bF_buf117), .B(u2__abc_44228_n3972), .Y(u2__abc_44228_n8985) );
  AND2X2 AND2X2_3423 ( .A(u2__abc_44228_n8986), .B(u2__abc_44228_n2972_bF_buf21), .Y(u2__abc_44228_n8987) );
  AND2X2 AND2X2_3424 ( .A(u2__abc_44228_n8984_1), .B(u2__abc_44228_n8987), .Y(u2__abc_44228_n8988) );
  AND2X2 AND2X2_3425 ( .A(u2__abc_44228_n8989_1), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_remHi_84__FF_INPUT) );
  AND2X2 AND2X2_3426 ( .A(u2__abc_44228_n3062_bF_buf7), .B(u2_remHi_85_), .Y(u2__abc_44228_n8991) );
  AND2X2 AND2X2_3427 ( .A(u2__abc_44228_n8979), .B(u2__abc_44228_n4188), .Y(u2__abc_44228_n8993) );
  AND2X2 AND2X2_3428 ( .A(u2__abc_44228_n8996), .B(u2__abc_44228_n8994_1), .Y(u2__abc_44228_n8997) );
  AND2X2 AND2X2_3429 ( .A(u2__abc_44228_n8998), .B(u2__abc_44228_n8999), .Y(u2__abc_44228_n9000_1) );
  AND2X2 AND2X2_343 ( .A(aNan_bF_buf0), .B(\a[119] ), .Y(_abc_64468_n1593) );
  AND2X2 AND2X2_3430 ( .A(u2__abc_44228_n2983_bF_buf115), .B(u2__abc_44228_n3966), .Y(u2__abc_44228_n9002) );
  AND2X2 AND2X2_3431 ( .A(u2__abc_44228_n9003), .B(u2__abc_44228_n2972_bF_buf20), .Y(u2__abc_44228_n9004) );
  AND2X2 AND2X2_3432 ( .A(u2__abc_44228_n9001), .B(u2__abc_44228_n9004), .Y(u2__abc_44228_n9005_1) );
  AND2X2 AND2X2_3433 ( .A(u2__abc_44228_n9006_1), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_remHi_85__FF_INPUT) );
  AND2X2 AND2X2_3434 ( .A(u2__abc_44228_n3062_bF_buf6), .B(u2_remHi_86_), .Y(u2__abc_44228_n9008) );
  AND2X2 AND2X2_3435 ( .A(u2__abc_44228_n8977), .B(u2__abc_44228_n3990), .Y(u2__abc_44228_n9009) );
  AND2X2 AND2X2_3436 ( .A(u2__abc_44228_n9010), .B(u2__abc_44228_n3975), .Y(u2__abc_44228_n9012) );
  AND2X2 AND2X2_3437 ( .A(u2__abc_44228_n9013), .B(u2__abc_44228_n9011_1), .Y(u2__abc_44228_n9014) );
  AND2X2 AND2X2_3438 ( .A(u2__abc_44228_n9015), .B(u2__abc_44228_n9016_1), .Y(u2__abc_44228_n9017_1) );
  AND2X2 AND2X2_3439 ( .A(u2__abc_44228_n2983_bF_buf113), .B(u2__abc_44228_n3949_1), .Y(u2__abc_44228_n9019) );
  AND2X2 AND2X2_344 ( .A(_abc_64468_n1581), .B(\a[119] ), .Y(_abc_64468_n1596) );
  AND2X2 AND2X2_3440 ( .A(u2__abc_44228_n9020), .B(u2__abc_44228_n2972_bF_buf19), .Y(u2__abc_44228_n9021) );
  AND2X2 AND2X2_3441 ( .A(u2__abc_44228_n9018), .B(u2__abc_44228_n9021), .Y(u2__abc_44228_n9022_1) );
  AND2X2 AND2X2_3442 ( .A(u2__abc_44228_n9023), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_remHi_86__FF_INPUT) );
  AND2X2 AND2X2_3443 ( .A(u2__abc_44228_n3062_bF_buf5), .B(u2_remHi_87_), .Y(u2__abc_44228_n9025) );
  AND2X2 AND2X2_3444 ( .A(u2__abc_44228_n9030), .B(u2__abc_44228_n9027_1), .Y(u2__abc_44228_n9031) );
  AND2X2 AND2X2_3445 ( .A(u2__abc_44228_n9031), .B(u2__abc_44228_n7547_bF_buf27), .Y(u2__abc_44228_n9032) );
  AND2X2 AND2X2_3446 ( .A(u2__abc_44228_n7548_1_bF_buf28), .B(u2_remHi_85_), .Y(u2__abc_44228_n9033_1) );
  AND2X2 AND2X2_3447 ( .A(u2__abc_44228_n2983_bF_buf111), .B(u2__abc_44228_n3956), .Y(u2__abc_44228_n9036) );
  AND2X2 AND2X2_3448 ( .A(u2__abc_44228_n9037), .B(u2__abc_44228_n2972_bF_buf18), .Y(u2__abc_44228_n9038_1) );
  AND2X2 AND2X2_3449 ( .A(u2__abc_44228_n9035), .B(u2__abc_44228_n9038_1), .Y(u2__abc_44228_n9039_1) );
  AND2X2 AND2X2_345 ( .A(_abc_64468_n1596), .B(_abc_64468_n1595), .Y(_abc_64468_n1598) );
  AND2X2 AND2X2_3450 ( .A(u2__abc_44228_n9040), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_remHi_87__FF_INPUT) );
  AND2X2 AND2X2_3451 ( .A(u2__abc_44228_n3062_bF_buf4), .B(u2_remHi_88_), .Y(u2__abc_44228_n9042) );
  AND2X2 AND2X2_3452 ( .A(u2__abc_44228_n7548_1_bF_buf27), .B(u2_remHi_86_), .Y(u2__abc_44228_n9043) );
  AND2X2 AND2X2_3453 ( .A(u2__abc_44228_n8907_1), .B(u2__abc_44228_n4021), .Y(u2__abc_44228_n9044_1) );
  AND2X2 AND2X2_3454 ( .A(u2__abc_44228_n9045), .B(u2__abc_44228_n3952), .Y(u2__abc_44228_n9047) );
  AND2X2 AND2X2_3455 ( .A(u2__abc_44228_n9048), .B(u2__abc_44228_n9046), .Y(u2__abc_44228_n9049_1) );
  AND2X2 AND2X2_3456 ( .A(u2__abc_44228_n7547_bF_buf26), .B(u2__abc_44228_n9049_1), .Y(u2__abc_44228_n9050_1) );
  AND2X2 AND2X2_3457 ( .A(u2__abc_44228_n2983_bF_buf109), .B(u2__abc_44228_n3942), .Y(u2__abc_44228_n9053) );
  AND2X2 AND2X2_3458 ( .A(u2__abc_44228_n9054), .B(u2__abc_44228_n2972_bF_buf17), .Y(u2__abc_44228_n9055_1) );
  AND2X2 AND2X2_3459 ( .A(u2__abc_44228_n9052), .B(u2__abc_44228_n9055_1), .Y(u2__abc_44228_n9056) );
  AND2X2 AND2X2_346 ( .A(_abc_64468_n1599), .B(_abc_64468_n1597), .Y(_abc_64468_n1600) );
  AND2X2 AND2X2_3460 ( .A(u2__abc_44228_n9057), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_remHi_88__FF_INPUT) );
  AND2X2 AND2X2_3461 ( .A(u2__abc_44228_n3062_bF_buf3), .B(u2_remHi_89_), .Y(u2__abc_44228_n9059) );
  AND2X2 AND2X2_3462 ( .A(u2__abc_44228_n7548_1_bF_buf26), .B(u2_remHi_87_), .Y(u2__abc_44228_n9060_1) );
  AND2X2 AND2X2_3463 ( .A(u2__abc_44228_n9048), .B(u2__abc_44228_n4198), .Y(u2__abc_44228_n9062) );
  AND2X2 AND2X2_3464 ( .A(u2__abc_44228_n9063), .B(u2__abc_44228_n9061_1), .Y(u2__abc_44228_n9064) );
  AND2X2 AND2X2_3465 ( .A(u2__abc_44228_n9062), .B(u2__abc_44228_n3959), .Y(u2__abc_44228_n9065) );
  AND2X2 AND2X2_3466 ( .A(u2__abc_44228_n7547_bF_buf25), .B(u2__abc_44228_n9066_1), .Y(u2__abc_44228_n9067) );
  AND2X2 AND2X2_3467 ( .A(u2__abc_44228_n2983_bF_buf107), .B(u2__abc_44228_n3936), .Y(u2__abc_44228_n9070) );
  AND2X2 AND2X2_3468 ( .A(u2__abc_44228_n9071_1), .B(u2__abc_44228_n2972_bF_buf16), .Y(u2__abc_44228_n9072_1) );
  AND2X2 AND2X2_3469 ( .A(u2__abc_44228_n9069), .B(u2__abc_44228_n9072_1), .Y(u2__abc_44228_n9073) );
  AND2X2 AND2X2_347 ( .A(_abc_64468_n1594), .B(_abc_64468_n1601), .Y(_abc_64468_n1602) );
  AND2X2 AND2X2_3470 ( .A(u2__abc_44228_n9074), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_remHi_89__FF_INPUT) );
  AND2X2 AND2X2_3471 ( .A(u2__abc_44228_n3062_bF_buf2), .B(u2_remHi_90_), .Y(u2__abc_44228_n9076) );
  AND2X2 AND2X2_3472 ( .A(u2__abc_44228_n9048), .B(u2__abc_44228_n4199), .Y(u2__abc_44228_n9077_1) );
  AND2X2 AND2X2_3473 ( .A(u2__abc_44228_n9079), .B(u2__abc_44228_n3945), .Y(u2__abc_44228_n9081) );
  AND2X2 AND2X2_3474 ( .A(u2__abc_44228_n9082_1), .B(u2__abc_44228_n9080), .Y(u2__abc_44228_n9083_1) );
  AND2X2 AND2X2_3475 ( .A(u2__abc_44228_n9084), .B(u2__abc_44228_n9085), .Y(u2__abc_44228_n9086) );
  AND2X2 AND2X2_3476 ( .A(u2__abc_44228_n2983_bF_buf105), .B(u2__abc_44228_n3920), .Y(u2__abc_44228_n9088_1) );
  AND2X2 AND2X2_3477 ( .A(u2__abc_44228_n9089), .B(u2__abc_44228_n2972_bF_buf15), .Y(u2__abc_44228_n9090) );
  AND2X2 AND2X2_3478 ( .A(u2__abc_44228_n9087), .B(u2__abc_44228_n9090), .Y(u2__abc_44228_n9091) );
  AND2X2 AND2X2_3479 ( .A(u2__abc_44228_n9092), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_remHi_90__FF_INPUT) );
  AND2X2 AND2X2_348 ( .A(_abc_64468_n1588), .B(_abc_64468_n1600), .Y(_abc_64468_n1603) );
  AND2X2 AND2X2_3480 ( .A(u2__abc_44228_n3062_bF_buf1), .B(u2_remHi_91_), .Y(u2__abc_44228_n9094_1) );
  AND2X2 AND2X2_3481 ( .A(u2__abc_44228_n9099_1), .B(u2__abc_44228_n7547_bF_buf23), .Y(u2__abc_44228_n9100) );
  AND2X2 AND2X2_3482 ( .A(u2__abc_44228_n9100), .B(u2__abc_44228_n9098), .Y(u2__abc_44228_n9101) );
  AND2X2 AND2X2_3483 ( .A(u2__abc_44228_n7548_1_bF_buf24), .B(u2_remHi_89_), .Y(u2__abc_44228_n9102) );
  AND2X2 AND2X2_3484 ( .A(u2__abc_44228_n2983_bF_buf103), .B(u2__abc_44228_n3927), .Y(u2__abc_44228_n9105_1) );
  AND2X2 AND2X2_3485 ( .A(u2__abc_44228_n9106), .B(u2__abc_44228_n2972_bF_buf14), .Y(u2__abc_44228_n9107) );
  AND2X2 AND2X2_3486 ( .A(u2__abc_44228_n9104_1), .B(u2__abc_44228_n9107), .Y(u2__abc_44228_n9108) );
  AND2X2 AND2X2_3487 ( .A(u2__abc_44228_n9109), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_remHi_91__FF_INPUT) );
  AND2X2 AND2X2_3488 ( .A(u2__abc_44228_n3062_bF_buf0), .B(u2_remHi_92_), .Y(u2__abc_44228_n9111) );
  AND2X2 AND2X2_3489 ( .A(u2__abc_44228_n9045), .B(u2__abc_44228_n3961), .Y(u2__abc_44228_n9112) );
  AND2X2 AND2X2_349 ( .A(_abc_64468_n1604), .B(_abc_64468_n753_bF_buf12), .Y(_abc_64468_n1605) );
  AND2X2 AND2X2_3490 ( .A(u2__abc_44228_n9113), .B(u2__abc_44228_n3923), .Y(u2__abc_44228_n9114) );
  AND2X2 AND2X2_3491 ( .A(u2__abc_44228_n9115_1), .B(u2__abc_44228_n9116_1), .Y(u2__abc_44228_n9117) );
  AND2X2 AND2X2_3492 ( .A(u2__abc_44228_n9118), .B(u2__abc_44228_n9119), .Y(u2__abc_44228_n9120) );
  AND2X2 AND2X2_3493 ( .A(u2__abc_44228_n2983_bF_buf101), .B(u2__abc_44228_n3913), .Y(u2__abc_44228_n9122) );
  AND2X2 AND2X2_3494 ( .A(u2__abc_44228_n9123), .B(u2__abc_44228_n2972_bF_buf13), .Y(u2__abc_44228_n9124) );
  AND2X2 AND2X2_3495 ( .A(u2__abc_44228_n9121_1), .B(u2__abc_44228_n9124), .Y(u2__abc_44228_n9125) );
  AND2X2 AND2X2_3496 ( .A(u2__abc_44228_n9126_1), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_remHi_92__FF_INPUT) );
  AND2X2 AND2X2_3497 ( .A(u2__abc_44228_n3062_bF_buf92), .B(u2_remHi_93_), .Y(u2__abc_44228_n9128) );
  AND2X2 AND2X2_3498 ( .A(u2__abc_44228_n9115_1), .B(u2__abc_44228_n4207), .Y(u2__abc_44228_n9129) );
  AND2X2 AND2X2_3499 ( .A(u2__abc_44228_n9129), .B(u2__abc_44228_n3930_1), .Y(u2__abc_44228_n9130) );
  AND2X2 AND2X2_35 ( .A(_abc_64468_n753_bF_buf7), .B(sqrto_34_), .Y(_auto_iopadmap_cc_313_execute_65414_70_) );
  AND2X2 AND2X2_350 ( .A(_abc_64468_n1596), .B(\a[120] ), .Y(_abc_64468_n1609) );
  AND2X2 AND2X2_3500 ( .A(u2__abc_44228_n9132_1), .B(u2__abc_44228_n9131), .Y(u2__abc_44228_n9133) );
  AND2X2 AND2X2_3501 ( .A(u2__abc_44228_n9134), .B(u2__abc_44228_n7547_bF_buf21), .Y(u2__abc_44228_n9135) );
  AND2X2 AND2X2_3502 ( .A(u2__abc_44228_n7548_1_bF_buf22), .B(u2_remHi_91_), .Y(u2__abc_44228_n9136) );
  AND2X2 AND2X2_3503 ( .A(u2__abc_44228_n2983_bF_buf99), .B(u2__abc_44228_n3907), .Y(u2__abc_44228_n9139) );
  AND2X2 AND2X2_3504 ( .A(u2__abc_44228_n9140), .B(u2__abc_44228_n2972_bF_buf12), .Y(u2__abc_44228_n9141) );
  AND2X2 AND2X2_3505 ( .A(u2__abc_44228_n9138_1), .B(u2__abc_44228_n9141), .Y(u2__abc_44228_n9142) );
  AND2X2 AND2X2_3506 ( .A(u2__abc_44228_n9143_1), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_remHi_93__FF_INPUT) );
  AND2X2 AND2X2_3507 ( .A(u2__abc_44228_n3062_bF_buf91), .B(u2_remHi_94_), .Y(u2__abc_44228_n9145) );
  AND2X2 AND2X2_3508 ( .A(u2__abc_44228_n9115_1), .B(u2__abc_44228_n4208), .Y(u2__abc_44228_n9146) );
  AND2X2 AND2X2_3509 ( .A(u2__abc_44228_n9148_1), .B(u2__abc_44228_n3916), .Y(u2__abc_44228_n9150) );
  AND2X2 AND2X2_351 ( .A(_abc_64468_n1609), .B(_abc_64468_n1608), .Y(_abc_64468_n1611) );
  AND2X2 AND2X2_3510 ( .A(u2__abc_44228_n9151), .B(u2__abc_44228_n9149_1), .Y(u2__abc_44228_n9152) );
  AND2X2 AND2X2_3511 ( .A(u2__abc_44228_n9152), .B(u2__abc_44228_n7547_bF_buf20), .Y(u2__abc_44228_n9153) );
  AND2X2 AND2X2_3512 ( .A(u2__abc_44228_n7548_1_bF_buf21), .B(u2_remHi_92_), .Y(u2__abc_44228_n9154_1) );
  AND2X2 AND2X2_3513 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n3888), .Y(u2__abc_44228_n9157) );
  AND2X2 AND2X2_3514 ( .A(u2__abc_44228_n9158), .B(u2__abc_44228_n2972_bF_buf11), .Y(u2__abc_44228_n9159_1) );
  AND2X2 AND2X2_3515 ( .A(u2__abc_44228_n9156), .B(u2__abc_44228_n9159_1), .Y(u2__abc_44228_n9160_1) );
  AND2X2 AND2X2_3516 ( .A(u2__abc_44228_n9161), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_remHi_94__FF_INPUT) );
  AND2X2 AND2X2_3517 ( .A(u2__abc_44228_n3062_bF_buf90), .B(u2_remHi_95_), .Y(u2__abc_44228_n9163) );
  AND2X2 AND2X2_3518 ( .A(u2__abc_44228_n9168), .B(u2__abc_44228_n7547_bF_buf19), .Y(u2__abc_44228_n9169) );
  AND2X2 AND2X2_3519 ( .A(u2__abc_44228_n9169), .B(u2__abc_44228_n9167), .Y(u2__abc_44228_n9170_1) );
  AND2X2 AND2X2_352 ( .A(_abc_64468_n1612), .B(_abc_64468_n1610), .Y(_abc_64468_n1613) );
  AND2X2 AND2X2_3520 ( .A(u2__abc_44228_n7548_1_bF_buf20), .B(u2_remHi_93_), .Y(u2__abc_44228_n9171_1) );
  AND2X2 AND2X2_3521 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n3895), .Y(u2__abc_44228_n9174) );
  AND2X2 AND2X2_3522 ( .A(u2__abc_44228_n9175), .B(u2__abc_44228_n2972_bF_buf10), .Y(u2__abc_44228_n9176_1) );
  AND2X2 AND2X2_3523 ( .A(u2__abc_44228_n9173), .B(u2__abc_44228_n9176_1), .Y(u2__abc_44228_n9177) );
  AND2X2 AND2X2_3524 ( .A(u2__abc_44228_n9178), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_remHi_95__FF_INPUT) );
  AND2X2 AND2X2_3525 ( .A(u2__abc_44228_n3062_bF_buf89), .B(u2_remHi_96_), .Y(u2__abc_44228_n9180) );
  AND2X2 AND2X2_3526 ( .A(u2__abc_44228_n3664), .B(u2__abc_44228_n4139), .Y(u2__abc_44228_n9181_1) );
  AND2X2 AND2X2_3527 ( .A(u2__abc_44228_n9182_1), .B(u2__abc_44228_n3891), .Y(u2__abc_44228_n9183) );
  AND2X2 AND2X2_3528 ( .A(u2__abc_44228_n9184), .B(u2__abc_44228_n9185), .Y(u2__abc_44228_n9186) );
  AND2X2 AND2X2_3529 ( .A(u2__abc_44228_n7547_bF_buf18), .B(u2__abc_44228_n9186), .Y(u2__abc_44228_n9187_1) );
  AND2X2 AND2X2_353 ( .A(_abc_64468_n1607), .B(_abc_64468_n1614), .Y(_abc_64468_n1615) );
  AND2X2 AND2X2_3530 ( .A(u2__abc_44228_n7548_1_bF_buf19), .B(u2_remHi_94_), .Y(u2__abc_44228_n9188) );
  AND2X2 AND2X2_3531 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n3881), .Y(u2__abc_44228_n9191) );
  AND2X2 AND2X2_3532 ( .A(u2__abc_44228_n9192_1), .B(u2__abc_44228_n2972_bF_buf9), .Y(u2__abc_44228_n9193_1) );
  AND2X2 AND2X2_3533 ( .A(u2__abc_44228_n9190), .B(u2__abc_44228_n9193_1), .Y(u2__abc_44228_n9194) );
  AND2X2 AND2X2_3534 ( .A(u2__abc_44228_n9195), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_remHi_96__FF_INPUT) );
  AND2X2 AND2X2_3535 ( .A(u2__abc_44228_n3062_bF_buf88), .B(u2_remHi_97_), .Y(u2__abc_44228_n9197) );
  AND2X2 AND2X2_3536 ( .A(u2__abc_44228_n9184), .B(u2__abc_44228_n4219), .Y(u2__abc_44228_n9198_1) );
  AND2X2 AND2X2_3537 ( .A(u2__abc_44228_n9198_1), .B(u2__abc_44228_n3898), .Y(u2__abc_44228_n9199) );
  AND2X2 AND2X2_3538 ( .A(u2__abc_44228_n9201), .B(u2__abc_44228_n9200), .Y(u2__abc_44228_n9202) );
  AND2X2 AND2X2_3539 ( .A(u2__abc_44228_n7547_bF_buf17), .B(u2__abc_44228_n9203_1), .Y(u2__abc_44228_n9204_1) );
  AND2X2 AND2X2_354 ( .A(_abc_64468_n1603), .B(_abc_64468_n1613), .Y(_abc_64468_n1616) );
  AND2X2 AND2X2_3540 ( .A(u2__abc_44228_n7548_1_bF_buf18), .B(u2_remHi_95_), .Y(u2__abc_44228_n9205) );
  AND2X2 AND2X2_3541 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n3875), .Y(u2__abc_44228_n9208) );
  AND2X2 AND2X2_3542 ( .A(u2__abc_44228_n9209_1), .B(u2__abc_44228_n2972_bF_buf8), .Y(u2__abc_44228_n9210) );
  AND2X2 AND2X2_3543 ( .A(u2__abc_44228_n9207), .B(u2__abc_44228_n9210), .Y(u2__abc_44228_n9211) );
  AND2X2 AND2X2_3544 ( .A(u2__abc_44228_n9212), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_remHi_97__FF_INPUT) );
  AND2X2 AND2X2_3545 ( .A(u2__abc_44228_n3062_bF_buf87), .B(u2_remHi_98_), .Y(u2__abc_44228_n9214_1) );
  AND2X2 AND2X2_3546 ( .A(u2__abc_44228_n9184), .B(u2__abc_44228_n4220), .Y(u2__abc_44228_n9215_1) );
  AND2X2 AND2X2_3547 ( .A(u2__abc_44228_n9217), .B(u2__abc_44228_n3884), .Y(u2__abc_44228_n9219) );
  AND2X2 AND2X2_3548 ( .A(u2__abc_44228_n9220_1), .B(u2__abc_44228_n9218), .Y(u2__abc_44228_n9221) );
  AND2X2 AND2X2_3549 ( .A(u2__abc_44228_n7547_bF_buf16), .B(u2__abc_44228_n9221), .Y(u2__abc_44228_n9222) );
  AND2X2 AND2X2_355 ( .A(_abc_64468_n1617), .B(_abc_64468_n753_bF_buf11), .Y(_abc_64468_n1618) );
  AND2X2 AND2X2_3550 ( .A(u2__abc_44228_n7548_1_bF_buf17), .B(u2_remHi_96_), .Y(u2__abc_44228_n9223) );
  AND2X2 AND2X2_3551 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n3859), .Y(u2__abc_44228_n9226_1) );
  AND2X2 AND2X2_3552 ( .A(u2__abc_44228_n9227), .B(u2__abc_44228_n2972_bF_buf7), .Y(u2__abc_44228_n9228) );
  AND2X2 AND2X2_3553 ( .A(u2__abc_44228_n9225_1), .B(u2__abc_44228_n9228), .Y(u2__abc_44228_n9229) );
  AND2X2 AND2X2_3554 ( .A(u2__abc_44228_n9230), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_remHi_98__FF_INPUT) );
  AND2X2 AND2X2_3555 ( .A(u2__abc_44228_n3062_bF_buf86), .B(u2_remHi_99_), .Y(u2__abc_44228_n9232) );
  AND2X2 AND2X2_3556 ( .A(u2__abc_44228_n9237_1), .B(u2__abc_44228_n9234), .Y(u2__abc_44228_n9238) );
  AND2X2 AND2X2_3557 ( .A(u2__abc_44228_n9239), .B(u2__abc_44228_n9240), .Y(u2__abc_44228_n9241) );
  AND2X2 AND2X2_3558 ( .A(u2__abc_44228_n2983_bF_buf88), .B(u2__abc_44228_n3866), .Y(u2__abc_44228_n9243) );
  AND2X2 AND2X2_3559 ( .A(u2__abc_44228_n9244), .B(u2__abc_44228_n2972_bF_buf6), .Y(u2__abc_44228_n9245) );
  AND2X2 AND2X2_356 ( .A(aNan_bF_buf10), .B(\a[120] ), .Y(_abc_64468_n1619) );
  AND2X2 AND2X2_3560 ( .A(u2__abc_44228_n9242_1), .B(u2__abc_44228_n9245), .Y(u2__abc_44228_n9246) );
  AND2X2 AND2X2_3561 ( .A(u2__abc_44228_n9247_1), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_remHi_99__FF_INPUT) );
  AND2X2 AND2X2_3562 ( .A(u2__abc_44228_n3062_bF_buf85), .B(u2_remHi_100_), .Y(u2__abc_44228_n9249) );
  AND2X2 AND2X2_3563 ( .A(u2__abc_44228_n7548_1_bF_buf15), .B(u2_remHi_98_), .Y(u2__abc_44228_n9250) );
  AND2X2 AND2X2_3564 ( .A(u2__abc_44228_n9182_1), .B(u2__abc_44228_n3900), .Y(u2__abc_44228_n9251) );
  AND2X2 AND2X2_3565 ( .A(u2__abc_44228_n9252), .B(u2__abc_44228_n3862), .Y(u2__abc_44228_n9253_1) );
  AND2X2 AND2X2_3566 ( .A(u2__abc_44228_n9254), .B(u2__abc_44228_n9255), .Y(u2__abc_44228_n9256) );
  AND2X2 AND2X2_3567 ( .A(u2__abc_44228_n7547_bF_buf14), .B(u2__abc_44228_n9256), .Y(u2__abc_44228_n9257) );
  AND2X2 AND2X2_3568 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n3852), .Y(u2__abc_44228_n9260) );
  AND2X2 AND2X2_3569 ( .A(u2__abc_44228_n9261), .B(u2__abc_44228_n2972_bF_buf5), .Y(u2__abc_44228_n9262) );
  AND2X2 AND2X2_357 ( .A(aNan_bF_buf9), .B(\a[121] ), .Y(_abc_64468_n1621) );
  AND2X2 AND2X2_3570 ( .A(u2__abc_44228_n9259_1), .B(u2__abc_44228_n9262), .Y(u2__abc_44228_n9263) );
  AND2X2 AND2X2_3571 ( .A(u2__abc_44228_n9264_1), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_remHi_100__FF_INPUT) );
  AND2X2 AND2X2_3572 ( .A(u2__abc_44228_n3062_bF_buf84), .B(u2_remHi_101_), .Y(u2__abc_44228_n9266) );
  AND2X2 AND2X2_3573 ( .A(u2__abc_44228_n9254), .B(u2__abc_44228_n4228), .Y(u2__abc_44228_n9268) );
  AND2X2 AND2X2_3574 ( .A(u2__abc_44228_n9271), .B(u2__abc_44228_n9269_1), .Y(u2__abc_44228_n9272) );
  AND2X2 AND2X2_3575 ( .A(u2__abc_44228_n9273), .B(u2__abc_44228_n9274), .Y(u2__abc_44228_n9275_1) );
  AND2X2 AND2X2_3576 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n3846), .Y(u2__abc_44228_n9277) );
  AND2X2 AND2X2_3577 ( .A(u2__abc_44228_n9278), .B(u2__abc_44228_n2972_bF_buf4), .Y(u2__abc_44228_n9279) );
  AND2X2 AND2X2_3578 ( .A(u2__abc_44228_n9276), .B(u2__abc_44228_n9279), .Y(u2__abc_44228_n9280_1) );
  AND2X2 AND2X2_3579 ( .A(u2__abc_44228_n9281_1), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_remHi_101__FF_INPUT) );
  AND2X2 AND2X2_358 ( .A(_abc_64468_n1609), .B(\a[121] ), .Y(_abc_64468_n1624) );
  AND2X2 AND2X2_3580 ( .A(u2__abc_44228_n3062_bF_buf83), .B(u2_remHi_102_), .Y(u2__abc_44228_n9283) );
  AND2X2 AND2X2_3581 ( .A(u2__abc_44228_n9252), .B(u2__abc_44228_n3870), .Y(u2__abc_44228_n9284) );
  AND2X2 AND2X2_3582 ( .A(u2__abc_44228_n9285), .B(u2__abc_44228_n3855), .Y(u2__abc_44228_n9287) );
  AND2X2 AND2X2_3583 ( .A(u2__abc_44228_n9288), .B(u2__abc_44228_n9286_1), .Y(u2__abc_44228_n9289) );
  AND2X2 AND2X2_3584 ( .A(u2__abc_44228_n9290), .B(u2__abc_44228_n9291_1), .Y(u2__abc_44228_n9292_1) );
  AND2X2 AND2X2_3585 ( .A(u2__abc_44228_n2983_bF_buf82), .B(u2__abc_44228_n3822), .Y(u2__abc_44228_n9294) );
  AND2X2 AND2X2_3586 ( .A(u2__abc_44228_n9295), .B(u2__abc_44228_n2972_bF_buf3), .Y(u2__abc_44228_n9296) );
  AND2X2 AND2X2_3587 ( .A(u2__abc_44228_n9293), .B(u2__abc_44228_n9296), .Y(u2__abc_44228_n9297_1) );
  AND2X2 AND2X2_3588 ( .A(u2__abc_44228_n9298), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_remHi_102__FF_INPUT) );
  AND2X2 AND2X2_3589 ( .A(u2__abc_44228_n3062_bF_buf82), .B(u2_remHi_103_), .Y(u2__abc_44228_n9300) );
  AND2X2 AND2X2_359 ( .A(_abc_64468_n1624), .B(_abc_64468_n1623), .Y(_abc_64468_n1626) );
  AND2X2 AND2X2_3590 ( .A(u2__abc_44228_n9305), .B(u2__abc_44228_n9302_1), .Y(u2__abc_44228_n9306) );
  AND2X2 AND2X2_3591 ( .A(u2__abc_44228_n9306), .B(u2__abc_44228_n7547_bF_buf11), .Y(u2__abc_44228_n9307) );
  AND2X2 AND2X2_3592 ( .A(u2__abc_44228_n7548_1_bF_buf12), .B(u2_remHi_101_), .Y(u2__abc_44228_n9308_1) );
  AND2X2 AND2X2_3593 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n3816_1), .Y(u2__abc_44228_n9311) );
  AND2X2 AND2X2_3594 ( .A(u2__abc_44228_n9312), .B(u2__abc_44228_n2972_bF_buf2), .Y(u2__abc_44228_n9313_1) );
  AND2X2 AND2X2_3595 ( .A(u2__abc_44228_n9310), .B(u2__abc_44228_n9313_1), .Y(u2__abc_44228_n9314_1) );
  AND2X2 AND2X2_3596 ( .A(u2__abc_44228_n9315), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_remHi_103__FF_INPUT) );
  AND2X2 AND2X2_3597 ( .A(u2__abc_44228_n3062_bF_buf81), .B(u2_remHi_104_), .Y(u2__abc_44228_n9317) );
  AND2X2 AND2X2_3598 ( .A(u2__abc_44228_n7548_1_bF_buf11), .B(u2_remHi_102_), .Y(u2__abc_44228_n9318) );
  AND2X2 AND2X2_3599 ( .A(u2__abc_44228_n9182_1), .B(u2__abc_44228_n3901), .Y(u2__abc_44228_n9319_1) );
  AND2X2 AND2X2_36 ( .A(_abc_64468_n753_bF_buf6), .B(sqrto_35_), .Y(_auto_iopadmap_cc_313_execute_65414_71_) );
  AND2X2 AND2X2_360 ( .A(_abc_64468_n1627), .B(_abc_64468_n1625), .Y(_abc_64468_n1628) );
  AND2X2 AND2X2_3600 ( .A(u2__abc_44228_n9320), .B(u2__abc_44228_n3825_1), .Y(u2__abc_44228_n9322) );
  AND2X2 AND2X2_3601 ( .A(u2__abc_44228_n9323), .B(u2__abc_44228_n9321), .Y(u2__abc_44228_n9324_1) );
  AND2X2 AND2X2_3602 ( .A(u2__abc_44228_n7547_bF_buf10), .B(u2__abc_44228_n9324_1), .Y(u2__abc_44228_n9325_1) );
  AND2X2 AND2X2_3603 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n3836), .Y(u2__abc_44228_n9328) );
  AND2X2 AND2X2_3604 ( .A(u2__abc_44228_n9329), .B(u2__abc_44228_n2972_bF_buf1), .Y(u2__abc_44228_n9330_1) );
  AND2X2 AND2X2_3605 ( .A(u2__abc_44228_n9327), .B(u2__abc_44228_n9330_1), .Y(u2__abc_44228_n9331) );
  AND2X2 AND2X2_3606 ( .A(u2__abc_44228_n9332), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_remHi_104__FF_INPUT) );
  AND2X2 AND2X2_3607 ( .A(u2__abc_44228_n3062_bF_buf80), .B(u2_remHi_105_), .Y(u2__abc_44228_n9334) );
  AND2X2 AND2X2_3608 ( .A(u2__abc_44228_n7548_1_bF_buf10), .B(u2_remHi_103_), .Y(u2__abc_44228_n9335_1) );
  AND2X2 AND2X2_3609 ( .A(u2__abc_44228_n9323), .B(u2__abc_44228_n4238), .Y(u2__abc_44228_n9337) );
  AND2X2 AND2X2_361 ( .A(_abc_64468_n1622), .B(_abc_64468_n1629), .Y(_abc_64468_n1630) );
  AND2X2 AND2X2_3610 ( .A(u2__abc_44228_n9338), .B(u2__abc_44228_n9336_1), .Y(u2__abc_44228_n9339) );
  AND2X2 AND2X2_3611 ( .A(u2__abc_44228_n9337), .B(u2__abc_44228_n3819), .Y(u2__abc_44228_n9340) );
  AND2X2 AND2X2_3612 ( .A(u2__abc_44228_n7547_bF_buf9), .B(u2__abc_44228_n9341_1), .Y(u2__abc_44228_n9342) );
  AND2X2 AND2X2_3613 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n3830), .Y(u2__abc_44228_n9345) );
  AND2X2 AND2X2_3614 ( .A(u2__abc_44228_n9346_1), .B(u2__abc_44228_n2972_bF_buf0), .Y(u2__abc_44228_n9347_1) );
  AND2X2 AND2X2_3615 ( .A(u2__abc_44228_n9344), .B(u2__abc_44228_n9347_1), .Y(u2__abc_44228_n9348) );
  AND2X2 AND2X2_3616 ( .A(u2__abc_44228_n9349), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_remHi_105__FF_INPUT) );
  AND2X2 AND2X2_3617 ( .A(u2__abc_44228_n3062_bF_buf79), .B(u2_remHi_106_), .Y(u2__abc_44228_n9351) );
  AND2X2 AND2X2_3618 ( .A(u2__abc_44228_n9320), .B(u2__abc_44228_n3826), .Y(u2__abc_44228_n9352_1) );
  AND2X2 AND2X2_3619 ( .A(u2__abc_44228_n9353), .B(u2__abc_44228_n3839), .Y(u2__abc_44228_n9355) );
  AND2X2 AND2X2_362 ( .A(_abc_64468_n1616), .B(_abc_64468_n1628), .Y(_abc_64468_n1631) );
  AND2X2 AND2X2_3620 ( .A(u2__abc_44228_n9356), .B(u2__abc_44228_n9354), .Y(u2__abc_44228_n9357_1) );
  AND2X2 AND2X2_3621 ( .A(u2__abc_44228_n9358_1), .B(u2__abc_44228_n9359), .Y(u2__abc_44228_n9360) );
  AND2X2 AND2X2_3622 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n3800), .Y(u2__abc_44228_n9362) );
  AND2X2 AND2X2_3623 ( .A(u2__abc_44228_n9363_1), .B(u2__abc_44228_n2972_bF_buf107), .Y(u2__abc_44228_n9364) );
  AND2X2 AND2X2_3624 ( .A(u2__abc_44228_n9361), .B(u2__abc_44228_n9364), .Y(u2__abc_44228_n9365) );
  AND2X2 AND2X2_3625 ( .A(u2__abc_44228_n9366), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_remHi_106__FF_INPUT) );
  AND2X2 AND2X2_3626 ( .A(u2__abc_44228_n3062_bF_buf78), .B(u2_remHi_107_), .Y(u2__abc_44228_n9368_1) );
  AND2X2 AND2X2_3627 ( .A(u2__abc_44228_n9356), .B(u2__abc_44228_n4243_1), .Y(u2__abc_44228_n9370) );
  AND2X2 AND2X2_3628 ( .A(u2__abc_44228_n9373), .B(u2__abc_44228_n9371), .Y(u2__abc_44228_n9374_1) );
  AND2X2 AND2X2_3629 ( .A(u2__abc_44228_n9374_1), .B(u2__abc_44228_n7547_bF_buf7), .Y(u2__abc_44228_n9375) );
  AND2X2 AND2X2_363 ( .A(_abc_64468_n1632), .B(_abc_64468_n753_bF_buf10), .Y(_abc_64468_n1633) );
  AND2X2 AND2X2_3630 ( .A(u2__abc_44228_n7548_1_bF_buf8), .B(u2_remHi_105_), .Y(u2__abc_44228_n9376) );
  AND2X2 AND2X2_3631 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n3807_1), .Y(u2__abc_44228_n9379_1) );
  AND2X2 AND2X2_3632 ( .A(u2__abc_44228_n9380_1), .B(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n9381) );
  AND2X2 AND2X2_3633 ( .A(u2__abc_44228_n9378), .B(u2__abc_44228_n9381), .Y(u2__abc_44228_n9382) );
  AND2X2 AND2X2_3634 ( .A(u2__abc_44228_n9383), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_remHi_107__FF_INPUT) );
  AND2X2 AND2X2_3635 ( .A(u2__abc_44228_n3062_bF_buf77), .B(u2_remHi_108_), .Y(u2__abc_44228_n9385_1) );
  AND2X2 AND2X2_3636 ( .A(u2__abc_44228_n9356), .B(u2__abc_44228_n4244), .Y(u2__abc_44228_n9386) );
  AND2X2 AND2X2_3637 ( .A(u2__abc_44228_n9388), .B(u2__abc_44228_n3803), .Y(u2__abc_44228_n9389) );
  AND2X2 AND2X2_3638 ( .A(u2__abc_44228_n9390_1), .B(u2__abc_44228_n9391_1), .Y(u2__abc_44228_n9392) );
  AND2X2 AND2X2_3639 ( .A(u2__abc_44228_n9393), .B(u2__abc_44228_n9394), .Y(u2__abc_44228_n9395) );
  AND2X2 AND2X2_364 ( .A(_abc_64468_n1624), .B(\a[122] ), .Y(_abc_64468_n1637) );
  AND2X2 AND2X2_3640 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n3793), .Y(u2__abc_44228_n9397) );
  AND2X2 AND2X2_3641 ( .A(u2__abc_44228_n9398), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n9399) );
  AND2X2 AND2X2_3642 ( .A(u2__abc_44228_n9396_1), .B(u2__abc_44228_n9399), .Y(u2__abc_44228_n9400) );
  AND2X2 AND2X2_3643 ( .A(u2__abc_44228_n9401_1), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_remHi_108__FF_INPUT) );
  AND2X2 AND2X2_3644 ( .A(u2__abc_44228_n3062_bF_buf76), .B(u2_remHi_109_), .Y(u2__abc_44228_n9403) );
  AND2X2 AND2X2_3645 ( .A(u2__abc_44228_n9390_1), .B(u2__abc_44228_n4249), .Y(u2__abc_44228_n9404) );
  AND2X2 AND2X2_3646 ( .A(u2__abc_44228_n9404), .B(u2__abc_44228_n3810), .Y(u2__abc_44228_n9405) );
  AND2X2 AND2X2_3647 ( .A(u2__abc_44228_n9407_1), .B(u2__abc_44228_n9406), .Y(u2__abc_44228_n9408) );
  AND2X2 AND2X2_3648 ( .A(u2__abc_44228_n9409), .B(u2__abc_44228_n7547_bF_buf5), .Y(u2__abc_44228_n9410) );
  AND2X2 AND2X2_3649 ( .A(u2__abc_44228_n7548_1_bF_buf6), .B(u2_remHi_107_), .Y(u2__abc_44228_n9411) );
  AND2X2 AND2X2_365 ( .A(_abc_64468_n1637), .B(_abc_64468_n1636), .Y(_abc_64468_n1639) );
  AND2X2 AND2X2_3650 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n3787), .Y(u2__abc_44228_n9414) );
  AND2X2 AND2X2_3651 ( .A(u2__abc_44228_n9415), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n9416) );
  AND2X2 AND2X2_3652 ( .A(u2__abc_44228_n9413_1), .B(u2__abc_44228_n9416), .Y(u2__abc_44228_n9417) );
  AND2X2 AND2X2_3653 ( .A(u2__abc_44228_n9418_1), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_remHi_109__FF_INPUT) );
  AND2X2 AND2X2_3654 ( .A(u2__abc_44228_n3062_bF_buf75), .B(u2_remHi_110_), .Y(u2__abc_44228_n9420) );
  AND2X2 AND2X2_3655 ( .A(u2__abc_44228_n9390_1), .B(u2__abc_44228_n4250), .Y(u2__abc_44228_n9421) );
  AND2X2 AND2X2_3656 ( .A(u2__abc_44228_n9423_1), .B(u2__abc_44228_n3796), .Y(u2__abc_44228_n9425) );
  AND2X2 AND2X2_3657 ( .A(u2__abc_44228_n9426), .B(u2__abc_44228_n9424_1), .Y(u2__abc_44228_n9427) );
  AND2X2 AND2X2_3658 ( .A(u2__abc_44228_n9427), .B(u2__abc_44228_n7547_bF_buf4), .Y(u2__abc_44228_n9428) );
  AND2X2 AND2X2_3659 ( .A(u2__abc_44228_n7548_1_bF_buf5), .B(u2_remHi_108_), .Y(u2__abc_44228_n9429_1) );
  AND2X2 AND2X2_366 ( .A(_abc_64468_n1640), .B(_abc_64468_n1638), .Y(_abc_64468_n1641) );
  AND2X2 AND2X2_3660 ( .A(u2__abc_44228_n2983_bF_buf67), .B(u2__abc_44228_n3769), .Y(u2__abc_44228_n9432) );
  AND2X2 AND2X2_3661 ( .A(u2__abc_44228_n9433), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n9434_1) );
  AND2X2 AND2X2_3662 ( .A(u2__abc_44228_n9431), .B(u2__abc_44228_n9434_1), .Y(u2__abc_44228_n9435_1) );
  AND2X2 AND2X2_3663 ( .A(u2__abc_44228_n9436), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_remHi_110__FF_INPUT) );
  AND2X2 AND2X2_3664 ( .A(u2__abc_44228_n3062_bF_buf74), .B(u2_remHi_111_), .Y(u2__abc_44228_n9438) );
  AND2X2 AND2X2_3665 ( .A(u2__abc_44228_n9443), .B(u2__abc_44228_n7547_bF_buf3), .Y(u2__abc_44228_n9444) );
  AND2X2 AND2X2_3666 ( .A(u2__abc_44228_n9444), .B(u2__abc_44228_n9442), .Y(u2__abc_44228_n9445_1) );
  AND2X2 AND2X2_3667 ( .A(u2__abc_44228_n7548_1_bF_buf4), .B(u2_remHi_109_), .Y(u2__abc_44228_n9446_1) );
  AND2X2 AND2X2_3668 ( .A(u2__abc_44228_n2983_bF_buf65), .B(u2__abc_44228_n3776), .Y(u2__abc_44228_n9449) );
  AND2X2 AND2X2_3669 ( .A(u2__abc_44228_n9450), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n9451_1) );
  AND2X2 AND2X2_367 ( .A(_abc_64468_n1635), .B(_abc_64468_n1642), .Y(_abc_64468_n1643) );
  AND2X2 AND2X2_3670 ( .A(u2__abc_44228_n9448), .B(u2__abc_44228_n9451_1), .Y(u2__abc_44228_n9452) );
  AND2X2 AND2X2_3671 ( .A(u2__abc_44228_n9453), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_remHi_111__FF_INPUT) );
  AND2X2 AND2X2_3672 ( .A(u2__abc_44228_n3062_bF_buf73), .B(u2_remHi_112_), .Y(u2__abc_44228_n9455) );
  AND2X2 AND2X2_3673 ( .A(u2__abc_44228_n7548_1_bF_buf3), .B(u2_remHi_110_), .Y(u2__abc_44228_n9456_1) );
  AND2X2 AND2X2_3674 ( .A(u2__abc_44228_n9182_1), .B(u2__abc_44228_n3902), .Y(u2__abc_44228_n9457_1) );
  AND2X2 AND2X2_3675 ( .A(u2__abc_44228_n9458), .B(u2__abc_44228_n3772), .Y(u2__abc_44228_n9459) );
  AND2X2 AND2X2_3676 ( .A(u2__abc_44228_n9460), .B(u2__abc_44228_n9461), .Y(u2__abc_44228_n9462_1) );
  AND2X2 AND2X2_3677 ( .A(u2__abc_44228_n7547_bF_buf2), .B(u2__abc_44228_n9462_1), .Y(u2__abc_44228_n9463) );
  AND2X2 AND2X2_3678 ( .A(u2__abc_44228_n2983_bF_buf63), .B(u2__abc_44228_n3762), .Y(u2__abc_44228_n9466) );
  AND2X2 AND2X2_3679 ( .A(u2__abc_44228_n9467_1), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n9468_1) );
  AND2X2 AND2X2_368 ( .A(_abc_64468_n1631), .B(_abc_64468_n1641), .Y(_abc_64468_n1644) );
  AND2X2 AND2X2_3680 ( .A(u2__abc_44228_n9465), .B(u2__abc_44228_n9468_1), .Y(u2__abc_44228_n9469) );
  AND2X2 AND2X2_3681 ( .A(u2__abc_44228_n9470), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_remHi_112__FF_INPUT) );
  AND2X2 AND2X2_3682 ( .A(u2__abc_44228_n3062_bF_buf72), .B(u2_remHi_113_), .Y(u2__abc_44228_n9472) );
  AND2X2 AND2X2_3683 ( .A(u2__abc_44228_n7548_1_bF_buf2), .B(u2_remHi_111_), .Y(u2__abc_44228_n9473_1) );
  AND2X2 AND2X2_3684 ( .A(u2__abc_44228_n9460), .B(u2__abc_44228_n4278), .Y(u2__abc_44228_n9475) );
  AND2X2 AND2X2_3685 ( .A(u2__abc_44228_n9476), .B(u2__abc_44228_n9474), .Y(u2__abc_44228_n9477) );
  AND2X2 AND2X2_3686 ( .A(u2__abc_44228_n9475), .B(u2__abc_44228_n3779_1), .Y(u2__abc_44228_n9478_1) );
  AND2X2 AND2X2_3687 ( .A(u2__abc_44228_n7547_bF_buf1), .B(u2__abc_44228_n9479_1), .Y(u2__abc_44228_n9480) );
  AND2X2 AND2X2_3688 ( .A(u2__abc_44228_n2983_bF_buf61), .B(u2__abc_44228_n3756), .Y(u2__abc_44228_n9483) );
  AND2X2 AND2X2_3689 ( .A(u2__abc_44228_n9484_1), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n9485) );
  AND2X2 AND2X2_369 ( .A(_abc_64468_n1645), .B(_abc_64468_n753_bF_buf9), .Y(_abc_64468_n1646) );
  AND2X2 AND2X2_3690 ( .A(u2__abc_44228_n9482), .B(u2__abc_44228_n9485), .Y(u2__abc_44228_n9486) );
  AND2X2 AND2X2_3691 ( .A(u2__abc_44228_n9487), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_remHi_113__FF_INPUT) );
  AND2X2 AND2X2_3692 ( .A(u2__abc_44228_n3062_bF_buf71), .B(u2_remHi_114_), .Y(u2__abc_44228_n9489_1) );
  AND2X2 AND2X2_3693 ( .A(u2__abc_44228_n9460), .B(u2__abc_44228_n4279), .Y(u2__abc_44228_n9490_1) );
  AND2X2 AND2X2_3694 ( .A(u2__abc_44228_n9492), .B(u2__abc_44228_n3765), .Y(u2__abc_44228_n9494) );
  AND2X2 AND2X2_3695 ( .A(u2__abc_44228_n9495_1), .B(u2__abc_44228_n9493), .Y(u2__abc_44228_n9496) );
  AND2X2 AND2X2_3696 ( .A(u2__abc_44228_n9497), .B(u2__abc_44228_n9498), .Y(u2__abc_44228_n9499) );
  AND2X2 AND2X2_3697 ( .A(u2__abc_44228_n2983_bF_buf59), .B(u2__abc_44228_n3747), .Y(u2__abc_44228_n9501_1) );
  AND2X2 AND2X2_3698 ( .A(u2__abc_44228_n9502), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n9503) );
  AND2X2 AND2X2_3699 ( .A(u2__abc_44228_n9500_1), .B(u2__abc_44228_n9503), .Y(u2__abc_44228_n9504) );
  AND2X2 AND2X2_37 ( .A(_abc_64468_n753_bF_buf5), .B(sqrto_36_), .Y(_auto_iopadmap_cc_313_execute_65414_72_) );
  AND2X2 AND2X2_370 ( .A(aNan_bF_buf8), .B(\a[122] ), .Y(_abc_64468_n1647) );
  AND2X2 AND2X2_3700 ( .A(u2__abc_44228_n9505), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_remHi_114__FF_INPUT) );
  AND2X2 AND2X2_3701 ( .A(u2__abc_44228_n3062_bF_buf70), .B(u2_remHi_115_), .Y(u2__abc_44228_n9507) );
  AND2X2 AND2X2_3702 ( .A(u2__abc_44228_n9512_1), .B(u2__abc_44228_n7547_bF_buf57), .Y(u2__abc_44228_n9513) );
  AND2X2 AND2X2_3703 ( .A(u2__abc_44228_n9513), .B(u2__abc_44228_n9511_1), .Y(u2__abc_44228_n9514) );
  AND2X2 AND2X2_3704 ( .A(u2__abc_44228_n7548_1_bF_buf0), .B(u2_remHi_113_), .Y(u2__abc_44228_n9515) );
  AND2X2 AND2X2_3705 ( .A(u2__abc_44228_n2983_bF_buf57), .B(u2__abc_44228_n3741), .Y(u2__abc_44228_n9518) );
  AND2X2 AND2X2_3706 ( .A(u2__abc_44228_n9519), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n9520) );
  AND2X2 AND2X2_3707 ( .A(u2__abc_44228_n9517_1), .B(u2__abc_44228_n9520), .Y(u2__abc_44228_n9521) );
  AND2X2 AND2X2_3708 ( .A(u2__abc_44228_n9522_1), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_remHi_115__FF_INPUT) );
  AND2X2 AND2X2_3709 ( .A(u2__abc_44228_n3062_bF_buf69), .B(u2_remHi_116_), .Y(u2__abc_44228_n9524) );
  AND2X2 AND2X2_371 ( .A(aNan_bF_buf7), .B(\a[123] ), .Y(_abc_64468_n1649) );
  AND2X2 AND2X2_3710 ( .A(u2__abc_44228_n9458), .B(u2__abc_44228_n3781), .Y(u2__abc_44228_n9525) );
  AND2X2 AND2X2_3711 ( .A(u2__abc_44228_n9526), .B(u2__abc_44228_n3750_1), .Y(u2__abc_44228_n9527) );
  AND2X2 AND2X2_3712 ( .A(u2__abc_44228_n9528_1), .B(u2__abc_44228_n9529), .Y(u2__abc_44228_n9530) );
  AND2X2 AND2X2_3713 ( .A(u2__abc_44228_n9531), .B(u2__abc_44228_n9532), .Y(u2__abc_44228_n9533_1) );
  AND2X2 AND2X2_3714 ( .A(u2__abc_44228_n2983_bF_buf55), .B(u2__abc_44228_n3733), .Y(u2__abc_44228_n9535) );
  AND2X2 AND2X2_3715 ( .A(u2__abc_44228_n9536), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n9537) );
  AND2X2 AND2X2_3716 ( .A(u2__abc_44228_n9534_1), .B(u2__abc_44228_n9537), .Y(u2__abc_44228_n9538) );
  AND2X2 AND2X2_3717 ( .A(u2__abc_44228_n9539_1), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_remHi_116__FF_INPUT) );
  AND2X2 AND2X2_3718 ( .A(u2__abc_44228_n3062_bF_buf68), .B(u2_remHi_117_), .Y(u2__abc_44228_n9541) );
  AND2X2 AND2X2_3719 ( .A(u2__abc_44228_n9528_1), .B(u2__abc_44228_n4287), .Y(u2__abc_44228_n9542) );
  AND2X2 AND2X2_372 ( .A(_abc_64468_n1637), .B(\a[123] ), .Y(_abc_64468_n1652) );
  AND2X2 AND2X2_3720 ( .A(u2__abc_44228_n7547_bF_buf55), .B(u2__abc_44228_n9546), .Y(u2__abc_44228_n9547) );
  AND2X2 AND2X2_3721 ( .A(u2__abc_44228_n9547), .B(u2__abc_44228_n9544_1), .Y(u2__abc_44228_n9548) );
  AND2X2 AND2X2_3722 ( .A(u2__abc_44228_n7548_1_bF_buf56), .B(u2_remHi_115_), .Y(u2__abc_44228_n9549) );
  AND2X2 AND2X2_3723 ( .A(u2__abc_44228_n2983_bF_buf53), .B(u2__abc_44228_n3727), .Y(u2__abc_44228_n9552) );
  AND2X2 AND2X2_3724 ( .A(u2__abc_44228_n9553), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n9554) );
  AND2X2 AND2X2_3725 ( .A(u2__abc_44228_n9551), .B(u2__abc_44228_n9554), .Y(u2__abc_44228_n9555_1) );
  AND2X2 AND2X2_3726 ( .A(u2__abc_44228_n9556_1), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_remHi_117__FF_INPUT) );
  AND2X2 AND2X2_3727 ( .A(u2__abc_44228_n3062_bF_buf67), .B(u2_remHi_118_), .Y(u2__abc_44228_n9558) );
  AND2X2 AND2X2_3728 ( .A(u2__abc_44228_n9526), .B(u2__abc_44228_n3751), .Y(u2__abc_44228_n9559) );
  AND2X2 AND2X2_3729 ( .A(u2__abc_44228_n9560), .B(u2__abc_44228_n3736), .Y(u2__abc_44228_n9562) );
  AND2X2 AND2X2_373 ( .A(_abc_64468_n1652), .B(_abc_64468_n1651), .Y(_abc_64468_n1654) );
  AND2X2 AND2X2_3730 ( .A(u2__abc_44228_n9563), .B(u2__abc_44228_n9561_1), .Y(u2__abc_44228_n9564) );
  AND2X2 AND2X2_3731 ( .A(u2__abc_44228_n9565), .B(u2__abc_44228_n9566_1), .Y(u2__abc_44228_n9567_1) );
  AND2X2 AND2X2_3732 ( .A(u2__abc_44228_n2983_bF_buf51), .B(u2__abc_44228_n3703), .Y(u2__abc_44228_n9569) );
  AND2X2 AND2X2_3733 ( .A(u2__abc_44228_n9570), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n9571) );
  AND2X2 AND2X2_3734 ( .A(u2__abc_44228_n9568), .B(u2__abc_44228_n9571), .Y(u2__abc_44228_n9572_1) );
  AND2X2 AND2X2_3735 ( .A(u2__abc_44228_n9573), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_remHi_118__FF_INPUT) );
  AND2X2 AND2X2_3736 ( .A(u2__abc_44228_n3062_bF_buf66), .B(u2_remHi_119_), .Y(u2__abc_44228_n9575) );
  AND2X2 AND2X2_3737 ( .A(u2__abc_44228_n9580), .B(u2__abc_44228_n7547_bF_buf53), .Y(u2__abc_44228_n9581) );
  AND2X2 AND2X2_3738 ( .A(u2__abc_44228_n9581), .B(u2__abc_44228_n9579), .Y(u2__abc_44228_n9582) );
  AND2X2 AND2X2_3739 ( .A(u2__abc_44228_n7548_1_bF_buf54), .B(u2_remHi_117_), .Y(u2__abc_44228_n9583_1) );
  AND2X2 AND2X2_374 ( .A(_abc_64468_n1655), .B(_abc_64468_n1653), .Y(_abc_64468_n1656) );
  AND2X2 AND2X2_3740 ( .A(u2__abc_44228_n2983_bF_buf49), .B(u2__abc_44228_n3697), .Y(u2__abc_44228_n9586) );
  AND2X2 AND2X2_3741 ( .A(u2__abc_44228_n9587), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n9588_1) );
  AND2X2 AND2X2_3742 ( .A(u2__abc_44228_n9585), .B(u2__abc_44228_n9588_1), .Y(u2__abc_44228_n9589_1) );
  AND2X2 AND2X2_3743 ( .A(u2__abc_44228_n9590), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_remHi_119__FF_INPUT) );
  AND2X2 AND2X2_3744 ( .A(u2__abc_44228_n3062_bF_buf65), .B(u2_remHi_120_), .Y(u2__abc_44228_n9592) );
  AND2X2 AND2X2_3745 ( .A(u2__abc_44228_n9458), .B(u2__abc_44228_n3782), .Y(u2__abc_44228_n9593) );
  AND2X2 AND2X2_3746 ( .A(u2__abc_44228_n9594_1), .B(u2__abc_44228_n3706), .Y(u2__abc_44228_n9596) );
  AND2X2 AND2X2_3747 ( .A(u2__abc_44228_n9597), .B(u2__abc_44228_n9595), .Y(u2__abc_44228_n9598) );
  AND2X2 AND2X2_3748 ( .A(u2__abc_44228_n9599_1), .B(u2__abc_44228_n9600_1), .Y(u2__abc_44228_n9601) );
  AND2X2 AND2X2_3749 ( .A(u2__abc_44228_n2983_bF_buf47), .B(u2__abc_44228_n3717), .Y(u2__abc_44228_n9603) );
  AND2X2 AND2X2_375 ( .A(_abc_64468_n1650), .B(_abc_64468_n1657), .Y(_abc_64468_n1658) );
  AND2X2 AND2X2_3750 ( .A(u2__abc_44228_n9604), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n9605_1) );
  AND2X2 AND2X2_3751 ( .A(u2__abc_44228_n9602), .B(u2__abc_44228_n9605_1), .Y(u2__abc_44228_n9606) );
  AND2X2 AND2X2_3752 ( .A(u2__abc_44228_n9607), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_remHi_120__FF_INPUT) );
  AND2X2 AND2X2_3753 ( .A(u2__abc_44228_n3062_bF_buf64), .B(u2_remHi_121_), .Y(u2__abc_44228_n9609) );
  AND2X2 AND2X2_3754 ( .A(u2__abc_44228_n9597), .B(u2__abc_44228_n4260), .Y(u2__abc_44228_n9611_1) );
  AND2X2 AND2X2_3755 ( .A(u2__abc_44228_n9614), .B(u2__abc_44228_n9612), .Y(u2__abc_44228_n9615) );
  AND2X2 AND2X2_3756 ( .A(u2__abc_44228_n9615), .B(u2__abc_44228_n7547_bF_buf51), .Y(u2__abc_44228_n9616_1) );
  AND2X2 AND2X2_3757 ( .A(u2__abc_44228_n7548_1_bF_buf52), .B(u2_remHi_119_), .Y(u2__abc_44228_n9617) );
  AND2X2 AND2X2_3758 ( .A(u2__abc_44228_n2983_bF_buf45), .B(u2__abc_44228_n3711), .Y(u2__abc_44228_n9620) );
  AND2X2 AND2X2_3759 ( .A(u2__abc_44228_n9621_1), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n9622_1) );
  AND2X2 AND2X2_376 ( .A(_abc_64468_n1644), .B(_abc_64468_n1656), .Y(_abc_64468_n1659) );
  AND2X2 AND2X2_3760 ( .A(u2__abc_44228_n9619), .B(u2__abc_44228_n9622_1), .Y(u2__abc_44228_n9623) );
  AND2X2 AND2X2_3761 ( .A(u2__abc_44228_n9624), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_remHi_121__FF_INPUT) );
  AND2X2 AND2X2_3762 ( .A(u2__abc_44228_n3062_bF_buf63), .B(u2_remHi_122_), .Y(u2__abc_44228_n9626) );
  AND2X2 AND2X2_3763 ( .A(u2__abc_44228_n9594_1), .B(u2__abc_44228_n3707), .Y(u2__abc_44228_n9627_1) );
  AND2X2 AND2X2_3764 ( .A(u2__abc_44228_n9628), .B(u2__abc_44228_n3720), .Y(u2__abc_44228_n9630) );
  AND2X2 AND2X2_3765 ( .A(u2__abc_44228_n9631), .B(u2__abc_44228_n9629), .Y(u2__abc_44228_n9632_1) );
  AND2X2 AND2X2_3766 ( .A(u2__abc_44228_n9633_1), .B(u2__abc_44228_n9634), .Y(u2__abc_44228_n9635) );
  AND2X2 AND2X2_3767 ( .A(u2__abc_44228_n2983_bF_buf43), .B(u2__abc_44228_n3681), .Y(u2__abc_44228_n9637) );
  AND2X2 AND2X2_3768 ( .A(u2__abc_44228_n9638_1), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n9639) );
  AND2X2 AND2X2_3769 ( .A(u2__abc_44228_n9636), .B(u2__abc_44228_n9639), .Y(u2__abc_44228_n9640) );
  AND2X2 AND2X2_377 ( .A(_abc_64468_n1660), .B(_abc_64468_n753_bF_buf8), .Y(_abc_64468_n1661) );
  AND2X2 AND2X2_3770 ( .A(u2__abc_44228_n9641), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_remHi_122__FF_INPUT) );
  AND2X2 AND2X2_3771 ( .A(u2__abc_44228_n3062_bF_buf62), .B(u2_remHi_123_), .Y(u2__abc_44228_n9643_1) );
  AND2X2 AND2X2_3772 ( .A(u2__abc_44228_n9648), .B(u2__abc_44228_n7547_bF_buf49), .Y(u2__abc_44228_n9649_1) );
  AND2X2 AND2X2_3773 ( .A(u2__abc_44228_n9649_1), .B(u2__abc_44228_n9647), .Y(u2__abc_44228_n9650) );
  AND2X2 AND2X2_3774 ( .A(u2__abc_44228_n7548_1_bF_buf50), .B(u2_remHi_121_), .Y(u2__abc_44228_n9651) );
  AND2X2 AND2X2_3775 ( .A(u2__abc_44228_n2983_bF_buf41), .B(u2__abc_44228_n3688), .Y(u2__abc_44228_n9654_1) );
  AND2X2 AND2X2_3776 ( .A(u2__abc_44228_n9655_1), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n9656) );
  AND2X2 AND2X2_3777 ( .A(u2__abc_44228_n9653), .B(u2__abc_44228_n9656), .Y(u2__abc_44228_n9657) );
  AND2X2 AND2X2_3778 ( .A(u2__abc_44228_n9658), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_remHi_123__FF_INPUT) );
  AND2X2 AND2X2_3779 ( .A(u2__abc_44228_n3062_bF_buf61), .B(u2_remHi_124_), .Y(u2__abc_44228_n9660_1) );
  AND2X2 AND2X2_378 ( .A(_abc_64468_n1652), .B(\a[124] ), .Y(_abc_64468_n1665) );
  AND2X2 AND2X2_3780 ( .A(u2__abc_44228_n9594_1), .B(u2__abc_44228_n3722), .Y(u2__abc_44228_n9661) );
  AND2X2 AND2X2_3781 ( .A(u2__abc_44228_n9662), .B(u2__abc_44228_n3684), .Y(u2__abc_44228_n9663) );
  AND2X2 AND2X2_3782 ( .A(u2__abc_44228_n9664), .B(u2__abc_44228_n9665_1), .Y(u2__abc_44228_n9666_1) );
  AND2X2 AND2X2_3783 ( .A(u2__abc_44228_n9667), .B(u2__abc_44228_n9668), .Y(u2__abc_44228_n9669) );
  AND2X2 AND2X2_3784 ( .A(u2__abc_44228_n2983_bF_buf39), .B(u2__abc_44228_n3674), .Y(u2__abc_44228_n9671_1) );
  AND2X2 AND2X2_3785 ( .A(u2__abc_44228_n9672), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n9673) );
  AND2X2 AND2X2_3786 ( .A(u2__abc_44228_n9670), .B(u2__abc_44228_n9673), .Y(u2__abc_44228_n9674) );
  AND2X2 AND2X2_3787 ( .A(u2__abc_44228_n9675), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_remHi_124__FF_INPUT) );
  AND2X2 AND2X2_3788 ( .A(u2__abc_44228_n3062_bF_buf60), .B(u2_remHi_125_), .Y(u2__abc_44228_n9677_1) );
  AND2X2 AND2X2_3789 ( .A(u2__abc_44228_n9664), .B(u2__abc_44228_n4269), .Y(u2__abc_44228_n9678) );
  AND2X2 AND2X2_379 ( .A(_abc_64468_n1665), .B(_abc_64468_n1664), .Y(_abc_64468_n1667) );
  AND2X2 AND2X2_3790 ( .A(u2__abc_44228_n9678), .B(u2__abc_44228_n3691), .Y(u2__abc_44228_n9679) );
  AND2X2 AND2X2_3791 ( .A(u2__abc_44228_n9681), .B(u2__abc_44228_n9680), .Y(u2__abc_44228_n9682_1) );
  AND2X2 AND2X2_3792 ( .A(u2__abc_44228_n9683), .B(u2__abc_44228_n7547_bF_buf47), .Y(u2__abc_44228_n9684) );
  AND2X2 AND2X2_3793 ( .A(u2__abc_44228_n7548_1_bF_buf48), .B(u2_remHi_123_), .Y(u2__abc_44228_n9685) );
  AND2X2 AND2X2_3794 ( .A(u2__abc_44228_n2983_bF_buf37), .B(u2__abc_44228_n3668), .Y(u2__abc_44228_n9688_1) );
  AND2X2 AND2X2_3795 ( .A(u2__abc_44228_n9689), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n9690) );
  AND2X2 AND2X2_3796 ( .A(u2__abc_44228_n9687_1), .B(u2__abc_44228_n9690), .Y(u2__abc_44228_n9691) );
  AND2X2 AND2X2_3797 ( .A(u2__abc_44228_n9692), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_remHi_125__FF_INPUT) );
  AND2X2 AND2X2_3798 ( .A(u2__abc_44228_n3062_bF_buf59), .B(u2_remHi_126_), .Y(u2__abc_44228_n9694) );
  AND2X2 AND2X2_3799 ( .A(u2__abc_44228_n9664), .B(u2__abc_44228_n4270), .Y(u2__abc_44228_n9695) );
  AND2X2 AND2X2_38 ( .A(_abc_64468_n753_bF_buf4), .B(sqrto_37_), .Y(_auto_iopadmap_cc_313_execute_65414_73_) );
  AND2X2 AND2X2_380 ( .A(_abc_64468_n1668), .B(_abc_64468_n1666), .Y(_abc_64468_n1669) );
  AND2X2 AND2X2_3800 ( .A(u2__abc_44228_n9697), .B(u2__abc_44228_n3677), .Y(u2__abc_44228_n9699_1) );
  AND2X2 AND2X2_3801 ( .A(u2__abc_44228_n9700), .B(u2__abc_44228_n9698_1), .Y(u2__abc_44228_n9701) );
  AND2X2 AND2X2_3802 ( .A(u2__abc_44228_n9701), .B(u2__abc_44228_n7547_bF_buf46), .Y(u2__abc_44228_n9702) );
  AND2X2 AND2X2_3803 ( .A(u2__abc_44228_n7548_1_bF_buf47), .B(u2_remHi_124_), .Y(u2__abc_44228_n9703) );
  AND2X2 AND2X2_3804 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n5246), .Y(u2__abc_44228_n9706) );
  AND2X2 AND2X2_3805 ( .A(u2__abc_44228_n9707), .B(u2__abc_44228_n2972_bF_buf87), .Y(u2__abc_44228_n9708) );
  AND2X2 AND2X2_3806 ( .A(u2__abc_44228_n9705), .B(u2__abc_44228_n9708), .Y(u2__abc_44228_n9709_1) );
  AND2X2 AND2X2_3807 ( .A(u2__abc_44228_n9710_1), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_remHi_126__FF_INPUT) );
  AND2X2 AND2X2_3808 ( .A(u2__abc_44228_n3062_bF_buf58), .B(u2_remHi_127_), .Y(u2__abc_44228_n9712) );
  AND2X2 AND2X2_3809 ( .A(u2__abc_44228_n9717), .B(u2__abc_44228_n7547_bF_buf45), .Y(u2__abc_44228_n9718) );
  AND2X2 AND2X2_381 ( .A(_abc_64468_n1663), .B(_abc_64468_n1670), .Y(_abc_64468_n1671) );
  AND2X2 AND2X2_3810 ( .A(u2__abc_44228_n9718), .B(u2__abc_44228_n9716), .Y(u2__abc_44228_n9719) );
  AND2X2 AND2X2_3811 ( .A(u2__abc_44228_n7548_1_bF_buf46), .B(u2_remHi_125_), .Y(u2__abc_44228_n9720_1) );
  AND2X2 AND2X2_3812 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n5240), .Y(u2__abc_44228_n9723) );
  AND2X2 AND2X2_3813 ( .A(u2__abc_44228_n9724), .B(u2__abc_44228_n2972_bF_buf86), .Y(u2__abc_44228_n9725) );
  AND2X2 AND2X2_3814 ( .A(u2__abc_44228_n9722), .B(u2__abc_44228_n9725), .Y(u2__abc_44228_n9726_1) );
  AND2X2 AND2X2_3815 ( .A(u2__abc_44228_n9727), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_remHi_127__FF_INPUT) );
  AND2X2 AND2X2_3816 ( .A(u2__abc_44228_n3062_bF_buf57), .B(u2_remHi_128_), .Y(u2__abc_44228_n9729) );
  AND2X2 AND2X2_3817 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5249), .Y(u2__abc_44228_n9730) );
  AND2X2 AND2X2_3818 ( .A(u2__abc_44228_n9731_1), .B(u2__abc_44228_n9732_1), .Y(u2__abc_44228_n9733) );
  AND2X2 AND2X2_3819 ( .A(u2__abc_44228_n7547_bF_buf44), .B(u2__abc_44228_n9733), .Y(u2__abc_44228_n9734) );
  AND2X2 AND2X2_382 ( .A(_abc_64468_n1659), .B(_abc_64468_n1669), .Y(_abc_64468_n1672) );
  AND2X2 AND2X2_3820 ( .A(u2__abc_44228_n7548_1_bF_buf45), .B(u2_remHi_126_), .Y(u2__abc_44228_n9735) );
  AND2X2 AND2X2_3821 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n5231), .Y(u2__abc_44228_n9738) );
  AND2X2 AND2X2_3822 ( .A(u2__abc_44228_n9739), .B(u2__abc_44228_n2972_bF_buf85), .Y(u2__abc_44228_n9740) );
  AND2X2 AND2X2_3823 ( .A(u2__abc_44228_n9737_1), .B(u2__abc_44228_n9740), .Y(u2__abc_44228_n9741) );
  AND2X2 AND2X2_3824 ( .A(u2__abc_44228_n9742_1), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_remHi_128__FF_INPUT) );
  AND2X2 AND2X2_3825 ( .A(u2__abc_44228_n3062_bF_buf56), .B(u2_remHi_129_), .Y(u2__abc_44228_n9744) );
  AND2X2 AND2X2_3826 ( .A(u2__abc_44228_n9746), .B(u2__abc_44228_n9745), .Y(u2__abc_44228_n9747) );
  AND2X2 AND2X2_3827 ( .A(u2__abc_44228_n9748_1), .B(u2__abc_44228_n5243), .Y(u2__abc_44228_n9749) );
  AND2X2 AND2X2_3828 ( .A(u2__abc_44228_n7547_bF_buf43), .B(u2__abc_44228_n9750), .Y(u2__abc_44228_n9751) );
  AND2X2 AND2X2_3829 ( .A(u2__abc_44228_n7548_1_bF_buf44), .B(u2_remHi_127_), .Y(u2__abc_44228_n9752) );
  AND2X2 AND2X2_383 ( .A(_abc_64468_n1673), .B(_abc_64468_n753_bF_buf7), .Y(_abc_64468_n1674) );
  AND2X2 AND2X2_3830 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n5226), .Y(u2__abc_44228_n9755) );
  AND2X2 AND2X2_3831 ( .A(u2__abc_44228_n9756), .B(u2__abc_44228_n2972_bF_buf84), .Y(u2__abc_44228_n9757) );
  AND2X2 AND2X2_3832 ( .A(u2__abc_44228_n9754_1), .B(u2__abc_44228_n9757), .Y(u2__abc_44228_n9758) );
  AND2X2 AND2X2_3833 ( .A(u2__abc_44228_n9759_1), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_remHi_129__FF_INPUT) );
  AND2X2 AND2X2_3834 ( .A(u2__abc_44228_n3062_bF_buf55), .B(u2_remHi_130_), .Y(u2__abc_44228_n9761) );
  AND2X2 AND2X2_3835 ( .A(u2__abc_44228_n7548_1_bF_buf43), .B(u2_remHi_128_), .Y(u2__abc_44228_n9762) );
  AND2X2 AND2X2_3836 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5250_1), .Y(u2__abc_44228_n9763) );
  AND2X2 AND2X2_3837 ( .A(u2__abc_44228_n9764_1), .B(u2__abc_44228_n5235), .Y(u2__abc_44228_n9766) );
  AND2X2 AND2X2_3838 ( .A(u2__abc_44228_n9767), .B(u2__abc_44228_n9765_1), .Y(u2__abc_44228_n9768) );
  AND2X2 AND2X2_3839 ( .A(u2__abc_44228_n7547_bF_buf42), .B(u2__abc_44228_n9768), .Y(u2__abc_44228_n9769) );
  AND2X2 AND2X2_384 ( .A(aNan_bF_buf6), .B(\a[124] ), .Y(_abc_64468_n1675) );
  AND2X2 AND2X2_3840 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n5220), .Y(u2__abc_44228_n9772) );
  AND2X2 AND2X2_3841 ( .A(u2__abc_44228_n9773), .B(u2__abc_44228_n2972_bF_buf83), .Y(u2__abc_44228_n9774) );
  AND2X2 AND2X2_3842 ( .A(u2__abc_44228_n9771), .B(u2__abc_44228_n9774), .Y(u2__abc_44228_n9775_1) );
  AND2X2 AND2X2_3843 ( .A(u2__abc_44228_n9776_1), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_remHi_130__FF_INPUT) );
  AND2X2 AND2X2_3844 ( .A(u2__abc_44228_n3062_bF_buf54), .B(u2_remHi_131_), .Y(u2__abc_44228_n9778) );
  AND2X2 AND2X2_3845 ( .A(u2__abc_44228_n7548_1_bF_buf42), .B(u2_remHi_129_), .Y(u2__abc_44228_n9779) );
  AND2X2 AND2X2_3846 ( .A(u2__abc_44228_n9767), .B(u2__abc_44228_n5232), .Y(u2__abc_44228_n9781_1) );
  AND2X2 AND2X2_3847 ( .A(u2__abc_44228_n9782), .B(u2__abc_44228_n9780), .Y(u2__abc_44228_n9783) );
  AND2X2 AND2X2_3848 ( .A(u2__abc_44228_n9781_1), .B(u2__abc_44228_n5230_1), .Y(u2__abc_44228_n9784) );
  AND2X2 AND2X2_3849 ( .A(u2__abc_44228_n7547_bF_buf41), .B(u2__abc_44228_n9785), .Y(u2__abc_44228_n9786_1) );
  AND2X2 AND2X2_385 ( .A(_abc_64468_n1665), .B(\a[125] ), .Y(_abc_64468_n1679) );
  AND2X2 AND2X2_3850 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n5214), .Y(u2__abc_44228_n9789) );
  AND2X2 AND2X2_3851 ( .A(u2__abc_44228_n9790), .B(u2__abc_44228_n2972_bF_buf82), .Y(u2__abc_44228_n9791) );
  AND2X2 AND2X2_3852 ( .A(u2__abc_44228_n9788), .B(u2__abc_44228_n9791), .Y(u2__abc_44228_n9792_1) );
  AND2X2 AND2X2_3853 ( .A(u2__abc_44228_n9793), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_remHi_131__FF_INPUT) );
  AND2X2 AND2X2_3854 ( .A(u2__abc_44228_n3062_bF_buf53), .B(u2_remHi_132_), .Y(u2__abc_44228_n9795) );
  AND2X2 AND2X2_3855 ( .A(u2__abc_44228_n7548_1_bF_buf41), .B(u2_remHi_130_), .Y(u2__abc_44228_n9796) );
  AND2X2 AND2X2_3856 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5251), .Y(u2__abc_44228_n9797_1) );
  AND2X2 AND2X2_3857 ( .A(u2__abc_44228_n9798_1), .B(u2__abc_44228_n5223), .Y(u2__abc_44228_n9799) );
  AND2X2 AND2X2_3858 ( .A(u2__abc_44228_n9800), .B(u2__abc_44228_n9801), .Y(u2__abc_44228_n9802) );
  AND2X2 AND2X2_3859 ( .A(u2__abc_44228_n7547_bF_buf40), .B(u2__abc_44228_n9802), .Y(u2__abc_44228_n9803_1) );
  AND2X2 AND2X2_386 ( .A(_abc_64468_n1679), .B(_abc_64468_n1678), .Y(_abc_64468_n1681) );
  AND2X2 AND2X2_3860 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n5206), .Y(u2__abc_44228_n9806) );
  AND2X2 AND2X2_3861 ( .A(u2__abc_44228_n9807), .B(u2__abc_44228_n2972_bF_buf81), .Y(u2__abc_44228_n9808_1) );
  AND2X2 AND2X2_3862 ( .A(u2__abc_44228_n9805), .B(u2__abc_44228_n9808_1), .Y(u2__abc_44228_n9809_1) );
  AND2X2 AND2X2_3863 ( .A(u2__abc_44228_n9810), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_remHi_132__FF_INPUT) );
  AND2X2 AND2X2_3864 ( .A(u2__abc_44228_n3062_bF_buf52), .B(u2_remHi_133_), .Y(u2__abc_44228_n9812) );
  AND2X2 AND2X2_3865 ( .A(u2__abc_44228_n7548_1_bF_buf40), .B(u2_remHi_131_), .Y(u2__abc_44228_n9813) );
  AND2X2 AND2X2_3866 ( .A(u2__abc_44228_n9815), .B(u2__abc_44228_n9814_1), .Y(u2__abc_44228_n9816) );
  AND2X2 AND2X2_3867 ( .A(u2__abc_44228_n9817), .B(u2__abc_44228_n5217), .Y(u2__abc_44228_n9818) );
  AND2X2 AND2X2_3868 ( .A(u2__abc_44228_n7547_bF_buf39), .B(u2__abc_44228_n9819_1), .Y(u2__abc_44228_n9820_1) );
  AND2X2 AND2X2_3869 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n5200), .Y(u2__abc_44228_n9823) );
  AND2X2 AND2X2_387 ( .A(_abc_64468_n1682), .B(_abc_64468_n1680), .Y(_abc_64468_n1683) );
  AND2X2 AND2X2_3870 ( .A(u2__abc_44228_n9824), .B(u2__abc_44228_n2972_bF_buf80), .Y(u2__abc_44228_n9825_1) );
  AND2X2 AND2X2_3871 ( .A(u2__abc_44228_n9822), .B(u2__abc_44228_n9825_1), .Y(u2__abc_44228_n9826) );
  AND2X2 AND2X2_3872 ( .A(u2__abc_44228_n9827), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_remHi_133__FF_INPUT) );
  AND2X2 AND2X2_3873 ( .A(u2__abc_44228_n3062_bF_buf51), .B(u2_remHi_134_), .Y(u2__abc_44228_n9829) );
  AND2X2 AND2X2_3874 ( .A(u2__abc_44228_n9798_1), .B(u2__abc_44228_n5224), .Y(u2__abc_44228_n9830_1) );
  AND2X2 AND2X2_3875 ( .A(u2__abc_44228_n9831_1), .B(u2__abc_44228_n5209), .Y(u2__abc_44228_n9833) );
  AND2X2 AND2X2_3876 ( .A(u2__abc_44228_n9834), .B(u2__abc_44228_n9832), .Y(u2__abc_44228_n9835) );
  AND2X2 AND2X2_3877 ( .A(u2__abc_44228_n9836_1), .B(u2__abc_44228_n9837), .Y(u2__abc_44228_n9838) );
  AND2X2 AND2X2_3878 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n5176), .Y(u2__abc_44228_n9840) );
  AND2X2 AND2X2_3879 ( .A(u2__abc_44228_n9841_1), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n9842_1) );
  AND2X2 AND2X2_388 ( .A(_abc_64468_n1672), .B(_abc_64468_n1683), .Y(_abc_64468_n1685) );
  AND2X2 AND2X2_3880 ( .A(u2__abc_44228_n9839), .B(u2__abc_44228_n9842_1), .Y(u2__abc_44228_n9843) );
  AND2X2 AND2X2_3881 ( .A(u2__abc_44228_n9844), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_remHi_134__FF_INPUT) );
  AND2X2 AND2X2_3882 ( .A(u2__abc_44228_n3062_bF_buf50), .B(u2_remHi_135_), .Y(u2__abc_44228_n9846) );
  AND2X2 AND2X2_3883 ( .A(u2__abc_44228_n9851), .B(u2__abc_44228_n9848), .Y(u2__abc_44228_n9852_1) );
  AND2X2 AND2X2_3884 ( .A(u2__abc_44228_n9852_1), .B(u2__abc_44228_n7547_bF_buf37), .Y(u2__abc_44228_n9853_1) );
  AND2X2 AND2X2_3885 ( .A(u2__abc_44228_n7548_1_bF_buf38), .B(u2_remHi_133_), .Y(u2__abc_44228_n9854) );
  AND2X2 AND2X2_3886 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n5170), .Y(u2__abc_44228_n9857) );
  AND2X2 AND2X2_3887 ( .A(u2__abc_44228_n9858_1), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n9859) );
  AND2X2 AND2X2_3888 ( .A(u2__abc_44228_n9856), .B(u2__abc_44228_n9859), .Y(u2__abc_44228_n9860) );
  AND2X2 AND2X2_3889 ( .A(u2__abc_44228_n9861), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_remHi_135__FF_INPUT) );
  AND2X2 AND2X2_389 ( .A(_abc_64468_n1686), .B(_abc_64468_n1684), .Y(_abc_64468_n1687) );
  AND2X2 AND2X2_3890 ( .A(u2__abc_44228_n3062_bF_buf49), .B(u2_remHi_136_), .Y(u2__abc_44228_n9863_1) );
  AND2X2 AND2X2_3891 ( .A(u2__abc_44228_n7548_1_bF_buf37), .B(u2_remHi_134_), .Y(u2__abc_44228_n9864_1) );
  AND2X2 AND2X2_3892 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5252), .Y(u2__abc_44228_n9865) );
  AND2X2 AND2X2_3893 ( .A(u2__abc_44228_n9866), .B(u2__abc_44228_n5179), .Y(u2__abc_44228_n9868) );
  AND2X2 AND2X2_3894 ( .A(u2__abc_44228_n9869_1), .B(u2__abc_44228_n9867), .Y(u2__abc_44228_n9870) );
  AND2X2 AND2X2_3895 ( .A(u2__abc_44228_n7547_bF_buf36), .B(u2__abc_44228_n9870), .Y(u2__abc_44228_n9871) );
  AND2X2 AND2X2_3896 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n5190), .Y(u2__abc_44228_n9874_1) );
  AND2X2 AND2X2_3897 ( .A(u2__abc_44228_n9875_1), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n9876) );
  AND2X2 AND2X2_3898 ( .A(u2__abc_44228_n9873), .B(u2__abc_44228_n9876), .Y(u2__abc_44228_n9877) );
  AND2X2 AND2X2_3899 ( .A(u2__abc_44228_n9878), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_remHi_136__FF_INPUT) );
  AND2X2 AND2X2_39 ( .A(_abc_64468_n753_bF_buf3), .B(sqrto_38_), .Y(_auto_iopadmap_cc_313_execute_65414_74_) );
  AND2X2 AND2X2_390 ( .A(_abc_64468_n1688), .B(_abc_64468_n1677), .Y(_auto_iopadmap_cc_313_execute_65414_239_) );
  AND2X2 AND2X2_3900 ( .A(u2__abc_44228_n3062_bF_buf48), .B(u2_remHi_137_), .Y(u2__abc_44228_n9880_1) );
  AND2X2 AND2X2_3901 ( .A(u2__abc_44228_n7548_1_bF_buf36), .B(u2_remHi_135_), .Y(u2__abc_44228_n9881) );
  AND2X2 AND2X2_3902 ( .A(u2__abc_44228_n9883), .B(u2__abc_44228_n9882), .Y(u2__abc_44228_n9884) );
  AND2X2 AND2X2_3903 ( .A(u2__abc_44228_n9885_1), .B(u2__abc_44228_n5173_1), .Y(u2__abc_44228_n9886_1) );
  AND2X2 AND2X2_3904 ( .A(u2__abc_44228_n7547_bF_buf35), .B(u2__abc_44228_n9887), .Y(u2__abc_44228_n9888) );
  AND2X2 AND2X2_3905 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n5184), .Y(u2__abc_44228_n9891_1) );
  AND2X2 AND2X2_3906 ( .A(u2__abc_44228_n9892), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n9893) );
  AND2X2 AND2X2_3907 ( .A(u2__abc_44228_n9890), .B(u2__abc_44228_n9893), .Y(u2__abc_44228_n9894) );
  AND2X2 AND2X2_3908 ( .A(u2__abc_44228_n9895), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_remHi_137__FF_INPUT) );
  AND2X2 AND2X2_3909 ( .A(u2__abc_44228_n3062_bF_buf47), .B(u2_remHi_138_), .Y(u2__abc_44228_n9897_1) );
  AND2X2 AND2X2_391 ( .A(_abc_64468_n1690), .B(\a[126] ), .Y(_abc_64468_n1691) );
  AND2X2 AND2X2_3910 ( .A(u2__abc_44228_n9866), .B(u2__abc_44228_n5180), .Y(u2__abc_44228_n9898) );
  AND2X2 AND2X2_3911 ( .A(u2__abc_44228_n9899), .B(u2__abc_44228_n5193), .Y(u2__abc_44228_n9901) );
  AND2X2 AND2X2_3912 ( .A(u2__abc_44228_n9902_1), .B(u2__abc_44228_n9900), .Y(u2__abc_44228_n9903) );
  AND2X2 AND2X2_3913 ( .A(u2__abc_44228_n9904), .B(u2__abc_44228_n9905), .Y(u2__abc_44228_n9906) );
  AND2X2 AND2X2_3914 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n5161), .Y(u2__abc_44228_n9908_1) );
  AND2X2 AND2X2_3915 ( .A(u2__abc_44228_n9909), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n9910) );
  AND2X2 AND2X2_3916 ( .A(u2__abc_44228_n9907_1), .B(u2__abc_44228_n9910), .Y(u2__abc_44228_n9911) );
  AND2X2 AND2X2_3917 ( .A(u2__abc_44228_n9912), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_remHi_138__FF_INPUT) );
  AND2X2 AND2X2_3918 ( .A(u2__abc_44228_n3062_bF_buf46), .B(u2_remHi_139_), .Y(u2__abc_44228_n9914) );
  AND2X2 AND2X2_3919 ( .A(u2__abc_44228_n9918_1), .B(u2__abc_44228_n9919_1), .Y(u2__abc_44228_n9920) );
  AND2X2 AND2X2_392 ( .A(_abc_64468_n1692), .B(_abc_64468_n753_bF_buf5), .Y(_abc_64468_n1693) );
  AND2X2 AND2X2_3920 ( .A(u2__abc_44228_n9920), .B(u2__abc_44228_n7547_bF_buf33), .Y(u2__abc_44228_n9921) );
  AND2X2 AND2X2_3921 ( .A(u2__abc_44228_n7548_1_bF_buf34), .B(u2_remHi_137_), .Y(u2__abc_44228_n9922) );
  AND2X2 AND2X2_3922 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n5155_1), .Y(u2__abc_44228_n9925) );
  AND2X2 AND2X2_3923 ( .A(u2__abc_44228_n9926), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n9927) );
  AND2X2 AND2X2_3924 ( .A(u2__abc_44228_n9924_1), .B(u2__abc_44228_n9927), .Y(u2__abc_44228_n9928) );
  AND2X2 AND2X2_3925 ( .A(u2__abc_44228_n9929_1), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_remHi_139__FF_INPUT) );
  AND2X2 AND2X2_3926 ( .A(u2__abc_44228_n3062_bF_buf45), .B(u2_remHi_140_), .Y(u2__abc_44228_n9931) );
  AND2X2 AND2X2_3927 ( .A(u2__abc_44228_n9866), .B(u2__abc_44228_n5195), .Y(u2__abc_44228_n9932) );
  AND2X2 AND2X2_3928 ( .A(u2__abc_44228_n9933), .B(u2__abc_44228_n5164_1), .Y(u2__abc_44228_n9934) );
  AND2X2 AND2X2_3929 ( .A(u2__abc_44228_n9935_1), .B(u2__abc_44228_n9936), .Y(u2__abc_44228_n9937) );
  AND2X2 AND2X2_393 ( .A(aNan_bF_buf3), .B(\a[127] ), .Y(_auto_iopadmap_cc_313_execute_65414_241_) );
  AND2X2 AND2X2_3930 ( .A(u2__abc_44228_n9938), .B(u2__abc_44228_n9939), .Y(u2__abc_44228_n9940_1) );
  AND2X2 AND2X2_3931 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n5147), .Y(u2__abc_44228_n9942) );
  AND2X2 AND2X2_3932 ( .A(u2__abc_44228_n9943), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n9944) );
  AND2X2 AND2X2_3933 ( .A(u2__abc_44228_n9941_1), .B(u2__abc_44228_n9944), .Y(u2__abc_44228_n9945) );
  AND2X2 AND2X2_3934 ( .A(u2__abc_44228_n9946_1), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_remHi_140__FF_INPUT) );
  AND2X2 AND2X2_3935 ( .A(u2__abc_44228_n3062_bF_buf44), .B(u2_remHi_141_), .Y(u2__abc_44228_n9948) );
  AND2X2 AND2X2_3936 ( .A(u2__abc_44228_n9935_1), .B(u2__abc_44228_n5282), .Y(u2__abc_44228_n9949) );
  AND2X2 AND2X2_3937 ( .A(u2__abc_44228_n9949), .B(u2__abc_44228_n5158), .Y(u2__abc_44228_n9950) );
  AND2X2 AND2X2_3938 ( .A(u2__abc_44228_n9952_1), .B(u2__abc_44228_n9951_1), .Y(u2__abc_44228_n9953) );
  AND2X2 AND2X2_3939 ( .A(u2__abc_44228_n9954), .B(u2__abc_44228_n7547_bF_buf31), .Y(u2__abc_44228_n9955) );
  AND2X2 AND2X2_394 ( .A(\a[125] ), .B(\a[126] ), .Y(u1__abc_43968_n152) );
  AND2X2 AND2X2_3940 ( .A(u2__abc_44228_n7548_1_bF_buf32), .B(u2_remHi_139_), .Y(u2__abc_44228_n9956) );
  AND2X2 AND2X2_3941 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n5141), .Y(u2__abc_44228_n9959) );
  AND2X2 AND2X2_3942 ( .A(u2__abc_44228_n9960), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n9961) );
  AND2X2 AND2X2_3943 ( .A(u2__abc_44228_n9958), .B(u2__abc_44228_n9961), .Y(u2__abc_44228_n9962_1) );
  AND2X2 AND2X2_3944 ( .A(u2__abc_44228_n9963_1), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_remHi_141__FF_INPUT) );
  AND2X2 AND2X2_3945 ( .A(u2__abc_44228_n3062_bF_buf43), .B(u2_remHi_142_), .Y(u2__abc_44228_n9965) );
  AND2X2 AND2X2_3946 ( .A(u2__abc_44228_n9935_1), .B(u2__abc_44228_n5283), .Y(u2__abc_44228_n9966) );
  AND2X2 AND2X2_3947 ( .A(u2__abc_44228_n9968_1), .B(u2__abc_44228_n5150), .Y(u2__abc_44228_n9970) );
  AND2X2 AND2X2_3948 ( .A(u2__abc_44228_n9971), .B(u2__abc_44228_n9969), .Y(u2__abc_44228_n9972) );
  AND2X2 AND2X2_3949 ( .A(u2__abc_44228_n9972), .B(u2__abc_44228_n7547_bF_buf30), .Y(u2__abc_44228_n9973_1) );
  AND2X2 AND2X2_395 ( .A(\a[123] ), .B(\a[124] ), .Y(u1__abc_43968_n153) );
  AND2X2 AND2X2_3950 ( .A(u2__abc_44228_n7548_1_bF_buf31), .B(u2_remHi_140_), .Y(u2__abc_44228_n9974_1) );
  AND2X2 AND2X2_3951 ( .A(u2__abc_44228_n2983_bF_buf5), .B(u2__abc_44228_n5130), .Y(u2__abc_44228_n9977) );
  AND2X2 AND2X2_3952 ( .A(u2__abc_44228_n9978), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n9979_1) );
  AND2X2 AND2X2_3953 ( .A(u2__abc_44228_n9976), .B(u2__abc_44228_n9979_1), .Y(u2__abc_44228_n9980) );
  AND2X2 AND2X2_3954 ( .A(u2__abc_44228_n9981), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_remHi_142__FF_INPUT) );
  AND2X2 AND2X2_3955 ( .A(u2__abc_44228_n3062_bF_buf42), .B(u2_remHi_143_), .Y(u2__abc_44228_n9983) );
  AND2X2 AND2X2_3956 ( .A(u2__abc_44228_n9988), .B(u2__abc_44228_n7547_bF_buf29), .Y(u2__abc_44228_n9989) );
  AND2X2 AND2X2_3957 ( .A(u2__abc_44228_n9989), .B(u2__abc_44228_n9987), .Y(u2__abc_44228_n9990_1) );
  AND2X2 AND2X2_3958 ( .A(u2__abc_44228_n7548_1_bF_buf30), .B(u2_remHi_141_), .Y(u2__abc_44228_n9991) );
  AND2X2 AND2X2_3959 ( .A(u2__abc_44228_n2983_bF_buf3), .B(u2__abc_44228_n5124), .Y(u2__abc_44228_n9994) );
  AND2X2 AND2X2_396 ( .A(u1__abc_43968_n152), .B(u1__abc_43968_n153), .Y(u1__abc_43968_n154_1) );
  AND2X2 AND2X2_3960 ( .A(u2__abc_44228_n9995_1), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n9996_1) );
  AND2X2 AND2X2_3961 ( .A(u2__abc_44228_n9993), .B(u2__abc_44228_n9996_1), .Y(u2__abc_44228_n9997) );
  AND2X2 AND2X2_3962 ( .A(u2__abc_44228_n9998), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_remHi_143__FF_INPUT) );
  AND2X2 AND2X2_3963 ( .A(u2__abc_44228_n3062_bF_buf41), .B(u2_remHi_144_), .Y(u2__abc_44228_n10000) );
  AND2X2 AND2X2_3964 ( .A(u2__abc_44228_n7548_1_bF_buf29), .B(u2_remHi_142_), .Y(u2__abc_44228_n10001_1) );
  AND2X2 AND2X2_3965 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5253), .Y(u2__abc_44228_n10002) );
  AND2X2 AND2X2_3966 ( .A(u2__abc_44228_n10003), .B(u2__abc_44228_n5133), .Y(u2__abc_44228_n10004) );
  AND2X2 AND2X2_3967 ( .A(u2__abc_44228_n10005), .B(u2__abc_44228_n10006_1), .Y(u2__abc_44228_n10007_1) );
  AND2X2 AND2X2_3968 ( .A(u2__abc_44228_n7547_bF_buf28), .B(u2__abc_44228_n10007_1), .Y(u2__abc_44228_n10008) );
  AND2X2 AND2X2_3969 ( .A(u2__abc_44228_n2983_bF_buf1), .B(u2__abc_44228_n5116), .Y(u2__abc_44228_n10011) );
  AND2X2 AND2X2_397 ( .A(\a[121] ), .B(\a[122] ), .Y(u1__abc_43968_n155_1) );
  AND2X2 AND2X2_3970 ( .A(u2__abc_44228_n10012_1), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n10013) );
  AND2X2 AND2X2_3971 ( .A(u2__abc_44228_n10010), .B(u2__abc_44228_n10013), .Y(u2__abc_44228_n10014) );
  AND2X2 AND2X2_3972 ( .A(u2__abc_44228_n10015), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_remHi_144__FF_INPUT) );
  AND2X2 AND2X2_3973 ( .A(u2__abc_44228_n3062_bF_buf40), .B(u2_remHi_145_), .Y(u2__abc_44228_n10017_1) );
  AND2X2 AND2X2_3974 ( .A(u2__abc_44228_n10021), .B(u2__abc_44228_n10022), .Y(u2__abc_44228_n10023_1) );
  AND2X2 AND2X2_3975 ( .A(u2__abc_44228_n7547_bF_buf27), .B(u2__abc_44228_n10023_1), .Y(u2__abc_44228_n10024) );
  AND2X2 AND2X2_3976 ( .A(u2__abc_44228_n7548_1_bF_buf28), .B(u2_remHi_143_), .Y(u2__abc_44228_n10025) );
  AND2X2 AND2X2_3977 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n5110), .Y(u2__abc_44228_n10028_1) );
  AND2X2 AND2X2_3978 ( .A(u2__abc_44228_n10029_1), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n10030) );
  AND2X2 AND2X2_3979 ( .A(u2__abc_44228_n10027), .B(u2__abc_44228_n10030), .Y(u2__abc_44228_n10031) );
  AND2X2 AND2X2_398 ( .A(\a[119] ), .B(\a[120] ), .Y(u1__abc_43968_n156) );
  AND2X2 AND2X2_3980 ( .A(u2__abc_44228_n10032), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_remHi_145__FF_INPUT) );
  AND2X2 AND2X2_3981 ( .A(u2__abc_44228_n3062_bF_buf39), .B(u2_remHi_146_), .Y(u2__abc_44228_n10034_1) );
  AND2X2 AND2X2_3982 ( .A(u2__abc_44228_n10003), .B(u2__abc_44228_n5134), .Y(u2__abc_44228_n10035) );
  AND2X2 AND2X2_3983 ( .A(u2__abc_44228_n10036), .B(u2__abc_44228_n5119), .Y(u2__abc_44228_n10038) );
  AND2X2 AND2X2_3984 ( .A(u2__abc_44228_n10039_1), .B(u2__abc_44228_n10037), .Y(u2__abc_44228_n10040_1) );
  AND2X2 AND2X2_3985 ( .A(u2__abc_44228_n10041), .B(u2__abc_44228_n10042), .Y(u2__abc_44228_n10043) );
  AND2X2 AND2X2_3986 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n5094), .Y(u2__abc_44228_n10045_1) );
  AND2X2 AND2X2_3987 ( .A(u2__abc_44228_n10046), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n10047) );
  AND2X2 AND2X2_3988 ( .A(u2__abc_44228_n10044), .B(u2__abc_44228_n10047), .Y(u2__abc_44228_n10048) );
  AND2X2 AND2X2_3989 ( .A(u2__abc_44228_n10049), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_remHi_146__FF_INPUT) );
  AND2X2 AND2X2_399 ( .A(u1__abc_43968_n155_1), .B(u1__abc_43968_n156), .Y(u1__abc_43968_n157_1) );
  AND2X2 AND2X2_3990 ( .A(u2__abc_44228_n3062_bF_buf38), .B(u2_remHi_147_), .Y(u2__abc_44228_n10051_1) );
  AND2X2 AND2X2_3991 ( .A(u2__abc_44228_n10039_1), .B(u2__abc_44228_n5296), .Y(u2__abc_44228_n10052) );
  AND2X2 AND2X2_3992 ( .A(u2__abc_44228_n10052), .B(u2__abc_44228_n5113), .Y(u2__abc_44228_n10053) );
  AND2X2 AND2X2_3993 ( .A(u2__abc_44228_n10055), .B(u2__abc_44228_n10054), .Y(u2__abc_44228_n10056_1) );
  AND2X2 AND2X2_3994 ( .A(u2__abc_44228_n10057), .B(u2__abc_44228_n7547_bF_buf25), .Y(u2__abc_44228_n10058) );
  AND2X2 AND2X2_3995 ( .A(u2__abc_44228_n7548_1_bF_buf26), .B(u2_remHi_145_), .Y(u2__abc_44228_n10059) );
  AND2X2 AND2X2_3996 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n5101), .Y(u2__abc_44228_n10062_1) );
  AND2X2 AND2X2_3997 ( .A(u2__abc_44228_n10063), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n10064) );
  AND2X2 AND2X2_3998 ( .A(u2__abc_44228_n10061_1), .B(u2__abc_44228_n10064), .Y(u2__abc_44228_n10065) );
  AND2X2 AND2X2_3999 ( .A(u2__abc_44228_n10066), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_remHi_147__FF_INPUT) );
  AND2X2 AND2X2_4 ( .A(_abc_64468_n753_bF_buf10), .B(sqrto_3_), .Y(_auto_iopadmap_cc_313_execute_65414_39_) );
  AND2X2 AND2X2_40 ( .A(_abc_64468_n753_bF_buf2), .B(sqrto_39_), .Y(_auto_iopadmap_cc_313_execute_65414_75_) );
  AND2X2 AND2X2_400 ( .A(u1__abc_43968_n154_1), .B(u1__abc_43968_n157_1), .Y(u1__abc_43968_n158_1) );
  AND2X2 AND2X2_4000 ( .A(u2__abc_44228_n3062_bF_buf37), .B(u2_remHi_148_), .Y(u2__abc_44228_n10068) );
  AND2X2 AND2X2_4001 ( .A(u2__abc_44228_n10039_1), .B(u2__abc_44228_n5297_1), .Y(u2__abc_44228_n10069) );
  AND2X2 AND2X2_4002 ( .A(u2__abc_44228_n10071), .B(u2__abc_44228_n5097), .Y(u2__abc_44228_n10072_1) );
  AND2X2 AND2X2_4003 ( .A(u2__abc_44228_n10073_1), .B(u2__abc_44228_n10074), .Y(u2__abc_44228_n10075) );
  AND2X2 AND2X2_4004 ( .A(u2__abc_44228_n10076), .B(u2__abc_44228_n10077), .Y(u2__abc_44228_n10078_1) );
  AND2X2 AND2X2_4005 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n5087), .Y(u2__abc_44228_n10080) );
  AND2X2 AND2X2_4006 ( .A(u2__abc_44228_n10081), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n10082) );
  AND2X2 AND2X2_4007 ( .A(u2__abc_44228_n10079), .B(u2__abc_44228_n10082), .Y(u2__abc_44228_n10083_1) );
  AND2X2 AND2X2_4008 ( .A(u2__abc_44228_n10084_1), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_remHi_148__FF_INPUT) );
  AND2X2 AND2X2_4009 ( .A(u2__abc_44228_n3062_bF_buf36), .B(u2_remHi_149_), .Y(u2__abc_44228_n10086) );
  AND2X2 AND2X2_401 ( .A(\a[118] ), .B(\a[115] ), .Y(u1__abc_43968_n159) );
  AND2X2 AND2X2_4010 ( .A(u2__abc_44228_n10073_1), .B(u2__abc_44228_n5302), .Y(u2__abc_44228_n10087) );
  AND2X2 AND2X2_4011 ( .A(u2__abc_44228_n10091), .B(u2__abc_44228_n7547_bF_buf23), .Y(u2__abc_44228_n10092) );
  AND2X2 AND2X2_4012 ( .A(u2__abc_44228_n10092), .B(u2__abc_44228_n10089_1), .Y(u2__abc_44228_n10093) );
  AND2X2 AND2X2_4013 ( .A(u2__abc_44228_n7548_1_bF_buf24), .B(u2_remHi_147_), .Y(u2__abc_44228_n10094_1) );
  AND2X2 AND2X2_4014 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n5081), .Y(u2__abc_44228_n10097) );
  AND2X2 AND2X2_4015 ( .A(u2__abc_44228_n10098), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n10099) );
  AND2X2 AND2X2_4016 ( .A(u2__abc_44228_n10096), .B(u2__abc_44228_n10099), .Y(u2__abc_44228_n10100_1) );
  AND2X2 AND2X2_4017 ( .A(u2__abc_44228_n10101), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_remHi_149__FF_INPUT) );
  AND2X2 AND2X2_4018 ( .A(u2__abc_44228_n3062_bF_buf35), .B(u2_remHi_150_), .Y(u2__abc_44228_n10103) );
  AND2X2 AND2X2_4019 ( .A(u2__abc_44228_n10073_1), .B(u2__abc_44228_n5303), .Y(u2__abc_44228_n10104) );
  AND2X2 AND2X2_402 ( .A(u1__abc_43968_n159), .B(\a[116] ), .Y(u1__abc_43968_n160) );
  AND2X2 AND2X2_4020 ( .A(u2__abc_44228_n10106_1), .B(u2__abc_44228_n5090), .Y(u2__abc_44228_n10108) );
  AND2X2 AND2X2_4021 ( .A(u2__abc_44228_n10109), .B(u2__abc_44228_n10107), .Y(u2__abc_44228_n10110) );
  AND2X2 AND2X2_4022 ( .A(u2__abc_44228_n10110), .B(u2__abc_44228_n7547_bF_buf22), .Y(u2__abc_44228_n10111_1) );
  AND2X2 AND2X2_4023 ( .A(u2__abc_44228_n7548_1_bF_buf23), .B(u2_remHi_148_), .Y(u2__abc_44228_n10112) );
  AND2X2 AND2X2_4024 ( .A(u2__abc_44228_n2983_bF_buf133), .B(u2__abc_44228_n5064), .Y(u2__abc_44228_n10115) );
  AND2X2 AND2X2_4025 ( .A(u2__abc_44228_n10116_1), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n10117_1) );
  AND2X2 AND2X2_4026 ( .A(u2__abc_44228_n10114), .B(u2__abc_44228_n10117_1), .Y(u2__abc_44228_n10118) );
  AND2X2 AND2X2_4027 ( .A(u2__abc_44228_n10119), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_remHi_150__FF_INPUT) );
  AND2X2 AND2X2_4028 ( .A(u2__abc_44228_n3062_bF_buf34), .B(u2_remHi_151_), .Y(u2__abc_44228_n10121) );
  AND2X2 AND2X2_4029 ( .A(u2__abc_44228_n10126), .B(u2__abc_44228_n7547_bF_buf21), .Y(u2__abc_44228_n10127_1) );
  AND2X2 AND2X2_403 ( .A(\a[113] ), .B(\a[114] ), .Y(u1__abc_43968_n161_1) );
  AND2X2 AND2X2_4030 ( .A(u2__abc_44228_n10127_1), .B(u2__abc_44228_n10125), .Y(u2__abc_44228_n10128_1) );
  AND2X2 AND2X2_4031 ( .A(u2__abc_44228_n7548_1_bF_buf22), .B(u2_remHi_149_), .Y(u2__abc_44228_n10129) );
  AND2X2 AND2X2_4032 ( .A(u2__abc_44228_n2983_bF_buf131), .B(u2__abc_44228_n5071_1), .Y(u2__abc_44228_n10132) );
  AND2X2 AND2X2_4033 ( .A(u2__abc_44228_n10133_1), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n10134) );
  AND2X2 AND2X2_4034 ( .A(u2__abc_44228_n10131), .B(u2__abc_44228_n10134), .Y(u2__abc_44228_n10135) );
  AND2X2 AND2X2_4035 ( .A(u2__abc_44228_n10136), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_remHi_151__FF_INPUT) );
  AND2X2 AND2X2_4036 ( .A(u2__abc_44228_n3062_bF_buf33), .B(u2_remHi_152_), .Y(u2__abc_44228_n10138_1) );
  AND2X2 AND2X2_4037 ( .A(u2__abc_44228_n10003), .B(u2__abc_44228_n5136_1), .Y(u2__abc_44228_n10139_1) );
  AND2X2 AND2X2_4038 ( .A(u2__abc_44228_n10140), .B(u2__abc_44228_n5067), .Y(u2__abc_44228_n10142) );
  AND2X2 AND2X2_4039 ( .A(u2__abc_44228_n10143), .B(u2__abc_44228_n10141), .Y(u2__abc_44228_n10144_1) );
  AND2X2 AND2X2_404 ( .A(a_112_bF_buf1), .B(\a[117] ), .Y(u1__abc_43968_n162_1) );
  AND2X2 AND2X2_4040 ( .A(u2__abc_44228_n10145), .B(u2__abc_44228_n10146), .Y(u2__abc_44228_n10147) );
  AND2X2 AND2X2_4041 ( .A(u2__abc_44228_n2983_bF_buf129), .B(u2__abc_44228_n5057), .Y(u2__abc_44228_n10149_1) );
  AND2X2 AND2X2_4042 ( .A(u2__abc_44228_n10150_1), .B(u2__abc_44228_n2972_bF_buf61), .Y(u2__abc_44228_n10151) );
  AND2X2 AND2X2_4043 ( .A(u2__abc_44228_n10148), .B(u2__abc_44228_n10151), .Y(u2__abc_44228_n10152) );
  AND2X2 AND2X2_4044 ( .A(u2__abc_44228_n10153), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_remHi_152__FF_INPUT) );
  AND2X2 AND2X2_4045 ( .A(u2__abc_44228_n3062_bF_buf32), .B(u2_remHi_153_), .Y(u2__abc_44228_n10155_1) );
  AND2X2 AND2X2_4046 ( .A(u2__abc_44228_n10143), .B(u2__abc_44228_n5314), .Y(u2__abc_44228_n10156) );
  AND2X2 AND2X2_4047 ( .A(u2__abc_44228_n10156), .B(u2__abc_44228_n5074), .Y(u2__abc_44228_n10157) );
  AND2X2 AND2X2_4048 ( .A(u2__abc_44228_n10159), .B(u2__abc_44228_n10158), .Y(u2__abc_44228_n10160_1) );
  AND2X2 AND2X2_4049 ( .A(u2__abc_44228_n10161_1), .B(u2__abc_44228_n7547_bF_buf19), .Y(u2__abc_44228_n10162) );
  AND2X2 AND2X2_405 ( .A(u1__abc_43968_n161_1), .B(u1__abc_43968_n162_1), .Y(u1__abc_43968_n163) );
  AND2X2 AND2X2_4050 ( .A(u2__abc_44228_n7548_1_bF_buf20), .B(u2_remHi_151_), .Y(u2__abc_44228_n10163) );
  AND2X2 AND2X2_4051 ( .A(u2__abc_44228_n2983_bF_buf127), .B(u2__abc_44228_n5051_1), .Y(u2__abc_44228_n10166_1) );
  AND2X2 AND2X2_4052 ( .A(u2__abc_44228_n10167), .B(u2__abc_44228_n2972_bF_buf60), .Y(u2__abc_44228_n10168) );
  AND2X2 AND2X2_4053 ( .A(u2__abc_44228_n10165), .B(u2__abc_44228_n10168), .Y(u2__abc_44228_n10169) );
  AND2X2 AND2X2_4054 ( .A(u2__abc_44228_n10170), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_remHi_153__FF_INPUT) );
  AND2X2 AND2X2_4055 ( .A(u2__abc_44228_n3062_bF_buf31), .B(u2_remHi_154_), .Y(u2__abc_44228_n10172_1) );
  AND2X2 AND2X2_4056 ( .A(u2__abc_44228_n10143), .B(u2__abc_44228_n5315_1), .Y(u2__abc_44228_n10173) );
  AND2X2 AND2X2_4057 ( .A(u2__abc_44228_n10175), .B(u2__abc_44228_n5060), .Y(u2__abc_44228_n10177_1) );
  AND2X2 AND2X2_4058 ( .A(u2__abc_44228_n10178), .B(u2__abc_44228_n10176), .Y(u2__abc_44228_n10179) );
  AND2X2 AND2X2_4059 ( .A(u2__abc_44228_n10179), .B(u2__abc_44228_n7547_bF_buf18), .Y(u2__abc_44228_n10180) );
  AND2X2 AND2X2_406 ( .A(u1__abc_43968_n163), .B(u1__abc_43968_n160), .Y(u1__abc_43968_n164_1) );
  AND2X2 AND2X2_4060 ( .A(u2__abc_44228_n7548_1_bF_buf19), .B(u2_remHi_152_), .Y(u2__abc_44228_n10181) );
  AND2X2 AND2X2_4061 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n5042_1), .Y(u2__abc_44228_n10184) );
  AND2X2 AND2X2_4062 ( .A(u2__abc_44228_n10185), .B(u2__abc_44228_n2972_bF_buf59), .Y(u2__abc_44228_n10186) );
  AND2X2 AND2X2_4063 ( .A(u2__abc_44228_n10183_1), .B(u2__abc_44228_n10186), .Y(u2__abc_44228_n10187) );
  AND2X2 AND2X2_4064 ( .A(u2__abc_44228_n10188_1), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_remHi_154__FF_INPUT) );
  AND2X2 AND2X2_4065 ( .A(u2__abc_44228_n3062_bF_buf30), .B(u2_remHi_155_), .Y(u2__abc_44228_n10190) );
  AND2X2 AND2X2_4066 ( .A(u2__abc_44228_n10195), .B(u2__abc_44228_n7547_bF_buf17), .Y(u2__abc_44228_n10196) );
  AND2X2 AND2X2_4067 ( .A(u2__abc_44228_n10196), .B(u2__abc_44228_n10194_1), .Y(u2__abc_44228_n10197) );
  AND2X2 AND2X2_4068 ( .A(u2__abc_44228_n7548_1_bF_buf18), .B(u2_remHi_153_), .Y(u2__abc_44228_n10198) );
  AND2X2 AND2X2_4069 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n5036), .Y(u2__abc_44228_n10201) );
  AND2X2 AND2X2_407 ( .A(u1__abc_43968_n158_1), .B(u1__abc_43968_n164_1), .Y(u1_xinf) );
  AND2X2 AND2X2_4070 ( .A(u2__abc_44228_n10202), .B(u2__abc_44228_n2972_bF_buf58), .Y(u2__abc_44228_n10203) );
  AND2X2 AND2X2_4071 ( .A(u2__abc_44228_n10200), .B(u2__abc_44228_n10203), .Y(u2__abc_44228_n10204_1) );
  AND2X2 AND2X2_4072 ( .A(u2__abc_44228_n10205_1), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_remHi_155__FF_INPUT) );
  AND2X2 AND2X2_4073 ( .A(u2__abc_44228_n3062_bF_buf29), .B(u2_remHi_156_), .Y(u2__abc_44228_n10207) );
  AND2X2 AND2X2_4074 ( .A(u2__abc_44228_n10140), .B(u2__abc_44228_n5076), .Y(u2__abc_44228_n10208) );
  AND2X2 AND2X2_4075 ( .A(u2__abc_44228_n10209), .B(u2__abc_44228_n5045), .Y(u2__abc_44228_n10210_1) );
  AND2X2 AND2X2_4076 ( .A(u2__abc_44228_n10211), .B(u2__abc_44228_n10212), .Y(u2__abc_44228_n10213) );
  AND2X2 AND2X2_4077 ( .A(u2__abc_44228_n10214), .B(u2__abc_44228_n10215_1), .Y(u2__abc_44228_n10216_1) );
  AND2X2 AND2X2_4078 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n5028), .Y(u2__abc_44228_n10218) );
  AND2X2 AND2X2_4079 ( .A(u2__abc_44228_n10219), .B(u2__abc_44228_n2972_bF_buf57), .Y(u2__abc_44228_n10220) );
  AND2X2 AND2X2_408 ( .A(u1__abc_43968_n166), .B(u1__abc_43968_n167), .Y(u1__abc_43968_n168) );
  AND2X2 AND2X2_4080 ( .A(u2__abc_44228_n10217), .B(u2__abc_44228_n10220), .Y(u2__abc_44228_n10221_1) );
  AND2X2 AND2X2_4081 ( .A(u2__abc_44228_n10222), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_remHi_156__FF_INPUT) );
  AND2X2 AND2X2_4082 ( .A(u2__abc_44228_n3062_bF_buf28), .B(u2_remHi_157_), .Y(u2__abc_44228_n10224) );
  AND2X2 AND2X2_4083 ( .A(u2__abc_44228_n10211), .B(u2__abc_44228_n5323), .Y(u2__abc_44228_n10226_1) );
  AND2X2 AND2X2_4084 ( .A(u2__abc_44228_n10229), .B(u2__abc_44228_n10227_1), .Y(u2__abc_44228_n10230) );
  AND2X2 AND2X2_4085 ( .A(u2__abc_44228_n10230), .B(u2__abc_44228_n7547_bF_buf15), .Y(u2__abc_44228_n10231) );
  AND2X2 AND2X2_4086 ( .A(u2__abc_44228_n7548_1_bF_buf16), .B(u2_remHi_155_), .Y(u2__abc_44228_n10232_1) );
  AND2X2 AND2X2_4087 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n5022), .Y(u2__abc_44228_n10235) );
  AND2X2 AND2X2_4088 ( .A(u2__abc_44228_n10236), .B(u2__abc_44228_n2972_bF_buf56), .Y(u2__abc_44228_n10237_1) );
  AND2X2 AND2X2_4089 ( .A(u2__abc_44228_n10234), .B(u2__abc_44228_n10237_1), .Y(u2__abc_44228_n10238_1) );
  AND2X2 AND2X2_409 ( .A(u1__abc_43968_n169), .B(u1__abc_43968_n170_1), .Y(u1__abc_43968_n171_1) );
  AND2X2 AND2X2_4090 ( .A(u2__abc_44228_n10239), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_remHi_157__FF_INPUT) );
  AND2X2 AND2X2_4091 ( .A(u2__abc_44228_n3062_bF_buf27), .B(u2_remHi_158_), .Y(u2__abc_44228_n10241) );
  AND2X2 AND2X2_4092 ( .A(u2__abc_44228_n10209), .B(u2__abc_44228_n5046), .Y(u2__abc_44228_n10242) );
  AND2X2 AND2X2_4093 ( .A(u2__abc_44228_n10243_1), .B(u2__abc_44228_n5031), .Y(u2__abc_44228_n10245) );
  AND2X2 AND2X2_4094 ( .A(u2__abc_44228_n10246), .B(u2__abc_44228_n10244), .Y(u2__abc_44228_n10247) );
  AND2X2 AND2X2_4095 ( .A(u2__abc_44228_n10247), .B(u2__abc_44228_n7547_bF_buf14), .Y(u2__abc_44228_n10248_1) );
  AND2X2 AND2X2_4096 ( .A(u2__abc_44228_n7548_1_bF_buf15), .B(u2_remHi_156_), .Y(u2__abc_44228_n10249_1) );
  AND2X2 AND2X2_4097 ( .A(u2__abc_44228_n2983_bF_buf119), .B(u2__abc_44228_n5003), .Y(u2__abc_44228_n10252) );
  AND2X2 AND2X2_4098 ( .A(u2__abc_44228_n10253), .B(u2__abc_44228_n2972_bF_buf55), .Y(u2__abc_44228_n10254_1) );
  AND2X2 AND2X2_4099 ( .A(u2__abc_44228_n10251), .B(u2__abc_44228_n10254_1), .Y(u2__abc_44228_n10255) );
  AND2X2 AND2X2_41 ( .A(_abc_64468_n753_bF_buf1), .B(sqrto_40_), .Y(_auto_iopadmap_cc_313_execute_65414_76_) );
  AND2X2 AND2X2_410 ( .A(u1__abc_43968_n168), .B(u1__abc_43968_n171_1), .Y(u1__abc_43968_n172) );
  AND2X2 AND2X2_4100 ( .A(u2__abc_44228_n10256), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_remHi_158__FF_INPUT) );
  AND2X2 AND2X2_4101 ( .A(u2__abc_44228_n3062_bF_buf26), .B(u2_remHi_159_), .Y(u2__abc_44228_n10258) );
  AND2X2 AND2X2_4102 ( .A(u2__abc_44228_n10263), .B(u2__abc_44228_n7547_bF_buf13), .Y(u2__abc_44228_n10264) );
  AND2X2 AND2X2_4103 ( .A(u2__abc_44228_n10264), .B(u2__abc_44228_n10262), .Y(u2__abc_44228_n10265_1) );
  AND2X2 AND2X2_4104 ( .A(u2__abc_44228_n7548_1_bF_buf14), .B(u2_remHi_157_), .Y(u2__abc_44228_n10266) );
  AND2X2 AND2X2_4105 ( .A(u2__abc_44228_n2983_bF_buf117), .B(u2__abc_44228_n5010), .Y(u2__abc_44228_n10269) );
  AND2X2 AND2X2_4106 ( .A(u2__abc_44228_n10270_1), .B(u2__abc_44228_n2972_bF_buf54), .Y(u2__abc_44228_n10271_1) );
  AND2X2 AND2X2_4107 ( .A(u2__abc_44228_n10268), .B(u2__abc_44228_n10271_1), .Y(u2__abc_44228_n10272) );
  AND2X2 AND2X2_4108 ( .A(u2__abc_44228_n10273), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_remHi_159__FF_INPUT) );
  AND2X2 AND2X2_4109 ( .A(u2__abc_44228_n3062_bF_buf25), .B(u2_remHi_160_), .Y(u2__abc_44228_n10275) );
  AND2X2 AND2X2_411 ( .A(u1__abc_43968_n173_1), .B(u1__abc_43968_n174_1), .Y(u1__abc_43968_n175) );
  AND2X2 AND2X2_4110 ( .A(u2__abc_44228_n7548_1_bF_buf13), .B(u2_remHi_158_), .Y(u2__abc_44228_n10276_1) );
  AND2X2 AND2X2_4111 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5254), .Y(u2__abc_44228_n10277) );
  AND2X2 AND2X2_4112 ( .A(u2__abc_44228_n10278), .B(u2__abc_44228_n5006), .Y(u2__abc_44228_n10280) );
  AND2X2 AND2X2_4113 ( .A(u2__abc_44228_n10281_1), .B(u2__abc_44228_n10279), .Y(u2__abc_44228_n10282_1) );
  AND2X2 AND2X2_4114 ( .A(u2__abc_44228_n7547_bF_buf12), .B(u2__abc_44228_n10282_1), .Y(u2__abc_44228_n10283) );
  AND2X2 AND2X2_4115 ( .A(u2__abc_44228_n2983_bF_buf115), .B(u2__abc_44228_n4996_1), .Y(u2__abc_44228_n10286) );
  AND2X2 AND2X2_4116 ( .A(u2__abc_44228_n10287_1), .B(u2__abc_44228_n2972_bF_buf53), .Y(u2__abc_44228_n10288) );
  AND2X2 AND2X2_4117 ( .A(u2__abc_44228_n10285), .B(u2__abc_44228_n10288), .Y(u2__abc_44228_n10289) );
  AND2X2 AND2X2_4118 ( .A(u2__abc_44228_n10290), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_remHi_160__FF_INPUT) );
  AND2X2 AND2X2_4119 ( .A(u2__abc_44228_n3062_bF_buf24), .B(u2_remHi_161_), .Y(u2__abc_44228_n10292_1) );
  AND2X2 AND2X2_412 ( .A(u1__abc_43968_n176), .B(u1__abc_43968_n177_1), .Y(u1__abc_43968_n178_1) );
  AND2X2 AND2X2_4120 ( .A(u2__abc_44228_n10296), .B(u2__abc_44228_n10297), .Y(u2__abc_44228_n10298_1) );
  AND2X2 AND2X2_4121 ( .A(u2__abc_44228_n7547_bF_buf11), .B(u2__abc_44228_n10298_1), .Y(u2__abc_44228_n10299) );
  AND2X2 AND2X2_4122 ( .A(u2__abc_44228_n7548_1_bF_buf12), .B(u2_remHi_159_), .Y(u2__abc_44228_n10300) );
  AND2X2 AND2X2_4123 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n4990), .Y(u2__abc_44228_n10303_1) );
  AND2X2 AND2X2_4124 ( .A(u2__abc_44228_n10304_1), .B(u2__abc_44228_n2972_bF_buf52), .Y(u2__abc_44228_n10305) );
  AND2X2 AND2X2_4125 ( .A(u2__abc_44228_n10302), .B(u2__abc_44228_n10305), .Y(u2__abc_44228_n10306) );
  AND2X2 AND2X2_4126 ( .A(u2__abc_44228_n10307), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_remHi_161__FF_INPUT) );
  AND2X2 AND2X2_4127 ( .A(u2__abc_44228_n3062_bF_buf23), .B(u2_remHi_162_), .Y(u2__abc_44228_n10309_1) );
  AND2X2 AND2X2_4128 ( .A(u2__abc_44228_n10278), .B(u2__abc_44228_n5014_1), .Y(u2__abc_44228_n10310) );
  AND2X2 AND2X2_4129 ( .A(u2__abc_44228_n10311), .B(u2__abc_44228_n4999), .Y(u2__abc_44228_n10313) );
  AND2X2 AND2X2_413 ( .A(u1__abc_43968_n175), .B(u1__abc_43968_n178_1), .Y(u1__abc_43968_n179) );
  AND2X2 AND2X2_4130 ( .A(u2__abc_44228_n10314_1), .B(u2__abc_44228_n10312), .Y(u2__abc_44228_n10315_1) );
  AND2X2 AND2X2_4131 ( .A(u2__abc_44228_n10316), .B(u2__abc_44228_n10317), .Y(u2__abc_44228_n10318) );
  AND2X2 AND2X2_4132 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n4974), .Y(u2__abc_44228_n10320_1) );
  AND2X2 AND2X2_4133 ( .A(u2__abc_44228_n10321), .B(u2__abc_44228_n2972_bF_buf51), .Y(u2__abc_44228_n10322) );
  AND2X2 AND2X2_4134 ( .A(u2__abc_44228_n10319), .B(u2__abc_44228_n10322), .Y(u2__abc_44228_n10323) );
  AND2X2 AND2X2_4135 ( .A(u2__abc_44228_n10324), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_remHi_162__FF_INPUT) );
  AND2X2 AND2X2_4136 ( .A(u2__abc_44228_n3062_bF_buf22), .B(u2_remHi_163_), .Y(u2__abc_44228_n10326_1) );
  AND2X2 AND2X2_4137 ( .A(u2__abc_44228_n10331), .B(u2__abc_44228_n10328), .Y(u2__abc_44228_n10332_1) );
  AND2X2 AND2X2_4138 ( .A(u2__abc_44228_n10332_1), .B(u2__abc_44228_n7547_bF_buf9), .Y(u2__abc_44228_n10333_1) );
  AND2X2 AND2X2_4139 ( .A(u2__abc_44228_n7548_1_bF_buf10), .B(u2_remHi_161_), .Y(u2__abc_44228_n10334) );
  AND2X2 AND2X2_414 ( .A(u1__abc_43968_n172), .B(u1__abc_43968_n179), .Y(u1__abc_43968_n180_1) );
  AND2X2 AND2X2_4140 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n4981), .Y(u2__abc_44228_n10337) );
  AND2X2 AND2X2_4141 ( .A(u2__abc_44228_n10338), .B(u2__abc_44228_n2972_bF_buf50), .Y(u2__abc_44228_n10339_1) );
  AND2X2 AND2X2_4142 ( .A(u2__abc_44228_n10336), .B(u2__abc_44228_n10339_1), .Y(u2__abc_44228_n10340_1) );
  AND2X2 AND2X2_4143 ( .A(u2__abc_44228_n10341), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_remHi_163__FF_INPUT) );
  AND2X2 AND2X2_4144 ( .A(u2__abc_44228_n3062_bF_buf21), .B(u2_remHi_164_), .Y(u2__abc_44228_n10343) );
  AND2X2 AND2X2_4145 ( .A(u2__abc_44228_n10278), .B(u2__abc_44228_n5015), .Y(u2__abc_44228_n10344) );
  AND2X2 AND2X2_4146 ( .A(u2__abc_44228_n10345), .B(u2__abc_44228_n4977), .Y(u2__abc_44228_n10346_1) );
  AND2X2 AND2X2_4147 ( .A(u2__abc_44228_n10347_1), .B(u2__abc_44228_n10348), .Y(u2__abc_44228_n10349) );
  AND2X2 AND2X2_4148 ( .A(u2__abc_44228_n10350), .B(u2__abc_44228_n10351), .Y(u2__abc_44228_n10352) );
  AND2X2 AND2X2_4149 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n4967_1), .Y(u2__abc_44228_n10354_1) );
  AND2X2 AND2X2_415 ( .A(u1__abc_43968_n181_1), .B(u1__abc_43968_n182), .Y(u1__abc_43968_n183) );
  AND2X2 AND2X2_4150 ( .A(u2__abc_44228_n10355), .B(u2__abc_44228_n2972_bF_buf49), .Y(u2__abc_44228_n10356) );
  AND2X2 AND2X2_4151 ( .A(u2__abc_44228_n10353_1), .B(u2__abc_44228_n10356), .Y(u2__abc_44228_n10357) );
  AND2X2 AND2X2_4152 ( .A(u2__abc_44228_n10358), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_remHi_164__FF_INPUT) );
  AND2X2 AND2X2_4153 ( .A(u2__abc_44228_n3062_bF_buf20), .B(u2_remHi_165_), .Y(u2__abc_44228_n10360_1) );
  AND2X2 AND2X2_4154 ( .A(u2__abc_44228_n10347_1), .B(u2__abc_44228_n5340), .Y(u2__abc_44228_n10361_1) );
  AND2X2 AND2X2_4155 ( .A(u2__abc_44228_n10361_1), .B(u2__abc_44228_n4984), .Y(u2__abc_44228_n10362) );
  AND2X2 AND2X2_4156 ( .A(u2__abc_44228_n10364), .B(u2__abc_44228_n10363), .Y(u2__abc_44228_n10365) );
  AND2X2 AND2X2_4157 ( .A(u2__abc_44228_n10366), .B(u2__abc_44228_n7547_bF_buf7), .Y(u2__abc_44228_n10367_1) );
  AND2X2 AND2X2_4158 ( .A(u2__abc_44228_n7548_1_bF_buf8), .B(u2_remHi_163_), .Y(u2__abc_44228_n10368_1) );
  AND2X2 AND2X2_4159 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n4961), .Y(u2__abc_44228_n10371) );
  AND2X2 AND2X2_416 ( .A(u1__abc_43968_n184), .B(u1__abc_43968_n185_1), .Y(u1__abc_43968_n186_1) );
  AND2X2 AND2X2_4160 ( .A(u2__abc_44228_n10372), .B(u2__abc_44228_n2972_bF_buf48), .Y(u2__abc_44228_n10373) );
  AND2X2 AND2X2_4161 ( .A(u2__abc_44228_n10370), .B(u2__abc_44228_n10373), .Y(u2__abc_44228_n10374_1) );
  AND2X2 AND2X2_4162 ( .A(u2__abc_44228_n10375_1), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_remHi_165__FF_INPUT) );
  AND2X2 AND2X2_4163 ( .A(u2__abc_44228_n3062_bF_buf19), .B(u2_remHi_166_), .Y(u2__abc_44228_n10377) );
  AND2X2 AND2X2_4164 ( .A(u2__abc_44228_n10347_1), .B(u2__abc_44228_n5341), .Y(u2__abc_44228_n10378) );
  AND2X2 AND2X2_4165 ( .A(u2__abc_44228_n10380), .B(u2__abc_44228_n4970), .Y(u2__abc_44228_n10382_1) );
  AND2X2 AND2X2_4166 ( .A(u2__abc_44228_n10383), .B(u2__abc_44228_n10381_1), .Y(u2__abc_44228_n10384) );
  AND2X2 AND2X2_4167 ( .A(u2__abc_44228_n10384), .B(u2__abc_44228_n7547_bF_buf6), .Y(u2__abc_44228_n10385) );
  AND2X2 AND2X2_4168 ( .A(u2__abc_44228_n7548_1_bF_buf7), .B(u2_remHi_164_), .Y(u2__abc_44228_n10386) );
  AND2X2 AND2X2_4169 ( .A(u2__abc_44228_n2983_bF_buf105), .B(u2__abc_44228_n4944), .Y(u2__abc_44228_n10389_1) );
  AND2X2 AND2X2_417 ( .A(u1__abc_43968_n183), .B(u1__abc_43968_n186_1), .Y(u1__abc_43968_n187) );
  AND2X2 AND2X2_4170 ( .A(u2__abc_44228_n10390), .B(u2__abc_44228_n2972_bF_buf47), .Y(u2__abc_44228_n10391) );
  AND2X2 AND2X2_4171 ( .A(u2__abc_44228_n10388_1), .B(u2__abc_44228_n10391), .Y(u2__abc_44228_n10392) );
  AND2X2 AND2X2_4172 ( .A(u2__abc_44228_n10393), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_remHi_166__FF_INPUT) );
  AND2X2 AND2X2_4173 ( .A(u2__abc_44228_n3062_bF_buf18), .B(u2_remHi_167_), .Y(u2__abc_44228_n10395_1) );
  AND2X2 AND2X2_4174 ( .A(u2__abc_44228_n10400), .B(u2__abc_44228_n7547_bF_buf5), .Y(u2__abc_44228_n10401) );
  AND2X2 AND2X2_4175 ( .A(u2__abc_44228_n10401), .B(u2__abc_44228_n10399), .Y(u2__abc_44228_n10402_1) );
  AND2X2 AND2X2_4176 ( .A(u2__abc_44228_n7548_1_bF_buf6), .B(u2_remHi_165_), .Y(u2__abc_44228_n10403_1) );
  AND2X2 AND2X2_4177 ( .A(u2__abc_44228_n2983_bF_buf103), .B(u2__abc_44228_n4951), .Y(u2__abc_44228_n10406) );
  AND2X2 AND2X2_4178 ( .A(u2__abc_44228_n10407), .B(u2__abc_44228_n2972_bF_buf46), .Y(u2__abc_44228_n10408) );
  AND2X2 AND2X2_4179 ( .A(u2__abc_44228_n10405), .B(u2__abc_44228_n10408), .Y(u2__abc_44228_n10409_1) );
  AND2X2 AND2X2_418 ( .A(u1__abc_43968_n188_1), .B(u1__abc_43968_n189_1), .Y(u1__abc_43968_n190) );
  AND2X2 AND2X2_4180 ( .A(u2__abc_44228_n10410_1), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_remHi_167__FF_INPUT) );
  AND2X2 AND2X2_4181 ( .A(u2__abc_44228_n3062_bF_buf17), .B(u2_remHi_168_), .Y(u2__abc_44228_n10412) );
  AND2X2 AND2X2_4182 ( .A(u2__abc_44228_n10278), .B(u2__abc_44228_n5016), .Y(u2__abc_44228_n10413) );
  AND2X2 AND2X2_4183 ( .A(u2__abc_44228_n10414), .B(u2__abc_44228_n4947), .Y(u2__abc_44228_n10416_1) );
  AND2X2 AND2X2_4184 ( .A(u2__abc_44228_n10417_1), .B(u2__abc_44228_n10415), .Y(u2__abc_44228_n10418) );
  AND2X2 AND2X2_4185 ( .A(u2__abc_44228_n10419), .B(u2__abc_44228_n10420), .Y(u2__abc_44228_n10421) );
  AND2X2 AND2X2_4186 ( .A(u2__abc_44228_n2983_bF_buf101), .B(u2__abc_44228_n4937), .Y(u2__abc_44228_n10423_1) );
  AND2X2 AND2X2_4187 ( .A(u2__abc_44228_n10424_1), .B(u2__abc_44228_n2972_bF_buf45), .Y(u2__abc_44228_n10425) );
  AND2X2 AND2X2_4188 ( .A(u2__abc_44228_n10422), .B(u2__abc_44228_n10425), .Y(u2__abc_44228_n10426) );
  AND2X2 AND2X2_4189 ( .A(u2__abc_44228_n10427), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_remHi_168__FF_INPUT) );
  AND2X2 AND2X2_419 ( .A(u1__abc_43968_n191), .B(u1__abc_43968_n192_1), .Y(u1__abc_43968_n193_1) );
  AND2X2 AND2X2_4190 ( .A(u2__abc_44228_n3062_bF_buf16), .B(u2_remHi_169_), .Y(u2__abc_44228_n10429) );
  AND2X2 AND2X2_4191 ( .A(u2__abc_44228_n10417_1), .B(u2__abc_44228_n5352_1), .Y(u2__abc_44228_n10430_1) );
  AND2X2 AND2X2_4192 ( .A(u2__abc_44228_n10430_1), .B(u2__abc_44228_n4954), .Y(u2__abc_44228_n10431_1) );
  AND2X2 AND2X2_4193 ( .A(u2__abc_44228_n10433), .B(u2__abc_44228_n10432), .Y(u2__abc_44228_n10434) );
  AND2X2 AND2X2_4194 ( .A(u2__abc_44228_n10435), .B(u2__abc_44228_n7547_bF_buf3), .Y(u2__abc_44228_n10436) );
  AND2X2 AND2X2_4195 ( .A(u2__abc_44228_n7548_1_bF_buf4), .B(u2_remHi_167_), .Y(u2__abc_44228_n10437_1) );
  AND2X2 AND2X2_4196 ( .A(u2__abc_44228_n2983_bF_buf99), .B(u2__abc_44228_n4931), .Y(u2__abc_44228_n10440) );
  AND2X2 AND2X2_4197 ( .A(u2__abc_44228_n10441), .B(u2__abc_44228_n2972_bF_buf44), .Y(u2__abc_44228_n10442) );
  AND2X2 AND2X2_4198 ( .A(u2__abc_44228_n10439), .B(u2__abc_44228_n10442), .Y(u2__abc_44228_n10443) );
  AND2X2 AND2X2_4199 ( .A(u2__abc_44228_n10444_1), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_remHi_169__FF_INPUT) );
  AND2X2 AND2X2_42 ( .A(_abc_64468_n753_bF_buf0), .B(sqrto_41_), .Y(_auto_iopadmap_cc_313_execute_65414_77_) );
  AND2X2 AND2X2_420 ( .A(u1__abc_43968_n190), .B(u1__abc_43968_n193_1), .Y(u1__abc_43968_n194) );
  AND2X2 AND2X2_4200 ( .A(u2__abc_44228_n3062_bF_buf15), .B(u2_remHi_170_), .Y(u2__abc_44228_n10446) );
  AND2X2 AND2X2_4201 ( .A(u2__abc_44228_n10417_1), .B(u2__abc_44228_n5353), .Y(u2__abc_44228_n10447) );
  AND2X2 AND2X2_4202 ( .A(u2__abc_44228_n10449), .B(u2__abc_44228_n4940), .Y(u2__abc_44228_n10451_1) );
  AND2X2 AND2X2_4203 ( .A(u2__abc_44228_n10452_1), .B(u2__abc_44228_n10450), .Y(u2__abc_44228_n10453) );
  AND2X2 AND2X2_4204 ( .A(u2__abc_44228_n10453), .B(u2__abc_44228_n7547_bF_buf2), .Y(u2__abc_44228_n10454) );
  AND2X2 AND2X2_4205 ( .A(u2__abc_44228_n7548_1_bF_buf3), .B(u2_remHi_168_), .Y(u2__abc_44228_n10455) );
  AND2X2 AND2X2_4206 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n4915), .Y(u2__abc_44228_n10458_1) );
  AND2X2 AND2X2_4207 ( .A(u2__abc_44228_n10459_1), .B(u2__abc_44228_n2972_bF_buf43), .Y(u2__abc_44228_n10460) );
  AND2X2 AND2X2_4208 ( .A(u2__abc_44228_n10457), .B(u2__abc_44228_n10460), .Y(u2__abc_44228_n10461) );
  AND2X2 AND2X2_4209 ( .A(u2__abc_44228_n10462), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_remHi_170__FF_INPUT) );
  AND2X2 AND2X2_421 ( .A(u1__abc_43968_n187), .B(u1__abc_43968_n194), .Y(u1__abc_43968_n195_1) );
  AND2X2 AND2X2_4210 ( .A(u2__abc_44228_n3062_bF_buf14), .B(u2_remHi_171_), .Y(u2__abc_44228_n10464) );
  AND2X2 AND2X2_4211 ( .A(u2__abc_44228_n10469), .B(u2__abc_44228_n7547_bF_buf1), .Y(u2__abc_44228_n10470) );
  AND2X2 AND2X2_4212 ( .A(u2__abc_44228_n10470), .B(u2__abc_44228_n10468), .Y(u2__abc_44228_n10471) );
  AND2X2 AND2X2_4213 ( .A(u2__abc_44228_n7548_1_bF_buf2), .B(u2_remHi_169_), .Y(u2__abc_44228_n10472_1) );
  AND2X2 AND2X2_4214 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n4922), .Y(u2__abc_44228_n10475) );
  AND2X2 AND2X2_4215 ( .A(u2__abc_44228_n10476), .B(u2__abc_44228_n2972_bF_buf42), .Y(u2__abc_44228_n10477) );
  AND2X2 AND2X2_4216 ( .A(u2__abc_44228_n10474), .B(u2__abc_44228_n10477), .Y(u2__abc_44228_n10478) );
  AND2X2 AND2X2_4217 ( .A(u2__abc_44228_n10479_1), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_remHi_171__FF_INPUT) );
  AND2X2 AND2X2_4218 ( .A(u2__abc_44228_n3062_bF_buf13), .B(u2_remHi_172_), .Y(u2__abc_44228_n10481) );
  AND2X2 AND2X2_4219 ( .A(u2__abc_44228_n10414), .B(u2__abc_44228_n4956), .Y(u2__abc_44228_n10482) );
  AND2X2 AND2X2_422 ( .A(u1__abc_43968_n180_1), .B(u1__abc_43968_n195_1), .Y(u1__abc_43968_n196_1) );
  AND2X2 AND2X2_4220 ( .A(u2__abc_44228_n10483), .B(u2__abc_44228_n4918), .Y(u2__abc_44228_n10484) );
  AND2X2 AND2X2_4221 ( .A(u2__abc_44228_n10485), .B(u2__abc_44228_n10486_1), .Y(u2__abc_44228_n10487_1) );
  AND2X2 AND2X2_4222 ( .A(u2__abc_44228_n10488), .B(u2__abc_44228_n10489), .Y(u2__abc_44228_n10490) );
  AND2X2 AND2X2_4223 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n4908), .Y(u2__abc_44228_n10492) );
  AND2X2 AND2X2_4224 ( .A(u2__abc_44228_n10493_1), .B(u2__abc_44228_n2972_bF_buf41), .Y(u2__abc_44228_n10494_1) );
  AND2X2 AND2X2_4225 ( .A(u2__abc_44228_n10491), .B(u2__abc_44228_n10494_1), .Y(u2__abc_44228_n10495) );
  AND2X2 AND2X2_4226 ( .A(u2__abc_44228_n10496), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_remHi_172__FF_INPUT) );
  AND2X2 AND2X2_4227 ( .A(u2__abc_44228_n3062_bF_buf12), .B(u2_remHi_173_), .Y(u2__abc_44228_n10498) );
  AND2X2 AND2X2_4228 ( .A(u2__abc_44228_n10485), .B(u2__abc_44228_n5359), .Y(u2__abc_44228_n10499) );
  AND2X2 AND2X2_4229 ( .A(u2__abc_44228_n10503), .B(u2__abc_44228_n7547_bF_buf57), .Y(u2__abc_44228_n10504) );
  AND2X2 AND2X2_423 ( .A(u1__abc_43968_n197), .B(u1__abc_43968_n198), .Y(u1__abc_43968_n199) );
  AND2X2 AND2X2_4230 ( .A(u2__abc_44228_n10504), .B(u2__abc_44228_n10501_1), .Y(u2__abc_44228_n10505) );
  AND2X2 AND2X2_4231 ( .A(u2__abc_44228_n7548_1_bF_buf0), .B(u2_remHi_171_), .Y(u2__abc_44228_n10506) );
  AND2X2 AND2X2_4232 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n4902), .Y(u2__abc_44228_n10509) );
  AND2X2 AND2X2_4233 ( .A(u2__abc_44228_n10510), .B(u2__abc_44228_n2972_bF_buf40), .Y(u2__abc_44228_n10511) );
  AND2X2 AND2X2_4234 ( .A(u2__abc_44228_n10508_1), .B(u2__abc_44228_n10511), .Y(u2__abc_44228_n10512) );
  AND2X2 AND2X2_4235 ( .A(u2__abc_44228_n10513), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_remHi_173__FF_INPUT) );
  AND2X2 AND2X2_4236 ( .A(u2__abc_44228_n3062_bF_buf11), .B(u2_remHi_174_), .Y(u2__abc_44228_n10515_1) );
  AND2X2 AND2X2_4237 ( .A(u2__abc_44228_n10485), .B(u2__abc_44228_n5360), .Y(u2__abc_44228_n10516) );
  AND2X2 AND2X2_4238 ( .A(u2__abc_44228_n10518), .B(u2__abc_44228_n4911_1), .Y(u2__abc_44228_n10520) );
  AND2X2 AND2X2_4239 ( .A(u2__abc_44228_n10521_1), .B(u2__abc_44228_n10519), .Y(u2__abc_44228_n10522_1) );
  AND2X2 AND2X2_424 ( .A(u1__abc_43968_n200), .B(u1__abc_43968_n201), .Y(u1__abc_43968_n202_1) );
  AND2X2 AND2X2_4240 ( .A(u2__abc_44228_n10522_1), .B(u2__abc_44228_n7547_bF_buf56), .Y(u2__abc_44228_n10523) );
  AND2X2 AND2X2_4241 ( .A(u2__abc_44228_n7548_1_bF_buf57), .B(u2_remHi_172_), .Y(u2__abc_44228_n10524) );
  AND2X2 AND2X2_4242 ( .A(u2__abc_44228_n2983_bF_buf91), .B(u2__abc_44228_n4891), .Y(u2__abc_44228_n10527) );
  AND2X2 AND2X2_4243 ( .A(u2__abc_44228_n10528_1), .B(u2__abc_44228_n2972_bF_buf39), .Y(u2__abc_44228_n10529_1) );
  AND2X2 AND2X2_4244 ( .A(u2__abc_44228_n10526), .B(u2__abc_44228_n10529_1), .Y(u2__abc_44228_n10530) );
  AND2X2 AND2X2_4245 ( .A(u2__abc_44228_n10531), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_remHi_174__FF_INPUT) );
  AND2X2 AND2X2_4246 ( .A(u2__abc_44228_n3062_bF_buf10), .B(u2_remHi_175_), .Y(u2__abc_44228_n10533) );
  AND2X2 AND2X2_4247 ( .A(u2__abc_44228_n10538), .B(u2__abc_44228_n7547_bF_buf55), .Y(u2__abc_44228_n10539) );
  AND2X2 AND2X2_4248 ( .A(u2__abc_44228_n10539), .B(u2__abc_44228_n10537), .Y(u2__abc_44228_n10540) );
  AND2X2 AND2X2_4249 ( .A(u2__abc_44228_n7548_1_bF_buf56), .B(u2_remHi_173_), .Y(u2__abc_44228_n10541) );
  AND2X2 AND2X2_425 ( .A(u1__abc_43968_n199), .B(u1__abc_43968_n202_1), .Y(u1__abc_43968_n203_1) );
  AND2X2 AND2X2_4250 ( .A(u2__abc_44228_n2983_bF_buf89), .B(u2__abc_44228_n4885), .Y(u2__abc_44228_n10544) );
  AND2X2 AND2X2_4251 ( .A(u2__abc_44228_n10545), .B(u2__abc_44228_n2972_bF_buf38), .Y(u2__abc_44228_n10546) );
  AND2X2 AND2X2_4252 ( .A(u2__abc_44228_n10543_1), .B(u2__abc_44228_n10546), .Y(u2__abc_44228_n10547) );
  AND2X2 AND2X2_4253 ( .A(u2__abc_44228_n10548), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_remHi_175__FF_INPUT) );
  AND2X2 AND2X2_4254 ( .A(u2__abc_44228_n3062_bF_buf9), .B(u2_remHi_176_), .Y(u2__abc_44228_n10550_1) );
  AND2X2 AND2X2_4255 ( .A(u2__abc_44228_n10278), .B(u2__abc_44228_n5017), .Y(u2__abc_44228_n10551) );
  AND2X2 AND2X2_4256 ( .A(u2__abc_44228_n10552), .B(u2__abc_44228_n4894), .Y(u2__abc_44228_n10553) );
  AND2X2 AND2X2_4257 ( .A(u2__abc_44228_n10554), .B(u2__abc_44228_n10555), .Y(u2__abc_44228_n10556_1) );
  AND2X2 AND2X2_4258 ( .A(u2__abc_44228_n10557_1), .B(u2__abc_44228_n10558), .Y(u2__abc_44228_n10559) );
  AND2X2 AND2X2_4259 ( .A(u2__abc_44228_n2983_bF_buf87), .B(u2__abc_44228_n4877), .Y(u2__abc_44228_n10561) );
  AND2X2 AND2X2_426 ( .A(u1__abc_43968_n204), .B(u1__abc_43968_n205_1), .Y(u1__abc_43968_n206_1) );
  AND2X2 AND2X2_4260 ( .A(u2__abc_44228_n10562), .B(u2__abc_44228_n2972_bF_buf37), .Y(u2__abc_44228_n10563_1) );
  AND2X2 AND2X2_4261 ( .A(u2__abc_44228_n10560), .B(u2__abc_44228_n10563_1), .Y(u2__abc_44228_n10564_1) );
  AND2X2 AND2X2_4262 ( .A(u2__abc_44228_n10565), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_remHi_176__FF_INPUT) );
  AND2X2 AND2X2_4263 ( .A(u2__abc_44228_n3062_bF_buf8), .B(u2_remHi_177_), .Y(u2__abc_44228_n10567) );
  AND2X2 AND2X2_4264 ( .A(u2__abc_44228_n10554), .B(u2__abc_44228_n5370), .Y(u2__abc_44228_n10568) );
  AND2X2 AND2X2_4265 ( .A(u2__abc_44228_n10570_1), .B(u2__abc_44228_n10572), .Y(u2__abc_44228_n10573) );
  AND2X2 AND2X2_4266 ( .A(u2__abc_44228_n10573), .B(u2__abc_44228_n7547_bF_buf53), .Y(u2__abc_44228_n10574) );
  AND2X2 AND2X2_4267 ( .A(u2__abc_44228_n7548_1_bF_buf54), .B(u2_remHi_175_), .Y(u2__abc_44228_n10575) );
  AND2X2 AND2X2_4268 ( .A(u2__abc_44228_n2983_bF_buf85), .B(u2__abc_44228_n4871), .Y(u2__abc_44228_n10578_1) );
  AND2X2 AND2X2_4269 ( .A(u2__abc_44228_n10579), .B(u2__abc_44228_n2972_bF_buf36), .Y(u2__abc_44228_n10580) );
  AND2X2 AND2X2_427 ( .A(u1__abc_43968_n207), .B(u1__abc_43968_n208), .Y(u1__abc_43968_n209_1) );
  AND2X2 AND2X2_4270 ( .A(u2__abc_44228_n10577_1), .B(u2__abc_44228_n10580), .Y(u2__abc_44228_n10581) );
  AND2X2 AND2X2_4271 ( .A(u2__abc_44228_n10582), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_remHi_177__FF_INPUT) );
  AND2X2 AND2X2_4272 ( .A(u2__abc_44228_n3062_bF_buf7), .B(u2_remHi_178_), .Y(u2__abc_44228_n10584_1) );
  AND2X2 AND2X2_4273 ( .A(u2__abc_44228_n10552), .B(u2__abc_44228_n4895), .Y(u2__abc_44228_n10585_1) );
  AND2X2 AND2X2_4274 ( .A(u2__abc_44228_n10586), .B(u2__abc_44228_n4880), .Y(u2__abc_44228_n10588) );
  AND2X2 AND2X2_4275 ( .A(u2__abc_44228_n10589), .B(u2__abc_44228_n10587), .Y(u2__abc_44228_n10590) );
  AND2X2 AND2X2_4276 ( .A(u2__abc_44228_n10591_1), .B(u2__abc_44228_n10592_1), .Y(u2__abc_44228_n10593) );
  AND2X2 AND2X2_4277 ( .A(u2__abc_44228_n2983_bF_buf83), .B(u2__abc_44228_n4862), .Y(u2__abc_44228_n10595) );
  AND2X2 AND2X2_4278 ( .A(u2__abc_44228_n10596), .B(u2__abc_44228_n2972_bF_buf35), .Y(u2__abc_44228_n10597) );
  AND2X2 AND2X2_4279 ( .A(u2__abc_44228_n10594), .B(u2__abc_44228_n10597), .Y(u2__abc_44228_n10598_1) );
  AND2X2 AND2X2_428 ( .A(u1__abc_43968_n206_1), .B(u1__abc_43968_n209_1), .Y(u1__abc_43968_n210_1) );
  AND2X2 AND2X2_4280 ( .A(u2__abc_44228_n10599_1), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_remHi_178__FF_INPUT) );
  AND2X2 AND2X2_4281 ( .A(u2__abc_44228_n3062_bF_buf6), .B(u2_remHi_179_), .Y(u2__abc_44228_n10601) );
  AND2X2 AND2X2_4282 ( .A(u2__abc_44228_n10606_1), .B(u2__abc_44228_n7547_bF_buf51), .Y(u2__abc_44228_n10607) );
  AND2X2 AND2X2_4283 ( .A(u2__abc_44228_n10607), .B(u2__abc_44228_n10605_1), .Y(u2__abc_44228_n10608) );
  AND2X2 AND2X2_4284 ( .A(u2__abc_44228_n7548_1_bF_buf52), .B(u2_remHi_177_), .Y(u2__abc_44228_n10609) );
  AND2X2 AND2X2_4285 ( .A(u2__abc_44228_n2983_bF_buf81), .B(u2__abc_44228_n4856), .Y(u2__abc_44228_n10612_1) );
  AND2X2 AND2X2_4286 ( .A(u2__abc_44228_n10613_1), .B(u2__abc_44228_n2972_bF_buf34), .Y(u2__abc_44228_n10614) );
  AND2X2 AND2X2_4287 ( .A(u2__abc_44228_n10611), .B(u2__abc_44228_n10614), .Y(u2__abc_44228_n10615) );
  AND2X2 AND2X2_4288 ( .A(u2__abc_44228_n10616), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_remHi_179__FF_INPUT) );
  AND2X2 AND2X2_4289 ( .A(u2__abc_44228_n3062_bF_buf5), .B(u2_remHi_180_), .Y(u2__abc_44228_n10618) );
  AND2X2 AND2X2_429 ( .A(u1__abc_43968_n203_1), .B(u1__abc_43968_n210_1), .Y(u1__abc_43968_n211) );
  AND2X2 AND2X2_4290 ( .A(u2__abc_44228_n10552), .B(u2__abc_44228_n4896), .Y(u2__abc_44228_n10619_1) );
  AND2X2 AND2X2_4291 ( .A(u2__abc_44228_n10620_1), .B(u2__abc_44228_n4865), .Y(u2__abc_44228_n10621) );
  AND2X2 AND2X2_4292 ( .A(u2__abc_44228_n10622), .B(u2__abc_44228_n10623), .Y(u2__abc_44228_n10624) );
  AND2X2 AND2X2_4293 ( .A(u2__abc_44228_n10625), .B(u2__abc_44228_n10626_1), .Y(u2__abc_44228_n10627_1) );
  AND2X2 AND2X2_4294 ( .A(u2__abc_44228_n2983_bF_buf79), .B(u2__abc_44228_n4848), .Y(u2__abc_44228_n10629) );
  AND2X2 AND2X2_4295 ( .A(u2__abc_44228_n10630), .B(u2__abc_44228_n2972_bF_buf33), .Y(u2__abc_44228_n10631) );
  AND2X2 AND2X2_4296 ( .A(u2__abc_44228_n10628), .B(u2__abc_44228_n10631), .Y(u2__abc_44228_n10632) );
  AND2X2 AND2X2_4297 ( .A(u2__abc_44228_n10633_1), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_remHi_180__FF_INPUT) );
  AND2X2 AND2X2_4298 ( .A(u2__abc_44228_n3062_bF_buf4), .B(u2_remHi_181_), .Y(u2__abc_44228_n10635) );
  AND2X2 AND2X2_4299 ( .A(u2__abc_44228_n10622), .B(u2__abc_44228_n5379), .Y(u2__abc_44228_n10637) );
  AND2X2 AND2X2_43 ( .A(_abc_64468_n753_bF_buf13), .B(sqrto_42_), .Y(_auto_iopadmap_cc_313_execute_65414_78_) );
  AND2X2 AND2X2_430 ( .A(u1__abc_43968_n212_1), .B(u1__abc_43968_n213_1), .Y(u1__abc_43968_n214) );
  AND2X2 AND2X2_4300 ( .A(u2__abc_44228_n10640_1), .B(u2__abc_44228_n10638), .Y(u2__abc_44228_n10641_1) );
  AND2X2 AND2X2_4301 ( .A(u2__abc_44228_n10641_1), .B(u2__abc_44228_n7547_bF_buf49), .Y(u2__abc_44228_n10642) );
  AND2X2 AND2X2_4302 ( .A(u2__abc_44228_n7548_1_bF_buf50), .B(u2_remHi_179_), .Y(u2__abc_44228_n10643) );
  AND2X2 AND2X2_4303 ( .A(u2__abc_44228_n2983_bF_buf77), .B(u2__abc_44228_n4842), .Y(u2__abc_44228_n10646) );
  AND2X2 AND2X2_4304 ( .A(u2__abc_44228_n10647_1), .B(u2__abc_44228_n2972_bF_buf32), .Y(u2__abc_44228_n10648_1) );
  AND2X2 AND2X2_4305 ( .A(u2__abc_44228_n10645), .B(u2__abc_44228_n10648_1), .Y(u2__abc_44228_n10649) );
  AND2X2 AND2X2_4306 ( .A(u2__abc_44228_n10650), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_remHi_181__FF_INPUT) );
  AND2X2 AND2X2_4307 ( .A(u2__abc_44228_n3062_bF_buf3), .B(u2_remHi_182_), .Y(u2__abc_44228_n10652) );
  AND2X2 AND2X2_4308 ( .A(u2__abc_44228_n10620_1), .B(u2__abc_44228_n4866), .Y(u2__abc_44228_n10653) );
  AND2X2 AND2X2_4309 ( .A(u2__abc_44228_n10654_1), .B(u2__abc_44228_n4851), .Y(u2__abc_44228_n10656) );
  AND2X2 AND2X2_431 ( .A(u1__abc_43968_n215), .B(u1__abc_43968_n216), .Y(u1__abc_43968_n217_1) );
  AND2X2 AND2X2_4310 ( .A(u2__abc_44228_n10657), .B(u2__abc_44228_n10655_1), .Y(u2__abc_44228_n10658) );
  AND2X2 AND2X2_4311 ( .A(u2__abc_44228_n10658), .B(u2__abc_44228_n7547_bF_buf48), .Y(u2__abc_44228_n10659) );
  AND2X2 AND2X2_4312 ( .A(u2__abc_44228_n7548_1_bF_buf49), .B(u2_remHi_180_), .Y(u2__abc_44228_n10660) );
  AND2X2 AND2X2_4313 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n4818_1), .Y(u2__abc_44228_n10663) );
  AND2X2 AND2X2_4314 ( .A(u2__abc_44228_n10664), .B(u2__abc_44228_n2972_bF_buf31), .Y(u2__abc_44228_n10665) );
  AND2X2 AND2X2_4315 ( .A(u2__abc_44228_n10662_1), .B(u2__abc_44228_n10665), .Y(u2__abc_44228_n10666) );
  AND2X2 AND2X2_4316 ( .A(u2__abc_44228_n10667), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_remHi_182__FF_INPUT) );
  AND2X2 AND2X2_4317 ( .A(u2__abc_44228_n3062_bF_buf2), .B(u2_remHi_183_), .Y(u2__abc_44228_n10669_1) );
  AND2X2 AND2X2_4318 ( .A(u2__abc_44228_n10674), .B(u2__abc_44228_n7547_bF_buf47), .Y(u2__abc_44228_n10675_1) );
  AND2X2 AND2X2_4319 ( .A(u2__abc_44228_n10675_1), .B(u2__abc_44228_n10673), .Y(u2__abc_44228_n10676_1) );
  AND2X2 AND2X2_432 ( .A(u1__abc_43968_n214), .B(u1__abc_43968_n217_1), .Y(u1__abc_43968_n218_1) );
  AND2X2 AND2X2_4320 ( .A(u2__abc_44228_n7548_1_bF_buf48), .B(u2_remHi_181_), .Y(u2__abc_44228_n10677) );
  AND2X2 AND2X2_4321 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n4812), .Y(u2__abc_44228_n10680) );
  AND2X2 AND2X2_4322 ( .A(u2__abc_44228_n10681), .B(u2__abc_44228_n2972_bF_buf30), .Y(u2__abc_44228_n10682_1) );
  AND2X2 AND2X2_4323 ( .A(u2__abc_44228_n10679), .B(u2__abc_44228_n10682_1), .Y(u2__abc_44228_n10683_1) );
  AND2X2 AND2X2_4324 ( .A(u2__abc_44228_n10684), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_remHi_183__FF_INPUT) );
  AND2X2 AND2X2_4325 ( .A(u2__abc_44228_n3062_bF_buf1), .B(u2_remHi_184_), .Y(u2__abc_44228_n10686) );
  AND2X2 AND2X2_4326 ( .A(u2__abc_44228_n10552), .B(u2__abc_44228_n4897), .Y(u2__abc_44228_n10687) );
  AND2X2 AND2X2_4327 ( .A(u2__abc_44228_n10688), .B(u2__abc_44228_n4821), .Y(u2__abc_44228_n10690_1) );
  AND2X2 AND2X2_4328 ( .A(u2__abc_44228_n10691), .B(u2__abc_44228_n10689_1), .Y(u2__abc_44228_n10692) );
  AND2X2 AND2X2_4329 ( .A(u2__abc_44228_n10693), .B(u2__abc_44228_n10694), .Y(u2__abc_44228_n10695) );
  AND2X2 AND2X2_433 ( .A(u1__abc_43968_n219), .B(u1__abc_43968_n220_1), .Y(u1__abc_43968_n221_1) );
  AND2X2 AND2X2_4330 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n4832), .Y(u2__abc_44228_n10697_1) );
  AND2X2 AND2X2_4331 ( .A(u2__abc_44228_n10698), .B(u2__abc_44228_n2972_bF_buf29), .Y(u2__abc_44228_n10699) );
  AND2X2 AND2X2_4332 ( .A(u2__abc_44228_n10696_1), .B(u2__abc_44228_n10699), .Y(u2__abc_44228_n10700) );
  AND2X2 AND2X2_4333 ( .A(u2__abc_44228_n10701), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_remHi_184__FF_INPUT) );
  AND2X2 AND2X2_4334 ( .A(u2__abc_44228_n3062_bF_buf0), .B(u2_remHi_185_), .Y(u2__abc_44228_n10703_1) );
  AND2X2 AND2X2_4335 ( .A(u2__abc_44228_n10691), .B(u2__abc_44228_n5397), .Y(u2__abc_44228_n10705) );
  AND2X2 AND2X2_4336 ( .A(u2__abc_44228_n10708), .B(u2__abc_44228_n10706), .Y(u2__abc_44228_n10709) );
  AND2X2 AND2X2_4337 ( .A(u2__abc_44228_n10709), .B(u2__abc_44228_n7547_bF_buf45), .Y(u2__abc_44228_n10710_1) );
  AND2X2 AND2X2_4338 ( .A(u2__abc_44228_n7548_1_bF_buf46), .B(u2_remHi_183_), .Y(u2__abc_44228_n10711_1) );
  AND2X2 AND2X2_4339 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n4826), .Y(u2__abc_44228_n10714) );
  AND2X2 AND2X2_434 ( .A(u1__abc_43968_n222), .B(u1__abc_43968_n223), .Y(u1__abc_43968_n224_1) );
  AND2X2 AND2X2_4340 ( .A(u2__abc_44228_n10715), .B(u2__abc_44228_n2972_bF_buf28), .Y(u2__abc_44228_n10716) );
  AND2X2 AND2X2_4341 ( .A(u2__abc_44228_n10713), .B(u2__abc_44228_n10716), .Y(u2__abc_44228_n10717_1) );
  AND2X2 AND2X2_4342 ( .A(u2__abc_44228_n10718_1), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_remHi_185__FF_INPUT) );
  AND2X2 AND2X2_4343 ( .A(u2__abc_44228_n3062_bF_buf92), .B(u2_remHi_186_), .Y(u2__abc_44228_n10720) );
  AND2X2 AND2X2_4344 ( .A(u2__abc_44228_n10688), .B(u2__abc_44228_n4822), .Y(u2__abc_44228_n10721) );
  AND2X2 AND2X2_4345 ( .A(u2__abc_44228_n10722), .B(u2__abc_44228_n4835), .Y(u2__abc_44228_n10724_1) );
  AND2X2 AND2X2_4346 ( .A(u2__abc_44228_n10725_1), .B(u2__abc_44228_n10723), .Y(u2__abc_44228_n10726) );
  AND2X2 AND2X2_4347 ( .A(u2__abc_44228_n10726), .B(u2__abc_44228_n7547_bF_buf44), .Y(u2__abc_44228_n10727) );
  AND2X2 AND2X2_4348 ( .A(u2__abc_44228_n7548_1_bF_buf45), .B(u2_remHi_184_), .Y(u2__abc_44228_n10728) );
  AND2X2 AND2X2_4349 ( .A(u2__abc_44228_n2983_bF_buf69), .B(u2__abc_44228_n4803), .Y(u2__abc_44228_n10731_1) );
  AND2X2 AND2X2_435 ( .A(u1__abc_43968_n221_1), .B(u1__abc_43968_n224_1), .Y(u1__abc_43968_n225_1) );
  AND2X2 AND2X2_4350 ( .A(u2__abc_44228_n10732_1), .B(u2__abc_44228_n2972_bF_buf27), .Y(u2__abc_44228_n10733) );
  AND2X2 AND2X2_4351 ( .A(u2__abc_44228_n10730), .B(u2__abc_44228_n10733), .Y(u2__abc_44228_n10734) );
  AND2X2 AND2X2_4352 ( .A(u2__abc_44228_n10735), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_remHi_186__FF_INPUT) );
  AND2X2 AND2X2_4353 ( .A(u2__abc_44228_n3062_bF_buf91), .B(u2_remHi_187_), .Y(u2__abc_44228_n10737) );
  AND2X2 AND2X2_4354 ( .A(u2__abc_44228_n10725_1), .B(u2__abc_44228_n5402), .Y(u2__abc_44228_n10739_1) );
  AND2X2 AND2X2_4355 ( .A(u2__abc_44228_n10742), .B(u2__abc_44228_n10740), .Y(u2__abc_44228_n10743) );
  AND2X2 AND2X2_4356 ( .A(u2__abc_44228_n10743), .B(u2__abc_44228_n7547_bF_buf43), .Y(u2__abc_44228_n10744) );
  AND2X2 AND2X2_4357 ( .A(u2__abc_44228_n7548_1_bF_buf44), .B(u2_remHi_185_), .Y(u2__abc_44228_n10745_1) );
  AND2X2 AND2X2_4358 ( .A(u2__abc_44228_n2983_bF_buf67), .B(u2__abc_44228_n4797), .Y(u2__abc_44228_n10748) );
  AND2X2 AND2X2_4359 ( .A(u2__abc_44228_n10749), .B(u2__abc_44228_n2972_bF_buf26), .Y(u2__abc_44228_n10750) );
  AND2X2 AND2X2_436 ( .A(u1__abc_43968_n218_1), .B(u1__abc_43968_n225_1), .Y(u1__abc_43968_n226) );
  AND2X2 AND2X2_4360 ( .A(u2__abc_44228_n10747), .B(u2__abc_44228_n10750), .Y(u2__abc_44228_n10751) );
  AND2X2 AND2X2_4361 ( .A(u2__abc_44228_n10752_1), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_remHi_187__FF_INPUT) );
  AND2X2 AND2X2_4362 ( .A(u2__abc_44228_n3062_bF_buf90), .B(u2_remHi_188_), .Y(u2__abc_44228_n10754) );
  AND2X2 AND2X2_4363 ( .A(u2__abc_44228_n10725_1), .B(u2__abc_44228_n5403), .Y(u2__abc_44228_n10755) );
  AND2X2 AND2X2_4364 ( .A(u2__abc_44228_n10757), .B(u2__abc_44228_n4806), .Y(u2__abc_44228_n10758) );
  AND2X2 AND2X2_4365 ( .A(u2__abc_44228_n10759_1), .B(u2__abc_44228_n10760_1), .Y(u2__abc_44228_n10761) );
  AND2X2 AND2X2_4366 ( .A(u2__abc_44228_n10761), .B(u2__abc_44228_n7547_bF_buf42), .Y(u2__abc_44228_n10762) );
  AND2X2 AND2X2_4367 ( .A(u2__abc_44228_n7548_1_bF_buf43), .B(u2_remHi_186_), .Y(u2__abc_44228_n10763) );
  AND2X2 AND2X2_4368 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n4789), .Y(u2__abc_44228_n10766_1) );
  AND2X2 AND2X2_4369 ( .A(u2__abc_44228_n10767_1), .B(u2__abc_44228_n2972_bF_buf25), .Y(u2__abc_44228_n10768) );
  AND2X2 AND2X2_437 ( .A(u1__abc_43968_n211), .B(u1__abc_43968_n226), .Y(u1__abc_43968_n227_1) );
  AND2X2 AND2X2_4370 ( .A(u2__abc_44228_n10765), .B(u2__abc_44228_n10768), .Y(u2__abc_44228_n10769) );
  AND2X2 AND2X2_4371 ( .A(u2__abc_44228_n10770), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_remHi_188__FF_INPUT) );
  AND2X2 AND2X2_4372 ( .A(u2__abc_44228_n3062_bF_buf89), .B(u2_remHi_189_), .Y(u2__abc_44228_n10772) );
  AND2X2 AND2X2_4373 ( .A(u2__abc_44228_n10759_1), .B(u2__abc_44228_n5389), .Y(u2__abc_44228_n10774_1) );
  AND2X2 AND2X2_4374 ( .A(u2__abc_44228_n10777), .B(u2__abc_44228_n10775), .Y(u2__abc_44228_n10778) );
  AND2X2 AND2X2_4375 ( .A(u2__abc_44228_n10778), .B(u2__abc_44228_n7547_bF_buf41), .Y(u2__abc_44228_n10779) );
  AND2X2 AND2X2_4376 ( .A(u2__abc_44228_n7548_1_bF_buf42), .B(u2_remHi_187_), .Y(u2__abc_44228_n10780_1) );
  AND2X2 AND2X2_4377 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n4783), .Y(u2__abc_44228_n10783) );
  AND2X2 AND2X2_4378 ( .A(u2__abc_44228_n10784), .B(u2__abc_44228_n2972_bF_buf24), .Y(u2__abc_44228_n10785) );
  AND2X2 AND2X2_4379 ( .A(u2__abc_44228_n10782), .B(u2__abc_44228_n10785), .Y(u2__abc_44228_n10786) );
  AND2X2 AND2X2_438 ( .A(u1__abc_43968_n228_1), .B(u1__abc_43968_n229), .Y(u1__abc_43968_n230) );
  AND2X2 AND2X2_4380 ( .A(u2__abc_44228_n10787_1), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_remHi_189__FF_INPUT) );
  AND2X2 AND2X2_4381 ( .A(u2__abc_44228_n3062_bF_buf88), .B(u2_remHi_190_), .Y(u2__abc_44228_n10789) );
  AND2X2 AND2X2_4382 ( .A(u2__abc_44228_n10757), .B(u2__abc_44228_n4807), .Y(u2__abc_44228_n10790) );
  AND2X2 AND2X2_4383 ( .A(u2__abc_44228_n10791), .B(u2__abc_44228_n4792), .Y(u2__abc_44228_n10793) );
  AND2X2 AND2X2_4384 ( .A(u2__abc_44228_n10794_1), .B(u2__abc_44228_n10792), .Y(u2__abc_44228_n10795_1) );
  AND2X2 AND2X2_4385 ( .A(u2__abc_44228_n10795_1), .B(u2__abc_44228_n7547_bF_buf40), .Y(u2__abc_44228_n10796) );
  AND2X2 AND2X2_4386 ( .A(u2__abc_44228_n7548_1_bF_buf41), .B(u2_remHi_188_), .Y(u2__abc_44228_n10797) );
  AND2X2 AND2X2_4387 ( .A(u2__abc_44228_n2983_bF_buf63), .B(u2__abc_44228_n4763), .Y(u2__abc_44228_n10800) );
  AND2X2 AND2X2_4388 ( .A(u2__abc_44228_n10801_1), .B(u2__abc_44228_n2972_bF_buf23), .Y(u2__abc_44228_n10802_1) );
  AND2X2 AND2X2_4389 ( .A(u2__abc_44228_n10799), .B(u2__abc_44228_n10802_1), .Y(u2__abc_44228_n10803) );
  AND2X2 AND2X2_439 ( .A(u1__abc_43968_n231), .B(u1__abc_43968_n232), .Y(u1__abc_43968_n233_1) );
  AND2X2 AND2X2_4390 ( .A(u2__abc_44228_n10804), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_remHi_190__FF_INPUT) );
  AND2X2 AND2X2_4391 ( .A(u2__abc_44228_n3062_bF_buf87), .B(u2_remHi_191_), .Y(u2__abc_44228_n10806) );
  AND2X2 AND2X2_4392 ( .A(u2__abc_44228_n10811), .B(u2__abc_44228_n7547_bF_buf39), .Y(u2__abc_44228_n10812) );
  AND2X2 AND2X2_4393 ( .A(u2__abc_44228_n10812), .B(u2__abc_44228_n10810), .Y(u2__abc_44228_n10813) );
  AND2X2 AND2X2_4394 ( .A(u2__abc_44228_n7548_1_bF_buf40), .B(u2_remHi_189_), .Y(u2__abc_44228_n10814) );
  AND2X2 AND2X2_4395 ( .A(u2__abc_44228_n2983_bF_buf61), .B(u2__abc_44228_n4770_1), .Y(u2__abc_44228_n10817) );
  AND2X2 AND2X2_4396 ( .A(u2__abc_44228_n10818), .B(u2__abc_44228_n2972_bF_buf22), .Y(u2__abc_44228_n10819) );
  AND2X2 AND2X2_4397 ( .A(u2__abc_44228_n10816_1), .B(u2__abc_44228_n10819), .Y(u2__abc_44228_n10820) );
  AND2X2 AND2X2_4398 ( .A(u2__abc_44228_n10821), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_remHi_191__FF_INPUT) );
  AND2X2 AND2X2_4399 ( .A(u2__abc_44228_n3062_bF_buf86), .B(u2_remHi_192_), .Y(u2__abc_44228_n10823_1) );
  AND2X2 AND2X2_44 ( .A(_abc_64468_n753_bF_buf12), .B(sqrto_43_), .Y(_auto_iopadmap_cc_313_execute_65414_79_) );
  AND2X2 AND2X2_440 ( .A(u1__abc_43968_n230), .B(u1__abc_43968_n233_1), .Y(u1__abc_43968_n234_1) );
  AND2X2 AND2X2_4400 ( .A(u2__abc_44228_n7548_1_bF_buf39), .B(u2_remHi_190_), .Y(u2__abc_44228_n10824) );
  AND2X2 AND2X2_4401 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5255), .Y(u2__abc_44228_n10825) );
  AND2X2 AND2X2_4402 ( .A(u2__abc_44228_n10826), .B(u2__abc_44228_n4766), .Y(u2__abc_44228_n10827) );
  AND2X2 AND2X2_4403 ( .A(u2__abc_44228_n10828), .B(u2__abc_44228_n10829_1), .Y(u2__abc_44228_n10830_1) );
  AND2X2 AND2X2_4404 ( .A(u2__abc_44228_n7547_bF_buf38), .B(u2__abc_44228_n10830_1), .Y(u2__abc_44228_n10831) );
  AND2X2 AND2X2_4405 ( .A(u2__abc_44228_n2983_bF_buf59), .B(u2__abc_44228_n4756), .Y(u2__abc_44228_n10834) );
  AND2X2 AND2X2_4406 ( .A(u2__abc_44228_n10835), .B(u2__abc_44228_n2972_bF_buf21), .Y(u2__abc_44228_n10836_1) );
  AND2X2 AND2X2_4407 ( .A(u2__abc_44228_n10833), .B(u2__abc_44228_n10836_1), .Y(u2__abc_44228_n10837_1) );
  AND2X2 AND2X2_4408 ( .A(u2__abc_44228_n10838), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_remHi_192__FF_INPUT) );
  AND2X2 AND2X2_4409 ( .A(u2__abc_44228_n3062_bF_buf85), .B(u2_remHi_193_), .Y(u2__abc_44228_n10840) );
  AND2X2 AND2X2_441 ( .A(u1__abc_43968_n235), .B(u1__abc_43968_n236_1), .Y(u1__abc_43968_n237_1) );
  AND2X2 AND2X2_4410 ( .A(u2__abc_44228_n10844_1), .B(u2__abc_44228_n10845), .Y(u2__abc_44228_n10846) );
  AND2X2 AND2X2_4411 ( .A(u2__abc_44228_n7547_bF_buf37), .B(u2__abc_44228_n10846), .Y(u2__abc_44228_n10847) );
  AND2X2 AND2X2_4412 ( .A(u2__abc_44228_n7548_1_bF_buf38), .B(u2_remHi_191_), .Y(u2__abc_44228_n10848) );
  AND2X2 AND2X2_4413 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n4750_1), .Y(u2__abc_44228_n10851_1) );
  AND2X2 AND2X2_4414 ( .A(u2__abc_44228_n10852), .B(u2__abc_44228_n2972_bF_buf20), .Y(u2__abc_44228_n10853) );
  AND2X2 AND2X2_4415 ( .A(u2__abc_44228_n10850_1), .B(u2__abc_44228_n10853), .Y(u2__abc_44228_n10854) );
  AND2X2 AND2X2_4416 ( .A(u2__abc_44228_n10855), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_remHi_193__FF_INPUT) );
  AND2X2 AND2X2_4417 ( .A(u2__abc_44228_n3062_bF_buf84), .B(u2_remHi_194_), .Y(u2__abc_44228_n10857_1) );
  AND2X2 AND2X2_4418 ( .A(u2__abc_44228_n10826), .B(u2__abc_44228_n4774), .Y(u2__abc_44228_n10858_1) );
  AND2X2 AND2X2_4419 ( .A(u2__abc_44228_n10859), .B(u2__abc_44228_n4759), .Y(u2__abc_44228_n10861) );
  AND2X2 AND2X2_442 ( .A(u1__abc_43968_n238), .B(u1__abc_43968_n239), .Y(u1__abc_43968_n240_1) );
  AND2X2 AND2X2_4420 ( .A(u2__abc_44228_n10862), .B(u2__abc_44228_n10860), .Y(u2__abc_44228_n10863) );
  AND2X2 AND2X2_4421 ( .A(u2__abc_44228_n10864_1), .B(u2__abc_44228_n10865_1), .Y(u2__abc_44228_n10866) );
  AND2X2 AND2X2_4422 ( .A(u2__abc_44228_n2983_bF_buf56), .B(u2__abc_44228_n4741_1), .Y(u2__abc_44228_n10868) );
  AND2X2 AND2X2_4423 ( .A(u2__abc_44228_n10869), .B(u2__abc_44228_n2972_bF_buf19), .Y(u2__abc_44228_n10870) );
  AND2X2 AND2X2_4424 ( .A(u2__abc_44228_n10867), .B(u2__abc_44228_n10870), .Y(u2__abc_44228_n10871_1) );
  AND2X2 AND2X2_4425 ( .A(u2__abc_44228_n10872_1), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_remHi_194__FF_INPUT) );
  AND2X2 AND2X2_4426 ( .A(u2__abc_44228_n3062_bF_buf83), .B(u2_remHi_195_), .Y(u2__abc_44228_n10874) );
  AND2X2 AND2X2_4427 ( .A(u2__abc_44228_n10876), .B(u2__abc_44228_n4753), .Y(u2__abc_44228_n10877) );
  AND2X2 AND2X2_4428 ( .A(u2__abc_44228_n10875), .B(u2__abc_44228_n10878_1), .Y(u2__abc_44228_n10879_1) );
  AND2X2 AND2X2_4429 ( .A(u2__abc_44228_n10880), .B(u2__abc_44228_n7547_bF_buf35), .Y(u2__abc_44228_n10881) );
  AND2X2 AND2X2_443 ( .A(u1__abc_43968_n237_1), .B(u1__abc_43968_n240_1), .Y(u1__abc_43968_n241_1) );
  AND2X2 AND2X2_4430 ( .A(u2__abc_44228_n7548_1_bF_buf36), .B(u2_remHi_193_), .Y(u2__abc_44228_n10882) );
  AND2X2 AND2X2_4431 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n4735), .Y(u2__abc_44228_n10885_1) );
  AND2X2 AND2X2_4432 ( .A(u2__abc_44228_n10886_1), .B(u2__abc_44228_n2972_bF_buf18), .Y(u2__abc_44228_n10887) );
  AND2X2 AND2X2_4433 ( .A(u2__abc_44228_n10884), .B(u2__abc_44228_n10887), .Y(u2__abc_44228_n10888) );
  AND2X2 AND2X2_4434 ( .A(u2__abc_44228_n10889), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_remHi_195__FF_INPUT) );
  AND2X2 AND2X2_4435 ( .A(u2__abc_44228_n3062_bF_buf82), .B(u2_remHi_196_), .Y(u2__abc_44228_n10891) );
  AND2X2 AND2X2_4436 ( .A(u2__abc_44228_n10826), .B(u2__abc_44228_n4775), .Y(u2__abc_44228_n10892_1) );
  AND2X2 AND2X2_4437 ( .A(u2__abc_44228_n10893_1), .B(u2__abc_44228_n4744), .Y(u2__abc_44228_n10894) );
  AND2X2 AND2X2_4438 ( .A(u2__abc_44228_n10895), .B(u2__abc_44228_n10896), .Y(u2__abc_44228_n10897) );
  AND2X2 AND2X2_4439 ( .A(u2__abc_44228_n10898), .B(u2__abc_44228_n10899_1), .Y(u2__abc_44228_n10900_1) );
  AND2X2 AND2X2_444 ( .A(u1__abc_43968_n234_1), .B(u1__abc_43968_n241_1), .Y(u1__abc_43968_n242) );
  AND2X2 AND2X2_4440 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n4727), .Y(u2__abc_44228_n10902) );
  AND2X2 AND2X2_4441 ( .A(u2__abc_44228_n10903), .B(u2__abc_44228_n2972_bF_buf17), .Y(u2__abc_44228_n10904) );
  AND2X2 AND2X2_4442 ( .A(u2__abc_44228_n10901), .B(u2__abc_44228_n10904), .Y(u2__abc_44228_n10905) );
  AND2X2 AND2X2_4443 ( .A(u2__abc_44228_n10906_1), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_remHi_196__FF_INPUT) );
  AND2X2 AND2X2_4444 ( .A(u2__abc_44228_n3062_bF_buf81), .B(u2_remHi_197_), .Y(u2__abc_44228_n10908) );
  AND2X2 AND2X2_4445 ( .A(u2__abc_44228_n10895), .B(u2__abc_44228_n5420), .Y(u2__abc_44228_n10910) );
  AND2X2 AND2X2_4446 ( .A(u2__abc_44228_n10913_1), .B(u2__abc_44228_n10911), .Y(u2__abc_44228_n10914_1) );
  AND2X2 AND2X2_4447 ( .A(u2__abc_44228_n10914_1), .B(u2__abc_44228_n7547_bF_buf33), .Y(u2__abc_44228_n10915) );
  AND2X2 AND2X2_4448 ( .A(u2__abc_44228_n7548_1_bF_buf34), .B(u2_remHi_195_), .Y(u2__abc_44228_n10916) );
  AND2X2 AND2X2_4449 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2__abc_44228_n4721), .Y(u2__abc_44228_n10919) );
  AND2X2 AND2X2_445 ( .A(u1__abc_43968_n243_1), .B(u1__abc_43968_n244_1), .Y(u1__abc_43968_n245) );
  AND2X2 AND2X2_4450 ( .A(u2__abc_44228_n10920_1), .B(u2__abc_44228_n2972_bF_buf16), .Y(u2__abc_44228_n10921_1) );
  AND2X2 AND2X2_4451 ( .A(u2__abc_44228_n10918), .B(u2__abc_44228_n10921_1), .Y(u2__abc_44228_n10922) );
  AND2X2 AND2X2_4452 ( .A(u2__abc_44228_n10923), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_remHi_197__FF_INPUT) );
  AND2X2 AND2X2_4453 ( .A(u2__abc_44228_n3062_bF_buf80), .B(u2_remHi_198_), .Y(u2__abc_44228_n10925) );
  AND2X2 AND2X2_4454 ( .A(u2__abc_44228_n10893_1), .B(u2__abc_44228_n4745), .Y(u2__abc_44228_n10926) );
  AND2X2 AND2X2_4455 ( .A(u2__abc_44228_n10927_1), .B(u2__abc_44228_n4730), .Y(u2__abc_44228_n10929) );
  AND2X2 AND2X2_4456 ( .A(u2__abc_44228_n10930), .B(u2__abc_44228_n10928_1), .Y(u2__abc_44228_n10931) );
  AND2X2 AND2X2_4457 ( .A(u2__abc_44228_n10932), .B(u2__abc_44228_n10933), .Y(u2__abc_44228_n10934_1) );
  AND2X2 AND2X2_4458 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n4704_1), .Y(u2__abc_44228_n10936) );
  AND2X2 AND2X2_4459 ( .A(u2__abc_44228_n10937), .B(u2__abc_44228_n2972_bF_buf15), .Y(u2__abc_44228_n10938) );
  AND2X2 AND2X2_446 ( .A(u1__abc_43968_n246), .B(u1__abc_43968_n247), .Y(u1__abc_43968_n248_1) );
  AND2X2 AND2X2_4460 ( .A(u2__abc_44228_n10935_1), .B(u2__abc_44228_n10938), .Y(u2__abc_44228_n10939) );
  AND2X2 AND2X2_4461 ( .A(u2__abc_44228_n10940), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_remHi_198__FF_INPUT) );
  AND2X2 AND2X2_4462 ( .A(u2__abc_44228_n3062_bF_buf79), .B(u2_remHi_199_), .Y(u2__abc_44228_n10942_1) );
  AND2X2 AND2X2_4463 ( .A(u2__abc_44228_n10947), .B(u2__abc_44228_n7547_bF_buf31), .Y(u2__abc_44228_n10948_1) );
  AND2X2 AND2X2_4464 ( .A(u2__abc_44228_n10948_1), .B(u2__abc_44228_n10946), .Y(u2__abc_44228_n10949_1) );
  AND2X2 AND2X2_4465 ( .A(u2__abc_44228_n7548_1_bF_buf32), .B(u2_remHi_197_), .Y(u2__abc_44228_n10950) );
  AND2X2 AND2X2_4466 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n4711), .Y(u2__abc_44228_n10953) );
  AND2X2 AND2X2_4467 ( .A(u2__abc_44228_n10954), .B(u2__abc_44228_n2972_bF_buf14), .Y(u2__abc_44228_n10955_1) );
  AND2X2 AND2X2_4468 ( .A(u2__abc_44228_n10952), .B(u2__abc_44228_n10955_1), .Y(u2__abc_44228_n10956_1) );
  AND2X2 AND2X2_4469 ( .A(u2__abc_44228_n10957), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_remHi_199__FF_INPUT) );
  AND2X2 AND2X2_447 ( .A(u1__abc_43968_n245), .B(u1__abc_43968_n248_1), .Y(u1__abc_43968_n249_1) );
  AND2X2 AND2X2_4470 ( .A(u2__abc_44228_n3062_bF_buf78), .B(u2_remHi_200_), .Y(u2__abc_44228_n10959) );
  AND2X2 AND2X2_4471 ( .A(u2__abc_44228_n10826), .B(u2__abc_44228_n4776), .Y(u2__abc_44228_n10960) );
  AND2X2 AND2X2_4472 ( .A(u2__abc_44228_n10961), .B(u2__abc_44228_n4707), .Y(u2__abc_44228_n10963_1) );
  AND2X2 AND2X2_4473 ( .A(u2__abc_44228_n10964), .B(u2__abc_44228_n10962_1), .Y(u2__abc_44228_n10965) );
  AND2X2 AND2X2_4474 ( .A(u2__abc_44228_n10966), .B(u2__abc_44228_n10967), .Y(u2__abc_44228_n10968) );
  AND2X2 AND2X2_4475 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n4697), .Y(u2__abc_44228_n10970_1) );
  AND2X2 AND2X2_4476 ( .A(u2__abc_44228_n10971), .B(u2__abc_44228_n2972_bF_buf13), .Y(u2__abc_44228_n10972) );
  AND2X2 AND2X2_4477 ( .A(u2__abc_44228_n10969_1), .B(u2__abc_44228_n10972), .Y(u2__abc_44228_n10973) );
  AND2X2 AND2X2_4478 ( .A(u2__abc_44228_n10974), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_remHi_200__FF_INPUT) );
  AND2X2 AND2X2_4479 ( .A(u2__abc_44228_n3062_bF_buf77), .B(u2_remHi_201_), .Y(u2__abc_44228_n10976_1) );
  AND2X2 AND2X2_448 ( .A(u1__abc_43968_n250), .B(u1__abc_43968_n251_1), .Y(u1__abc_43968_n252_1) );
  AND2X2 AND2X2_4480 ( .A(u2__abc_44228_n10964), .B(u2__abc_44228_n5430), .Y(u2__abc_44228_n10977_1) );
  AND2X2 AND2X2_4481 ( .A(u2__abc_44228_n10979), .B(u2__abc_44228_n10981), .Y(u2__abc_44228_n10982) );
  AND2X2 AND2X2_4482 ( .A(u2__abc_44228_n10982), .B(u2__abc_44228_n7547_bF_buf29), .Y(u2__abc_44228_n10983_1) );
  AND2X2 AND2X2_4483 ( .A(u2__abc_44228_n7548_1_bF_buf30), .B(u2_remHi_199_), .Y(u2__abc_44228_n10984_1) );
  AND2X2 AND2X2_4484 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n4691), .Y(u2__abc_44228_n10987) );
  AND2X2 AND2X2_4485 ( .A(u2__abc_44228_n10988), .B(u2__abc_44228_n2972_bF_buf12), .Y(u2__abc_44228_n10989) );
  AND2X2 AND2X2_4486 ( .A(u2__abc_44228_n10986), .B(u2__abc_44228_n10989), .Y(u2__abc_44228_n10990_1) );
  AND2X2 AND2X2_4487 ( .A(u2__abc_44228_n10991_1), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_remHi_201__FF_INPUT) );
  AND2X2 AND2X2_4488 ( .A(u2__abc_44228_n3062_bF_buf76), .B(u2_remHi_202_), .Y(u2__abc_44228_n10993) );
  AND2X2 AND2X2_4489 ( .A(u2__abc_44228_n10964), .B(u2__abc_44228_n5431), .Y(u2__abc_44228_n10994) );
  AND2X2 AND2X2_449 ( .A(u1__abc_43968_n253), .B(u1__abc_43968_n254), .Y(u1__abc_43968_n255_1) );
  AND2X2 AND2X2_4490 ( .A(u2__abc_44228_n10996), .B(u2__abc_44228_n4700), .Y(u2__abc_44228_n10998_1) );
  AND2X2 AND2X2_4491 ( .A(u2__abc_44228_n10999), .B(u2__abc_44228_n10997_1), .Y(u2__abc_44228_n11000) );
  AND2X2 AND2X2_4492 ( .A(u2__abc_44228_n11000), .B(u2__abc_44228_n7547_bF_buf28), .Y(u2__abc_44228_n11001) );
  AND2X2 AND2X2_4493 ( .A(u2__abc_44228_n7548_1_bF_buf29), .B(u2_remHi_200_), .Y(u2__abc_44228_n11002) );
  AND2X2 AND2X2_4494 ( .A(u2__abc_44228_n2983_bF_buf41), .B(u2__abc_44228_n4682), .Y(u2__abc_44228_n11005_1) );
  AND2X2 AND2X2_4495 ( .A(u2__abc_44228_n11006), .B(u2__abc_44228_n2972_bF_buf11), .Y(u2__abc_44228_n11007) );
  AND2X2 AND2X2_4496 ( .A(u2__abc_44228_n11004_1), .B(u2__abc_44228_n11007), .Y(u2__abc_44228_n11008) );
  AND2X2 AND2X2_4497 ( .A(u2__abc_44228_n11009), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_remHi_202__FF_INPUT) );
  AND2X2 AND2X2_4498 ( .A(u2__abc_44228_n3062_bF_buf75), .B(u2_remHi_203_), .Y(u2__abc_44228_n11011_1) );
  AND2X2 AND2X2_4499 ( .A(u2__abc_44228_n11016), .B(u2__abc_44228_n7547_bF_buf27), .Y(u2__abc_44228_n11017) );
  AND2X2 AND2X2_45 ( .A(_abc_64468_n753_bF_buf11), .B(sqrto_44_), .Y(_auto_iopadmap_cc_313_execute_65414_80_) );
  AND2X2 AND2X2_450 ( .A(u1__abc_43968_n252_1), .B(u1__abc_43968_n255_1), .Y(u1__abc_43968_n256_1) );
  AND2X2 AND2X2_4500 ( .A(u2__abc_44228_n11017), .B(u2__abc_44228_n11015), .Y(u2__abc_44228_n11018_1) );
  AND2X2 AND2X2_4501 ( .A(u2__abc_44228_n7548_1_bF_buf28), .B(u2_remHi_201_), .Y(u2__abc_44228_n11019_1) );
  AND2X2 AND2X2_4502 ( .A(u2__abc_44228_n2983_bF_buf39), .B(u2__abc_44228_n4676), .Y(u2__abc_44228_n11022) );
  AND2X2 AND2X2_4503 ( .A(u2__abc_44228_n11023), .B(u2__abc_44228_n2972_bF_buf10), .Y(u2__abc_44228_n11024) );
  AND2X2 AND2X2_4504 ( .A(u2__abc_44228_n11021), .B(u2__abc_44228_n11024), .Y(u2__abc_44228_n11025_1) );
  AND2X2 AND2X2_4505 ( .A(u2__abc_44228_n11026_1), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_remHi_203__FF_INPUT) );
  AND2X2 AND2X2_4506 ( .A(u2__abc_44228_n3062_bF_buf74), .B(u2_remHi_204_), .Y(u2__abc_44228_n11028) );
  AND2X2 AND2X2_4507 ( .A(u2__abc_44228_n10961), .B(u2__abc_44228_n4716), .Y(u2__abc_44228_n11029) );
  AND2X2 AND2X2_4508 ( .A(u2__abc_44228_n11030), .B(u2__abc_44228_n4685_1), .Y(u2__abc_44228_n11031) );
  AND2X2 AND2X2_4509 ( .A(u2__abc_44228_n11032_1), .B(u2__abc_44228_n11033_1), .Y(u2__abc_44228_n11034) );
  AND2X2 AND2X2_451 ( .A(u1__abc_43968_n249_1), .B(u1__abc_43968_n256_1), .Y(u1__abc_43968_n257) );
  AND2X2 AND2X2_4510 ( .A(u2__abc_44228_n11035), .B(u2__abc_44228_n11036), .Y(u2__abc_44228_n11037) );
  AND2X2 AND2X2_4511 ( .A(u2__abc_44228_n2983_bF_buf37), .B(u2__abc_44228_n4668), .Y(u2__abc_44228_n11039_1) );
  AND2X2 AND2X2_4512 ( .A(u2__abc_44228_n11040_1), .B(u2__abc_44228_n2972_bF_buf9), .Y(u2__abc_44228_n11041) );
  AND2X2 AND2X2_4513 ( .A(u2__abc_44228_n11038), .B(u2__abc_44228_n11041), .Y(u2__abc_44228_n11042) );
  AND2X2 AND2X2_4514 ( .A(u2__abc_44228_n11043), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_remHi_204__FF_INPUT) );
  AND2X2 AND2X2_4515 ( .A(u2__abc_44228_n3062_bF_buf73), .B(u2_remHi_205_), .Y(u2__abc_44228_n11045) );
  AND2X2 AND2X2_4516 ( .A(u2__abc_44228_n11032_1), .B(u2__abc_44228_n5439), .Y(u2__abc_44228_n11047_1) );
  AND2X2 AND2X2_4517 ( .A(u2__abc_44228_n11050), .B(u2__abc_44228_n11048), .Y(u2__abc_44228_n11051) );
  AND2X2 AND2X2_4518 ( .A(u2__abc_44228_n11051), .B(u2__abc_44228_n7547_bF_buf25), .Y(u2__abc_44228_n11052) );
  AND2X2 AND2X2_4519 ( .A(u2__abc_44228_n7548_1_bF_buf26), .B(u2_remHi_203_), .Y(u2__abc_44228_n11053_1) );
  AND2X2 AND2X2_452 ( .A(u1__abc_43968_n242), .B(u1__abc_43968_n257), .Y(u1__abc_43968_n258_1) );
  AND2X2 AND2X2_4520 ( .A(u2__abc_44228_n2983_bF_buf35), .B(u2__abc_44228_n4662), .Y(u2__abc_44228_n11056) );
  AND2X2 AND2X2_4521 ( .A(u2__abc_44228_n11057), .B(u2__abc_44228_n2972_bF_buf8), .Y(u2__abc_44228_n11058) );
  AND2X2 AND2X2_4522 ( .A(u2__abc_44228_n11055), .B(u2__abc_44228_n11058), .Y(u2__abc_44228_n11059) );
  AND2X2 AND2X2_4523 ( .A(u2__abc_44228_n11060_1), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_remHi_205__FF_INPUT) );
  AND2X2 AND2X2_4524 ( .A(u2__abc_44228_n3062_bF_buf72), .B(u2_remHi_206_), .Y(u2__abc_44228_n11062) );
  AND2X2 AND2X2_4525 ( .A(u2__abc_44228_n11030), .B(u2__abc_44228_n4686), .Y(u2__abc_44228_n11063) );
  AND2X2 AND2X2_4526 ( .A(u2__abc_44228_n11064), .B(u2__abc_44228_n4671), .Y(u2__abc_44228_n11066) );
  AND2X2 AND2X2_4527 ( .A(u2__abc_44228_n11067_1), .B(u2__abc_44228_n11065), .Y(u2__abc_44228_n11068_1) );
  AND2X2 AND2X2_4528 ( .A(u2__abc_44228_n11068_1), .B(u2__abc_44228_n7547_bF_buf24), .Y(u2__abc_44228_n11069) );
  AND2X2 AND2X2_4529 ( .A(u2__abc_44228_n7548_1_bF_buf25), .B(u2_remHi_204_), .Y(u2__abc_44228_n11070) );
  AND2X2 AND2X2_453 ( .A(u1__abc_43968_n227_1), .B(u1__abc_43968_n258_1), .Y(u1__abc_43968_n259_1) );
  AND2X2 AND2X2_4530 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n4651), .Y(u2__abc_44228_n11073) );
  AND2X2 AND2X2_4531 ( .A(u2__abc_44228_n11074_1), .B(u2__abc_44228_n2972_bF_buf7), .Y(u2__abc_44228_n11075_1) );
  AND2X2 AND2X2_4532 ( .A(u2__abc_44228_n11072), .B(u2__abc_44228_n11075_1), .Y(u2__abc_44228_n11076) );
  AND2X2 AND2X2_4533 ( .A(u2__abc_44228_n11077), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_remHi_206__FF_INPUT) );
  AND2X2 AND2X2_4534 ( .A(u2__abc_44228_n3062_bF_buf71), .B(u2_remHi_207_), .Y(u2__abc_44228_n11079) );
  AND2X2 AND2X2_4535 ( .A(u2__abc_44228_n11084), .B(u2__abc_44228_n7547_bF_buf23), .Y(u2__abc_44228_n11085) );
  AND2X2 AND2X2_4536 ( .A(u2__abc_44228_n11085), .B(u2__abc_44228_n11083), .Y(u2__abc_44228_n11086) );
  AND2X2 AND2X2_4537 ( .A(u2__abc_44228_n7548_1_bF_buf24), .B(u2_remHi_205_), .Y(u2__abc_44228_n11087) );
  AND2X2 AND2X2_4538 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n4645), .Y(u2__abc_44228_n11090) );
  AND2X2 AND2X2_4539 ( .A(u2__abc_44228_n11091), .B(u2__abc_44228_n2972_bF_buf6), .Y(u2__abc_44228_n11092) );
  AND2X2 AND2X2_454 ( .A(u1__abc_43968_n259_1), .B(u1__abc_43968_n196_1), .Y(u1__abc_43968_n260) );
  AND2X2 AND2X2_4540 ( .A(u2__abc_44228_n11089_1), .B(u2__abc_44228_n11092), .Y(u2__abc_44228_n11093) );
  AND2X2 AND2X2_4541 ( .A(u2__abc_44228_n11094), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_remHi_207__FF_INPUT) );
  AND2X2 AND2X2_4542 ( .A(u2__abc_44228_n3062_bF_buf70), .B(u2_remHi_208_), .Y(u2__abc_44228_n11096_1) );
  AND2X2 AND2X2_4543 ( .A(u2__abc_44228_n10826), .B(u2__abc_44228_n4777), .Y(u2__abc_44228_n11097) );
  AND2X2 AND2X2_4544 ( .A(u2__abc_44228_n11098), .B(u2__abc_44228_n4654), .Y(u2__abc_44228_n11099) );
  AND2X2 AND2X2_4545 ( .A(u2__abc_44228_n11100), .B(u2__abc_44228_n11101), .Y(u2__abc_44228_n11102_1) );
  AND2X2 AND2X2_4546 ( .A(u2__abc_44228_n11103_1), .B(u2__abc_44228_n11104), .Y(u2__abc_44228_n11105) );
  AND2X2 AND2X2_4547 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n4637), .Y(u2__abc_44228_n11107) );
  AND2X2 AND2X2_4548 ( .A(u2__abc_44228_n11108), .B(u2__abc_44228_n2972_bF_buf5), .Y(u2__abc_44228_n11109_1) );
  AND2X2 AND2X2_4549 ( .A(u2__abc_44228_n11106), .B(u2__abc_44228_n11109_1), .Y(u2__abc_44228_n11110_1) );
  AND2X2 AND2X2_455 ( .A(u1__abc_43968_n261), .B(u1__abc_43968_n262), .Y(u1__abc_43968_n263) );
  AND2X2 AND2X2_4550 ( .A(u2__abc_44228_n11111), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_remHi_208__FF_INPUT) );
  AND2X2 AND2X2_4551 ( .A(u2__abc_44228_n3062_bF_buf69), .B(u2_remHi_209_), .Y(u2__abc_44228_n11113) );
  AND2X2 AND2X2_4552 ( .A(u2__abc_44228_n11100), .B(u2__abc_44228_n5450), .Y(u2__abc_44228_n11114) );
  AND2X2 AND2X2_4553 ( .A(u2__abc_44228_n11116_1), .B(u2__abc_44228_n11118), .Y(u2__abc_44228_n11119) );
  AND2X2 AND2X2_4554 ( .A(u2__abc_44228_n11119), .B(u2__abc_44228_n7547_bF_buf21), .Y(u2__abc_44228_n11120) );
  AND2X2 AND2X2_4555 ( .A(u2__abc_44228_n7548_1_bF_buf22), .B(u2_remHi_207_), .Y(u2__abc_44228_n11121) );
  AND2X2 AND2X2_4556 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n4631), .Y(u2__abc_44228_n11124_1) );
  AND2X2 AND2X2_4557 ( .A(u2__abc_44228_n11125), .B(u2__abc_44228_n2972_bF_buf4), .Y(u2__abc_44228_n11126) );
  AND2X2 AND2X2_4558 ( .A(u2__abc_44228_n11123_1), .B(u2__abc_44228_n11126), .Y(u2__abc_44228_n11127) );
  AND2X2 AND2X2_4559 ( .A(u2__abc_44228_n11128), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_remHi_209__FF_INPUT) );
  AND2X2 AND2X2_456 ( .A(u1__abc_43968_n264), .B(u1__abc_43968_n265), .Y(u1__abc_43968_n266_1) );
  AND2X2 AND2X2_4560 ( .A(u2__abc_44228_n3062_bF_buf68), .B(u2_remHi_210_), .Y(u2__abc_44228_n11130_1) );
  AND2X2 AND2X2_4561 ( .A(u2__abc_44228_n11098), .B(u2__abc_44228_n4655), .Y(u2__abc_44228_n11131_1) );
  AND2X2 AND2X2_4562 ( .A(u2__abc_44228_n11132), .B(u2__abc_44228_n4640), .Y(u2__abc_44228_n11134) );
  AND2X2 AND2X2_4563 ( .A(u2__abc_44228_n11135), .B(u2__abc_44228_n11133), .Y(u2__abc_44228_n11136) );
  AND2X2 AND2X2_4564 ( .A(u2__abc_44228_n11137_1), .B(u2__abc_44228_n11138_1), .Y(u2__abc_44228_n11139) );
  AND2X2 AND2X2_4565 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n4615), .Y(u2__abc_44228_n11141) );
  AND2X2 AND2X2_4566 ( .A(u2__abc_44228_n11142), .B(u2__abc_44228_n2972_bF_buf3), .Y(u2__abc_44228_n11143) );
  AND2X2 AND2X2_4567 ( .A(u2__abc_44228_n11140), .B(u2__abc_44228_n11143), .Y(u2__abc_44228_n11144_1) );
  AND2X2 AND2X2_4568 ( .A(u2__abc_44228_n11145_1), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_remHi_210__FF_INPUT) );
  AND2X2 AND2X2_4569 ( .A(u2__abc_44228_n3062_bF_buf67), .B(u2_remHi_211_), .Y(u2__abc_44228_n11147) );
  AND2X2 AND2X2_457 ( .A(u1__abc_43968_n263), .B(u1__abc_43968_n266_1), .Y(u1__abc_43968_n267_1) );
  AND2X2 AND2X2_4570 ( .A(u2__abc_44228_n11152_1), .B(u2__abc_44228_n7547_bF_buf19), .Y(u2__abc_44228_n11153) );
  AND2X2 AND2X2_4571 ( .A(u2__abc_44228_n11153), .B(u2__abc_44228_n11151_1), .Y(u2__abc_44228_n11154) );
  AND2X2 AND2X2_4572 ( .A(u2__abc_44228_n7548_1_bF_buf20), .B(u2_remHi_209_), .Y(u2__abc_44228_n11155) );
  AND2X2 AND2X2_4573 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n4622), .Y(u2__abc_44228_n11158_1) );
  AND2X2 AND2X2_4574 ( .A(u2__abc_44228_n11159_1), .B(u2__abc_44228_n2972_bF_buf2), .Y(u2__abc_44228_n11160) );
  AND2X2 AND2X2_4575 ( .A(u2__abc_44228_n11157), .B(u2__abc_44228_n11160), .Y(u2__abc_44228_n11161) );
  AND2X2 AND2X2_4576 ( .A(u2__abc_44228_n11162), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_remHi_211__FF_INPUT) );
  AND2X2 AND2X2_4577 ( .A(u2__abc_44228_n3062_bF_buf66), .B(u2_remHi_212_), .Y(u2__abc_44228_n11164) );
  AND2X2 AND2X2_4578 ( .A(u2__abc_44228_n11098), .B(u2__abc_44228_n4656_1), .Y(u2__abc_44228_n11165_1) );
  AND2X2 AND2X2_4579 ( .A(u2__abc_44228_n11166_1), .B(u2__abc_44228_n4618), .Y(u2__abc_44228_n11167) );
  AND2X2 AND2X2_458 ( .A(u1__abc_43968_n268_1), .B(u1__abc_43968_n269_1), .Y(u1__abc_43968_n270) );
  AND2X2 AND2X2_4580 ( .A(u2__abc_44228_n11168), .B(u2__abc_44228_n11169), .Y(u2__abc_44228_n11170) );
  AND2X2 AND2X2_4581 ( .A(u2__abc_44228_n11171), .B(u2__abc_44228_n11172_1), .Y(u2__abc_44228_n11173_1) );
  AND2X2 AND2X2_4582 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n4608), .Y(u2__abc_44228_n11175) );
  AND2X2 AND2X2_4583 ( .A(u2__abc_44228_n11176), .B(u2__abc_44228_n2972_bF_buf1), .Y(u2__abc_44228_n11177) );
  AND2X2 AND2X2_4584 ( .A(u2__abc_44228_n11174), .B(u2__abc_44228_n11177), .Y(u2__abc_44228_n11178) );
  AND2X2 AND2X2_4585 ( .A(u2__abc_44228_n11179_1), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_remHi_212__FF_INPUT) );
  AND2X2 AND2X2_4586 ( .A(u2__abc_44228_n3062_bF_buf65), .B(u2_remHi_213_), .Y(u2__abc_44228_n11181) );
  AND2X2 AND2X2_4587 ( .A(u2__abc_44228_n11168), .B(u2__abc_44228_n5459), .Y(u2__abc_44228_n11182) );
  AND2X2 AND2X2_4588 ( .A(u2__abc_44228_n11182), .B(u2__abc_44228_n4625), .Y(u2__abc_44228_n11183) );
  AND2X2 AND2X2_4589 ( .A(u2__abc_44228_n11185), .B(u2__abc_44228_n11184), .Y(u2__abc_44228_n11186_1) );
  AND2X2 AND2X2_459 ( .A(u1__abc_43968_n271), .B(u1__abc_43968_n272_1), .Y(u1__abc_43968_n273_1) );
  AND2X2 AND2X2_4590 ( .A(u2__abc_44228_n11187_1), .B(u2__abc_44228_n7547_bF_buf17), .Y(u2__abc_44228_n11188) );
  AND2X2 AND2X2_4591 ( .A(u2__abc_44228_n7548_1_bF_buf18), .B(u2_remHi_211_), .Y(u2__abc_44228_n11189) );
  AND2X2 AND2X2_4592 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n4602), .Y(u2__abc_44228_n11192) );
  AND2X2 AND2X2_4593 ( .A(u2__abc_44228_n11193_1), .B(u2__abc_44228_n2972_bF_buf0), .Y(u2__abc_44228_n11194_1) );
  AND2X2 AND2X2_4594 ( .A(u2__abc_44228_n11191), .B(u2__abc_44228_n11194_1), .Y(u2__abc_44228_n11195) );
  AND2X2 AND2X2_4595 ( .A(u2__abc_44228_n11196), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_remHi_213__FF_INPUT) );
  AND2X2 AND2X2_4596 ( .A(u2__abc_44228_n3062_bF_buf64), .B(u2_remHi_214_), .Y(u2__abc_44228_n11198) );
  AND2X2 AND2X2_4597 ( .A(u2__abc_44228_n11168), .B(u2__abc_44228_n5460), .Y(u2__abc_44228_n11199) );
  AND2X2 AND2X2_4598 ( .A(u2__abc_44228_n11201_1), .B(u2__abc_44228_n4611), .Y(u2__abc_44228_n11203) );
  AND2X2 AND2X2_4599 ( .A(u2__abc_44228_n11204), .B(u2__abc_44228_n11202), .Y(u2__abc_44228_n11205) );
  AND2X2 AND2X2_46 ( .A(_abc_64468_n753_bF_buf10), .B(sqrto_45_), .Y(_auto_iopadmap_cc_313_execute_65414_81_) );
  AND2X2 AND2X2_460 ( .A(u1__abc_43968_n270), .B(u1__abc_43968_n273_1), .Y(u1__abc_43968_n274) );
  AND2X2 AND2X2_4600 ( .A(u2__abc_44228_n11205), .B(u2__abc_44228_n7547_bF_buf16), .Y(u2__abc_44228_n11206) );
  AND2X2 AND2X2_4601 ( .A(u2__abc_44228_n7548_1_bF_buf17), .B(u2_remHi_212_), .Y(u2__abc_44228_n11207_1) );
  AND2X2 AND2X2_4602 ( .A(u2__abc_44228_n2983_bF_buf19), .B(u2__abc_44228_n4585), .Y(u2__abc_44228_n11210) );
  AND2X2 AND2X2_4603 ( .A(u2__abc_44228_n11211), .B(u2__abc_44228_n2972_bF_buf107), .Y(u2__abc_44228_n11212) );
  AND2X2 AND2X2_4604 ( .A(u2__abc_44228_n11209), .B(u2__abc_44228_n11212), .Y(u2__abc_44228_n11213) );
  AND2X2 AND2X2_4605 ( .A(u2__abc_44228_n11214_1), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_remHi_214__FF_INPUT) );
  AND2X2 AND2X2_4606 ( .A(u2__abc_44228_n3062_bF_buf63), .B(u2_remHi_215_), .Y(u2__abc_44228_n11216) );
  AND2X2 AND2X2_4607 ( .A(u2__abc_44228_n11221_1), .B(u2__abc_44228_n7547_bF_buf15), .Y(u2__abc_44228_n11222_1) );
  AND2X2 AND2X2_4608 ( .A(u2__abc_44228_n11222_1), .B(u2__abc_44228_n11220), .Y(u2__abc_44228_n11223) );
  AND2X2 AND2X2_4609 ( .A(u2__abc_44228_n7548_1_bF_buf16), .B(u2_remHi_213_), .Y(u2__abc_44228_n11224) );
  AND2X2 AND2X2_461 ( .A(u1__abc_43968_n267_1), .B(u1__abc_43968_n274), .Y(u1__abc_43968_n275) );
  AND2X2 AND2X2_4610 ( .A(u2__abc_44228_n2983_bF_buf17), .B(u2__abc_44228_n4592), .Y(u2__abc_44228_n11227) );
  AND2X2 AND2X2_4611 ( .A(u2__abc_44228_n11228_1), .B(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n11229_1) );
  AND2X2 AND2X2_4612 ( .A(u2__abc_44228_n11226), .B(u2__abc_44228_n11229_1), .Y(u2__abc_44228_n11230) );
  AND2X2 AND2X2_4613 ( .A(u2__abc_44228_n11231), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_remHi_215__FF_INPUT) );
  AND2X2 AND2X2_4614 ( .A(u2__abc_44228_n3062_bF_buf62), .B(u2_remHi_216_), .Y(u2__abc_44228_n11233) );
  AND2X2 AND2X2_4615 ( .A(u2__abc_44228_n11098), .B(u2__abc_44228_n4657), .Y(u2__abc_44228_n11234) );
  AND2X2 AND2X2_4616 ( .A(u2__abc_44228_n11235_1), .B(u2__abc_44228_n4588), .Y(u2__abc_44228_n11237) );
  AND2X2 AND2X2_4617 ( .A(u2__abc_44228_n11238), .B(u2__abc_44228_n11236_1), .Y(u2__abc_44228_n11239) );
  AND2X2 AND2X2_4618 ( .A(u2__abc_44228_n11240), .B(u2__abc_44228_n11241), .Y(u2__abc_44228_n11242_1) );
  AND2X2 AND2X2_4619 ( .A(u2__abc_44228_n2983_bF_buf15), .B(u2__abc_44228_n4578), .Y(u2__abc_44228_n11244) );
  AND2X2 AND2X2_462 ( .A(u1__abc_43968_n276), .B(u1__abc_43968_n277), .Y(u1__abc_43968_n278) );
  AND2X2 AND2X2_4620 ( .A(u2__abc_44228_n11245), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n11246) );
  AND2X2 AND2X2_4621 ( .A(u2__abc_44228_n11243_1), .B(u2__abc_44228_n11246), .Y(u2__abc_44228_n11247) );
  AND2X2 AND2X2_4622 ( .A(u2__abc_44228_n11248), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_remHi_216__FF_INPUT) );
  AND2X2 AND2X2_4623 ( .A(u2__abc_44228_n3062_bF_buf61), .B(u2_remHi_217_), .Y(u2__abc_44228_n11250_1) );
  AND2X2 AND2X2_4624 ( .A(u2__abc_44228_n11238), .B(u2__abc_44228_n5469), .Y(u2__abc_44228_n11251) );
  AND2X2 AND2X2_4625 ( .A(u2__abc_44228_n11251), .B(u2__abc_44228_n4595), .Y(u2__abc_44228_n11252) );
  AND2X2 AND2X2_4626 ( .A(u2__abc_44228_n11254), .B(u2__abc_44228_n11253), .Y(u2__abc_44228_n11255) );
  AND2X2 AND2X2_4627 ( .A(u2__abc_44228_n11256_1), .B(u2__abc_44228_n7547_bF_buf13), .Y(u2__abc_44228_n11257_1) );
  AND2X2 AND2X2_4628 ( .A(u2__abc_44228_n7548_1_bF_buf14), .B(u2_remHi_215_), .Y(u2__abc_44228_n11258) );
  AND2X2 AND2X2_4629 ( .A(u2__abc_44228_n2983_bF_buf13), .B(u2__abc_44228_n4572_1), .Y(u2__abc_44228_n11261) );
  AND2X2 AND2X2_463 ( .A(u1__abc_43968_n279), .B(u1__abc_43968_n280), .Y(u1__abc_43968_n281) );
  AND2X2 AND2X2_4630 ( .A(u2__abc_44228_n11262), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n11263_1) );
  AND2X2 AND2X2_4631 ( .A(u2__abc_44228_n11260), .B(u2__abc_44228_n11263_1), .Y(u2__abc_44228_n11264_1) );
  AND2X2 AND2X2_4632 ( .A(u2__abc_44228_n11265), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_remHi_217__FF_INPUT) );
  AND2X2 AND2X2_4633 ( .A(u2__abc_44228_n3062_bF_buf60), .B(u2_remHi_218_), .Y(u2__abc_44228_n11267) );
  AND2X2 AND2X2_4634 ( .A(u2__abc_44228_n11238), .B(u2__abc_44228_n5470), .Y(u2__abc_44228_n11268) );
  AND2X2 AND2X2_4635 ( .A(u2__abc_44228_n11270_1), .B(u2__abc_44228_n4581_1), .Y(u2__abc_44228_n11272) );
  AND2X2 AND2X2_4636 ( .A(u2__abc_44228_n11273), .B(u2__abc_44228_n11271_1), .Y(u2__abc_44228_n11274) );
  AND2X2 AND2X2_4637 ( .A(u2__abc_44228_n11274), .B(u2__abc_44228_n7547_bF_buf12), .Y(u2__abc_44228_n11275) );
  AND2X2 AND2X2_4638 ( .A(u2__abc_44228_n7548_1_bF_buf13), .B(u2_remHi_216_), .Y(u2__abc_44228_n11276) );
  AND2X2 AND2X2_4639 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n4556), .Y(u2__abc_44228_n11279) );
  AND2X2 AND2X2_464 ( .A(u1__abc_43968_n278), .B(u1__abc_43968_n281), .Y(u1__abc_43968_n282) );
  AND2X2 AND2X2_4640 ( .A(u2__abc_44228_n11280), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n11281) );
  AND2X2 AND2X2_4641 ( .A(u2__abc_44228_n11278_1), .B(u2__abc_44228_n11281), .Y(u2__abc_44228_n11282) );
  AND2X2 AND2X2_4642 ( .A(u2__abc_44228_n11283), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_remHi_218__FF_INPUT) );
  AND2X2 AND2X2_4643 ( .A(u2__abc_44228_n3062_bF_buf59), .B(u2_remHi_219_), .Y(u2__abc_44228_n11285_1) );
  AND2X2 AND2X2_4644 ( .A(u2__abc_44228_n11290), .B(u2__abc_44228_n7547_bF_buf11), .Y(u2__abc_44228_n11291_1) );
  AND2X2 AND2X2_4645 ( .A(u2__abc_44228_n11291_1), .B(u2__abc_44228_n11289), .Y(u2__abc_44228_n11292_1) );
  AND2X2 AND2X2_4646 ( .A(u2__abc_44228_n7548_1_bF_buf12), .B(u2_remHi_217_), .Y(u2__abc_44228_n11293) );
  AND2X2 AND2X2_4647 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n4563_1), .Y(u2__abc_44228_n11296) );
  AND2X2 AND2X2_4648 ( .A(u2__abc_44228_n11297), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n11298_1) );
  AND2X2 AND2X2_4649 ( .A(u2__abc_44228_n11295), .B(u2__abc_44228_n11298_1), .Y(u2__abc_44228_n11299_1) );
  AND2X2 AND2X2_465 ( .A(u1__abc_43968_n283), .B(u1__abc_43968_n284), .Y(u1__abc_43968_n285) );
  AND2X2 AND2X2_4650 ( .A(u2__abc_44228_n11300), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_remHi_219__FF_INPUT) );
  AND2X2 AND2X2_4651 ( .A(u2__abc_44228_n3062_bF_buf58), .B(u2_remHi_220_), .Y(u2__abc_44228_n11302) );
  AND2X2 AND2X2_4652 ( .A(u2__abc_44228_n11235_1), .B(u2__abc_44228_n4597), .Y(u2__abc_44228_n11303) );
  AND2X2 AND2X2_4653 ( .A(u2__abc_44228_n11304), .B(u2__abc_44228_n4559), .Y(u2__abc_44228_n11305_1) );
  AND2X2 AND2X2_4654 ( .A(u2__abc_44228_n11306_1), .B(u2__abc_44228_n11307), .Y(u2__abc_44228_n11308) );
  AND2X2 AND2X2_4655 ( .A(u2__abc_44228_n11308), .B(u2__abc_44228_n7547_bF_buf10), .Y(u2__abc_44228_n11309) );
  AND2X2 AND2X2_4656 ( .A(u2__abc_44228_n7548_1_bF_buf11), .B(u2_remHi_218_), .Y(u2__abc_44228_n11310) );
  AND2X2 AND2X2_4657 ( .A(u2__abc_44228_n2983_bF_buf9), .B(u2__abc_44228_n4549), .Y(u2__abc_44228_n11313_1) );
  AND2X2 AND2X2_4658 ( .A(u2__abc_44228_n11314), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n11315) );
  AND2X2 AND2X2_4659 ( .A(u2__abc_44228_n11312_1), .B(u2__abc_44228_n11315), .Y(u2__abc_44228_n11316) );
  AND2X2 AND2X2_466 ( .A(u1__abc_43968_n286), .B(u1__abc_43968_n287), .Y(u1__abc_43968_n288) );
  AND2X2 AND2X2_4660 ( .A(u2__abc_44228_n11317), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_remHi_220__FF_INPUT) );
  AND2X2 AND2X2_4661 ( .A(u2__abc_44228_n3062_bF_buf57), .B(u2_remHi_221_), .Y(u2__abc_44228_n11319_1) );
  AND2X2 AND2X2_4662 ( .A(u2__abc_44228_n11306_1), .B(u2__abc_44228_n5480), .Y(u2__abc_44228_n11320_1) );
  AND2X2 AND2X2_4663 ( .A(u2__abc_44228_n11324), .B(u2__abc_44228_n7547_bF_buf9), .Y(u2__abc_44228_n11325) );
  AND2X2 AND2X2_4664 ( .A(u2__abc_44228_n11325), .B(u2__abc_44228_n11322), .Y(u2__abc_44228_n11326_1) );
  AND2X2 AND2X2_4665 ( .A(u2__abc_44228_n7548_1_bF_buf10), .B(u2_remHi_219_), .Y(u2__abc_44228_n11327_1) );
  AND2X2 AND2X2_4666 ( .A(u2__abc_44228_n2983_bF_buf7), .B(u2__abc_44228_n4543), .Y(u2__abc_44228_n11330) );
  AND2X2 AND2X2_4667 ( .A(u2__abc_44228_n11331), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n11332) );
  AND2X2 AND2X2_4668 ( .A(u2__abc_44228_n11329), .B(u2__abc_44228_n11332), .Y(u2__abc_44228_n11333_1) );
  AND2X2 AND2X2_4669 ( .A(u2__abc_44228_n11334_1), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_remHi_221__FF_INPUT) );
  AND2X2 AND2X2_467 ( .A(u1__abc_43968_n285), .B(u1__abc_43968_n288), .Y(u1__abc_43968_n289) );
  AND2X2 AND2X2_4670 ( .A(u2__abc_44228_n3062_bF_buf56), .B(u2_remHi_222_), .Y(u2__abc_44228_n11336) );
  AND2X2 AND2X2_4671 ( .A(u2__abc_44228_n11306_1), .B(u2__abc_44228_n5481), .Y(u2__abc_44228_n11337) );
  AND2X2 AND2X2_4672 ( .A(u2__abc_44228_n11339), .B(u2__abc_44228_n4552), .Y(u2__abc_44228_n11341_1) );
  AND2X2 AND2X2_4673 ( .A(u2__abc_44228_n11342), .B(u2__abc_44228_n11340_1), .Y(u2__abc_44228_n11343) );
  AND2X2 AND2X2_4674 ( .A(u2__abc_44228_n11343), .B(u2__abc_44228_n7547_bF_buf8), .Y(u2__abc_44228_n11344) );
  AND2X2 AND2X2_4675 ( .A(u2__abc_44228_n7548_1_bF_buf9), .B(u2_remHi_220_), .Y(u2__abc_44228_n11345) );
  AND2X2 AND2X2_4676 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n4524), .Y(u2__abc_44228_n11348_1) );
  AND2X2 AND2X2_4677 ( .A(u2__abc_44228_n11349), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n11350) );
  AND2X2 AND2X2_4678 ( .A(u2__abc_44228_n11347_1), .B(u2__abc_44228_n11350), .Y(u2__abc_44228_n11351) );
  AND2X2 AND2X2_4679 ( .A(u2__abc_44228_n11352), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_remHi_222__FF_INPUT) );
  AND2X2 AND2X2_468 ( .A(u1__abc_43968_n282), .B(u1__abc_43968_n289), .Y(u1__abc_43968_n290) );
  AND2X2 AND2X2_4680 ( .A(u2__abc_44228_n3062_bF_buf55), .B(u2_remHi_223_), .Y(u2__abc_44228_n11354_1) );
  AND2X2 AND2X2_4681 ( .A(u2__abc_44228_n11359), .B(u2__abc_44228_n7547_bF_buf7), .Y(u2__abc_44228_n11360) );
  AND2X2 AND2X2_4682 ( .A(u2__abc_44228_n11360), .B(u2__abc_44228_n11358), .Y(u2__abc_44228_n11361_1) );
  AND2X2 AND2X2_4683 ( .A(u2__abc_44228_n7548_1_bF_buf8), .B(u2_remHi_221_), .Y(u2__abc_44228_n11362_1) );
  AND2X2 AND2X2_4684 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n4531), .Y(u2__abc_44228_n11365) );
  AND2X2 AND2X2_4685 ( .A(u2__abc_44228_n11366), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n11367) );
  AND2X2 AND2X2_4686 ( .A(u2__abc_44228_n11364), .B(u2__abc_44228_n11367), .Y(u2__abc_44228_n11368_1) );
  AND2X2 AND2X2_4687 ( .A(u2__abc_44228_n11369_1), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_remHi_223__FF_INPUT) );
  AND2X2 AND2X2_4688 ( .A(u2__abc_44228_n3062_bF_buf54), .B(u2_remHi_224_), .Y(u2__abc_44228_n11371) );
  AND2X2 AND2X2_4689 ( .A(u2__abc_44228_n10826), .B(u2__abc_44228_n4778), .Y(u2__abc_44228_n11372) );
  AND2X2 AND2X2_469 ( .A(u1__abc_43968_n275), .B(u1__abc_43968_n290), .Y(u1__abc_43968_n291) );
  AND2X2 AND2X2_4690 ( .A(u2__abc_44228_n11373), .B(u2__abc_44228_n4527), .Y(u2__abc_44228_n11375_1) );
  AND2X2 AND2X2_4691 ( .A(u2__abc_44228_n11376_1), .B(u2__abc_44228_n11374), .Y(u2__abc_44228_n11377) );
  AND2X2 AND2X2_4692 ( .A(u2__abc_44228_n11378), .B(u2__abc_44228_n11379), .Y(u2__abc_44228_n11380) );
  AND2X2 AND2X2_4693 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n4517_1), .Y(u2__abc_44228_n11382_1) );
  AND2X2 AND2X2_4694 ( .A(u2__abc_44228_n11383_1), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n11384) );
  AND2X2 AND2X2_4695 ( .A(u2__abc_44228_n11381), .B(u2__abc_44228_n11384), .Y(u2__abc_44228_n11385) );
  AND2X2 AND2X2_4696 ( .A(u2__abc_44228_n11386), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_remHi_224__FF_INPUT) );
  AND2X2 AND2X2_4697 ( .A(u2__abc_44228_n3062_bF_buf53), .B(u2_remHi_225_), .Y(u2__abc_44228_n11388) );
  AND2X2 AND2X2_4698 ( .A(u2__abc_44228_n11376_1), .B(u2__abc_44228_n5490), .Y(u2__abc_44228_n11390_1) );
  AND2X2 AND2X2_4699 ( .A(u2__abc_44228_n11393), .B(u2__abc_44228_n11391), .Y(u2__abc_44228_n11394) );
  AND2X2 AND2X2_47 ( .A(_abc_64468_n753_bF_buf9), .B(sqrto_46_), .Y(_auto_iopadmap_cc_313_execute_65414_82_) );
  AND2X2 AND2X2_470 ( .A(u1__abc_43968_n292), .B(u1__abc_43968_n293), .Y(u1__abc_43968_n294) );
  AND2X2 AND2X2_4700 ( .A(u2__abc_44228_n11394), .B(u2__abc_44228_n7547_bF_buf5), .Y(u2__abc_44228_n11395) );
  AND2X2 AND2X2_4701 ( .A(u2__abc_44228_n7548_1_bF_buf6), .B(u2_remHi_223_), .Y(u2__abc_44228_n11396_1) );
  AND2X2 AND2X2_4702 ( .A(u2__abc_44228_n2983_bF_buf1), .B(u2__abc_44228_n4511), .Y(u2__abc_44228_n11399) );
  AND2X2 AND2X2_4703 ( .A(u2__abc_44228_n11400), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n11401) );
  AND2X2 AND2X2_4704 ( .A(u2__abc_44228_n11398), .B(u2__abc_44228_n11401), .Y(u2__abc_44228_n11402) );
  AND2X2 AND2X2_4705 ( .A(u2__abc_44228_n11403_1), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_remHi_225__FF_INPUT) );
  AND2X2 AND2X2_4706 ( .A(u2__abc_44228_n3062_bF_buf52), .B(u2_remHi_226_), .Y(u2__abc_44228_n11405) );
  AND2X2 AND2X2_4707 ( .A(u2__abc_44228_n11373), .B(u2__abc_44228_n4535_1), .Y(u2__abc_44228_n11406) );
  AND2X2 AND2X2_4708 ( .A(u2__abc_44228_n11407), .B(u2__abc_44228_n4520), .Y(u2__abc_44228_n11409) );
  AND2X2 AND2X2_4709 ( .A(u2__abc_44228_n11410_1), .B(u2__abc_44228_n11408), .Y(u2__abc_44228_n11411_1) );
  AND2X2 AND2X2_471 ( .A(u1__abc_43968_n295), .B(u1__abc_43968_n296), .Y(u1__abc_43968_n297) );
  AND2X2 AND2X2_4710 ( .A(u2__abc_44228_n11412), .B(u2__abc_44228_n11413), .Y(u2__abc_44228_n11414) );
  AND2X2 AND2X2_4711 ( .A(u2__abc_44228_n2983_bF_buf141), .B(u2__abc_44228_n4495), .Y(u2__abc_44228_n11416) );
  AND2X2 AND2X2_4712 ( .A(u2__abc_44228_n11417_1), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n11418_1) );
  AND2X2 AND2X2_4713 ( .A(u2__abc_44228_n11415), .B(u2__abc_44228_n11418_1), .Y(u2__abc_44228_n11419) );
  AND2X2 AND2X2_4714 ( .A(u2__abc_44228_n11420), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_remHi_226__FF_INPUT) );
  AND2X2 AND2X2_4715 ( .A(u2__abc_44228_n3062_bF_buf51), .B(u2_remHi_227_), .Y(u2__abc_44228_n11422) );
  AND2X2 AND2X2_4716 ( .A(u2__abc_44228_n11427), .B(u2__abc_44228_n7547_bF_buf3), .Y(u2__abc_44228_n11428) );
  AND2X2 AND2X2_4717 ( .A(u2__abc_44228_n11428), .B(u2__abc_44228_n11426), .Y(u2__abc_44228_n11429) );
  AND2X2 AND2X2_4718 ( .A(u2__abc_44228_n7548_1_bF_buf4), .B(u2_remHi_225_), .Y(u2__abc_44228_n11430) );
  AND2X2 AND2X2_4719 ( .A(u2__abc_44228_n2983_bF_buf139), .B(u2__abc_44228_n4502), .Y(u2__abc_44228_n11433) );
  AND2X2 AND2X2_472 ( .A(u1__abc_43968_n294), .B(u1__abc_43968_n297), .Y(u1__abc_43968_n298) );
  AND2X2 AND2X2_4720 ( .A(u2__abc_44228_n11434), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n11435) );
  AND2X2 AND2X2_4721 ( .A(u2__abc_44228_n11432_1), .B(u2__abc_44228_n11435), .Y(u2__abc_44228_n11436) );
  AND2X2 AND2X2_4722 ( .A(u2__abc_44228_n11437), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_remHi_227__FF_INPUT) );
  AND2X2 AND2X2_4723 ( .A(u2__abc_44228_n3062_bF_buf50), .B(u2_remHi_228_), .Y(u2__abc_44228_n11439_1) );
  AND2X2 AND2X2_4724 ( .A(u2__abc_44228_n11373), .B(u2__abc_44228_n4536), .Y(u2__abc_44228_n11440) );
  AND2X2 AND2X2_4725 ( .A(u2__abc_44228_n11441), .B(u2__abc_44228_n4498_1), .Y(u2__abc_44228_n11442) );
  AND2X2 AND2X2_4726 ( .A(u2__abc_44228_n11443), .B(u2__abc_44228_n11444), .Y(u2__abc_44228_n11445_1) );
  AND2X2 AND2X2_4727 ( .A(u2__abc_44228_n11446_1), .B(u2__abc_44228_n11447), .Y(u2__abc_44228_n11448) );
  AND2X2 AND2X2_4728 ( .A(u2__abc_44228_n2983_bF_buf137), .B(u2__abc_44228_n4488), .Y(u2__abc_44228_n11450) );
  AND2X2 AND2X2_4729 ( .A(u2__abc_44228_n11451), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n11452_1) );
  AND2X2 AND2X2_473 ( .A(u1__abc_43968_n299), .B(u1__abc_43968_n300), .Y(u1__abc_43968_n301) );
  AND2X2 AND2X2_4730 ( .A(u2__abc_44228_n11449), .B(u2__abc_44228_n11452_1), .Y(u2__abc_44228_n11453_1) );
  AND2X2 AND2X2_4731 ( .A(u2__abc_44228_n11454), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_remHi_228__FF_INPUT) );
  AND2X2 AND2X2_4732 ( .A(u2__abc_44228_n3062_bF_buf49), .B(u2_remHi_229_), .Y(u2__abc_44228_n11456) );
  AND2X2 AND2X2_4733 ( .A(u2__abc_44228_n11443), .B(u2__abc_44228_n5499), .Y(u2__abc_44228_n11457) );
  AND2X2 AND2X2_4734 ( .A(u2__abc_44228_n11461), .B(u2__abc_44228_n7547_bF_buf1), .Y(u2__abc_44228_n11462) );
  AND2X2 AND2X2_4735 ( .A(u2__abc_44228_n11462), .B(u2__abc_44228_n11459_1), .Y(u2__abc_44228_n11463) );
  AND2X2 AND2X2_4736 ( .A(u2__abc_44228_n7548_1_bF_buf2), .B(u2_remHi_227_), .Y(u2__abc_44228_n11464) );
  AND2X2 AND2X2_4737 ( .A(u2__abc_44228_n2983_bF_buf135), .B(u2__abc_44228_n4482), .Y(u2__abc_44228_n11467_1) );
  AND2X2 AND2X2_4738 ( .A(u2__abc_44228_n11468), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n11469) );
  AND2X2 AND2X2_4739 ( .A(u2__abc_44228_n11466_1), .B(u2__abc_44228_n11469), .Y(u2__abc_44228_n11470) );
  AND2X2 AND2X2_474 ( .A(u1__abc_43968_n302), .B(u1__abc_43968_n303), .Y(u1__abc_43968_n304) );
  AND2X2 AND2X2_4740 ( .A(u2__abc_44228_n11471), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_remHi_229__FF_INPUT) );
  AND2X2 AND2X2_4741 ( .A(u2__abc_44228_n3062_bF_buf48), .B(u2_remHi_230_), .Y(u2__abc_44228_n11473_1) );
  AND2X2 AND2X2_4742 ( .A(u2__abc_44228_n11443), .B(u2__abc_44228_n5500), .Y(u2__abc_44228_n11474_1) );
  AND2X2 AND2X2_4743 ( .A(u2__abc_44228_n11476), .B(u2__abc_44228_n4491), .Y(u2__abc_44228_n11478) );
  AND2X2 AND2X2_4744 ( .A(u2__abc_44228_n11479), .B(u2__abc_44228_n11477), .Y(u2__abc_44228_n11480_1) );
  AND2X2 AND2X2_4745 ( .A(u2__abc_44228_n11480_1), .B(u2__abc_44228_n7547_bF_buf0), .Y(u2__abc_44228_n11481_1) );
  AND2X2 AND2X2_4746 ( .A(u2__abc_44228_n7548_1_bF_buf1), .B(u2_remHi_228_), .Y(u2__abc_44228_n11482) );
  AND2X2 AND2X2_4747 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n4458), .Y(u2__abc_44228_n11485) );
  AND2X2 AND2X2_4748 ( .A(u2__abc_44228_n11486), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n11487_1) );
  AND2X2 AND2X2_4749 ( .A(u2__abc_44228_n11484), .B(u2__abc_44228_n11487_1), .Y(u2__abc_44228_n11488_1) );
  AND2X2 AND2X2_475 ( .A(u1__abc_43968_n301), .B(u1__abc_43968_n304), .Y(u1__abc_43968_n305) );
  AND2X2 AND2X2_4750 ( .A(u2__abc_44228_n11489), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_remHi_230__FF_INPUT) );
  AND2X2 AND2X2_4751 ( .A(u2__abc_44228_n3062_bF_buf47), .B(u2_remHi_231_), .Y(u2__abc_44228_n11491) );
  AND2X2 AND2X2_4752 ( .A(u2__abc_44228_n11496), .B(u2__abc_44228_n7547_bF_buf57), .Y(u2__abc_44228_n11497) );
  AND2X2 AND2X2_4753 ( .A(u2__abc_44228_n11497), .B(u2__abc_44228_n11495_1), .Y(u2__abc_44228_n11498) );
  AND2X2 AND2X2_4754 ( .A(u2__abc_44228_n7548_1_bF_buf0), .B(u2_remHi_229_), .Y(u2__abc_44228_n11499) );
  AND2X2 AND2X2_4755 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n4452), .Y(u2__abc_44228_n11502_1) );
  AND2X2 AND2X2_4756 ( .A(u2__abc_44228_n11503), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n11504) );
  AND2X2 AND2X2_4757 ( .A(u2__abc_44228_n11501_1), .B(u2__abc_44228_n11504), .Y(u2__abc_44228_n11505) );
  AND2X2 AND2X2_4758 ( .A(u2__abc_44228_n11506), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_remHi_231__FF_INPUT) );
  AND2X2 AND2X2_4759 ( .A(u2__abc_44228_n3062_bF_buf46), .B(u2_remHi_232_), .Y(u2__abc_44228_n11508_1) );
  AND2X2 AND2X2_476 ( .A(u1__abc_43968_n298), .B(u1__abc_43968_n305), .Y(u1__abc_43968_n306) );
  AND2X2 AND2X2_4760 ( .A(u2__abc_44228_n11373), .B(u2__abc_44228_n4537), .Y(u2__abc_44228_n11509_1) );
  AND2X2 AND2X2_4761 ( .A(u2__abc_44228_n11510), .B(u2__abc_44228_n4461_1), .Y(u2__abc_44228_n11512) );
  AND2X2 AND2X2_4762 ( .A(u2__abc_44228_n11513), .B(u2__abc_44228_n11511), .Y(u2__abc_44228_n11514) );
  AND2X2 AND2X2_4763 ( .A(u2__abc_44228_n11515_1), .B(u2__abc_44228_n11516_1), .Y(u2__abc_44228_n11517) );
  AND2X2 AND2X2_4764 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n4472), .Y(u2__abc_44228_n11519) );
  AND2X2 AND2X2_4765 ( .A(u2__abc_44228_n11520), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n11521) );
  AND2X2 AND2X2_4766 ( .A(u2__abc_44228_n11518), .B(u2__abc_44228_n11521), .Y(u2__abc_44228_n11522_1) );
  AND2X2 AND2X2_4767 ( .A(u2__abc_44228_n11523_1), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_remHi_232__FF_INPUT) );
  AND2X2 AND2X2_4768 ( .A(u2__abc_44228_n3062_bF_buf45), .B(u2_remHi_233_), .Y(u2__abc_44228_n11525) );
  AND2X2 AND2X2_4769 ( .A(u2__abc_44228_n11513), .B(u2__abc_44228_n5509), .Y(u2__abc_44228_n11527) );
  AND2X2 AND2X2_477 ( .A(u1__abc_43968_n307), .B(u1__abc_43968_n308), .Y(u1__abc_43968_n309) );
  AND2X2 AND2X2_4770 ( .A(u2__abc_44228_n11530_1), .B(u2__abc_44228_n11528), .Y(u2__abc_44228_n11531) );
  AND2X2 AND2X2_4771 ( .A(u2__abc_44228_n11531), .B(u2__abc_44228_n7547_bF_buf55), .Y(u2__abc_44228_n11532) );
  AND2X2 AND2X2_4772 ( .A(u2__abc_44228_n7548_1_bF_buf56), .B(u2_remHi_231_), .Y(u2__abc_44228_n11533) );
  AND2X2 AND2X2_4773 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n4466), .Y(u2__abc_44228_n11536_1) );
  AND2X2 AND2X2_4774 ( .A(u2__abc_44228_n11537_1), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n11538) );
  AND2X2 AND2X2_4775 ( .A(u2__abc_44228_n11535), .B(u2__abc_44228_n11538), .Y(u2__abc_44228_n11539) );
  AND2X2 AND2X2_4776 ( .A(u2__abc_44228_n11540), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_remHi_233__FF_INPUT) );
  AND2X2 AND2X2_4777 ( .A(u2__abc_44228_n3062_bF_buf44), .B(u2_remHi_234_), .Y(u2__abc_44228_n11542) );
  AND2X2 AND2X2_4778 ( .A(u2__abc_44228_n11510), .B(u2__abc_44228_n4462), .Y(u2__abc_44228_n11543_1) );
  AND2X2 AND2X2_4779 ( .A(u2__abc_44228_n11544_1), .B(u2__abc_44228_n4475), .Y(u2__abc_44228_n11546) );
  AND2X2 AND2X2_478 ( .A(u1__abc_43968_n310), .B(u1__abc_43968_n311), .Y(u1__abc_43968_n312) );
  AND2X2 AND2X2_4780 ( .A(u2__abc_44228_n11547), .B(u2__abc_44228_n11545), .Y(u2__abc_44228_n11548) );
  AND2X2 AND2X2_4781 ( .A(u2__abc_44228_n11548), .B(u2__abc_44228_n7547_bF_buf54), .Y(u2__abc_44228_n11549) );
  AND2X2 AND2X2_4782 ( .A(u2__abc_44228_n7548_1_bF_buf55), .B(u2_remHi_232_), .Y(u2__abc_44228_n11550_1) );
  AND2X2 AND2X2_4783 ( .A(u2__abc_44228_n2983_bF_buf127), .B(u2__abc_44228_n4436), .Y(u2__abc_44228_n11553) );
  AND2X2 AND2X2_4784 ( .A(u2__abc_44228_n11554), .B(u2__abc_44228_n2972_bF_buf87), .Y(u2__abc_44228_n11555) );
  AND2X2 AND2X2_4785 ( .A(u2__abc_44228_n11552), .B(u2__abc_44228_n11555), .Y(u2__abc_44228_n11556) );
  AND2X2 AND2X2_4786 ( .A(u2__abc_44228_n11557_1), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_remHi_234__FF_INPUT) );
  AND2X2 AND2X2_4787 ( .A(u2__abc_44228_n3062_bF_buf43), .B(u2_remHi_235_), .Y(u2__abc_44228_n11559) );
  AND2X2 AND2X2_4788 ( .A(u2__abc_44228_n11547), .B(u2__abc_44228_n5514), .Y(u2__abc_44228_n11561) );
  AND2X2 AND2X2_4789 ( .A(u2__abc_44228_n11564_1), .B(u2__abc_44228_n11562), .Y(u2__abc_44228_n11565_1) );
  AND2X2 AND2X2_479 ( .A(u1__abc_43968_n309), .B(u1__abc_43968_n312), .Y(u1__abc_43968_n313) );
  AND2X2 AND2X2_4790 ( .A(u2__abc_44228_n11565_1), .B(u2__abc_44228_n7547_bF_buf53), .Y(u2__abc_44228_n11566) );
  AND2X2 AND2X2_4791 ( .A(u2__abc_44228_n7548_1_bF_buf54), .B(u2_remHi_233_), .Y(u2__abc_44228_n11567) );
  AND2X2 AND2X2_4792 ( .A(u2__abc_44228_n2983_bF_buf125), .B(u2__abc_44228_n4443), .Y(u2__abc_44228_n11570) );
  AND2X2 AND2X2_4793 ( .A(u2__abc_44228_n11571_1), .B(u2__abc_44228_n2972_bF_buf86), .Y(u2__abc_44228_n11572_1) );
  AND2X2 AND2X2_4794 ( .A(u2__abc_44228_n11569), .B(u2__abc_44228_n11572_1), .Y(u2__abc_44228_n11573) );
  AND2X2 AND2X2_4795 ( .A(u2__abc_44228_n11574), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_remHi_235__FF_INPUT) );
  AND2X2 AND2X2_4796 ( .A(u2__abc_44228_n3062_bF_buf42), .B(u2_remHi_236_), .Y(u2__abc_44228_n11576) );
  AND2X2 AND2X2_4797 ( .A(u2__abc_44228_n11547), .B(u2__abc_44228_n5515), .Y(u2__abc_44228_n11577) );
  AND2X2 AND2X2_4798 ( .A(u2__abc_44228_n11579_1), .B(u2__abc_44228_n4439), .Y(u2__abc_44228_n11580) );
  AND2X2 AND2X2_4799 ( .A(u2__abc_44228_n11581), .B(u2__abc_44228_n11582), .Y(u2__abc_44228_n11583) );
  AND2X2 AND2X2_48 ( .A(_abc_64468_n753_bF_buf8), .B(sqrto_47_), .Y(_auto_iopadmap_cc_313_execute_65414_83_) );
  AND2X2 AND2X2_480 ( .A(u1__abc_43968_n314), .B(u1__abc_43968_n315), .Y(u1__abc_43968_n316) );
  AND2X2 AND2X2_4800 ( .A(u2__abc_44228_n11583), .B(u2__abc_44228_n7547_bF_buf52), .Y(u2__abc_44228_n11584) );
  AND2X2 AND2X2_4801 ( .A(u2__abc_44228_n7548_1_bF_buf53), .B(u2_remHi_234_), .Y(u2__abc_44228_n11585_1) );
  AND2X2 AND2X2_4802 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n4429), .Y(u2__abc_44228_n11588) );
  AND2X2 AND2X2_4803 ( .A(u2__abc_44228_n11589), .B(u2__abc_44228_n2972_bF_buf85), .Y(u2__abc_44228_n11590) );
  AND2X2 AND2X2_4804 ( .A(u2__abc_44228_n11587), .B(u2__abc_44228_n11590), .Y(u2__abc_44228_n11591) );
  AND2X2 AND2X2_4805 ( .A(u2__abc_44228_n11592_1), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_remHi_236__FF_INPUT) );
  AND2X2 AND2X2_4806 ( .A(u2__abc_44228_n3062_bF_buf41), .B(u2_remHi_237_), .Y(u2__abc_44228_n11594) );
  AND2X2 AND2X2_4807 ( .A(u2__abc_44228_n11581), .B(u2__abc_44228_n5520), .Y(u2__abc_44228_n11595) );
  AND2X2 AND2X2_4808 ( .A(u2__abc_44228_n11599_1), .B(u2__abc_44228_n7547_bF_buf51), .Y(u2__abc_44228_n11600_1) );
  AND2X2 AND2X2_4809 ( .A(u2__abc_44228_n11600_1), .B(u2__abc_44228_n11597), .Y(u2__abc_44228_n11601) );
  AND2X2 AND2X2_481 ( .A(u1__abc_43968_n317), .B(u1__abc_43968_n318), .Y(u1__abc_43968_n319) );
  AND2X2 AND2X2_4810 ( .A(u2__abc_44228_n7548_1_bF_buf52), .B(u2_remHi_235_), .Y(u2__abc_44228_n11602) );
  AND2X2 AND2X2_4811 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n4423_1), .Y(u2__abc_44228_n11605) );
  AND2X2 AND2X2_4812 ( .A(u2__abc_44228_n11606_1), .B(u2__abc_44228_n2972_bF_buf84), .Y(u2__abc_44228_n11607_1) );
  AND2X2 AND2X2_4813 ( .A(u2__abc_44228_n11604), .B(u2__abc_44228_n11607_1), .Y(u2__abc_44228_n11608) );
  AND2X2 AND2X2_4814 ( .A(u2__abc_44228_n11609), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_remHi_237__FF_INPUT) );
  AND2X2 AND2X2_4815 ( .A(u2__abc_44228_n3062_bF_buf40), .B(u2_remHi_238_), .Y(u2__abc_44228_n11611) );
  AND2X2 AND2X2_4816 ( .A(u2__abc_44228_n11581), .B(u2__abc_44228_n5521), .Y(u2__abc_44228_n11612) );
  AND2X2 AND2X2_4817 ( .A(u2__abc_44228_n11614_1), .B(u2__abc_44228_n4432_1), .Y(u2__abc_44228_n11615) );
  AND2X2 AND2X2_4818 ( .A(u2__abc_44228_n11617), .B(u2__abc_44228_n7547_bF_buf50), .Y(u2__abc_44228_n11618) );
  AND2X2 AND2X2_4819 ( .A(u2__abc_44228_n11618), .B(u2__abc_44228_n11616), .Y(u2__abc_44228_n11619) );
  AND2X2 AND2X2_482 ( .A(u1__abc_43968_n316), .B(u1__abc_43968_n319), .Y(u1__abc_43968_n320) );
  AND2X2 AND2X2_4820 ( .A(u2__abc_44228_n7548_1_bF_buf51), .B(u2_remHi_236_), .Y(u2__abc_44228_n11620_1) );
  AND2X2 AND2X2_4821 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n4405_1), .Y(u2__abc_44228_n11623) );
  AND2X2 AND2X2_4822 ( .A(u2__abc_44228_n11624), .B(u2__abc_44228_n2972_bF_buf83), .Y(u2__abc_44228_n11625) );
  AND2X2 AND2X2_4823 ( .A(u2__abc_44228_n11622), .B(u2__abc_44228_n11625), .Y(u2__abc_44228_n11626) );
  AND2X2 AND2X2_4824 ( .A(u2__abc_44228_n11627_1), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_remHi_238__FF_INPUT) );
  AND2X2 AND2X2_4825 ( .A(u2__abc_44228_n3062_bF_buf39), .B(u2_remHi_239_), .Y(u2__abc_44228_n11629) );
  AND2X2 AND2X2_4826 ( .A(u2__abc_44228_n11634_1), .B(u2__abc_44228_n7547_bF_buf49), .Y(u2__abc_44228_n11635_1) );
  AND2X2 AND2X2_4827 ( .A(u2__abc_44228_n11635_1), .B(u2__abc_44228_n11633), .Y(u2__abc_44228_n11636) );
  AND2X2 AND2X2_4828 ( .A(u2__abc_44228_n7548_1_bF_buf50), .B(u2_remHi_237_), .Y(u2__abc_44228_n11637) );
  AND2X2 AND2X2_4829 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n4412), .Y(u2__abc_44228_n11640) );
  AND2X2 AND2X2_483 ( .A(u1__abc_43968_n313), .B(u1__abc_43968_n320), .Y(u1__abc_43968_n321) );
  AND2X2 AND2X2_4830 ( .A(u2__abc_44228_n11641_1), .B(u2__abc_44228_n2972_bF_buf82), .Y(u2__abc_44228_n11642_1) );
  AND2X2 AND2X2_4831 ( .A(u2__abc_44228_n11639), .B(u2__abc_44228_n11642_1), .Y(u2__abc_44228_n11643) );
  AND2X2 AND2X2_4832 ( .A(u2__abc_44228_n11644), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_remHi_239__FF_INPUT) );
  AND2X2 AND2X2_4833 ( .A(u2__abc_44228_n3062_bF_buf38), .B(u2_remHi_240_), .Y(u2__abc_44228_n11646) );
  AND2X2 AND2X2_4834 ( .A(u2__abc_44228_n11373), .B(u2__abc_44228_n4538), .Y(u2__abc_44228_n11647) );
  AND2X2 AND2X2_4835 ( .A(u2__abc_44228_n11648_1), .B(u2__abc_44228_n4408), .Y(u2__abc_44228_n11649_1) );
  AND2X2 AND2X2_4836 ( .A(u2__abc_44228_n11650), .B(u2__abc_44228_n11651), .Y(u2__abc_44228_n11652) );
  AND2X2 AND2X2_4837 ( .A(u2__abc_44228_n11653), .B(u2__abc_44228_n11654), .Y(u2__abc_44228_n11655_1) );
  AND2X2 AND2X2_4838 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n4398), .Y(u2__abc_44228_n11657) );
  AND2X2 AND2X2_4839 ( .A(u2__abc_44228_n11658), .B(u2__abc_44228_n2972_bF_buf81), .Y(u2__abc_44228_n11659) );
  AND2X2 AND2X2_484 ( .A(u1__abc_43968_n306), .B(u1__abc_43968_n321), .Y(u1__abc_43968_n322) );
  AND2X2 AND2X2_4840 ( .A(u2__abc_44228_n11656_1), .B(u2__abc_44228_n11659), .Y(u2__abc_44228_n11660) );
  AND2X2 AND2X2_4841 ( .A(u2__abc_44228_n11661), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_remHi_240__FF_INPUT) );
  AND2X2 AND2X2_4842 ( .A(u2__abc_44228_n3062_bF_buf37), .B(u2_remHi_241_), .Y(u2__abc_44228_n11663_1) );
  AND2X2 AND2X2_4843 ( .A(u2__abc_44228_n11650), .B(u2__abc_44228_n5549_1), .Y(u2__abc_44228_n11665) );
  AND2X2 AND2X2_4844 ( .A(u2__abc_44228_n11668), .B(u2__abc_44228_n11666), .Y(u2__abc_44228_n11669_1) );
  AND2X2 AND2X2_4845 ( .A(u2__abc_44228_n11669_1), .B(u2__abc_44228_n7547_bF_buf47), .Y(u2__abc_44228_n11670) );
  AND2X2 AND2X2_4846 ( .A(u2__abc_44228_n7548_1_bF_buf48), .B(u2_remHi_239_), .Y(u2__abc_44228_n11671) );
  AND2X2 AND2X2_4847 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n4392), .Y(u2__abc_44228_n11674_1) );
  AND2X2 AND2X2_4848 ( .A(u2__abc_44228_n11675), .B(u2__abc_44228_n2972_bF_buf80), .Y(u2__abc_44228_n11676) );
  AND2X2 AND2X2_4849 ( .A(u2__abc_44228_n11673), .B(u2__abc_44228_n11676), .Y(u2__abc_44228_n11677) );
  AND2X2 AND2X2_485 ( .A(u1__abc_43968_n291), .B(u1__abc_43968_n322), .Y(u1__abc_43968_n323) );
  AND2X2 AND2X2_4850 ( .A(u2__abc_44228_n11678), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_remHi_241__FF_INPUT) );
  AND2X2 AND2X2_4851 ( .A(u2__abc_44228_n3062_bF_buf36), .B(u2_remHi_242_), .Y(u2__abc_44228_n11680) );
  AND2X2 AND2X2_4852 ( .A(u2__abc_44228_n11650), .B(u2__abc_44228_n5550), .Y(u2__abc_44228_n11681) );
  AND2X2 AND2X2_4853 ( .A(u2__abc_44228_n11683), .B(u2__abc_44228_n4401), .Y(u2__abc_44228_n11685) );
  AND2X2 AND2X2_4854 ( .A(u2__abc_44228_n11686), .B(u2__abc_44228_n11684_1), .Y(u2__abc_44228_n11687) );
  AND2X2 AND2X2_4855 ( .A(u2__abc_44228_n11687), .B(u2__abc_44228_n7547_bF_buf46), .Y(u2__abc_44228_n11688) );
  AND2X2 AND2X2_4856 ( .A(u2__abc_44228_n7548_1_bF_buf47), .B(u2_remHi_240_), .Y(u2__abc_44228_n11689) );
  AND2X2 AND2X2_4857 ( .A(u2__abc_44228_n2983_bF_buf113), .B(u2__abc_44228_n4376), .Y(u2__abc_44228_n11692) );
  AND2X2 AND2X2_4858 ( .A(u2__abc_44228_n11693), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n11694) );
  AND2X2 AND2X2_4859 ( .A(u2__abc_44228_n11691), .B(u2__abc_44228_n11694), .Y(u2__abc_44228_n11695) );
  AND2X2 AND2X2_486 ( .A(u1__abc_43968_n324), .B(u1__abc_43968_n325), .Y(u1__abc_43968_n326) );
  AND2X2 AND2X2_4860 ( .A(u2__abc_44228_n11696), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_remHi_242__FF_INPUT) );
  AND2X2 AND2X2_4861 ( .A(u2__abc_44228_n3062_bF_buf35), .B(u2_remHi_243_), .Y(u2__abc_44228_n11698) );
  AND2X2 AND2X2_4862 ( .A(u2__abc_44228_n11703), .B(u2__abc_44228_n7547_bF_buf45), .Y(u2__abc_44228_n11704_1) );
  AND2X2 AND2X2_4863 ( .A(u2__abc_44228_n11704_1), .B(u2__abc_44228_n11702), .Y(u2__abc_44228_n11705) );
  AND2X2 AND2X2_4864 ( .A(u2__abc_44228_n7548_1_bF_buf46), .B(u2_remHi_241_), .Y(u2__abc_44228_n11706) );
  AND2X2 AND2X2_4865 ( .A(u2__abc_44228_n2983_bF_buf111), .B(u2__abc_44228_n4383), .Y(u2__abc_44228_n11709) );
  AND2X2 AND2X2_4866 ( .A(u2__abc_44228_n11710), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n11711_1) );
  AND2X2 AND2X2_4867 ( .A(u2__abc_44228_n11708), .B(u2__abc_44228_n11711_1), .Y(u2__abc_44228_n11712) );
  AND2X2 AND2X2_4868 ( .A(u2__abc_44228_n11713), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_remHi_243__FF_INPUT) );
  AND2X2 AND2X2_4869 ( .A(u2__abc_44228_n3062_bF_buf34), .B(u2_remHi_244_), .Y(u2__abc_44228_n11715) );
  AND2X2 AND2X2_487 ( .A(u1__abc_43968_n327), .B(u1__abc_43968_n328), .Y(u1__abc_43968_n329) );
  AND2X2 AND2X2_4870 ( .A(u2__abc_44228_n11648_1), .B(u2__abc_44228_n4417), .Y(u2__abc_44228_n11716) );
  AND2X2 AND2X2_4871 ( .A(u2__abc_44228_n11717), .B(u2__abc_44228_n4379), .Y(u2__abc_44228_n11718) );
  AND2X2 AND2X2_4872 ( .A(u2__abc_44228_n11719_1), .B(u2__abc_44228_n11720), .Y(u2__abc_44228_n11721) );
  AND2X2 AND2X2_4873 ( .A(u2__abc_44228_n11721), .B(u2__abc_44228_n7547_bF_buf44), .Y(u2__abc_44228_n11722) );
  AND2X2 AND2X2_4874 ( .A(u2__abc_44228_n7548_1_bF_buf45), .B(u2_remHi_242_), .Y(u2__abc_44228_n11723) );
  AND2X2 AND2X2_4875 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n4369), .Y(u2__abc_44228_n11726_1) );
  AND2X2 AND2X2_4876 ( .A(u2__abc_44228_n11727), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n11728) );
  AND2X2 AND2X2_4877 ( .A(u2__abc_44228_n11725), .B(u2__abc_44228_n11728), .Y(u2__abc_44228_n11729) );
  AND2X2 AND2X2_4878 ( .A(u2__abc_44228_n11730), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_remHi_244__FF_INPUT) );
  AND2X2 AND2X2_4879 ( .A(u2__abc_44228_n3062_bF_buf33), .B(u2_remHi_245_), .Y(u2__abc_44228_n11732) );
  AND2X2 AND2X2_488 ( .A(u1__abc_43968_n326), .B(u1__abc_43968_n329), .Y(u1__abc_43968_n330) );
  AND2X2 AND2X2_4880 ( .A(u2__abc_44228_n11719_1), .B(u2__abc_44228_n5558_1), .Y(u2__abc_44228_n11733) );
  AND2X2 AND2X2_4881 ( .A(u2__abc_44228_n11737), .B(u2__abc_44228_n7547_bF_buf43), .Y(u2__abc_44228_n11738) );
  AND2X2 AND2X2_4882 ( .A(u2__abc_44228_n11738), .B(u2__abc_44228_n11735), .Y(u2__abc_44228_n11739) );
  AND2X2 AND2X2_4883 ( .A(u2__abc_44228_n7548_1_bF_buf44), .B(u2_remHi_243_), .Y(u2__abc_44228_n11740) );
  AND2X2 AND2X2_4884 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n4363), .Y(u2__abc_44228_n11743) );
  AND2X2 AND2X2_4885 ( .A(u2__abc_44228_n11744), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n11745) );
  AND2X2 AND2X2_4886 ( .A(u2__abc_44228_n11742), .B(u2__abc_44228_n11745), .Y(u2__abc_44228_n11746) );
  AND2X2 AND2X2_4887 ( .A(u2__abc_44228_n11747), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_remHi_245__FF_INPUT) );
  AND2X2 AND2X2_4888 ( .A(u2__abc_44228_n3062_bF_buf32), .B(u2_remHi_246_), .Y(u2__abc_44228_n11749) );
  AND2X2 AND2X2_4889 ( .A(u2__abc_44228_n11719_1), .B(u2__abc_44228_n5559), .Y(u2__abc_44228_n11750_1) );
  AND2X2 AND2X2_489 ( .A(u1__abc_43968_n331), .B(u1__abc_43968_n332), .Y(u1__abc_43968_n333) );
  AND2X2 AND2X2_4890 ( .A(u2__abc_44228_n11752), .B(u2__abc_44228_n4372), .Y(u2__abc_44228_n11754) );
  AND2X2 AND2X2_4891 ( .A(u2__abc_44228_n11755), .B(u2__abc_44228_n11753), .Y(u2__abc_44228_n11756) );
  AND2X2 AND2X2_4892 ( .A(u2__abc_44228_n11756), .B(u2__abc_44228_n7547_bF_buf42), .Y(u2__abc_44228_n11757_1) );
  AND2X2 AND2X2_4893 ( .A(u2__abc_44228_n7548_1_bF_buf43), .B(u2_remHi_244_), .Y(u2__abc_44228_n11758) );
  AND2X2 AND2X2_4894 ( .A(u2__abc_44228_n2983_bF_buf107), .B(u2__abc_44228_n4346), .Y(u2__abc_44228_n11761) );
  AND2X2 AND2X2_4895 ( .A(u2__abc_44228_n11762), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n11763) );
  AND2X2 AND2X2_4896 ( .A(u2__abc_44228_n11760), .B(u2__abc_44228_n11763), .Y(u2__abc_44228_n11764) );
  AND2X2 AND2X2_4897 ( .A(u2__abc_44228_n11765_1), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_remHi_246__FF_INPUT) );
  AND2X2 AND2X2_4898 ( .A(u2__abc_44228_n3062_bF_buf31), .B(u2_remHi_247_), .Y(u2__abc_44228_n11767) );
  AND2X2 AND2X2_4899 ( .A(u2__abc_44228_n11772_1), .B(u2__abc_44228_n7547_bF_buf41), .Y(u2__abc_44228_n11773) );
  AND2X2 AND2X2_49 ( .A(_abc_64468_n753_bF_buf7), .B(sqrto_48_), .Y(_auto_iopadmap_cc_313_execute_65414_84_) );
  AND2X2 AND2X2_490 ( .A(u1__abc_43968_n334), .B(u1__abc_43968_n335), .Y(u1__abc_43968_n336) );
  AND2X2 AND2X2_4900 ( .A(u2__abc_44228_n11773), .B(u2__abc_44228_n11771), .Y(u2__abc_44228_n11774) );
  AND2X2 AND2X2_4901 ( .A(u2__abc_44228_n7548_1_bF_buf42), .B(u2_remHi_245_), .Y(u2__abc_44228_n11775) );
  AND2X2 AND2X2_4902 ( .A(u2__abc_44228_n2983_bF_buf105), .B(u2__abc_44228_n4353), .Y(u2__abc_44228_n11778) );
  AND2X2 AND2X2_4903 ( .A(u2__abc_44228_n11779), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n11780) );
  AND2X2 AND2X2_4904 ( .A(u2__abc_44228_n11777), .B(u2__abc_44228_n11780), .Y(u2__abc_44228_n11781_1) );
  AND2X2 AND2X2_4905 ( .A(u2__abc_44228_n11782), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_remHi_247__FF_INPUT) );
  AND2X2 AND2X2_4906 ( .A(u2__abc_44228_n3062_bF_buf30), .B(u2_remHi_248_), .Y(u2__abc_44228_n11784) );
  AND2X2 AND2X2_4907 ( .A(u2__abc_44228_n11648_1), .B(u2__abc_44228_n4418), .Y(u2__abc_44228_n11785) );
  AND2X2 AND2X2_4908 ( .A(u2__abc_44228_n11786), .B(u2__abc_44228_n4349_1), .Y(u2__abc_44228_n11788_1) );
  AND2X2 AND2X2_4909 ( .A(u2__abc_44228_n11789), .B(u2__abc_44228_n11787), .Y(u2__abc_44228_n11790) );
  AND2X2 AND2X2_491 ( .A(u1__abc_43968_n333), .B(u1__abc_43968_n336), .Y(u1__abc_43968_n337) );
  AND2X2 AND2X2_4910 ( .A(u2__abc_44228_n11790), .B(u2__abc_44228_n7547_bF_buf40), .Y(u2__abc_44228_n11791) );
  AND2X2 AND2X2_4911 ( .A(u2__abc_44228_n7548_1_bF_buf41), .B(u2_remHi_246_), .Y(u2__abc_44228_n11792) );
  AND2X2 AND2X2_4912 ( .A(u2__abc_44228_n2983_bF_buf104), .B(u2__abc_44228_n4339), .Y(u2__abc_44228_n11795) );
  AND2X2 AND2X2_4913 ( .A(u2__abc_44228_n11796_1), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n11797) );
  AND2X2 AND2X2_4914 ( .A(u2__abc_44228_n11794), .B(u2__abc_44228_n11797), .Y(u2__abc_44228_n11798) );
  AND2X2 AND2X2_4915 ( .A(u2__abc_44228_n11799), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_remHi_248__FF_INPUT) );
  AND2X2 AND2X2_4916 ( .A(u2__abc_44228_n3062_bF_buf29), .B(u2_remHi_249_), .Y(u2__abc_44228_n11801) );
  AND2X2 AND2X2_4917 ( .A(u2__abc_44228_n11789), .B(u2__abc_44228_n5531_1), .Y(u2__abc_44228_n11802) );
  AND2X2 AND2X2_4918 ( .A(u2__abc_44228_n11802), .B(u2__abc_44228_n4356), .Y(u2__abc_44228_n11803_1) );
  AND2X2 AND2X2_4919 ( .A(u2__abc_44228_n11805), .B(u2__abc_44228_n11804), .Y(u2__abc_44228_n11806) );
  AND2X2 AND2X2_492 ( .A(u1__abc_43968_n330), .B(u1__abc_43968_n337), .Y(u1__abc_43968_n338) );
  AND2X2 AND2X2_4920 ( .A(u2__abc_44228_n11807), .B(u2__abc_44228_n7547_bF_buf39), .Y(u2__abc_44228_n11808) );
  AND2X2 AND2X2_4921 ( .A(u2__abc_44228_n7548_1_bF_buf40), .B(u2_remHi_247_), .Y(u2__abc_44228_n11809) );
  AND2X2 AND2X2_4922 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n4333), .Y(u2__abc_44228_n11812) );
  AND2X2 AND2X2_4923 ( .A(u2__abc_44228_n11813_1), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n11814) );
  AND2X2 AND2X2_4924 ( .A(u2__abc_44228_n11811), .B(u2__abc_44228_n11814), .Y(u2__abc_44228_n11815) );
  AND2X2 AND2X2_4925 ( .A(u2__abc_44228_n11816), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_remHi_249__FF_INPUT) );
  AND2X2 AND2X2_4926 ( .A(u2__abc_44228_n3062_bF_buf28), .B(u2_remHi_250_), .Y(u2__abc_44228_n11818) );
  AND2X2 AND2X2_4927 ( .A(u2__abc_44228_n11789), .B(u2__abc_44228_n5532), .Y(u2__abc_44228_n11819) );
  AND2X2 AND2X2_4928 ( .A(u2__abc_44228_n11821), .B(u2__abc_44228_n4342), .Y(u2__abc_44228_n11823) );
  AND2X2 AND2X2_4929 ( .A(u2__abc_44228_n11824), .B(u2__abc_44228_n11822), .Y(u2__abc_44228_n11825) );
  AND2X2 AND2X2_493 ( .A(u1__abc_43968_n339), .B(u1__abc_43968_n340), .Y(u1__abc_43968_n341) );
  AND2X2 AND2X2_4930 ( .A(u2__abc_44228_n11825), .B(u2__abc_44228_n7547_bF_buf38), .Y(u2__abc_44228_n11826) );
  AND2X2 AND2X2_4931 ( .A(u2__abc_44228_n7548_1_bF_buf39), .B(u2_remHi_248_), .Y(u2__abc_44228_n11827) );
  AND2X2 AND2X2_4932 ( .A(u2__abc_44228_n2983_bF_buf101), .B(u2__abc_44228_n4317), .Y(u2__abc_44228_n11830) );
  AND2X2 AND2X2_4933 ( .A(u2__abc_44228_n11831), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n11832) );
  AND2X2 AND2X2_4934 ( .A(u2__abc_44228_n11829), .B(u2__abc_44228_n11832), .Y(u2__abc_44228_n11833) );
  AND2X2 AND2X2_4935 ( .A(u2__abc_44228_n11834), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_remHi_250__FF_INPUT) );
  AND2X2 AND2X2_4936 ( .A(u2__abc_44228_n3062_bF_buf27), .B(u2_remHi_251_), .Y(u2__abc_44228_n11836) );
  AND2X2 AND2X2_4937 ( .A(u2__abc_44228_n11841), .B(u2__abc_44228_n7547_bF_buf37), .Y(u2__abc_44228_n11842) );
  AND2X2 AND2X2_4938 ( .A(u2__abc_44228_n11842), .B(u2__abc_44228_n11840), .Y(u2__abc_44228_n11843) );
  AND2X2 AND2X2_4939 ( .A(u2__abc_44228_n7548_1_bF_buf38), .B(u2_remHi_249_), .Y(u2__abc_44228_n11844_1) );
  AND2X2 AND2X2_494 ( .A(u1__abc_43968_n342), .B(u1__abc_43968_n343), .Y(u1__abc_43968_n344) );
  AND2X2 AND2X2_4940 ( .A(u2__abc_44228_n2983_bF_buf99), .B(u2__abc_44228_n4324), .Y(u2__abc_44228_n11847) );
  AND2X2 AND2X2_4941 ( .A(u2__abc_44228_n11848), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n11849) );
  AND2X2 AND2X2_4942 ( .A(u2__abc_44228_n11846), .B(u2__abc_44228_n11849), .Y(u2__abc_44228_n11850) );
  AND2X2 AND2X2_4943 ( .A(u2__abc_44228_n11851_1), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_remHi_251__FF_INPUT) );
  AND2X2 AND2X2_4944 ( .A(u2__abc_44228_n3062_bF_buf26), .B(u2_remHi_252_), .Y(u2__abc_44228_n11853) );
  AND2X2 AND2X2_4945 ( .A(u2__abc_44228_n11786), .B(u2__abc_44228_n4358), .Y(u2__abc_44228_n11854) );
  AND2X2 AND2X2_4946 ( .A(u2__abc_44228_n11855), .B(u2__abc_44228_n4320_1), .Y(u2__abc_44228_n11856) );
  AND2X2 AND2X2_4947 ( .A(u2__abc_44228_n11857), .B(u2__abc_44228_n11858), .Y(u2__abc_44228_n11859_1) );
  AND2X2 AND2X2_4948 ( .A(u2__abc_44228_n11859_1), .B(u2__abc_44228_n7547_bF_buf36), .Y(u2__abc_44228_n11860) );
  AND2X2 AND2X2_4949 ( .A(u2__abc_44228_n7548_1_bF_buf37), .B(u2_remHi_250_), .Y(u2__abc_44228_n11861) );
  AND2X2 AND2X2_495 ( .A(u1__abc_43968_n341), .B(u1__abc_43968_n344), .Y(u1__abc_43968_n345) );
  AND2X2 AND2X2_4950 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n4310_1), .Y(u2__abc_44228_n11864) );
  AND2X2 AND2X2_4951 ( .A(u2__abc_44228_n11865), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n11866_1) );
  AND2X2 AND2X2_4952 ( .A(u2__abc_44228_n11863), .B(u2__abc_44228_n11866_1), .Y(u2__abc_44228_n11867) );
  AND2X2 AND2X2_4953 ( .A(u2__abc_44228_n11868), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_remHi_252__FF_INPUT) );
  AND2X2 AND2X2_4954 ( .A(u2__abc_44228_n3062_bF_buf25), .B(u2_remHi_253_), .Y(u2__abc_44228_n11870) );
  AND2X2 AND2X2_4955 ( .A(u2__abc_44228_n11857), .B(u2__abc_44228_n5542), .Y(u2__abc_44228_n11871) );
  AND2X2 AND2X2_4956 ( .A(u2__abc_44228_n11871), .B(u2__abc_44228_n4327), .Y(u2__abc_44228_n11872) );
  AND2X2 AND2X2_4957 ( .A(u2__abc_44228_n11874), .B(u2__abc_44228_n11873), .Y(u2__abc_44228_n11875) );
  AND2X2 AND2X2_4958 ( .A(u2__abc_44228_n11876_1), .B(u2__abc_44228_n7547_bF_buf35), .Y(u2__abc_44228_n11877) );
  AND2X2 AND2X2_4959 ( .A(u2__abc_44228_n7548_1_bF_buf36), .B(u2_remHi_251_), .Y(u2__abc_44228_n11878) );
  AND2X2 AND2X2_496 ( .A(u1__abc_43968_n346), .B(u1__abc_43968_n347), .Y(u1__abc_43968_n348) );
  AND2X2 AND2X2_4960 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n4304), .Y(u2__abc_44228_n11881) );
  AND2X2 AND2X2_4961 ( .A(u2__abc_44228_n11882), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n11883_1) );
  AND2X2 AND2X2_4962 ( .A(u2__abc_44228_n11880), .B(u2__abc_44228_n11883_1), .Y(u2__abc_44228_n11884) );
  AND2X2 AND2X2_4963 ( .A(u2__abc_44228_n11885), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_remHi_253__FF_INPUT) );
  AND2X2 AND2X2_4964 ( .A(u2__abc_44228_n3062_bF_buf24), .B(u2_remHi_254_), .Y(u2__abc_44228_n11887) );
  AND2X2 AND2X2_4965 ( .A(u2__abc_44228_n11857), .B(u2__abc_44228_n5543), .Y(u2__abc_44228_n11888) );
  AND2X2 AND2X2_4966 ( .A(u2__abc_44228_n11890), .B(u2__abc_44228_n4313), .Y(u2__abc_44228_n11892) );
  AND2X2 AND2X2_4967 ( .A(u2__abc_44228_n11893), .B(u2__abc_44228_n11891_1), .Y(u2__abc_44228_n11894) );
  AND2X2 AND2X2_4968 ( .A(u2__abc_44228_n11894), .B(u2__abc_44228_n7547_bF_buf34), .Y(u2__abc_44228_n11895) );
  AND2X2 AND2X2_4969 ( .A(u2__abc_44228_n7548_1_bF_buf35), .B(u2_remHi_252_), .Y(u2__abc_44228_n11896) );
  AND2X2 AND2X2_497 ( .A(u1__abc_43968_n349), .B(u1__abc_43968_n350), .Y(u1__abc_43968_n351) );
  AND2X2 AND2X2_4970 ( .A(u2__abc_44228_n2983_bF_buf95), .B(u2__abc_44228_n6521), .Y(u2__abc_44228_n11899) );
  AND2X2 AND2X2_4971 ( .A(u2__abc_44228_n11900), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n11901) );
  AND2X2 AND2X2_4972 ( .A(u2__abc_44228_n11898_1), .B(u2__abc_44228_n11901), .Y(u2__abc_44228_n11902) );
  AND2X2 AND2X2_4973 ( .A(u2__abc_44228_n11903), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_remHi_254__FF_INPUT) );
  AND2X2 AND2X2_4974 ( .A(u2__abc_44228_n3062_bF_buf23), .B(u2_remHi_255_), .Y(u2__abc_44228_n11905) );
  AND2X2 AND2X2_4975 ( .A(u2__abc_44228_n11910), .B(u2__abc_44228_n7547_bF_buf33), .Y(u2__abc_44228_n11911) );
  AND2X2 AND2X2_4976 ( .A(u2__abc_44228_n11911), .B(u2__abc_44228_n11909), .Y(u2__abc_44228_n11912) );
  AND2X2 AND2X2_4977 ( .A(u2__abc_44228_n7548_1_bF_buf34), .B(u2_remHi_253_), .Y(u2__abc_44228_n11913) );
  AND2X2 AND2X2_4978 ( .A(u2__abc_44228_n2983_bF_buf93), .B(u2__abc_44228_n6515), .Y(u2__abc_44228_n11916) );
  AND2X2 AND2X2_4979 ( .A(u2__abc_44228_n11917), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n11918) );
  AND2X2 AND2X2_498 ( .A(u1__abc_43968_n348), .B(u1__abc_43968_n351), .Y(u1__abc_43968_n352) );
  AND2X2 AND2X2_4980 ( .A(u2__abc_44228_n11915), .B(u2__abc_44228_n11918), .Y(u2__abc_44228_n11919) );
  AND2X2 AND2X2_4981 ( .A(u2__abc_44228_n11920), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_remHi_255__FF_INPUT) );
  AND2X2 AND2X2_4982 ( .A(u2__abc_44228_n3062_bF_buf22), .B(u2_remHi_256_), .Y(u2__abc_44228_n11922_1) );
  AND2X2 AND2X2_4983 ( .A(u2__abc_44228_n7548_1_bF_buf33), .B(u2_remHi_254_), .Y(u2__abc_44228_n11923) );
  AND2X2 AND2X2_4984 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6524), .Y(u2__abc_44228_n11925) );
  AND2X2 AND2X2_4985 ( .A(u2__abc_44228_n11926), .B(u2__abc_44228_n11924), .Y(u2__abc_44228_n11927) );
  AND2X2 AND2X2_4986 ( .A(u2__abc_44228_n7547_bF_buf32), .B(u2__abc_44228_n11927), .Y(u2__abc_44228_n11928) );
  AND2X2 AND2X2_4987 ( .A(u2__abc_44228_n2983_bF_buf91), .B(u2__abc_44228_n6507_1), .Y(u2__abc_44228_n11931) );
  AND2X2 AND2X2_4988 ( .A(u2__abc_44228_n11932), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n11933) );
  AND2X2 AND2X2_4989 ( .A(u2__abc_44228_n11930), .B(u2__abc_44228_n11933), .Y(u2__abc_44228_n11934) );
  AND2X2 AND2X2_499 ( .A(u1__abc_43968_n345), .B(u1__abc_43968_n352), .Y(u1__abc_43968_n353) );
  AND2X2 AND2X2_4990 ( .A(u2__abc_44228_n11935), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_remHi_256__FF_INPUT) );
  AND2X2 AND2X2_4991 ( .A(u2__abc_44228_n3062_bF_buf21), .B(u2_remHi_257_), .Y(u2__abc_44228_n11937) );
  AND2X2 AND2X2_4992 ( .A(u2__abc_44228_n7548_1_bF_buf32), .B(u2_remHi_255_), .Y(u2__abc_44228_n11938) );
  AND2X2 AND2X2_4993 ( .A(u2__abc_44228_n11926), .B(u2__abc_44228_n6533), .Y(u2__abc_44228_n11940_1) );
  AND2X2 AND2X2_4994 ( .A(u2__abc_44228_n11941), .B(u2__abc_44228_n11939), .Y(u2__abc_44228_n11942) );
  AND2X2 AND2X2_4995 ( .A(u2__abc_44228_n11940_1), .B(u2__abc_44228_n6518), .Y(u2__abc_44228_n11943) );
  AND2X2 AND2X2_4996 ( .A(u2__abc_44228_n7547_bF_buf31), .B(u2__abc_44228_n11944), .Y(u2__abc_44228_n11945) );
  AND2X2 AND2X2_4997 ( .A(u2__abc_44228_n2983_bF_buf89), .B(u2__abc_44228_n6501), .Y(u2__abc_44228_n11948) );
  AND2X2 AND2X2_4998 ( .A(u2__abc_44228_n11949), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n11950) );
  AND2X2 AND2X2_4999 ( .A(u2__abc_44228_n11947_1), .B(u2__abc_44228_n11950), .Y(u2__abc_44228_n11951) );
  AND2X2 AND2X2_5 ( .A(_abc_64468_n753_bF_buf9), .B(sqrto_4_), .Y(_auto_iopadmap_cc_313_execute_65414_40_) );
  AND2X2 AND2X2_50 ( .A(_abc_64468_n753_bF_buf6), .B(sqrto_49_), .Y(_auto_iopadmap_cc_313_execute_65414_85_) );
  AND2X2 AND2X2_500 ( .A(u1__abc_43968_n338), .B(u1__abc_43968_n353), .Y(u1__abc_43968_n354) );
  AND2X2 AND2X2_5000 ( .A(u2__abc_44228_n11952), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_remHi_257__FF_INPUT) );
  AND2X2 AND2X2_5001 ( .A(u2__abc_44228_n3062_bF_buf20), .B(u2_remHi_258_), .Y(u2__abc_44228_n11954) );
  AND2X2 AND2X2_5002 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6525_1), .Y(u2__abc_44228_n11955_1) );
  AND2X2 AND2X2_5003 ( .A(u2__abc_44228_n11956), .B(u2__abc_44228_n6510), .Y(u2__abc_44228_n11957) );
  AND2X2 AND2X2_5004 ( .A(u2__abc_44228_n11958), .B(u2__abc_44228_n11959), .Y(u2__abc_44228_n11960) );
  AND2X2 AND2X2_5005 ( .A(u2__abc_44228_n11961), .B(u2__abc_44228_n11962_1), .Y(u2__abc_44228_n11963) );
  AND2X2 AND2X2_5006 ( .A(u2__abc_44228_n2983_bF_buf87), .B(u2__abc_44228_n6492), .Y(u2__abc_44228_n11965) );
  AND2X2 AND2X2_5007 ( .A(u2__abc_44228_n11966), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n11967) );
  AND2X2 AND2X2_5008 ( .A(u2__abc_44228_n11964), .B(u2__abc_44228_n11967), .Y(u2__abc_44228_n11968) );
  AND2X2 AND2X2_5009 ( .A(u2__abc_44228_n11969), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_remHi_258__FF_INPUT) );
  AND2X2 AND2X2_501 ( .A(u1__abc_43968_n355), .B(u1__abc_43968_n356), .Y(u1__abc_43968_n357) );
  AND2X2 AND2X2_5010 ( .A(u2__abc_44228_n3062_bF_buf19), .B(u2_remHi_259_), .Y(u2__abc_44228_n11971_1) );
  AND2X2 AND2X2_5011 ( .A(u2__abc_44228_n11976), .B(u2__abc_44228_n11973), .Y(u2__abc_44228_n11977) );
  AND2X2 AND2X2_5012 ( .A(u2__abc_44228_n11977), .B(u2__abc_44228_n7547_bF_buf29), .Y(u2__abc_44228_n11978_1) );
  AND2X2 AND2X2_5013 ( .A(u2__abc_44228_n7548_1_bF_buf30), .B(u2_remHi_257_), .Y(u2__abc_44228_n11979) );
  AND2X2 AND2X2_5014 ( .A(u2__abc_44228_n2983_bF_buf85), .B(u2__abc_44228_n6486), .Y(u2__abc_44228_n11982) );
  AND2X2 AND2X2_5015 ( .A(u2__abc_44228_n11983), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n11984) );
  AND2X2 AND2X2_5016 ( .A(u2__abc_44228_n11981), .B(u2__abc_44228_n11984), .Y(u2__abc_44228_n11985) );
  AND2X2 AND2X2_5017 ( .A(u2__abc_44228_n11986_1), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_remHi_259__FF_INPUT) );
  AND2X2 AND2X2_5018 ( .A(u2__abc_44228_n3062_bF_buf18), .B(u2_remHi_260_), .Y(u2__abc_44228_n11988) );
  AND2X2 AND2X2_5019 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6526), .Y(u2__abc_44228_n11989) );
  AND2X2 AND2X2_502 ( .A(u1__abc_43968_n358), .B(u1__abc_43968_n359), .Y(u1__abc_43968_n360) );
  AND2X2 AND2X2_5020 ( .A(u2__abc_44228_n11990), .B(u2__abc_44228_n6495), .Y(u2__abc_44228_n11992) );
  AND2X2 AND2X2_5021 ( .A(u2__abc_44228_n11993_1), .B(u2__abc_44228_n11991), .Y(u2__abc_44228_n11994) );
  AND2X2 AND2X2_5022 ( .A(u2__abc_44228_n11995), .B(u2__abc_44228_n11996), .Y(u2__abc_44228_n11997) );
  AND2X2 AND2X2_5023 ( .A(u2__abc_44228_n2983_bF_buf83), .B(u2__abc_44228_n6478), .Y(u2__abc_44228_n11999) );
  AND2X2 AND2X2_5024 ( .A(u2__abc_44228_n12000), .B(u2__abc_44228_n2972_bF_buf61), .Y(u2__abc_44228_n12001) );
  AND2X2 AND2X2_5025 ( .A(u2__abc_44228_n11998), .B(u2__abc_44228_n12001), .Y(u2__abc_44228_n12002) );
  AND2X2 AND2X2_5026 ( .A(u2__abc_44228_n12003_1), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_remHi_260__FF_INPUT) );
  AND2X2 AND2X2_5027 ( .A(u2__abc_44228_n3062_bF_buf17), .B(u2_remHi_261_), .Y(u2__abc_44228_n12005) );
  AND2X2 AND2X2_5028 ( .A(u2__abc_44228_n11993_1), .B(u2__abc_44228_n6542), .Y(u2__abc_44228_n12007) );
  AND2X2 AND2X2_5029 ( .A(u2__abc_44228_n12010_1), .B(u2__abc_44228_n12008), .Y(u2__abc_44228_n12011) );
  AND2X2 AND2X2_503 ( .A(u1__abc_43968_n357), .B(u1__abc_43968_n360), .Y(u1__abc_43968_n361) );
  AND2X2 AND2X2_5030 ( .A(u2__abc_44228_n12011), .B(u2__abc_44228_n7547_bF_buf27), .Y(u2__abc_44228_n12012) );
  AND2X2 AND2X2_5031 ( .A(u2__abc_44228_n7548_1_bF_buf28), .B(u2_remHi_259_), .Y(u2__abc_44228_n12013) );
  AND2X2 AND2X2_5032 ( .A(u2__abc_44228_n2983_bF_buf81), .B(u2__abc_44228_n6472), .Y(u2__abc_44228_n12016) );
  AND2X2 AND2X2_5033 ( .A(u2__abc_44228_n12017), .B(u2__abc_44228_n2972_bF_buf60), .Y(u2__abc_44228_n12018_1) );
  AND2X2 AND2X2_5034 ( .A(u2__abc_44228_n12015), .B(u2__abc_44228_n12018_1), .Y(u2__abc_44228_n12019) );
  AND2X2 AND2X2_5035 ( .A(u2__abc_44228_n12020), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_remHi_261__FF_INPUT) );
  AND2X2 AND2X2_5036 ( .A(u2__abc_44228_n3062_bF_buf16), .B(u2_remHi_262_), .Y(u2__abc_44228_n12022) );
  AND2X2 AND2X2_5037 ( .A(u2__abc_44228_n11990), .B(u2__abc_44228_n6496), .Y(u2__abc_44228_n12023) );
  AND2X2 AND2X2_5038 ( .A(u2__abc_44228_n12024), .B(u2__abc_44228_n6481), .Y(u2__abc_44228_n12025_1) );
  AND2X2 AND2X2_5039 ( .A(u2__abc_44228_n12026), .B(u2__abc_44228_n12027), .Y(u2__abc_44228_n12028) );
  AND2X2 AND2X2_504 ( .A(u1__abc_43968_n362), .B(u1__abc_43968_n363), .Y(u1__abc_43968_n364) );
  AND2X2 AND2X2_5040 ( .A(u2__abc_44228_n12029), .B(u2__abc_44228_n12030), .Y(u2__abc_44228_n12031) );
  AND2X2 AND2X2_5041 ( .A(u2__abc_44228_n2983_bF_buf79), .B(u2__abc_44228_n6462), .Y(u2__abc_44228_n12033) );
  AND2X2 AND2X2_5042 ( .A(u2__abc_44228_n12034_1), .B(u2__abc_44228_n2972_bF_buf59), .Y(u2__abc_44228_n12035) );
  AND2X2 AND2X2_5043 ( .A(u2__abc_44228_n12032), .B(u2__abc_44228_n12035), .Y(u2__abc_44228_n12036) );
  AND2X2 AND2X2_5044 ( .A(u2__abc_44228_n12037), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_remHi_262__FF_INPUT) );
  AND2X2 AND2X2_5045 ( .A(u2__abc_44228_n3062_bF_buf15), .B(u2_remHi_263_), .Y(u2__abc_44228_n12039) );
  AND2X2 AND2X2_5046 ( .A(u2__abc_44228_n12044), .B(u2__abc_44228_n7547_bF_buf25), .Y(u2__abc_44228_n12045) );
  AND2X2 AND2X2_5047 ( .A(u2__abc_44228_n12045), .B(u2__abc_44228_n12043), .Y(u2__abc_44228_n12046) );
  AND2X2 AND2X2_5048 ( .A(u2__abc_44228_n7548_1_bF_buf26), .B(u2_remHi_261_), .Y(u2__abc_44228_n12047) );
  AND2X2 AND2X2_5049 ( .A(u2__abc_44228_n2983_bF_buf77), .B(u2__abc_44228_n6456), .Y(u2__abc_44228_n12050) );
  AND2X2 AND2X2_505 ( .A(u1__abc_43968_n365), .B(u1__abc_43968_n366), .Y(u1__abc_43968_n367) );
  AND2X2 AND2X2_5050 ( .A(u2__abc_44228_n12051), .B(u2__abc_44228_n2972_bF_buf58), .Y(u2__abc_44228_n12052) );
  AND2X2 AND2X2_5051 ( .A(u2__abc_44228_n12049_1), .B(u2__abc_44228_n12052), .Y(u2__abc_44228_n12053) );
  AND2X2 AND2X2_5052 ( .A(u2__abc_44228_n12054), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_remHi_263__FF_INPUT) );
  AND2X2 AND2X2_5053 ( .A(u2__abc_44228_n3062_bF_buf14), .B(u2_remHi_264_), .Y(u2__abc_44228_n12056_1) );
  AND2X2 AND2X2_5054 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6527), .Y(u2__abc_44228_n12057) );
  AND2X2 AND2X2_5055 ( .A(u2__abc_44228_n12058), .B(u2__abc_44228_n6465), .Y(u2__abc_44228_n12059) );
  AND2X2 AND2X2_5056 ( .A(u2__abc_44228_n12060), .B(u2__abc_44228_n12061), .Y(u2__abc_44228_n12062) );
  AND2X2 AND2X2_5057 ( .A(u2__abc_44228_n12063), .B(u2__abc_44228_n12064), .Y(u2__abc_44228_n12065) );
  AND2X2 AND2X2_5058 ( .A(u2__abc_44228_n2983_bF_buf75), .B(u2__abc_44228_n6448), .Y(u2__abc_44228_n12067_1) );
  AND2X2 AND2X2_5059 ( .A(u2__abc_44228_n12068), .B(u2__abc_44228_n2972_bF_buf57), .Y(u2__abc_44228_n12069) );
  AND2X2 AND2X2_506 ( .A(u1__abc_43968_n364), .B(u1__abc_43968_n367), .Y(u1__abc_43968_n368) );
  AND2X2 AND2X2_5060 ( .A(u2__abc_44228_n12066), .B(u2__abc_44228_n12069), .Y(u2__abc_44228_n12070) );
  AND2X2 AND2X2_5061 ( .A(u2__abc_44228_n12071), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_remHi_264__FF_INPUT) );
  AND2X2 AND2X2_5062 ( .A(u2__abc_44228_n3062_bF_buf13), .B(u2_remHi_265_), .Y(u2__abc_44228_n12073) );
  AND2X2 AND2X2_5063 ( .A(u2__abc_44228_n12060), .B(u2__abc_44228_n6554), .Y(u2__abc_44228_n12075) );
  AND2X2 AND2X2_5064 ( .A(u2__abc_44228_n12078), .B(u2__abc_44228_n12076), .Y(u2__abc_44228_n12079) );
  AND2X2 AND2X2_5065 ( .A(u2__abc_44228_n12079), .B(u2__abc_44228_n7547_bF_buf23), .Y(u2__abc_44228_n12080) );
  AND2X2 AND2X2_5066 ( .A(u2__abc_44228_n7548_1_bF_buf24), .B(u2_remHi_263_), .Y(u2__abc_44228_n12081) );
  AND2X2 AND2X2_5067 ( .A(u2__abc_44228_n2983_bF_buf73), .B(u2__abc_44228_n6442), .Y(u2__abc_44228_n12084) );
  AND2X2 AND2X2_5068 ( .A(u2__abc_44228_n12085), .B(u2__abc_44228_n2972_bF_buf56), .Y(u2__abc_44228_n12086) );
  AND2X2 AND2X2_5069 ( .A(u2__abc_44228_n12083), .B(u2__abc_44228_n12086), .Y(u2__abc_44228_n12087) );
  AND2X2 AND2X2_507 ( .A(u1__abc_43968_n361), .B(u1__abc_43968_n368), .Y(u1__abc_43968_n369) );
  AND2X2 AND2X2_5070 ( .A(u2__abc_44228_n12088), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_remHi_265__FF_INPUT) );
  AND2X2 AND2X2_5071 ( .A(u2__abc_44228_n3062_bF_buf12), .B(u2_remHi_266_), .Y(u2__abc_44228_n12090) );
  AND2X2 AND2X2_5072 ( .A(u2__abc_44228_n12060), .B(u2__abc_44228_n6555), .Y(u2__abc_44228_n12091) );
  AND2X2 AND2X2_5073 ( .A(u2__abc_44228_n12093), .B(u2__abc_44228_n6451), .Y(u2__abc_44228_n12094) );
  AND2X2 AND2X2_5074 ( .A(u2__abc_44228_n12095), .B(u2__abc_44228_n12096), .Y(u2__abc_44228_n12097) );
  AND2X2 AND2X2_5075 ( .A(u2__abc_44228_n12097), .B(u2__abc_44228_n7547_bF_buf22), .Y(u2__abc_44228_n12098_1) );
  AND2X2 AND2X2_5076 ( .A(u2__abc_44228_n7548_1_bF_buf23), .B(u2_remHi_264_), .Y(u2__abc_44228_n12099) );
  AND2X2 AND2X2_5077 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n6433), .Y(u2__abc_44228_n12102) );
  AND2X2 AND2X2_5078 ( .A(u2__abc_44228_n12103), .B(u2__abc_44228_n2972_bF_buf55), .Y(u2__abc_44228_n12104) );
  AND2X2 AND2X2_5079 ( .A(u2__abc_44228_n12101), .B(u2__abc_44228_n12104), .Y(u2__abc_44228_n12105_1) );
  AND2X2 AND2X2_508 ( .A(u1__abc_43968_n370), .B(u1__abc_43968_n371), .Y(u1__abc_43968_n372) );
  AND2X2 AND2X2_5080 ( .A(u2__abc_44228_n12106), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_remHi_266__FF_INPUT) );
  AND2X2 AND2X2_5081 ( .A(u2__abc_44228_n3062_bF_buf11), .B(u2_remHi_267_), .Y(u2__abc_44228_n12108) );
  AND2X2 AND2X2_5082 ( .A(u2__abc_44228_n12113_1), .B(u2__abc_44228_n7547_bF_buf21), .Y(u2__abc_44228_n12114) );
  AND2X2 AND2X2_5083 ( .A(u2__abc_44228_n12114), .B(u2__abc_44228_n12112), .Y(u2__abc_44228_n12115) );
  AND2X2 AND2X2_5084 ( .A(u2__abc_44228_n7548_1_bF_buf22), .B(u2_remHi_265_), .Y(u2__abc_44228_n12116) );
  AND2X2 AND2X2_5085 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n6427), .Y(u2__abc_44228_n12119) );
  AND2X2 AND2X2_5086 ( .A(u2__abc_44228_n12120_1), .B(u2__abc_44228_n2972_bF_buf54), .Y(u2__abc_44228_n12121) );
  AND2X2 AND2X2_5087 ( .A(u2__abc_44228_n12118), .B(u2__abc_44228_n12121), .Y(u2__abc_44228_n12122) );
  AND2X2 AND2X2_5088 ( .A(u2__abc_44228_n12123), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_remHi_267__FF_INPUT) );
  AND2X2 AND2X2_5089 ( .A(u2__abc_44228_n3062_bF_buf10), .B(u2_remHi_268_), .Y(u2__abc_44228_n12125) );
  AND2X2 AND2X2_509 ( .A(u1__abc_43968_n373), .B(u1__abc_43968_n374), .Y(u1__abc_43968_n375) );
  AND2X2 AND2X2_5090 ( .A(u2__abc_44228_n12058), .B(u2__abc_44228_n6467), .Y(u2__abc_44228_n12126) );
  AND2X2 AND2X2_5091 ( .A(u2__abc_44228_n12127), .B(u2__abc_44228_n6436), .Y(u2__abc_44228_n12129) );
  AND2X2 AND2X2_5092 ( .A(u2__abc_44228_n12130_1), .B(u2__abc_44228_n12128), .Y(u2__abc_44228_n12131) );
  AND2X2 AND2X2_5093 ( .A(u2__abc_44228_n12132), .B(u2__abc_44228_n12133), .Y(u2__abc_44228_n12134) );
  AND2X2 AND2X2_5094 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n6419), .Y(u2__abc_44228_n12136) );
  AND2X2 AND2X2_5095 ( .A(u2__abc_44228_n12137_1), .B(u2__abc_44228_n2972_bF_buf53), .Y(u2__abc_44228_n12138) );
  AND2X2 AND2X2_5096 ( .A(u2__abc_44228_n12135), .B(u2__abc_44228_n12138), .Y(u2__abc_44228_n12139) );
  AND2X2 AND2X2_5097 ( .A(u2__abc_44228_n12140), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_remHi_268__FF_INPUT) );
  AND2X2 AND2X2_5098 ( .A(u2__abc_44228_n3062_bF_buf9), .B(u2_remHi_269_), .Y(u2__abc_44228_n12142) );
  AND2X2 AND2X2_5099 ( .A(u2__abc_44228_n12130_1), .B(u2__abc_44228_n6561_1), .Y(u2__abc_44228_n12144) );
  AND2X2 AND2X2_51 ( .A(_abc_64468_n753_bF_buf5), .B(sqrto_50_), .Y(_auto_iopadmap_cc_313_execute_65414_86_) );
  AND2X2 AND2X2_510 ( .A(u1__abc_43968_n372), .B(u1__abc_43968_n375), .Y(u1__abc_43968_n376) );
  AND2X2 AND2X2_5100 ( .A(u2__abc_44228_n12147), .B(u2__abc_44228_n12145_1), .Y(u2__abc_44228_n12148) );
  AND2X2 AND2X2_5101 ( .A(u2__abc_44228_n12148), .B(u2__abc_44228_n7547_bF_buf19), .Y(u2__abc_44228_n12149) );
  AND2X2 AND2X2_5102 ( .A(u2__abc_44228_n7548_1_bF_buf20), .B(u2_remHi_267_), .Y(u2__abc_44228_n12150) );
  AND2X2 AND2X2_5103 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n6413), .Y(u2__abc_44228_n12153) );
  AND2X2 AND2X2_5104 ( .A(u2__abc_44228_n12154), .B(u2__abc_44228_n2972_bF_buf52), .Y(u2__abc_44228_n12155) );
  AND2X2 AND2X2_5105 ( .A(u2__abc_44228_n12152_1), .B(u2__abc_44228_n12155), .Y(u2__abc_44228_n12156) );
  AND2X2 AND2X2_5106 ( .A(u2__abc_44228_n12157), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_remHi_269__FF_INPUT) );
  AND2X2 AND2X2_5107 ( .A(u2__abc_44228_n3062_bF_buf8), .B(u2_remHi_270_), .Y(u2__abc_44228_n12159) );
  AND2X2 AND2X2_5108 ( .A(u2__abc_44228_n12127), .B(u2__abc_44228_n6437), .Y(u2__abc_44228_n12160) );
  AND2X2 AND2X2_5109 ( .A(u2__abc_44228_n12161_1), .B(u2__abc_44228_n6422), .Y(u2__abc_44228_n12162) );
  AND2X2 AND2X2_511 ( .A(u1__abc_43968_n377), .B(u1__abc_43968_n378), .Y(u1__abc_43968_n379) );
  AND2X2 AND2X2_5110 ( .A(u2__abc_44228_n12163), .B(u2__abc_44228_n12164), .Y(u2__abc_44228_n12165) );
  AND2X2 AND2X2_5111 ( .A(u2__abc_44228_n12165), .B(u2__abc_44228_n7547_bF_buf18), .Y(u2__abc_44228_n12166) );
  AND2X2 AND2X2_5112 ( .A(u2__abc_44228_n7548_1_bF_buf19), .B(u2_remHi_268_), .Y(u2__abc_44228_n12167) );
  AND2X2 AND2X2_5113 ( .A(u2__abc_44228_n2983_bF_buf65), .B(u2__abc_44228_n6395), .Y(u2__abc_44228_n12170) );
  AND2X2 AND2X2_5114 ( .A(u2__abc_44228_n12171), .B(u2__abc_44228_n2972_bF_buf51), .Y(u2__abc_44228_n12172) );
  AND2X2 AND2X2_5115 ( .A(u2__abc_44228_n12169), .B(u2__abc_44228_n12172), .Y(u2__abc_44228_n12173) );
  AND2X2 AND2X2_5116 ( .A(u2__abc_44228_n12174), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_remHi_270__FF_INPUT) );
  AND2X2 AND2X2_5117 ( .A(u2__abc_44228_n3062_bF_buf7), .B(u2_remHi_271_), .Y(u2__abc_44228_n12176_1) );
  AND2X2 AND2X2_5118 ( .A(u2__abc_44228_n12181), .B(u2__abc_44228_n7547_bF_buf17), .Y(u2__abc_44228_n12182) );
  AND2X2 AND2X2_5119 ( .A(u2__abc_44228_n12182), .B(u2__abc_44228_n12180), .Y(u2__abc_44228_n12183_1) );
  AND2X2 AND2X2_512 ( .A(u1__abc_43968_n380), .B(u1__abc_43968_n381), .Y(u1__abc_43968_n382) );
  AND2X2 AND2X2_5120 ( .A(u2__abc_44228_n7548_1_bF_buf18), .B(u2_remHi_269_), .Y(u2__abc_44228_n12184) );
  AND2X2 AND2X2_5121 ( .A(u2__abc_44228_n2983_bF_buf63), .B(u2__abc_44228_n6402), .Y(u2__abc_44228_n12187) );
  AND2X2 AND2X2_5122 ( .A(u2__abc_44228_n12188), .B(u2__abc_44228_n2972_bF_buf50), .Y(u2__abc_44228_n12189) );
  AND2X2 AND2X2_5123 ( .A(u2__abc_44228_n12186), .B(u2__abc_44228_n12189), .Y(u2__abc_44228_n12190) );
  AND2X2 AND2X2_5124 ( .A(u2__abc_44228_n12191), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_remHi_271__FF_INPUT) );
  AND2X2 AND2X2_5125 ( .A(u2__abc_44228_n3062_bF_buf6), .B(u2_remHi_272_), .Y(u2__abc_44228_n12193) );
  AND2X2 AND2X2_5126 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6528), .Y(u2__abc_44228_n12194) );
  AND2X2 AND2X2_5127 ( .A(u2__abc_44228_n12195_1), .B(u2__abc_44228_n6398), .Y(u2__abc_44228_n12197) );
  AND2X2 AND2X2_5128 ( .A(u2__abc_44228_n12198), .B(u2__abc_44228_n12196), .Y(u2__abc_44228_n12199) );
  AND2X2 AND2X2_5129 ( .A(u2__abc_44228_n12200), .B(u2__abc_44228_n12201), .Y(u2__abc_44228_n12202_1) );
  AND2X2 AND2X2_513 ( .A(u1__abc_43968_n379), .B(u1__abc_43968_n382), .Y(u1__abc_43968_n383) );
  AND2X2 AND2X2_5130 ( .A(u2__abc_44228_n2983_bF_buf61), .B(u2__abc_44228_n6388), .Y(u2__abc_44228_n12204) );
  AND2X2 AND2X2_5131 ( .A(u2__abc_44228_n12205), .B(u2__abc_44228_n2972_bF_buf49), .Y(u2__abc_44228_n12206) );
  AND2X2 AND2X2_5132 ( .A(u2__abc_44228_n12203), .B(u2__abc_44228_n12206), .Y(u2__abc_44228_n12207) );
  AND2X2 AND2X2_5133 ( .A(u2__abc_44228_n12208), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_remHi_272__FF_INPUT) );
  AND2X2 AND2X2_5134 ( .A(u2__abc_44228_n3062_bF_buf5), .B(u2_remHi_273_), .Y(u2__abc_44228_n12210_1) );
  AND2X2 AND2X2_5135 ( .A(u2__abc_44228_n12198), .B(u2__abc_44228_n6572), .Y(u2__abc_44228_n12212) );
  AND2X2 AND2X2_5136 ( .A(u2__abc_44228_n12215), .B(u2__abc_44228_n12213), .Y(u2__abc_44228_n12216) );
  AND2X2 AND2X2_5137 ( .A(u2__abc_44228_n12216), .B(u2__abc_44228_n7547_bF_buf15), .Y(u2__abc_44228_n12217_1) );
  AND2X2 AND2X2_5138 ( .A(u2__abc_44228_n7548_1_bF_buf16), .B(u2_remHi_271_), .Y(u2__abc_44228_n12218) );
  AND2X2 AND2X2_5139 ( .A(u2__abc_44228_n2983_bF_buf59), .B(u2__abc_44228_n6382), .Y(u2__abc_44228_n12221) );
  AND2X2 AND2X2_514 ( .A(u1__abc_43968_n376), .B(u1__abc_43968_n383), .Y(u1__abc_43968_n384) );
  AND2X2 AND2X2_5140 ( .A(u2__abc_44228_n12222), .B(u2__abc_44228_n2972_bF_buf48), .Y(u2__abc_44228_n12223) );
  AND2X2 AND2X2_5141 ( .A(u2__abc_44228_n12220), .B(u2__abc_44228_n12223), .Y(u2__abc_44228_n12224) );
  AND2X2 AND2X2_5142 ( .A(u2__abc_44228_n12225), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_remHi_273__FF_INPUT) );
  AND2X2 AND2X2_5143 ( .A(u2__abc_44228_n3062_bF_buf4), .B(u2_remHi_274_), .Y(u2__abc_44228_n12227) );
  AND2X2 AND2X2_5144 ( .A(u2__abc_44228_n12198), .B(u2__abc_44228_n6573), .Y(u2__abc_44228_n12228) );
  AND2X2 AND2X2_5145 ( .A(u2__abc_44228_n12230), .B(u2__abc_44228_n6391), .Y(u2__abc_44228_n12231) );
  AND2X2 AND2X2_5146 ( .A(u2__abc_44228_n12232), .B(u2__abc_44228_n12233_1), .Y(u2__abc_44228_n12234) );
  AND2X2 AND2X2_5147 ( .A(u2__abc_44228_n12234), .B(u2__abc_44228_n7547_bF_buf14), .Y(u2__abc_44228_n12235) );
  AND2X2 AND2X2_5148 ( .A(u2__abc_44228_n7548_1_bF_buf15), .B(u2_remHi_272_), .Y(u2__abc_44228_n12236) );
  AND2X2 AND2X2_5149 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n6373), .Y(u2__abc_44228_n12239) );
  AND2X2 AND2X2_515 ( .A(u1__abc_43968_n369), .B(u1__abc_43968_n384), .Y(u1__abc_43968_n385) );
  AND2X2 AND2X2_5150 ( .A(u2__abc_44228_n12240), .B(u2__abc_44228_n2972_bF_buf47), .Y(u2__abc_44228_n12241_1) );
  AND2X2 AND2X2_5151 ( .A(u2__abc_44228_n12238), .B(u2__abc_44228_n12241_1), .Y(u2__abc_44228_n12242) );
  AND2X2 AND2X2_5152 ( .A(u2__abc_44228_n12243), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_remHi_274__FF_INPUT) );
  AND2X2 AND2X2_5153 ( .A(u2__abc_44228_n3062_bF_buf3), .B(u2_remHi_275_), .Y(u2__abc_44228_n12245) );
  AND2X2 AND2X2_5154 ( .A(u2__abc_44228_n12250), .B(u2__abc_44228_n7547_bF_buf13), .Y(u2__abc_44228_n12251) );
  AND2X2 AND2X2_5155 ( .A(u2__abc_44228_n12251), .B(u2__abc_44228_n12249), .Y(u2__abc_44228_n12252) );
  AND2X2 AND2X2_5156 ( .A(u2__abc_44228_n7548_1_bF_buf14), .B(u2_remHi_273_), .Y(u2__abc_44228_n12253) );
  AND2X2 AND2X2_5157 ( .A(u2__abc_44228_n2983_bF_buf56), .B(u2__abc_44228_n6367), .Y(u2__abc_44228_n12256) );
  AND2X2 AND2X2_5158 ( .A(u2__abc_44228_n12257), .B(u2__abc_44228_n2972_bF_buf46), .Y(u2__abc_44228_n12258_1) );
  AND2X2 AND2X2_5159 ( .A(u2__abc_44228_n12255), .B(u2__abc_44228_n12258_1), .Y(u2__abc_44228_n12259) );
  AND2X2 AND2X2_516 ( .A(u1__abc_43968_n354), .B(u1__abc_43968_n385), .Y(u1__abc_43968_n386) );
  AND2X2 AND2X2_5160 ( .A(u2__abc_44228_n12260), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_remHi_275__FF_INPUT) );
  AND2X2 AND2X2_5161 ( .A(u2__abc_44228_n3062_bF_buf2), .B(u2_remHi_276_), .Y(u2__abc_44228_n12262) );
  AND2X2 AND2X2_5162 ( .A(u2__abc_44228_n12195_1), .B(u2__abc_44228_n6407), .Y(u2__abc_44228_n12263) );
  AND2X2 AND2X2_5163 ( .A(u2__abc_44228_n12264), .B(u2__abc_44228_n6376), .Y(u2__abc_44228_n12266) );
  AND2X2 AND2X2_5164 ( .A(u2__abc_44228_n12267), .B(u2__abc_44228_n12265_1), .Y(u2__abc_44228_n12268) );
  AND2X2 AND2X2_5165 ( .A(u2__abc_44228_n12269), .B(u2__abc_44228_n12270), .Y(u2__abc_44228_n12271) );
  AND2X2 AND2X2_5166 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n6359), .Y(u2__abc_44228_n12273_1) );
  AND2X2 AND2X2_5167 ( .A(u2__abc_44228_n12274), .B(u2__abc_44228_n2972_bF_buf45), .Y(u2__abc_44228_n12275) );
  AND2X2 AND2X2_5168 ( .A(u2__abc_44228_n12272), .B(u2__abc_44228_n12275), .Y(u2__abc_44228_n12276) );
  AND2X2 AND2X2_5169 ( .A(u2__abc_44228_n12277), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_remHi_276__FF_INPUT) );
  AND2X2 AND2X2_517 ( .A(u1__abc_43968_n323), .B(u1__abc_43968_n386), .Y(u1__abc_43968_n387) );
  AND2X2 AND2X2_5170 ( .A(u2__abc_44228_n3062_bF_buf1), .B(u2_remHi_277_), .Y(u2__abc_44228_n12279) );
  AND2X2 AND2X2_5171 ( .A(u2__abc_44228_n12267), .B(u2__abc_44228_n6581), .Y(u2__abc_44228_n12281) );
  AND2X2 AND2X2_5172 ( .A(u2__abc_44228_n12284), .B(u2__abc_44228_n12282), .Y(u2__abc_44228_n12285) );
  AND2X2 AND2X2_5173 ( .A(u2__abc_44228_n12285), .B(u2__abc_44228_n7547_bF_buf11), .Y(u2__abc_44228_n12286) );
  AND2X2 AND2X2_5174 ( .A(u2__abc_44228_n7548_1_bF_buf12), .B(u2_remHi_275_), .Y(u2__abc_44228_n12287) );
  AND2X2 AND2X2_5175 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n6353), .Y(u2__abc_44228_n12290) );
  AND2X2 AND2X2_5176 ( .A(u2__abc_44228_n12291), .B(u2__abc_44228_n2972_bF_buf44), .Y(u2__abc_44228_n12292) );
  AND2X2 AND2X2_5177 ( .A(u2__abc_44228_n12289_1), .B(u2__abc_44228_n12292), .Y(u2__abc_44228_n12293) );
  AND2X2 AND2X2_5178 ( .A(u2__abc_44228_n12294), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_remHi_277__FF_INPUT) );
  AND2X2 AND2X2_5179 ( .A(u2__abc_44228_n3062_bF_buf0), .B(u2_remHi_278_), .Y(u2__abc_44228_n12296_1) );
  AND2X2 AND2X2_518 ( .A(u1__abc_43968_n387), .B(u1__abc_43968_n260), .Y(u1_mz) );
  AND2X2 AND2X2_5180 ( .A(u2__abc_44228_n12264), .B(u2__abc_44228_n6377), .Y(u2__abc_44228_n12297) );
  AND2X2 AND2X2_5181 ( .A(u2__abc_44228_n12298), .B(u2__abc_44228_n6362), .Y(u2__abc_44228_n12299) );
  AND2X2 AND2X2_5182 ( .A(u2__abc_44228_n12300), .B(u2__abc_44228_n12301), .Y(u2__abc_44228_n12302) );
  AND2X2 AND2X2_5183 ( .A(u2__abc_44228_n12302), .B(u2__abc_44228_n7547_bF_buf10), .Y(u2__abc_44228_n12303) );
  AND2X2 AND2X2_5184 ( .A(u2__abc_44228_n7548_1_bF_buf11), .B(u2_remHi_276_), .Y(u2__abc_44228_n12304_1) );
  AND2X2 AND2X2_5185 ( .A(u2__abc_44228_n2983_bF_buf51), .B(u2__abc_44228_n6329), .Y(u2__abc_44228_n12307) );
  AND2X2 AND2X2_5186 ( .A(u2__abc_44228_n12308), .B(u2__abc_44228_n2972_bF_buf43), .Y(u2__abc_44228_n12309) );
  AND2X2 AND2X2_5187 ( .A(u2__abc_44228_n12306), .B(u2__abc_44228_n12309), .Y(u2__abc_44228_n12310) );
  AND2X2 AND2X2_5188 ( .A(u2__abc_44228_n12311_1), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_remHi_278__FF_INPUT) );
  AND2X2 AND2X2_5189 ( .A(u2__abc_44228_n3062_bF_buf92), .B(u2_remHi_279_), .Y(u2__abc_44228_n12313) );
  AND2X2 AND2X2_519 ( .A(u1__abc_43968_n392), .B(u1_xinf), .Y(aNan) );
  AND2X2 AND2X2_5190 ( .A(u2__abc_44228_n12318), .B(u2__abc_44228_n7547_bF_buf9), .Y(u2__abc_44228_n12319) );
  AND2X2 AND2X2_5191 ( .A(u2__abc_44228_n12319), .B(u2__abc_44228_n12317), .Y(u2__abc_44228_n12320) );
  AND2X2 AND2X2_5192 ( .A(u2__abc_44228_n7548_1_bF_buf10), .B(u2_remHi_277_), .Y(u2__abc_44228_n12321) );
  AND2X2 AND2X2_5193 ( .A(u2__abc_44228_n2983_bF_buf49), .B(u2__abc_44228_n6323), .Y(u2__abc_44228_n12324) );
  AND2X2 AND2X2_5194 ( .A(u2__abc_44228_n12325), .B(u2__abc_44228_n2972_bF_buf42), .Y(u2__abc_44228_n12326) );
  AND2X2 AND2X2_5195 ( .A(u2__abc_44228_n12323), .B(u2__abc_44228_n12326), .Y(u2__abc_44228_n12327) );
  AND2X2 AND2X2_5196 ( .A(u2__abc_44228_n12328), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_remHi_279__FF_INPUT) );
  AND2X2 AND2X2_5197 ( .A(u2__abc_44228_n3062_bF_buf91), .B(u2_remHi_280_), .Y(u2__abc_44228_n12330) );
  AND2X2 AND2X2_5198 ( .A(u2__abc_44228_n12195_1), .B(u2__abc_44228_n6408), .Y(u2__abc_44228_n12331) );
  AND2X2 AND2X2_5199 ( .A(u2__abc_44228_n12332), .B(u2__abc_44228_n6332), .Y(u2__abc_44228_n12333) );
  AND2X2 AND2X2_52 ( .A(_abc_64468_n753_bF_buf4), .B(sqrto_51_), .Y(_auto_iopadmap_cc_313_execute_65414_87_) );
  AND2X2 AND2X2_520 ( .A(u2__abc_44228_n2962), .B(u2_state_0_), .Y(u2__abc_44228_n2963) );
  AND2X2 AND2X2_5200 ( .A(u2__abc_44228_n12334), .B(u2__abc_44228_n12335), .Y(u2__abc_44228_n12336) );
  AND2X2 AND2X2_5201 ( .A(u2__abc_44228_n12337_1), .B(u2__abc_44228_n12338), .Y(u2__abc_44228_n12339) );
  AND2X2 AND2X2_5202 ( .A(u2__abc_44228_n2983_bF_buf47), .B(u2__abc_44228_n6343), .Y(u2__abc_44228_n12341) );
  AND2X2 AND2X2_5203 ( .A(u2__abc_44228_n12342), .B(u2__abc_44228_n2972_bF_buf41), .Y(u2__abc_44228_n12343) );
  AND2X2 AND2X2_5204 ( .A(u2__abc_44228_n12340), .B(u2__abc_44228_n12343), .Y(u2__abc_44228_n12344_1) );
  AND2X2 AND2X2_5205 ( .A(u2__abc_44228_n12345), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_remHi_280__FF_INPUT) );
  AND2X2 AND2X2_5206 ( .A(u2__abc_44228_n3062_bF_buf90), .B(u2_remHi_281_), .Y(u2__abc_44228_n12347) );
  AND2X2 AND2X2_5207 ( .A(u2__abc_44228_n12334), .B(u2__abc_44228_n6591), .Y(u2__abc_44228_n12349) );
  AND2X2 AND2X2_5208 ( .A(u2__abc_44228_n12352), .B(u2__abc_44228_n12350), .Y(u2__abc_44228_n12353_1) );
  AND2X2 AND2X2_5209 ( .A(u2__abc_44228_n12353_1), .B(u2__abc_44228_n7547_bF_buf7), .Y(u2__abc_44228_n12354) );
  AND2X2 AND2X2_521 ( .A(u2__abc_44228_n2964), .B(ce), .Y(u2__abc_44228_n2965) );
  AND2X2 AND2X2_5210 ( .A(u2__abc_44228_n7548_1_bF_buf8), .B(u2_remHi_279_), .Y(u2__abc_44228_n12355) );
  AND2X2 AND2X2_5211 ( .A(u2__abc_44228_n2983_bF_buf45), .B(u2__abc_44228_n6337), .Y(u2__abc_44228_n12358) );
  AND2X2 AND2X2_5212 ( .A(u2__abc_44228_n12359), .B(u2__abc_44228_n2972_bF_buf40), .Y(u2__abc_44228_n12360_1) );
  AND2X2 AND2X2_5213 ( .A(u2__abc_44228_n12357), .B(u2__abc_44228_n12360_1), .Y(u2__abc_44228_n12361) );
  AND2X2 AND2X2_5214 ( .A(u2__abc_44228_n12362), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_remHi_281__FF_INPUT) );
  AND2X2 AND2X2_5215 ( .A(u2__abc_44228_n3062_bF_buf89), .B(u2_remHi_282_), .Y(u2__abc_44228_n12364) );
  AND2X2 AND2X2_5216 ( .A(u2__abc_44228_n12332), .B(u2__abc_44228_n6333_1), .Y(u2__abc_44228_n12365) );
  AND2X2 AND2X2_5217 ( .A(u2__abc_44228_n12366), .B(u2__abc_44228_n6346), .Y(u2__abc_44228_n12367) );
  AND2X2 AND2X2_5218 ( .A(u2__abc_44228_n12368_1), .B(u2__abc_44228_n12369), .Y(u2__abc_44228_n12370) );
  AND2X2 AND2X2_5219 ( .A(u2__abc_44228_n12370), .B(u2__abc_44228_n7547_bF_buf6), .Y(u2__abc_44228_n12371) );
  AND2X2 AND2X2_522 ( .A(u2__abc_44228_n2966_bF_buf107), .B(u2__abc_44228_n2967), .Y(u2__abc_44228_n2968) );
  AND2X2 AND2X2_5220 ( .A(u2__abc_44228_n7548_1_bF_buf7), .B(u2_remHi_280_), .Y(u2__abc_44228_n12372) );
  AND2X2 AND2X2_5221 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n6314), .Y(u2__abc_44228_n12375_1) );
  AND2X2 AND2X2_5222 ( .A(u2__abc_44228_n12376), .B(u2__abc_44228_n2972_bF_buf39), .Y(u2__abc_44228_n12377) );
  AND2X2 AND2X2_5223 ( .A(u2__abc_44228_n12374), .B(u2__abc_44228_n12377), .Y(u2__abc_44228_n12378) );
  AND2X2 AND2X2_5224 ( .A(u2__abc_44228_n12379), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_remHi_282__FF_INPUT) );
  AND2X2 AND2X2_5225 ( .A(u2__abc_44228_n3062_bF_buf88), .B(u2_remHi_283_), .Y(u2__abc_44228_n12381) );
  AND2X2 AND2X2_5226 ( .A(u2__abc_44228_n12368_1), .B(u2__abc_44228_n6596), .Y(u2__abc_44228_n12383) );
  AND2X2 AND2X2_5227 ( .A(u2__abc_44228_n12386), .B(u2__abc_44228_n12384), .Y(u2__abc_44228_n12387) );
  AND2X2 AND2X2_5228 ( .A(u2__abc_44228_n12387), .B(u2__abc_44228_n7547_bF_buf5), .Y(u2__abc_44228_n12388) );
  AND2X2 AND2X2_5229 ( .A(u2__abc_44228_n7548_1_bF_buf6), .B(u2_remHi_281_), .Y(u2__abc_44228_n12389) );
  AND2X2 AND2X2_523 ( .A(u2__abc_44228_n2968), .B(u2_state_0_), .Y(u2__abc_44228_n2969) );
  AND2X2 AND2X2_5230 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n6308), .Y(u2__abc_44228_n12392_1) );
  AND2X2 AND2X2_5231 ( .A(u2__abc_44228_n12393), .B(u2__abc_44228_n2972_bF_buf38), .Y(u2__abc_44228_n12394) );
  AND2X2 AND2X2_5232 ( .A(u2__abc_44228_n12391), .B(u2__abc_44228_n12394), .Y(u2__abc_44228_n12395) );
  AND2X2 AND2X2_5233 ( .A(u2__abc_44228_n12396), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_remHi_283__FF_INPUT) );
  AND2X2 AND2X2_5234 ( .A(u2__abc_44228_n3062_bF_buf87), .B(u2_remHi_284_), .Y(u2__abc_44228_n12398) );
  AND2X2 AND2X2_5235 ( .A(u2__abc_44228_n12368_1), .B(u2__abc_44228_n6597_1), .Y(u2__abc_44228_n12399) );
  AND2X2 AND2X2_5236 ( .A(u2__abc_44228_n12401), .B(u2__abc_44228_n6317), .Y(u2__abc_44228_n12403) );
  AND2X2 AND2X2_5237 ( .A(u2__abc_44228_n12404), .B(u2__abc_44228_n12402), .Y(u2__abc_44228_n12405) );
  AND2X2 AND2X2_5238 ( .A(u2__abc_44228_n12405), .B(u2__abc_44228_n7547_bF_buf4), .Y(u2__abc_44228_n12406) );
  AND2X2 AND2X2_5239 ( .A(u2__abc_44228_n7548_1_bF_buf5), .B(u2_remHi_282_), .Y(u2__abc_44228_n12407_1) );
  AND2X2 AND2X2_524 ( .A(ce), .B(u2_state_2_), .Y(u2__abc_44228_n2972) );
  AND2X2 AND2X2_5240 ( .A(u2__abc_44228_n2983_bF_buf41), .B(u2__abc_44228_n6300), .Y(u2__abc_44228_n12410) );
  AND2X2 AND2X2_5241 ( .A(u2__abc_44228_n12411), .B(u2__abc_44228_n2972_bF_buf37), .Y(u2__abc_44228_n12412) );
  AND2X2 AND2X2_5242 ( .A(u2__abc_44228_n12409), .B(u2__abc_44228_n12412), .Y(u2__abc_44228_n12413) );
  AND2X2 AND2X2_5243 ( .A(u2__abc_44228_n12414), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_remHi_284__FF_INPUT) );
  AND2X2 AND2X2_5244 ( .A(u2__abc_44228_n3062_bF_buf86), .B(u2_remHi_285_), .Y(u2__abc_44228_n12416_1) );
  AND2X2 AND2X2_5245 ( .A(u2__abc_44228_n12404), .B(u2__abc_44228_n6604), .Y(u2__abc_44228_n12417) );
  AND2X2 AND2X2_5246 ( .A(u2__abc_44228_n12417), .B(u2__abc_44228_n6311), .Y(u2__abc_44228_n12418) );
  AND2X2 AND2X2_5247 ( .A(u2__abc_44228_n12420), .B(u2__abc_44228_n12419), .Y(u2__abc_44228_n12421) );
  AND2X2 AND2X2_5248 ( .A(u2__abc_44228_n12422), .B(u2__abc_44228_n7547_bF_buf3), .Y(u2__abc_44228_n12423_1) );
  AND2X2 AND2X2_5249 ( .A(u2__abc_44228_n7548_1_bF_buf4), .B(u2_remHi_283_), .Y(u2__abc_44228_n12424) );
  AND2X2 AND2X2_525 ( .A(u2__abc_44228_n2972_bF_buf107), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2__abc_44228_n2973) );
  AND2X2 AND2X2_5250 ( .A(u2__abc_44228_n2983_bF_buf39), .B(u2__abc_44228_n6294), .Y(u2__abc_44228_n12427) );
  AND2X2 AND2X2_5251 ( .A(u2__abc_44228_n12428), .B(u2__abc_44228_n2972_bF_buf36), .Y(u2__abc_44228_n12429) );
  AND2X2 AND2X2_5252 ( .A(u2__abc_44228_n12426), .B(u2__abc_44228_n12429), .Y(u2__abc_44228_n12430) );
  AND2X2 AND2X2_5253 ( .A(u2__abc_44228_n12431_1), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_remHi_285__FF_INPUT) );
  AND2X2 AND2X2_5254 ( .A(u2__abc_44228_n3062_bF_buf85), .B(u2_remHi_286_), .Y(u2__abc_44228_n12433) );
  AND2X2 AND2X2_5255 ( .A(u2__abc_44228_n12404), .B(u2__abc_44228_n6605), .Y(u2__abc_44228_n12434) );
  AND2X2 AND2X2_5256 ( .A(u2__abc_44228_n12436), .B(u2__abc_44228_n6303), .Y(u2__abc_44228_n12437) );
  AND2X2 AND2X2_5257 ( .A(u2__abc_44228_n12439), .B(u2__abc_44228_n7547_bF_buf2), .Y(u2__abc_44228_n12440) );
  AND2X2 AND2X2_5258 ( .A(u2__abc_44228_n12440), .B(u2__abc_44228_n12438_1), .Y(u2__abc_44228_n12441) );
  AND2X2 AND2X2_5259 ( .A(u2__abc_44228_n7548_1_bF_buf3), .B(u2_remHi_284_), .Y(u2__abc_44228_n12442) );
  AND2X2 AND2X2_526 ( .A(u2__abc_44228_n2974), .B(u2_cnt_1_), .Y(u2__abc_44228_n2975) );
  AND2X2 AND2X2_5260 ( .A(u2__abc_44228_n2983_bF_buf37), .B(u2__abc_44228_n6282), .Y(u2__abc_44228_n12445) );
  AND2X2 AND2X2_5261 ( .A(u2__abc_44228_n12446), .B(u2__abc_44228_n2972_bF_buf35), .Y(u2__abc_44228_n12447) );
  AND2X2 AND2X2_5262 ( .A(u2__abc_44228_n12444), .B(u2__abc_44228_n12447), .Y(u2__abc_44228_n12448) );
  AND2X2 AND2X2_5263 ( .A(u2__abc_44228_n12449), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_remHi_286__FF_INPUT) );
  AND2X2 AND2X2_5264 ( .A(u2__abc_44228_n3062_bF_buf84), .B(u2_remHi_287_), .Y(u2__abc_44228_n12451) );
  AND2X2 AND2X2_5265 ( .A(u2__abc_44228_n12456), .B(u2__abc_44228_n7547_bF_buf1), .Y(u2__abc_44228_n12457_1) );
  AND2X2 AND2X2_5266 ( .A(u2__abc_44228_n12457_1), .B(u2__abc_44228_n12455), .Y(u2__abc_44228_n12458) );
  AND2X2 AND2X2_5267 ( .A(u2__abc_44228_n7548_1_bF_buf2), .B(u2_remHi_285_), .Y(u2__abc_44228_n12459) );
  AND2X2 AND2X2_5268 ( .A(u2__abc_44228_n2983_bF_buf35), .B(u2__abc_44228_n6276), .Y(u2__abc_44228_n12462) );
  AND2X2 AND2X2_5269 ( .A(u2__abc_44228_n12463), .B(u2__abc_44228_n2972_bF_buf34), .Y(u2__abc_44228_n12464) );
  AND2X2 AND2X2_527 ( .A(u2__abc_44228_n2977), .B(u2__abc_44228_n2975), .Y(u2__abc_44228_n2978) );
  AND2X2 AND2X2_5270 ( .A(u2__abc_44228_n12461), .B(u2__abc_44228_n12464), .Y(u2__abc_44228_n12465_1) );
  AND2X2 AND2X2_5271 ( .A(u2__abc_44228_n12466), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_remHi_287__FF_INPUT) );
  AND2X2 AND2X2_5272 ( .A(u2__abc_44228_n3062_bF_buf83), .B(u2_remHi_288_), .Y(u2__abc_44228_n12468) );
  AND2X2 AND2X2_5273 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6529), .Y(u2__abc_44228_n12469) );
  AND2X2 AND2X2_5274 ( .A(u2__abc_44228_n12470), .B(u2__abc_44228_n6285), .Y(u2__abc_44228_n12471) );
  AND2X2 AND2X2_5275 ( .A(u2__abc_44228_n12472_1), .B(u2__abc_44228_n12473), .Y(u2__abc_44228_n12474) );
  AND2X2 AND2X2_5276 ( .A(u2__abc_44228_n12475), .B(u2__abc_44228_n12476), .Y(u2__abc_44228_n12477) );
  AND2X2 AND2X2_5277 ( .A(u2__abc_44228_n2983_bF_buf33), .B(u2__abc_44228_n6268), .Y(u2__abc_44228_n12479) );
  AND2X2 AND2X2_5278 ( .A(u2__abc_44228_n12480), .B(u2__abc_44228_n2972_bF_buf33), .Y(u2__abc_44228_n12481_1) );
  AND2X2 AND2X2_5279 ( .A(u2__abc_44228_n12478), .B(u2__abc_44228_n12481_1), .Y(u2__abc_44228_n12482) );
  AND2X2 AND2X2_528 ( .A(u2__abc_44228_n2979), .B(u2_cnt_5_), .Y(u2__abc_44228_n2980) );
  AND2X2 AND2X2_5280 ( .A(u2__abc_44228_n12483), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_remHi_288__FF_INPUT) );
  AND2X2 AND2X2_5281 ( .A(u2__abc_44228_n3062_bF_buf82), .B(u2_remHi_289_), .Y(u2__abc_44228_n12485) );
  AND2X2 AND2X2_5282 ( .A(u2__abc_44228_n12472_1), .B(u2__abc_44228_n6614), .Y(u2__abc_44228_n12487) );
  AND2X2 AND2X2_5283 ( .A(u2__abc_44228_n12490), .B(u2__abc_44228_n12488_1), .Y(u2__abc_44228_n12491) );
  AND2X2 AND2X2_5284 ( .A(u2__abc_44228_n12491), .B(u2__abc_44228_n7547_bF_buf57), .Y(u2__abc_44228_n12492) );
  AND2X2 AND2X2_5285 ( .A(u2__abc_44228_n7548_1_bF_buf0), .B(u2_remHi_287_), .Y(u2__abc_44228_n12493) );
  AND2X2 AND2X2_5286 ( .A(u2__abc_44228_n2983_bF_buf31), .B(u2__abc_44228_n6262), .Y(u2__abc_44228_n12496_1) );
  AND2X2 AND2X2_5287 ( .A(u2__abc_44228_n12497), .B(u2__abc_44228_n2972_bF_buf32), .Y(u2__abc_44228_n12498) );
  AND2X2 AND2X2_5288 ( .A(u2__abc_44228_n12495), .B(u2__abc_44228_n12498), .Y(u2__abc_44228_n12499) );
  AND2X2 AND2X2_5289 ( .A(u2__abc_44228_n12500), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_remHi_289__FF_INPUT) );
  AND2X2 AND2X2_529 ( .A(u2_cnt_7_), .B(u2_cnt_6_), .Y(u2__abc_44228_n2981) );
  AND2X2 AND2X2_5290 ( .A(u2__abc_44228_n3062_bF_buf81), .B(u2_remHi_290_), .Y(u2__abc_44228_n12502) );
  AND2X2 AND2X2_5291 ( .A(u2__abc_44228_n12470), .B(u2__abc_44228_n6286), .Y(u2__abc_44228_n12503_1) );
  AND2X2 AND2X2_5292 ( .A(u2__abc_44228_n12504), .B(u2__abc_44228_n6271), .Y(u2__abc_44228_n12505) );
  AND2X2 AND2X2_5293 ( .A(u2__abc_44228_n12506), .B(u2__abc_44228_n12507), .Y(u2__abc_44228_n12508) );
  AND2X2 AND2X2_5294 ( .A(u2__abc_44228_n12509), .B(u2__abc_44228_n12510), .Y(u2__abc_44228_n12511) );
  AND2X2 AND2X2_5295 ( .A(u2__abc_44228_n2983_bF_buf29), .B(u2__abc_44228_n6253), .Y(u2__abc_44228_n12513_1) );
  AND2X2 AND2X2_5296 ( .A(u2__abc_44228_n12514), .B(u2__abc_44228_n2972_bF_buf31), .Y(u2__abc_44228_n12515) );
  AND2X2 AND2X2_5297 ( .A(u2__abc_44228_n12512), .B(u2__abc_44228_n12515), .Y(u2__abc_44228_n12516) );
  AND2X2 AND2X2_5298 ( .A(u2__abc_44228_n12517), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_remHi_290__FF_INPUT) );
  AND2X2 AND2X2_5299 ( .A(u2__abc_44228_n3062_bF_buf80), .B(u2_remHi_291_), .Y(u2__abc_44228_n12519) );
  AND2X2 AND2X2_53 ( .A(_abc_64468_n753_bF_buf3), .B(sqrto_52_), .Y(_auto_iopadmap_cc_313_execute_65414_88_) );
  AND2X2 AND2X2_530 ( .A(u2__abc_44228_n2980), .B(u2__abc_44228_n2981), .Y(u2__abc_44228_n2982) );
  AND2X2 AND2X2_5300 ( .A(u2__abc_44228_n12524), .B(u2__abc_44228_n7547_bF_buf55), .Y(u2__abc_44228_n12525) );
  AND2X2 AND2X2_5301 ( .A(u2__abc_44228_n12525), .B(u2__abc_44228_n12523), .Y(u2__abc_44228_n12526) );
  AND2X2 AND2X2_5302 ( .A(u2__abc_44228_n7548_1_bF_buf56), .B(u2_remHi_289_), .Y(u2__abc_44228_n12527) );
  AND2X2 AND2X2_5303 ( .A(u2__abc_44228_n2983_bF_buf27), .B(u2__abc_44228_n6247), .Y(u2__abc_44228_n12530) );
  AND2X2 AND2X2_5304 ( .A(u2__abc_44228_n12531), .B(u2__abc_44228_n2972_bF_buf30), .Y(u2__abc_44228_n12532) );
  AND2X2 AND2X2_5305 ( .A(u2__abc_44228_n12529), .B(u2__abc_44228_n12532), .Y(u2__abc_44228_n12533) );
  AND2X2 AND2X2_5306 ( .A(u2__abc_44228_n12534), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_remHi_291__FF_INPUT) );
  AND2X2 AND2X2_5307 ( .A(u2__abc_44228_n3062_bF_buf79), .B(u2_remHi_292_), .Y(u2__abc_44228_n12536) );
  AND2X2 AND2X2_5308 ( .A(u2__abc_44228_n12470), .B(u2__abc_44228_n6287_1), .Y(u2__abc_44228_n12537) );
  AND2X2 AND2X2_5309 ( .A(u2__abc_44228_n12538), .B(u2__abc_44228_n6256), .Y(u2__abc_44228_n12540) );
  AND2X2 AND2X2_531 ( .A(u2__abc_44228_n2978), .B(u2__abc_44228_n2982), .Y(u2__abc_44228_n2983) );
  AND2X2 AND2X2_5310 ( .A(u2__abc_44228_n12541), .B(u2__abc_44228_n12539), .Y(u2__abc_44228_n12542) );
  AND2X2 AND2X2_5311 ( .A(u2__abc_44228_n12543), .B(u2__abc_44228_n12544_1), .Y(u2__abc_44228_n12545) );
  AND2X2 AND2X2_5312 ( .A(u2__abc_44228_n2983_bF_buf25), .B(u2__abc_44228_n6239), .Y(u2__abc_44228_n12547) );
  AND2X2 AND2X2_5313 ( .A(u2__abc_44228_n12548), .B(u2__abc_44228_n2972_bF_buf29), .Y(u2__abc_44228_n12549) );
  AND2X2 AND2X2_5314 ( .A(u2__abc_44228_n12546), .B(u2__abc_44228_n12549), .Y(u2__abc_44228_n12550) );
  AND2X2 AND2X2_5315 ( .A(u2__abc_44228_n12551_1), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_remHi_292__FF_INPUT) );
  AND2X2 AND2X2_5316 ( .A(u2__abc_44228_n3062_bF_buf78), .B(u2_remHi_293_), .Y(u2__abc_44228_n12553) );
  AND2X2 AND2X2_5317 ( .A(u2__abc_44228_n12541), .B(u2__abc_44228_n6623), .Y(u2__abc_44228_n12555) );
  AND2X2 AND2X2_5318 ( .A(u2__abc_44228_n12558), .B(u2__abc_44228_n12556), .Y(u2__abc_44228_n12559_1) );
  AND2X2 AND2X2_5319 ( .A(u2__abc_44228_n12559_1), .B(u2__abc_44228_n7547_bF_buf53), .Y(u2__abc_44228_n12560) );
  AND2X2 AND2X2_532 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n2973), .Y(u2__abc_44228_n2985) );
  AND2X2 AND2X2_5320 ( .A(u2__abc_44228_n7548_1_bF_buf54), .B(u2_remHi_291_), .Y(u2__abc_44228_n12561) );
  AND2X2 AND2X2_5321 ( .A(u2__abc_44228_n2983_bF_buf23), .B(u2__abc_44228_n6233), .Y(u2__abc_44228_n12564) );
  AND2X2 AND2X2_5322 ( .A(u2__abc_44228_n12565), .B(u2__abc_44228_n2972_bF_buf28), .Y(u2__abc_44228_n12566_1) );
  AND2X2 AND2X2_5323 ( .A(u2__abc_44228_n12563), .B(u2__abc_44228_n12566_1), .Y(u2__abc_44228_n12567) );
  AND2X2 AND2X2_5324 ( .A(u2__abc_44228_n12568), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_remHi_293__FF_INPUT) );
  AND2X2 AND2X2_5325 ( .A(u2__abc_44228_n3062_bF_buf77), .B(u2_remHi_294_), .Y(u2__abc_44228_n12570) );
  AND2X2 AND2X2_5326 ( .A(u2__abc_44228_n12538), .B(u2__abc_44228_n6257), .Y(u2__abc_44228_n12571) );
  AND2X2 AND2X2_5327 ( .A(u2__abc_44228_n12572), .B(u2__abc_44228_n6242_1), .Y(u2__abc_44228_n12573) );
  AND2X2 AND2X2_5328 ( .A(u2__abc_44228_n12574), .B(u2__abc_44228_n12575), .Y(u2__abc_44228_n12576) );
  AND2X2 AND2X2_5329 ( .A(u2__abc_44228_n12576), .B(u2__abc_44228_n7547_bF_buf52), .Y(u2__abc_44228_n12577_1) );
  AND2X2 AND2X2_533 ( .A(u2__abc_44228_n2968), .B(u2_state_2_), .Y(u2__abc_44228_n2986) );
  AND2X2 AND2X2_5330 ( .A(u2__abc_44228_n7548_1_bF_buf53), .B(u2_remHi_292_), .Y(u2__abc_44228_n12578) );
  AND2X2 AND2X2_5331 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n6209), .Y(u2__abc_44228_n12581) );
  AND2X2 AND2X2_5332 ( .A(u2__abc_44228_n12582), .B(u2__abc_44228_n2972_bF_buf27), .Y(u2__abc_44228_n12583) );
  AND2X2 AND2X2_5333 ( .A(u2__abc_44228_n12580), .B(u2__abc_44228_n12583), .Y(u2__abc_44228_n12584_1) );
  AND2X2 AND2X2_5334 ( .A(u2__abc_44228_n12585), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_remHi_294__FF_INPUT) );
  AND2X2 AND2X2_5335 ( .A(u2__abc_44228_n3062_bF_buf76), .B(u2_remHi_295_), .Y(u2__abc_44228_n12587) );
  AND2X2 AND2X2_5336 ( .A(u2__abc_44228_n12592_1), .B(u2__abc_44228_n7547_bF_buf51), .Y(u2__abc_44228_n12593) );
  AND2X2 AND2X2_5337 ( .A(u2__abc_44228_n12593), .B(u2__abc_44228_n12591), .Y(u2__abc_44228_n12594) );
  AND2X2 AND2X2_5338 ( .A(u2__abc_44228_n7548_1_bF_buf52), .B(u2_remHi_293_), .Y(u2__abc_44228_n12595) );
  AND2X2 AND2X2_5339 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n6203), .Y(u2__abc_44228_n12598) );
  AND2X2 AND2X2_534 ( .A(u2__abc_44228_n2966_bF_buf105), .B(ce), .Y(u2__abc_44228_n2987) );
  AND2X2 AND2X2_5340 ( .A(u2__abc_44228_n12599_1), .B(u2__abc_44228_n2972_bF_buf26), .Y(u2__abc_44228_n12600) );
  AND2X2 AND2X2_5341 ( .A(u2__abc_44228_n12597), .B(u2__abc_44228_n12600), .Y(u2__abc_44228_n12601) );
  AND2X2 AND2X2_5342 ( .A(u2__abc_44228_n12602), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_remHi_295__FF_INPUT) );
  AND2X2 AND2X2_5343 ( .A(u2__abc_44228_n3062_bF_buf75), .B(u2_remHi_296_), .Y(u2__abc_44228_n12604) );
  AND2X2 AND2X2_5344 ( .A(u2__abc_44228_n12470), .B(u2__abc_44228_n6288), .Y(u2__abc_44228_n12605) );
  AND2X2 AND2X2_5345 ( .A(u2__abc_44228_n12606), .B(u2__abc_44228_n6212), .Y(u2__abc_44228_n12607) );
  AND2X2 AND2X2_5346 ( .A(u2__abc_44228_n12608_1), .B(u2__abc_44228_n12609), .Y(u2__abc_44228_n12610) );
  AND2X2 AND2X2_5347 ( .A(u2__abc_44228_n12611), .B(u2__abc_44228_n12612), .Y(u2__abc_44228_n12613) );
  AND2X2 AND2X2_5348 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n6223), .Y(u2__abc_44228_n12615_1) );
  AND2X2 AND2X2_5349 ( .A(u2__abc_44228_n12616), .B(u2__abc_44228_n2972_bF_buf25), .Y(u2__abc_44228_n12617) );
  AND2X2 AND2X2_535 ( .A(u2_state_0_), .B(ld), .Y(u2__abc_44228_n2988) );
  AND2X2 AND2X2_5350 ( .A(u2__abc_44228_n12614), .B(u2__abc_44228_n12617), .Y(u2__abc_44228_n12618) );
  AND2X2 AND2X2_5351 ( .A(u2__abc_44228_n12619), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_remHi_296__FF_INPUT) );
  AND2X2 AND2X2_5352 ( .A(u2__abc_44228_n3062_bF_buf74), .B(u2_remHi_297_), .Y(u2__abc_44228_n12621) );
  AND2X2 AND2X2_5353 ( .A(u2__abc_44228_n12608_1), .B(u2__abc_44228_n6633), .Y(u2__abc_44228_n12623_1) );
  AND2X2 AND2X2_5354 ( .A(u2__abc_44228_n12626), .B(u2__abc_44228_n12624), .Y(u2__abc_44228_n12627) );
  AND2X2 AND2X2_5355 ( .A(u2__abc_44228_n12627), .B(u2__abc_44228_n7547_bF_buf49), .Y(u2__abc_44228_n12628) );
  AND2X2 AND2X2_5356 ( .A(u2__abc_44228_n7548_1_bF_buf50), .B(u2_remHi_295_), .Y(u2__abc_44228_n12629) );
  AND2X2 AND2X2_5357 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n6217), .Y(u2__abc_44228_n12632) );
  AND2X2 AND2X2_5358 ( .A(u2__abc_44228_n12633), .B(u2__abc_44228_n2972_bF_buf24), .Y(u2__abc_44228_n12634) );
  AND2X2 AND2X2_5359 ( .A(u2__abc_44228_n12631), .B(u2__abc_44228_n12634), .Y(u2__abc_44228_n12635) );
  AND2X2 AND2X2_536 ( .A(u2__abc_44228_n2987_bF_buf14), .B(u2__abc_44228_n2988_bF_buf13), .Y(u2__abc_44228_n2989) );
  AND2X2 AND2X2_5360 ( .A(u2__abc_44228_n12636), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_remHi_297__FF_INPUT) );
  AND2X2 AND2X2_5361 ( .A(u2__abc_44228_n3062_bF_buf73), .B(u2_remHi_298_), .Y(u2__abc_44228_n12638) );
  AND2X2 AND2X2_5362 ( .A(u2__abc_44228_n12606), .B(u2__abc_44228_n6213), .Y(u2__abc_44228_n12639) );
  AND2X2 AND2X2_5363 ( .A(u2__abc_44228_n12640_1), .B(u2__abc_44228_n6226), .Y(u2__abc_44228_n12641) );
  AND2X2 AND2X2_5364 ( .A(u2__abc_44228_n12642), .B(u2__abc_44228_n12643), .Y(u2__abc_44228_n12644) );
  AND2X2 AND2X2_5365 ( .A(u2__abc_44228_n12644), .B(u2__abc_44228_n7547_bF_buf48), .Y(u2__abc_44228_n12645) );
  AND2X2 AND2X2_5366 ( .A(u2__abc_44228_n7548_1_bF_buf49), .B(u2_remHi_296_), .Y(u2__abc_44228_n12646) );
  AND2X2 AND2X2_5367 ( .A(u2__abc_44228_n2983_bF_buf15), .B(u2__abc_44228_n6194), .Y(u2__abc_44228_n12649) );
  AND2X2 AND2X2_5368 ( .A(u2__abc_44228_n12650), .B(u2__abc_44228_n2972_bF_buf23), .Y(u2__abc_44228_n12651) );
  AND2X2 AND2X2_5369 ( .A(u2__abc_44228_n12648), .B(u2__abc_44228_n12651), .Y(u2__abc_44228_n12652) );
  AND2X2 AND2X2_537 ( .A(u2__abc_44228_n2968), .B(_auto_iopadmap_cc_313_execute_65412), .Y(u2__abc_44228_n2992) );
  AND2X2 AND2X2_5370 ( .A(u2__abc_44228_n12653), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_remHi_298__FF_INPUT) );
  AND2X2 AND2X2_5371 ( .A(u2__abc_44228_n3062_bF_buf72), .B(u2_remHi_299_), .Y(u2__abc_44228_n12655_1) );
  AND2X2 AND2X2_5372 ( .A(u2__abc_44228_n12642), .B(u2__abc_44228_n6638), .Y(u2__abc_44228_n12657) );
  AND2X2 AND2X2_5373 ( .A(u2__abc_44228_n12660), .B(u2__abc_44228_n12658), .Y(u2__abc_44228_n12661) );
  AND2X2 AND2X2_5374 ( .A(u2__abc_44228_n12661), .B(u2__abc_44228_n7547_bF_buf47), .Y(u2__abc_44228_n12662_1) );
  AND2X2 AND2X2_5375 ( .A(u2__abc_44228_n7548_1_bF_buf48), .B(u2_remHi_297_), .Y(u2__abc_44228_n12663) );
  AND2X2 AND2X2_5376 ( .A(u2__abc_44228_n2983_bF_buf13), .B(u2__abc_44228_n6188), .Y(u2__abc_44228_n12666) );
  AND2X2 AND2X2_5377 ( .A(u2__abc_44228_n12667), .B(u2__abc_44228_n2972_bF_buf22), .Y(u2__abc_44228_n12668) );
  AND2X2 AND2X2_5378 ( .A(u2__abc_44228_n12665), .B(u2__abc_44228_n12668), .Y(u2__abc_44228_n12669) );
  AND2X2 AND2X2_5379 ( .A(u2__abc_44228_n12670), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_remHi_299__FF_INPUT) );
  AND2X2 AND2X2_538 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n2973), .Y(u2__abc_44228_n2993) );
  AND2X2 AND2X2_5380 ( .A(u2__abc_44228_n3062_bF_buf71), .B(u2_remHi_300_), .Y(u2__abc_44228_n12672) );
  AND2X2 AND2X2_5381 ( .A(u2__abc_44228_n12642), .B(u2__abc_44228_n6639), .Y(u2__abc_44228_n12673) );
  AND2X2 AND2X2_5382 ( .A(u2__abc_44228_n12675), .B(u2__abc_44228_n6197), .Y(u2__abc_44228_n12677) );
  AND2X2 AND2X2_5383 ( .A(u2__abc_44228_n12678_1), .B(u2__abc_44228_n12676), .Y(u2__abc_44228_n12679) );
  AND2X2 AND2X2_5384 ( .A(u2__abc_44228_n12679), .B(u2__abc_44228_n7547_bF_buf46), .Y(u2__abc_44228_n12680) );
  AND2X2 AND2X2_5385 ( .A(u2__abc_44228_n7548_1_bF_buf47), .B(u2_remHi_298_), .Y(u2__abc_44228_n12681) );
  AND2X2 AND2X2_5386 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n6180), .Y(u2__abc_44228_n12684) );
  AND2X2 AND2X2_5387 ( .A(u2__abc_44228_n12685), .B(u2__abc_44228_n2972_bF_buf21), .Y(u2__abc_44228_n12686_1) );
  AND2X2 AND2X2_5388 ( .A(u2__abc_44228_n12683), .B(u2__abc_44228_n12686_1), .Y(u2__abc_44228_n12687) );
  AND2X2 AND2X2_5389 ( .A(u2__abc_44228_n12688), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_remHi_300__FF_INPUT) );
  AND2X2 AND2X2_539 ( .A(u2__abc_44228_n2995), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n2996) );
  AND2X2 AND2X2_5390 ( .A(u2__abc_44228_n3062_bF_buf70), .B(u2_remHi_301_), .Y(u2__abc_44228_n12690) );
  AND2X2 AND2X2_5391 ( .A(u2__abc_44228_n12678_1), .B(u2__abc_44228_n6644_1), .Y(u2__abc_44228_n12691) );
  AND2X2 AND2X2_5392 ( .A(u2__abc_44228_n12695), .B(u2__abc_44228_n7547_bF_buf45), .Y(u2__abc_44228_n12696) );
  AND2X2 AND2X2_5393 ( .A(u2__abc_44228_n12696), .B(u2__abc_44228_n12693_1), .Y(u2__abc_44228_n12697) );
  AND2X2 AND2X2_5394 ( .A(u2__abc_44228_n7548_1_bF_buf46), .B(u2_remHi_299_), .Y(u2__abc_44228_n12698) );
  AND2X2 AND2X2_5395 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n6174), .Y(u2__abc_44228_n12701) );
  AND2X2 AND2X2_5396 ( .A(u2__abc_44228_n12702), .B(u2__abc_44228_n2972_bF_buf20), .Y(u2__abc_44228_n12703) );
  AND2X2 AND2X2_5397 ( .A(u2__abc_44228_n12700), .B(u2__abc_44228_n12703), .Y(u2__abc_44228_n12704) );
  AND2X2 AND2X2_5398 ( .A(u2__abc_44228_n12705), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_remHi_301__FF_INPUT) );
  AND2X2 AND2X2_5399 ( .A(u2__abc_44228_n3062_bF_buf69), .B(u2_remHi_302_), .Y(u2__abc_44228_n12707) );
  AND2X2 AND2X2_54 ( .A(_abc_64468_n753_bF_buf2), .B(sqrto_53_), .Y(_auto_iopadmap_cc_313_execute_65414_89_) );
  AND2X2 AND2X2_540 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n2996), .Y(u2__abc_44228_n2997) );
  AND2X2 AND2X2_5400 ( .A(u2__abc_44228_n12678_1), .B(u2__abc_44228_n6645), .Y(u2__abc_44228_n12708) );
  AND2X2 AND2X2_5401 ( .A(u2__abc_44228_n12710), .B(u2__abc_44228_n6183), .Y(u2__abc_44228_n12711) );
  AND2X2 AND2X2_5402 ( .A(u2__abc_44228_n12713_1), .B(u2__abc_44228_n7547_bF_buf44), .Y(u2__abc_44228_n12714) );
  AND2X2 AND2X2_5403 ( .A(u2__abc_44228_n12714), .B(u2__abc_44228_n12712), .Y(u2__abc_44228_n12715) );
  AND2X2 AND2X2_5404 ( .A(u2__abc_44228_n7548_1_bF_buf45), .B(u2_remHi_300_), .Y(u2__abc_44228_n12716) );
  AND2X2 AND2X2_5405 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n6156), .Y(u2__abc_44228_n12719) );
  AND2X2 AND2X2_5406 ( .A(u2__abc_44228_n12720), .B(u2__abc_44228_n2972_bF_buf19), .Y(u2__abc_44228_n12721_1) );
  AND2X2 AND2X2_5407 ( .A(u2__abc_44228_n12718), .B(u2__abc_44228_n12721_1), .Y(u2__abc_44228_n12722) );
  AND2X2 AND2X2_5408 ( .A(u2__abc_44228_n12723), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_remHi_302__FF_INPUT) );
  AND2X2 AND2X2_5409 ( .A(u2__abc_44228_n3062_bF_buf68), .B(u2_remHi_303_), .Y(u2__abc_44228_n12725) );
  AND2X2 AND2X2_541 ( .A(u2__abc_44228_n2998), .B(u2__abc_44228_n2999), .Y(u2_cnt_0__FF_INPUT) );
  AND2X2 AND2X2_5410 ( .A(u2__abc_44228_n12730), .B(u2__abc_44228_n7547_bF_buf43), .Y(u2__abc_44228_n12731) );
  AND2X2 AND2X2_5411 ( .A(u2__abc_44228_n12731), .B(u2__abc_44228_n12729), .Y(u2__abc_44228_n12732) );
  AND2X2 AND2X2_5412 ( .A(u2__abc_44228_n7548_1_bF_buf44), .B(u2_remHi_301_), .Y(u2__abc_44228_n12733) );
  AND2X2 AND2X2_5413 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n6163), .Y(u2__abc_44228_n12736) );
  AND2X2 AND2X2_5414 ( .A(u2__abc_44228_n12737_1), .B(u2__abc_44228_n2972_bF_buf18), .Y(u2__abc_44228_n12738) );
  AND2X2 AND2X2_5415 ( .A(u2__abc_44228_n12735), .B(u2__abc_44228_n12738), .Y(u2__abc_44228_n12739) );
  AND2X2 AND2X2_5416 ( .A(u2__abc_44228_n12740), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_remHi_303__FF_INPUT) );
  AND2X2 AND2X2_5417 ( .A(u2__abc_44228_n3062_bF_buf67), .B(u2_remHi_304_), .Y(u2__abc_44228_n12742) );
  AND2X2 AND2X2_5418 ( .A(u2__abc_44228_n12470), .B(u2__abc_44228_n6289), .Y(u2__abc_44228_n12743) );
  AND2X2 AND2X2_5419 ( .A(u2__abc_44228_n12744_1), .B(u2__abc_44228_n6159_1), .Y(u2__abc_44228_n12746) );
  AND2X2 AND2X2_542 ( .A(u2__abc_44228_n2968), .B(u2_cnt_1_), .Y(u2__abc_44228_n3001) );
  AND2X2 AND2X2_5420 ( .A(u2__abc_44228_n12747), .B(u2__abc_44228_n12745), .Y(u2__abc_44228_n12748) );
  AND2X2 AND2X2_5421 ( .A(u2__abc_44228_n12749), .B(u2__abc_44228_n12750), .Y(u2__abc_44228_n12751) );
  AND2X2 AND2X2_5422 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n6149), .Y(u2__abc_44228_n12753) );
  AND2X2 AND2X2_5423 ( .A(u2__abc_44228_n12754), .B(u2__abc_44228_n2972_bF_buf17), .Y(u2__abc_44228_n12755) );
  AND2X2 AND2X2_5424 ( .A(u2__abc_44228_n12752_1), .B(u2__abc_44228_n12755), .Y(u2__abc_44228_n12756) );
  AND2X2 AND2X2_5425 ( .A(u2__abc_44228_n12757), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_remHi_304__FF_INPUT) );
  AND2X2 AND2X2_5426 ( .A(u2__abc_44228_n3062_bF_buf66), .B(u2_remHi_305_), .Y(u2__abc_44228_n12759_1) );
  AND2X2 AND2X2_5427 ( .A(u2__abc_44228_n7548_1_bF_buf42), .B(u2_remHi_303_), .Y(u2__abc_44228_n12760) );
  AND2X2 AND2X2_5428 ( .A(u2__abc_44228_n12747), .B(u2__abc_44228_n6655), .Y(u2__abc_44228_n12763) );
  AND2X2 AND2X2_5429 ( .A(u2__abc_44228_n12766), .B(u2__abc_44228_n12764), .Y(u2__abc_44228_n12767) );
  AND2X2 AND2X2_543 ( .A(u2_cnt_1_), .B(u2_cnt_0_), .Y(u2__abc_44228_n3003) );
  AND2X2 AND2X2_5430 ( .A(u2__abc_44228_n12767), .B(u2__abc_44228_n7547_bF_buf41), .Y(u2__abc_44228_n12768) );
  AND2X2 AND2X2_5431 ( .A(u2__abc_44228_n2983_bF_buf3), .B(u2__abc_44228_n6143), .Y(u2__abc_44228_n12770) );
  AND2X2 AND2X2_5432 ( .A(u2__abc_44228_n12771), .B(u2__abc_44228_n2972_bF_buf16), .Y(u2__abc_44228_n12772) );
  AND2X2 AND2X2_5433 ( .A(u2__abc_44228_n12769_1), .B(u2__abc_44228_n12772), .Y(u2__abc_44228_n12773) );
  AND2X2 AND2X2_5434 ( .A(u2__abc_44228_n12774), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_remHi_305__FF_INPUT) );
  AND2X2 AND2X2_5435 ( .A(u2__abc_44228_n3062_bF_buf65), .B(u2_remHi_306_), .Y(u2__abc_44228_n12776_1) );
  AND2X2 AND2X2_5436 ( .A(u2__abc_44228_n12744_1), .B(u2__abc_44228_n6167), .Y(u2__abc_44228_n12777) );
  AND2X2 AND2X2_5437 ( .A(u2__abc_44228_n12778), .B(u2__abc_44228_n6152), .Y(u2__abc_44228_n12779) );
  AND2X2 AND2X2_5438 ( .A(u2__abc_44228_n12780), .B(u2__abc_44228_n12781), .Y(u2__abc_44228_n12782) );
  AND2X2 AND2X2_5439 ( .A(u2__abc_44228_n12782), .B(u2__abc_44228_n7547_bF_buf40), .Y(u2__abc_44228_n12783) );
  AND2X2 AND2X2_544 ( .A(u2__abc_44228_n3004), .B(u2__abc_44228_n3002), .Y(u2__abc_44228_n3005) );
  AND2X2 AND2X2_5440 ( .A(u2__abc_44228_n7548_1_bF_buf41), .B(u2_remHi_304_), .Y(u2__abc_44228_n12784_1) );
  AND2X2 AND2X2_5441 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n6127), .Y(u2__abc_44228_n12787) );
  AND2X2 AND2X2_5442 ( .A(u2__abc_44228_n12788), .B(u2__abc_44228_n2972_bF_buf15), .Y(u2__abc_44228_n12789) );
  AND2X2 AND2X2_5443 ( .A(u2__abc_44228_n12786), .B(u2__abc_44228_n12789), .Y(u2__abc_44228_n12790) );
  AND2X2 AND2X2_5444 ( .A(u2__abc_44228_n12791_1), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_remHi_306__FF_INPUT) );
  AND2X2 AND2X2_5445 ( .A(u2__abc_44228_n3062_bF_buf64), .B(u2_remHi_307_), .Y(u2__abc_44228_n12793) );
  AND2X2 AND2X2_5446 ( .A(u2__abc_44228_n12798), .B(u2__abc_44228_n7547_bF_buf39), .Y(u2__abc_44228_n12799) );
  AND2X2 AND2X2_5447 ( .A(u2__abc_44228_n12799), .B(u2__abc_44228_n12797), .Y(u2__abc_44228_n12800_1) );
  AND2X2 AND2X2_5448 ( .A(u2__abc_44228_n7548_1_bF_buf40), .B(u2_remHi_305_), .Y(u2__abc_44228_n12801) );
  AND2X2 AND2X2_5449 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n6134), .Y(u2__abc_44228_n12804) );
  AND2X2 AND2X2_545 ( .A(u2__abc_44228_n2996), .B(u2__abc_44228_n3005), .Y(u2__abc_44228_n3006) );
  AND2X2 AND2X2_5450 ( .A(u2__abc_44228_n12805), .B(u2__abc_44228_n2972_bF_buf14), .Y(u2__abc_44228_n12806) );
  AND2X2 AND2X2_5451 ( .A(u2__abc_44228_n12803), .B(u2__abc_44228_n12806), .Y(u2__abc_44228_n12807_1) );
  AND2X2 AND2X2_5452 ( .A(u2__abc_44228_n12808), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_remHi_307__FF_INPUT) );
  AND2X2 AND2X2_5453 ( .A(u2__abc_44228_n3062_bF_buf63), .B(u2_remHi_308_), .Y(u2__abc_44228_n12810) );
  AND2X2 AND2X2_5454 ( .A(u2__abc_44228_n12744_1), .B(u2__abc_44228_n6168), .Y(u2__abc_44228_n12811) );
  AND2X2 AND2X2_5455 ( .A(u2__abc_44228_n12812), .B(u2__abc_44228_n6130), .Y(u2__abc_44228_n12814) );
  AND2X2 AND2X2_5456 ( .A(u2__abc_44228_n12815_1), .B(u2__abc_44228_n12813), .Y(u2__abc_44228_n12816) );
  AND2X2 AND2X2_5457 ( .A(u2__abc_44228_n12816), .B(u2__abc_44228_n7547_bF_buf38), .Y(u2__abc_44228_n12817) );
  AND2X2 AND2X2_5458 ( .A(u2__abc_44228_n7548_1_bF_buf39), .B(u2_remHi_306_), .Y(u2__abc_44228_n12818) );
  AND2X2 AND2X2_5459 ( .A(u2__abc_44228_n2983_bF_buf141), .B(u2__abc_44228_n6120), .Y(u2__abc_44228_n12821) );
  AND2X2 AND2X2_546 ( .A(u2__abc_44228_n3003), .B(u2_cnt_2_), .Y(u2__abc_44228_n3011) );
  AND2X2 AND2X2_5460 ( .A(u2__abc_44228_n12822_1), .B(u2__abc_44228_n2972_bF_buf13), .Y(u2__abc_44228_n12823) );
  AND2X2 AND2X2_5461 ( .A(u2__abc_44228_n12820), .B(u2__abc_44228_n12823), .Y(u2__abc_44228_n12824) );
  AND2X2 AND2X2_5462 ( .A(u2__abc_44228_n12825), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_remHi_308__FF_INPUT) );
  AND2X2 AND2X2_5463 ( .A(u2__abc_44228_n3062_bF_buf62), .B(u2_remHi_309_), .Y(u2__abc_44228_n12827) );
  AND2X2 AND2X2_5464 ( .A(u2__abc_44228_n7548_1_bF_buf38), .B(u2_remHi_307_), .Y(u2__abc_44228_n12828) );
  AND2X2 AND2X2_5465 ( .A(u2__abc_44228_n12815_1), .B(u2__abc_44228_n6664), .Y(u2__abc_44228_n12831) );
  AND2X2 AND2X2_5466 ( .A(u2__abc_44228_n12834), .B(u2__abc_44228_n12832), .Y(u2__abc_44228_n12835) );
  AND2X2 AND2X2_5467 ( .A(u2__abc_44228_n12835), .B(u2__abc_44228_n7547_bF_buf37), .Y(u2__abc_44228_n12836) );
  AND2X2 AND2X2_5468 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n6114), .Y(u2__abc_44228_n12838) );
  AND2X2 AND2X2_5469 ( .A(u2__abc_44228_n12839), .B(u2__abc_44228_n2972_bF_buf12), .Y(u2__abc_44228_n12840_1) );
  AND2X2 AND2X2_547 ( .A(u2__abc_44228_n3013), .B(u2__abc_44228_n2995), .Y(u2__abc_44228_n3014) );
  AND2X2 AND2X2_5470 ( .A(u2__abc_44228_n12837), .B(u2__abc_44228_n12840_1), .Y(u2__abc_44228_n12841) );
  AND2X2 AND2X2_5471 ( .A(u2__abc_44228_n12842), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_remHi_309__FF_INPUT) );
  AND2X2 AND2X2_5472 ( .A(u2__abc_44228_n3062_bF_buf61), .B(u2_remHi_310_), .Y(u2__abc_44228_n12844) );
  AND2X2 AND2X2_5473 ( .A(u2__abc_44228_n12812), .B(u2__abc_44228_n6138), .Y(u2__abc_44228_n12845) );
  AND2X2 AND2X2_5474 ( .A(u2__abc_44228_n12846), .B(u2__abc_44228_n6123), .Y(u2__abc_44228_n12847) );
  AND2X2 AND2X2_5475 ( .A(u2__abc_44228_n12848_1), .B(u2__abc_44228_n12849), .Y(u2__abc_44228_n12850) );
  AND2X2 AND2X2_5476 ( .A(u2__abc_44228_n12850), .B(u2__abc_44228_n7547_bF_buf36), .Y(u2__abc_44228_n12851) );
  AND2X2 AND2X2_5477 ( .A(u2__abc_44228_n7548_1_bF_buf37), .B(u2_remHi_308_), .Y(u2__abc_44228_n12852) );
  AND2X2 AND2X2_5478 ( .A(u2__abc_44228_n2983_bF_buf139), .B(u2__abc_44228_n6104_1), .Y(u2__abc_44228_n12855_1) );
  AND2X2 AND2X2_5479 ( .A(u2__abc_44228_n12856), .B(u2__abc_44228_n2972_bF_buf11), .Y(u2__abc_44228_n12857) );
  AND2X2 AND2X2_548 ( .A(u2__abc_44228_n3014), .B(u2__abc_44228_n3012), .Y(u2__abc_44228_n3015) );
  AND2X2 AND2X2_5480 ( .A(u2__abc_44228_n12854), .B(u2__abc_44228_n12857), .Y(u2__abc_44228_n12858) );
  AND2X2 AND2X2_5481 ( .A(u2__abc_44228_n12859), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_remHi_310__FF_INPUT) );
  AND2X2 AND2X2_5482 ( .A(u2__abc_44228_n3062_bF_buf60), .B(u2_remHi_311_), .Y(u2__abc_44228_n12861) );
  AND2X2 AND2X2_5483 ( .A(u2__abc_44228_n12866), .B(u2__abc_44228_n7547_bF_buf35), .Y(u2__abc_44228_n12867) );
  AND2X2 AND2X2_5484 ( .A(u2__abc_44228_n12867), .B(u2__abc_44228_n12865), .Y(u2__abc_44228_n12868) );
  AND2X2 AND2X2_5485 ( .A(u2__abc_44228_n7548_1_bF_buf36), .B(u2_remHi_309_), .Y(u2__abc_44228_n12869) );
  AND2X2 AND2X2_5486 ( .A(u2__abc_44228_n2983_bF_buf137), .B(u2__abc_44228_n6098), .Y(u2__abc_44228_n12872) );
  AND2X2 AND2X2_5487 ( .A(u2__abc_44228_n12873), .B(u2__abc_44228_n2972_bF_buf10), .Y(u2__abc_44228_n12874) );
  AND2X2 AND2X2_5488 ( .A(u2__abc_44228_n12871_1), .B(u2__abc_44228_n12874), .Y(u2__abc_44228_n12875) );
  AND2X2 AND2X2_5489 ( .A(u2__abc_44228_n12876), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_remHi_311__FF_INPUT) );
  AND2X2 AND2X2_549 ( .A(u2__abc_44228_n3016), .B(u2__abc_44228_n3009), .Y(u2_cnt_2__FF_INPUT) );
  AND2X2 AND2X2_5490 ( .A(u2__abc_44228_n3062_bF_buf59), .B(u2_remHi_312_), .Y(u2__abc_44228_n12878) );
  AND2X2 AND2X2_5491 ( .A(u2__abc_44228_n12744_1), .B(u2__abc_44228_n6169_1), .Y(u2__abc_44228_n12879_1) );
  AND2X2 AND2X2_5492 ( .A(u2__abc_44228_n12880), .B(u2__abc_44228_n6107), .Y(u2__abc_44228_n12881) );
  AND2X2 AND2X2_5493 ( .A(u2__abc_44228_n12882), .B(u2__abc_44228_n12883), .Y(u2__abc_44228_n12884) );
  AND2X2 AND2X2_5494 ( .A(u2__abc_44228_n12884), .B(u2__abc_44228_n7547_bF_buf34), .Y(u2__abc_44228_n12885) );
  AND2X2 AND2X2_5495 ( .A(u2__abc_44228_n7548_1_bF_buf35), .B(u2_remHi_310_), .Y(u2__abc_44228_n12886_1) );
  AND2X2 AND2X2_5496 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n6090), .Y(u2__abc_44228_n12889) );
  AND2X2 AND2X2_5497 ( .A(u2__abc_44228_n12890), .B(u2__abc_44228_n2972_bF_buf9), .Y(u2__abc_44228_n12891) );
  AND2X2 AND2X2_5498 ( .A(u2__abc_44228_n12888), .B(u2__abc_44228_n12891), .Y(u2__abc_44228_n12892) );
  AND2X2 AND2X2_5499 ( .A(u2__abc_44228_n12893), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_remHi_312__FF_INPUT) );
  AND2X2 AND2X2_55 ( .A(_abc_64468_n753_bF_buf1), .B(sqrto_54_), .Y(_auto_iopadmap_cc_313_execute_65414_90_) );
  AND2X2 AND2X2_550 ( .A(u2__abc_44228_n2968), .B(u2_cnt_3_), .Y(u2__abc_44228_n3018) );
  AND2X2 AND2X2_5500 ( .A(u2__abc_44228_n3062_bF_buf58), .B(u2_remHi_313_), .Y(u2__abc_44228_n12895) );
  AND2X2 AND2X2_5501 ( .A(u2__abc_44228_n7548_1_bF_buf34), .B(u2_remHi_311_), .Y(u2__abc_44228_n12896_1) );
  AND2X2 AND2X2_5502 ( .A(u2__abc_44228_n12882), .B(u2__abc_44228_n6674), .Y(u2__abc_44228_n12899) );
  AND2X2 AND2X2_5503 ( .A(u2__abc_44228_n12902), .B(u2__abc_44228_n12900), .Y(u2__abc_44228_n12903_1) );
  AND2X2 AND2X2_5504 ( .A(u2__abc_44228_n12903_1), .B(u2__abc_44228_n7547_bF_buf33), .Y(u2__abc_44228_n12904) );
  AND2X2 AND2X2_5505 ( .A(u2__abc_44228_n2983_bF_buf135), .B(u2__abc_44228_n6084), .Y(u2__abc_44228_n12906) );
  AND2X2 AND2X2_5506 ( .A(u2__abc_44228_n12907), .B(u2__abc_44228_n2972_bF_buf8), .Y(u2__abc_44228_n12908) );
  AND2X2 AND2X2_5507 ( .A(u2__abc_44228_n12905), .B(u2__abc_44228_n12908), .Y(u2__abc_44228_n12909) );
  AND2X2 AND2X2_5508 ( .A(u2__abc_44228_n12910), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_remHi_313__FF_INPUT) );
  AND2X2 AND2X2_5509 ( .A(u2__abc_44228_n3062_bF_buf57), .B(u2_remHi_314_), .Y(u2__abc_44228_n12912) );
  AND2X2 AND2X2_551 ( .A(u2__abc_44228_n3011), .B(u2_cnt_3_), .Y(u2__abc_44228_n3020) );
  AND2X2 AND2X2_5510 ( .A(u2__abc_44228_n12880), .B(u2__abc_44228_n6108), .Y(u2__abc_44228_n12913) );
  AND2X2 AND2X2_5511 ( .A(u2__abc_44228_n12914), .B(u2__abc_44228_n6093), .Y(u2__abc_44228_n12915) );
  AND2X2 AND2X2_5512 ( .A(u2__abc_44228_n12916), .B(u2__abc_44228_n12917), .Y(u2__abc_44228_n12918_1) );
  AND2X2 AND2X2_5513 ( .A(u2__abc_44228_n12918_1), .B(u2__abc_44228_n7547_bF_buf32), .Y(u2__abc_44228_n12919) );
  AND2X2 AND2X2_5514 ( .A(u2__abc_44228_n7548_1_bF_buf33), .B(u2_remHi_312_), .Y(u2__abc_44228_n12920) );
  AND2X2 AND2X2_5515 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n6075), .Y(u2__abc_44228_n12923) );
  AND2X2 AND2X2_5516 ( .A(u2__abc_44228_n12924), .B(u2__abc_44228_n2972_bF_buf7), .Y(u2__abc_44228_n12925) );
  AND2X2 AND2X2_5517 ( .A(u2__abc_44228_n12922), .B(u2__abc_44228_n12925), .Y(u2__abc_44228_n12926) );
  AND2X2 AND2X2_5518 ( .A(u2__abc_44228_n12927_1), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_remHi_314__FF_INPUT) );
  AND2X2 AND2X2_5519 ( .A(u2__abc_44228_n3062_bF_buf56), .B(u2_remHi_315_), .Y(u2__abc_44228_n12929) );
  AND2X2 AND2X2_552 ( .A(u2__abc_44228_n3021), .B(u2__abc_44228_n3019), .Y(u2__abc_44228_n3022) );
  AND2X2 AND2X2_5520 ( .A(u2__abc_44228_n12916), .B(u2__abc_44228_n6679), .Y(u2__abc_44228_n12931) );
  AND2X2 AND2X2_5521 ( .A(u2__abc_44228_n12934_1), .B(u2__abc_44228_n12932), .Y(u2__abc_44228_n12935) );
  AND2X2 AND2X2_5522 ( .A(u2__abc_44228_n12935), .B(u2__abc_44228_n7547_bF_buf31), .Y(u2__abc_44228_n12936) );
  AND2X2 AND2X2_5523 ( .A(u2__abc_44228_n7548_1_bF_buf32), .B(u2_remHi_313_), .Y(u2__abc_44228_n12937) );
  AND2X2 AND2X2_5524 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n6069), .Y(u2__abc_44228_n12940) );
  AND2X2 AND2X2_5525 ( .A(u2__abc_44228_n12941), .B(u2__abc_44228_n2972_bF_buf6), .Y(u2__abc_44228_n12942_1) );
  AND2X2 AND2X2_5526 ( .A(u2__abc_44228_n12939), .B(u2__abc_44228_n12942_1), .Y(u2__abc_44228_n12943) );
  AND2X2 AND2X2_5527 ( .A(u2__abc_44228_n12944), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_remHi_315__FF_INPUT) );
  AND2X2 AND2X2_5528 ( .A(u2__abc_44228_n3062_bF_buf55), .B(u2_remHi_316_), .Y(u2__abc_44228_n12946) );
  AND2X2 AND2X2_5529 ( .A(u2__abc_44228_n12916), .B(u2__abc_44228_n6680), .Y(u2__abc_44228_n12947) );
  AND2X2 AND2X2_553 ( .A(u2__abc_44228_n3022), .B(u2__abc_44228_n2996), .Y(u2__abc_44228_n3023) );
  AND2X2 AND2X2_5530 ( .A(u2__abc_44228_n12949_1), .B(u2__abc_44228_n6078_1), .Y(u2__abc_44228_n12950) );
  AND2X2 AND2X2_5531 ( .A(u2__abc_44228_n12952), .B(u2__abc_44228_n7547_bF_buf30), .Y(u2__abc_44228_n12953) );
  AND2X2 AND2X2_5532 ( .A(u2__abc_44228_n12953), .B(u2__abc_44228_n12951), .Y(u2__abc_44228_n12954) );
  AND2X2 AND2X2_5533 ( .A(u2__abc_44228_n7548_1_bF_buf31), .B(u2_remHi_314_), .Y(u2__abc_44228_n12955) );
  AND2X2 AND2X2_5534 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n6061), .Y(u2__abc_44228_n12958) );
  AND2X2 AND2X2_5535 ( .A(u2__abc_44228_n12959), .B(u2__abc_44228_n2972_bF_buf5), .Y(u2__abc_44228_n12960) );
  AND2X2 AND2X2_5536 ( .A(u2__abc_44228_n12957), .B(u2__abc_44228_n12960), .Y(u2__abc_44228_n12961_1) );
  AND2X2 AND2X2_5537 ( .A(u2__abc_44228_n12962), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_remHi_316__FF_INPUT) );
  AND2X2 AND2X2_5538 ( .A(u2__abc_44228_n3062_bF_buf54), .B(u2_remHi_317_), .Y(u2__abc_44228_n12964) );
  AND2X2 AND2X2_5539 ( .A(u2__abc_44228_n12951), .B(u2__abc_44228_n6687), .Y(u2__abc_44228_n12966) );
  AND2X2 AND2X2_554 ( .A(u2__abc_44228_n2968), .B(u2_cnt_4_), .Y(u2__abc_44228_n3025) );
  AND2X2 AND2X2_5540 ( .A(u2__abc_44228_n12969), .B(u2__abc_44228_n12967), .Y(u2__abc_44228_n12970) );
  AND2X2 AND2X2_5541 ( .A(u2__abc_44228_n12970), .B(u2__abc_44228_n7547_bF_buf29), .Y(u2__abc_44228_n12971) );
  AND2X2 AND2X2_5542 ( .A(u2__abc_44228_n7548_1_bF_buf30), .B(u2_remHi_315_), .Y(u2__abc_44228_n12972) );
  AND2X2 AND2X2_5543 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n6055), .Y(u2__abc_44228_n12975) );
  AND2X2 AND2X2_5544 ( .A(u2__abc_44228_n12976_1), .B(u2__abc_44228_n2972_bF_buf4), .Y(u2__abc_44228_n12977) );
  AND2X2 AND2X2_5545 ( .A(u2__abc_44228_n12974), .B(u2__abc_44228_n12977), .Y(u2__abc_44228_n12978) );
  AND2X2 AND2X2_5546 ( .A(u2__abc_44228_n12979), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_remHi_317__FF_INPUT) );
  AND2X2 AND2X2_5547 ( .A(u2__abc_44228_n3062_bF_buf53), .B(u2_remHi_318_), .Y(u2__abc_44228_n12981) );
  AND2X2 AND2X2_5548 ( .A(u2__abc_44228_n12949_1), .B(u2__abc_44228_n6079), .Y(u2__abc_44228_n12982) );
  AND2X2 AND2X2_5549 ( .A(u2__abc_44228_n12983_1), .B(u2__abc_44228_n6064), .Y(u2__abc_44228_n12984) );
  AND2X2 AND2X2_555 ( .A(u2__abc_44228_n3020), .B(u2_cnt_4_), .Y(u2__abc_44228_n3026) );
  AND2X2 AND2X2_5550 ( .A(u2__abc_44228_n12986), .B(u2__abc_44228_n7547_bF_buf28), .Y(u2__abc_44228_n12987) );
  AND2X2 AND2X2_5551 ( .A(u2__abc_44228_n12987), .B(u2__abc_44228_n12985), .Y(u2__abc_44228_n12988) );
  AND2X2 AND2X2_5552 ( .A(u2__abc_44228_n7548_1_bF_buf29), .B(u2_remHi_316_), .Y(u2__abc_44228_n12989) );
  AND2X2 AND2X2_5553 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n6035), .Y(u2__abc_44228_n12992_1) );
  AND2X2 AND2X2_5554 ( .A(u2__abc_44228_n12993), .B(u2__abc_44228_n2972_bF_buf3), .Y(u2__abc_44228_n12994) );
  AND2X2 AND2X2_5555 ( .A(u2__abc_44228_n12991), .B(u2__abc_44228_n12994), .Y(u2__abc_44228_n12995) );
  AND2X2 AND2X2_5556 ( .A(u2__abc_44228_n12996), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_remHi_318__FF_INPUT) );
  AND2X2 AND2X2_5557 ( .A(u2__abc_44228_n3062_bF_buf52), .B(u2_remHi_319_), .Y(u2__abc_44228_n12998) );
  AND2X2 AND2X2_5558 ( .A(u2__abc_44228_n13003), .B(u2__abc_44228_n7547_bF_buf27), .Y(u2__abc_44228_n13004) );
  AND2X2 AND2X2_5559 ( .A(u2__abc_44228_n13004), .B(u2__abc_44228_n13002), .Y(u2__abc_44228_n13005) );
  AND2X2 AND2X2_556 ( .A(u2__abc_44228_n3028), .B(u2__abc_44228_n2996), .Y(u2__abc_44228_n3029) );
  AND2X2 AND2X2_5560 ( .A(u2__abc_44228_n7548_1_bF_buf28), .B(u2_remHi_317_), .Y(u2__abc_44228_n13006) );
  AND2X2 AND2X2_5561 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n6042), .Y(u2__abc_44228_n13009) );
  AND2X2 AND2X2_5562 ( .A(u2__abc_44228_n13010), .B(u2__abc_44228_n2972_bF_buf2), .Y(u2__abc_44228_n13011) );
  AND2X2 AND2X2_5563 ( .A(u2__abc_44228_n13008), .B(u2__abc_44228_n13011), .Y(u2__abc_44228_n13012) );
  AND2X2 AND2X2_5564 ( .A(u2__abc_44228_n13013), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_remHi_319__FF_INPUT) );
  AND2X2 AND2X2_5565 ( .A(u2__abc_44228_n3062_bF_buf51), .B(u2_remHi_320_), .Y(u2__abc_44228_n13015) );
  AND2X2 AND2X2_5566 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6530), .Y(u2__abc_44228_n13016) );
  AND2X2 AND2X2_5567 ( .A(u2__abc_44228_n13017), .B(u2__abc_44228_n6038), .Y(u2__abc_44228_n13018) );
  AND2X2 AND2X2_5568 ( .A(u2__abc_44228_n13019), .B(u2__abc_44228_n13020), .Y(u2__abc_44228_n13021) );
  AND2X2 AND2X2_5569 ( .A(u2__abc_44228_n13022), .B(u2__abc_44228_n13023), .Y(u2__abc_44228_n13024_1) );
  AND2X2 AND2X2_557 ( .A(u2__abc_44228_n3029), .B(u2__abc_44228_n3027), .Y(u2__abc_44228_n3030) );
  AND2X2 AND2X2_5570 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n6028), .Y(u2__abc_44228_n13026) );
  AND2X2 AND2X2_5571 ( .A(u2__abc_44228_n13027), .B(u2__abc_44228_n2972_bF_buf1), .Y(u2__abc_44228_n13028) );
  AND2X2 AND2X2_5572 ( .A(u2__abc_44228_n13025), .B(u2__abc_44228_n13028), .Y(u2__abc_44228_n13029) );
  AND2X2 AND2X2_5573 ( .A(u2__abc_44228_n13030), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_remHi_320__FF_INPUT) );
  AND2X2 AND2X2_5574 ( .A(u2__abc_44228_n3062_bF_buf50), .B(u2_remHi_321_), .Y(u2__abc_44228_n13032) );
  AND2X2 AND2X2_5575 ( .A(u2__abc_44228_n13019), .B(u2__abc_44228_n6698_1), .Y(u2__abc_44228_n13033) );
  AND2X2 AND2X2_5576 ( .A(u2__abc_44228_n13033), .B(u2__abc_44228_n6045), .Y(u2__abc_44228_n13034) );
  AND2X2 AND2X2_5577 ( .A(u2__abc_44228_n13036), .B(u2__abc_44228_n13035), .Y(u2__abc_44228_n13037) );
  AND2X2 AND2X2_5578 ( .A(u2__abc_44228_n13038), .B(u2__abc_44228_n7547_bF_buf25), .Y(u2__abc_44228_n13039_1) );
  AND2X2 AND2X2_5579 ( .A(u2__abc_44228_n7548_1_bF_buf26), .B(u2_remHi_319_), .Y(u2__abc_44228_n13040) );
  AND2X2 AND2X2_558 ( .A(u2__abc_44228_n2968), .B(u2_cnt_5_), .Y(u2__abc_44228_n3032) );
  AND2X2 AND2X2_5580 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n6022_1), .Y(u2__abc_44228_n13043) );
  AND2X2 AND2X2_5581 ( .A(u2__abc_44228_n13044), .B(u2__abc_44228_n2972_bF_buf0), .Y(u2__abc_44228_n13045) );
  AND2X2 AND2X2_5582 ( .A(u2__abc_44228_n13042), .B(u2__abc_44228_n13045), .Y(u2__abc_44228_n13046_1) );
  AND2X2 AND2X2_5583 ( .A(u2__abc_44228_n13047), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_remHi_321__FF_INPUT) );
  AND2X2 AND2X2_5584 ( .A(u2__abc_44228_n3062_bF_buf49), .B(u2_remHi_322_), .Y(u2__abc_44228_n13049) );
  AND2X2 AND2X2_5585 ( .A(u2__abc_44228_n13019), .B(u2__abc_44228_n6699), .Y(u2__abc_44228_n13050) );
  AND2X2 AND2X2_5586 ( .A(u2__abc_44228_n13052), .B(u2__abc_44228_n6031_1), .Y(u2__abc_44228_n13053) );
  AND2X2 AND2X2_5587 ( .A(u2__abc_44228_n13054), .B(u2__abc_44228_n13055_1), .Y(u2__abc_44228_n13056) );
  AND2X2 AND2X2_5588 ( .A(u2__abc_44228_n13056), .B(u2__abc_44228_n7547_bF_buf24), .Y(u2__abc_44228_n13057) );
  AND2X2 AND2X2_5589 ( .A(u2__abc_44228_n7548_1_bF_buf25), .B(u2_remHi_320_), .Y(u2__abc_44228_n13058) );
  AND2X2 AND2X2_559 ( .A(u2__abc_44228_n3026), .B(u2_cnt_5_), .Y(u2__abc_44228_n3034) );
  AND2X2 AND2X2_5590 ( .A(u2__abc_44228_n2983_bF_buf119), .B(u2__abc_44228_n6006), .Y(u2__abc_44228_n13061) );
  AND2X2 AND2X2_5591 ( .A(u2__abc_44228_n13062_1), .B(u2__abc_44228_n2972_bF_buf107), .Y(u2__abc_44228_n13063) );
  AND2X2 AND2X2_5592 ( .A(u2__abc_44228_n13060), .B(u2__abc_44228_n13063), .Y(u2__abc_44228_n13064) );
  AND2X2 AND2X2_5593 ( .A(u2__abc_44228_n13065), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_remHi_322__FF_INPUT) );
  AND2X2 AND2X2_5594 ( .A(u2__abc_44228_n3062_bF_buf48), .B(u2_remHi_323_), .Y(u2__abc_44228_n13067) );
  AND2X2 AND2X2_5595 ( .A(u2__abc_44228_n13072), .B(u2__abc_44228_n7547_bF_buf23), .Y(u2__abc_44228_n13073) );
  AND2X2 AND2X2_5596 ( .A(u2__abc_44228_n13073), .B(u2__abc_44228_n13071), .Y(u2__abc_44228_n13074) );
  AND2X2 AND2X2_5597 ( .A(u2__abc_44228_n7548_1_bF_buf24), .B(u2_remHi_321_), .Y(u2__abc_44228_n13075) );
  AND2X2 AND2X2_5598 ( .A(u2__abc_44228_n2983_bF_buf117), .B(u2__abc_44228_n6013), .Y(u2__abc_44228_n13078) );
  AND2X2 AND2X2_5599 ( .A(u2__abc_44228_n13079), .B(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n13080) );
  AND2X2 AND2X2_56 ( .A(_abc_64468_n753_bF_buf0), .B(sqrto_55_), .Y(_auto_iopadmap_cc_313_execute_65414_91_) );
  AND2X2 AND2X2_560 ( .A(u2__abc_44228_n3035), .B(u2__abc_44228_n3033), .Y(u2__abc_44228_n3036) );
  AND2X2 AND2X2_5600 ( .A(u2__abc_44228_n13077_1), .B(u2__abc_44228_n13080), .Y(u2__abc_44228_n13081) );
  AND2X2 AND2X2_5601 ( .A(u2__abc_44228_n13082), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_remHi_323__FF_INPUT) );
  AND2X2 AND2X2_5602 ( .A(u2__abc_44228_n3062_bF_buf47), .B(u2_remHi_324_), .Y(u2__abc_44228_n13084) );
  AND2X2 AND2X2_5603 ( .A(u2__abc_44228_n13017), .B(u2__abc_44228_n6047), .Y(u2__abc_44228_n13085) );
  AND2X2 AND2X2_5604 ( .A(u2__abc_44228_n13086), .B(u2__abc_44228_n6009), .Y(u2__abc_44228_n13088_1) );
  AND2X2 AND2X2_5605 ( .A(u2__abc_44228_n13089), .B(u2__abc_44228_n13087), .Y(u2__abc_44228_n13090) );
  AND2X2 AND2X2_5606 ( .A(u2__abc_44228_n13091), .B(u2__abc_44228_n13092), .Y(u2__abc_44228_n13093) );
  AND2X2 AND2X2_5607 ( .A(u2__abc_44228_n2983_bF_buf115), .B(u2__abc_44228_n5999), .Y(u2__abc_44228_n13095_1) );
  AND2X2 AND2X2_5608 ( .A(u2__abc_44228_n13096), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n13097) );
  AND2X2 AND2X2_5609 ( .A(u2__abc_44228_n13094), .B(u2__abc_44228_n13097), .Y(u2__abc_44228_n13098) );
  AND2X2 AND2X2_561 ( .A(u2__abc_44228_n3036), .B(u2__abc_44228_n2996), .Y(u2__abc_44228_n3037) );
  AND2X2 AND2X2_5610 ( .A(u2__abc_44228_n13099), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_remHi_324__FF_INPUT) );
  AND2X2 AND2X2_5611 ( .A(u2__abc_44228_n3062_bF_buf46), .B(u2_remHi_325_), .Y(u2__abc_44228_n13101) );
  AND2X2 AND2X2_5612 ( .A(u2__abc_44228_n13089), .B(u2__abc_44228_n6707_1), .Y(u2__abc_44228_n13102) );
  AND2X2 AND2X2_5613 ( .A(u2__abc_44228_n13106), .B(u2__abc_44228_n7547_bF_buf21), .Y(u2__abc_44228_n13107) );
  AND2X2 AND2X2_5614 ( .A(u2__abc_44228_n13107), .B(u2__abc_44228_n13104), .Y(u2__abc_44228_n13108) );
  AND2X2 AND2X2_5615 ( .A(u2__abc_44228_n7548_1_bF_buf22), .B(u2_remHi_323_), .Y(u2__abc_44228_n13109) );
  AND2X2 AND2X2_5616 ( .A(u2__abc_44228_n2983_bF_buf113), .B(u2__abc_44228_n5993), .Y(u2__abc_44228_n13112) );
  AND2X2 AND2X2_5617 ( .A(u2__abc_44228_n13113), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n13114) );
  AND2X2 AND2X2_5618 ( .A(u2__abc_44228_n13111), .B(u2__abc_44228_n13114), .Y(u2__abc_44228_n13115) );
  AND2X2 AND2X2_5619 ( .A(u2__abc_44228_n13116), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_remHi_325__FF_INPUT) );
  AND2X2 AND2X2_562 ( .A(u2__abc_44228_n3039), .B(u2__abc_44228_n3008), .Y(u2__abc_44228_n3040) );
  AND2X2 AND2X2_5620 ( .A(u2__abc_44228_n3062_bF_buf45), .B(u2_remHi_326_), .Y(u2__abc_44228_n13118) );
  AND2X2 AND2X2_5621 ( .A(u2__abc_44228_n13089), .B(u2__abc_44228_n6708), .Y(u2__abc_44228_n13119_1) );
  AND2X2 AND2X2_5622 ( .A(u2__abc_44228_n13121), .B(u2__abc_44228_n6002), .Y(u2__abc_44228_n13122) );
  AND2X2 AND2X2_5623 ( .A(u2__abc_44228_n13123), .B(u2__abc_44228_n13124), .Y(u2__abc_44228_n13125) );
  AND2X2 AND2X2_5624 ( .A(u2__abc_44228_n13125), .B(u2__abc_44228_n7547_bF_buf20), .Y(u2__abc_44228_n13126_1) );
  AND2X2 AND2X2_5625 ( .A(u2__abc_44228_n7548_1_bF_buf21), .B(u2_remHi_324_), .Y(u2__abc_44228_n13127) );
  AND2X2 AND2X2_5626 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n5983), .Y(u2__abc_44228_n13130) );
  AND2X2 AND2X2_5627 ( .A(u2__abc_44228_n13131), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n13132) );
  AND2X2 AND2X2_5628 ( .A(u2__abc_44228_n13129), .B(u2__abc_44228_n13132), .Y(u2__abc_44228_n13133) );
  AND2X2 AND2X2_5629 ( .A(u2__abc_44228_n13134_1), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_remHi_326__FF_INPUT) );
  AND2X2 AND2X2_563 ( .A(u2__abc_44228_n3034), .B(u2_cnt_6_), .Y(u2__abc_44228_n3042) );
  AND2X2 AND2X2_5630 ( .A(u2__abc_44228_n3062_bF_buf44), .B(u2_remHi_327_), .Y(u2__abc_44228_n13136) );
  AND2X2 AND2X2_5631 ( .A(u2__abc_44228_n13141_1), .B(u2__abc_44228_n7547_bF_buf19), .Y(u2__abc_44228_n13142) );
  AND2X2 AND2X2_5632 ( .A(u2__abc_44228_n13142), .B(u2__abc_44228_n13140), .Y(u2__abc_44228_n13143) );
  AND2X2 AND2X2_5633 ( .A(u2__abc_44228_n7548_1_bF_buf20), .B(u2_remHi_325_), .Y(u2__abc_44228_n13144) );
  AND2X2 AND2X2_5634 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n5977), .Y(u2__abc_44228_n13147) );
  AND2X2 AND2X2_5635 ( .A(u2__abc_44228_n13148), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n13149) );
  AND2X2 AND2X2_5636 ( .A(u2__abc_44228_n13146), .B(u2__abc_44228_n13149), .Y(u2__abc_44228_n13150) );
  AND2X2 AND2X2_5637 ( .A(u2__abc_44228_n13151_1), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_remHi_327__FF_INPUT) );
  AND2X2 AND2X2_5638 ( .A(u2__abc_44228_n3062_bF_buf43), .B(u2_remHi_328_), .Y(u2__abc_44228_n13153) );
  AND2X2 AND2X2_5639 ( .A(u2__abc_44228_n13017), .B(u2__abc_44228_n6048), .Y(u2__abc_44228_n13154) );
  AND2X2 AND2X2_564 ( .A(u2__abc_44228_n3043), .B(u2__abc_44228_n2995), .Y(u2__abc_44228_n3044) );
  AND2X2 AND2X2_5640 ( .A(u2__abc_44228_n13155), .B(u2__abc_44228_n5986), .Y(u2__abc_44228_n13156) );
  AND2X2 AND2X2_5641 ( .A(u2__abc_44228_n13157), .B(u2__abc_44228_n13158_1), .Y(u2__abc_44228_n13159) );
  AND2X2 AND2X2_5642 ( .A(u2__abc_44228_n13160), .B(u2__abc_44228_n13161), .Y(u2__abc_44228_n13162) );
  AND2X2 AND2X2_5643 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n5969), .Y(u2__abc_44228_n13164) );
  AND2X2 AND2X2_5644 ( .A(u2__abc_44228_n13165), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n13166_1) );
  AND2X2 AND2X2_5645 ( .A(u2__abc_44228_n13163), .B(u2__abc_44228_n13166_1), .Y(u2__abc_44228_n13167) );
  AND2X2 AND2X2_5646 ( .A(u2__abc_44228_n13168), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_remHi_328__FF_INPUT) );
  AND2X2 AND2X2_5647 ( .A(u2__abc_44228_n3062_bF_buf42), .B(u2_remHi_329_), .Y(u2__abc_44228_n13170) );
  AND2X2 AND2X2_5648 ( .A(u2__abc_44228_n13157), .B(u2__abc_44228_n6719), .Y(u2__abc_44228_n13171) );
  AND2X2 AND2X2_5649 ( .A(u2__abc_44228_n13171), .B(u2__abc_44228_n5980), .Y(u2__abc_44228_n13172) );
  AND2X2 AND2X2_565 ( .A(u2__abc_44228_n3045), .B(u2__abc_44228_n3041), .Y(u2_cnt_6__FF_INPUT) );
  AND2X2 AND2X2_5650 ( .A(u2__abc_44228_n13174), .B(u2__abc_44228_n13173_1), .Y(u2__abc_44228_n13175) );
  AND2X2 AND2X2_5651 ( .A(u2__abc_44228_n13176), .B(u2__abc_44228_n7547_bF_buf17), .Y(u2__abc_44228_n13177) );
  AND2X2 AND2X2_5652 ( .A(u2__abc_44228_n7548_1_bF_buf18), .B(u2_remHi_327_), .Y(u2__abc_44228_n13178) );
  AND2X2 AND2X2_5653 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n5963), .Y(u2__abc_44228_n13181) );
  AND2X2 AND2X2_5654 ( .A(u2__abc_44228_n13182_1), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n13183) );
  AND2X2 AND2X2_5655 ( .A(u2__abc_44228_n13180), .B(u2__abc_44228_n13183), .Y(u2__abc_44228_n13184) );
  AND2X2 AND2X2_5656 ( .A(u2__abc_44228_n13185), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_remHi_329__FF_INPUT) );
  AND2X2 AND2X2_5657 ( .A(u2__abc_44228_n3062_bF_buf41), .B(u2_remHi_330_), .Y(u2__abc_44228_n13187) );
  AND2X2 AND2X2_5658 ( .A(u2__abc_44228_n13157), .B(u2__abc_44228_n6720), .Y(u2__abc_44228_n13188) );
  AND2X2 AND2X2_5659 ( .A(u2__abc_44228_n13190), .B(u2__abc_44228_n5972), .Y(u2__abc_44228_n13191) );
  AND2X2 AND2X2_566 ( .A(u2_cnt_5_), .B(u2_cnt_6_), .Y(u2__abc_44228_n3048) );
  AND2X2 AND2X2_5660 ( .A(u2__abc_44228_n13192), .B(u2__abc_44228_n13193), .Y(u2__abc_44228_n13194) );
  AND2X2 AND2X2_5661 ( .A(u2__abc_44228_n13194), .B(u2__abc_44228_n7547_bF_buf16), .Y(u2__abc_44228_n13195) );
  AND2X2 AND2X2_5662 ( .A(u2__abc_44228_n7548_1_bF_buf17), .B(u2_remHi_328_), .Y(u2__abc_44228_n13196) );
  AND2X2 AND2X2_5663 ( .A(u2__abc_44228_n2983_bF_buf105), .B(u2__abc_44228_n5954), .Y(u2__abc_44228_n13199) );
  AND2X2 AND2X2_5664 ( .A(u2__abc_44228_n13200), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n13201) );
  AND2X2 AND2X2_5665 ( .A(u2__abc_44228_n13198), .B(u2__abc_44228_n13201), .Y(u2__abc_44228_n13202) );
  AND2X2 AND2X2_5666 ( .A(u2__abc_44228_n13203), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_remHi_330__FF_INPUT) );
  AND2X2 AND2X2_5667 ( .A(u2__abc_44228_n3062_bF_buf40), .B(u2_remHi_331_), .Y(u2__abc_44228_n13205) );
  AND2X2 AND2X2_5668 ( .A(u2__abc_44228_n13210), .B(u2__abc_44228_n7547_bF_buf15), .Y(u2__abc_44228_n13211) );
  AND2X2 AND2X2_5669 ( .A(u2__abc_44228_n13211), .B(u2__abc_44228_n13209), .Y(u2__abc_44228_n13212) );
  AND2X2 AND2X2_567 ( .A(u2__abc_44228_n3026), .B(u2__abc_44228_n3048), .Y(u2__abc_44228_n3049) );
  AND2X2 AND2X2_5670 ( .A(u2__abc_44228_n7548_1_bF_buf16), .B(u2_remHi_329_), .Y(u2__abc_44228_n13213) );
  AND2X2 AND2X2_5671 ( .A(u2__abc_44228_n2983_bF_buf103), .B(u2__abc_44228_n5948_1), .Y(u2__abc_44228_n13216) );
  AND2X2 AND2X2_5672 ( .A(u2__abc_44228_n13217_1), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n13218) );
  AND2X2 AND2X2_5673 ( .A(u2__abc_44228_n13215), .B(u2__abc_44228_n13218), .Y(u2__abc_44228_n13219) );
  AND2X2 AND2X2_5674 ( .A(u2__abc_44228_n13220), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_remHi_331__FF_INPUT) );
  AND2X2 AND2X2_5675 ( .A(u2__abc_44228_n3062_bF_buf39), .B(u2_remHi_332_), .Y(u2__abc_44228_n13222) );
  AND2X2 AND2X2_5676 ( .A(u2__abc_44228_n13155), .B(u2__abc_44228_n5988), .Y(u2__abc_44228_n13223) );
  AND2X2 AND2X2_5677 ( .A(u2__abc_44228_n13224_1), .B(u2__abc_44228_n5957_1), .Y(u2__abc_44228_n13226) );
  AND2X2 AND2X2_5678 ( .A(u2__abc_44228_n13227), .B(u2__abc_44228_n13225), .Y(u2__abc_44228_n13228) );
  AND2X2 AND2X2_5679 ( .A(u2__abc_44228_n13228), .B(u2__abc_44228_n7547_bF_buf14), .Y(u2__abc_44228_n13229) );
  AND2X2 AND2X2_568 ( .A(u2__abc_44228_n3049), .B(ce), .Y(u2__abc_44228_n3050) );
  AND2X2 AND2X2_5680 ( .A(u2__abc_44228_n7548_1_bF_buf15), .B(u2_remHi_330_), .Y(u2__abc_44228_n13230) );
  AND2X2 AND2X2_5681 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n5940), .Y(u2__abc_44228_n13233) );
  AND2X2 AND2X2_5682 ( .A(u2__abc_44228_n13234), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n13235) );
  AND2X2 AND2X2_5683 ( .A(u2__abc_44228_n13232_1), .B(u2__abc_44228_n13235), .Y(u2__abc_44228_n13236) );
  AND2X2 AND2X2_5684 ( .A(u2__abc_44228_n13237), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_remHi_332__FF_INPUT) );
  AND2X2 AND2X2_5685 ( .A(u2__abc_44228_n3062_bF_buf38), .B(u2_remHi_333_), .Y(u2__abc_44228_n13239_1) );
  AND2X2 AND2X2_5686 ( .A(u2__abc_44228_n13227), .B(u2__abc_44228_n6726), .Y(u2__abc_44228_n13240) );
  AND2X2 AND2X2_5687 ( .A(u2__abc_44228_n13240), .B(u2__abc_44228_n5951), .Y(u2__abc_44228_n13241) );
  AND2X2 AND2X2_5688 ( .A(u2__abc_44228_n13243), .B(u2__abc_44228_n13242), .Y(u2__abc_44228_n13244) );
  AND2X2 AND2X2_5689 ( .A(u2__abc_44228_n13245), .B(u2__abc_44228_n7547_bF_buf13), .Y(u2__abc_44228_n13246) );
  AND2X2 AND2X2_569 ( .A(u2__abc_44228_n3051), .B(u2_cnt_7_), .Y(u2__abc_44228_n3052) );
  AND2X2 AND2X2_5690 ( .A(u2__abc_44228_n7548_1_bF_buf14), .B(u2_remHi_331_), .Y(u2__abc_44228_n13247) );
  AND2X2 AND2X2_5691 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n5934), .Y(u2__abc_44228_n13250) );
  AND2X2 AND2X2_5692 ( .A(u2__abc_44228_n13251), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n13252) );
  AND2X2 AND2X2_5693 ( .A(u2__abc_44228_n13249), .B(u2__abc_44228_n13252), .Y(u2__abc_44228_n13253) );
  AND2X2 AND2X2_5694 ( .A(u2__abc_44228_n13254), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_remHi_333__FF_INPUT) );
  AND2X2 AND2X2_5695 ( .A(u2__abc_44228_n3062_bF_buf37), .B(u2_remHi_334_), .Y(u2__abc_44228_n13256) );
  AND2X2 AND2X2_5696 ( .A(u2__abc_44228_n13227), .B(u2__abc_44228_n6727), .Y(u2__abc_44228_n13257) );
  AND2X2 AND2X2_5697 ( .A(u2__abc_44228_n13259), .B(u2__abc_44228_n5943), .Y(u2__abc_44228_n13260) );
  AND2X2 AND2X2_5698 ( .A(u2__abc_44228_n13261), .B(u2__abc_44228_n13262), .Y(u2__abc_44228_n13263_1) );
  AND2X2 AND2X2_5699 ( .A(u2__abc_44228_n13263_1), .B(u2__abc_44228_n7547_bF_buf12), .Y(u2__abc_44228_n13264) );
  AND2X2 AND2X2_57 ( .A(_abc_64468_n753_bF_buf13), .B(sqrto_56_), .Y(_auto_iopadmap_cc_313_execute_65414_92_) );
  AND2X2 AND2X2_570 ( .A(u2__abc_44228_n3050), .B(u2__abc_44228_n3053), .Y(u2__abc_44228_n3054) );
  AND2X2 AND2X2_5700 ( .A(u2__abc_44228_n7548_1_bF_buf13), .B(u2_remHi_332_), .Y(u2__abc_44228_n13265) );
  AND2X2 AND2X2_5701 ( .A(u2__abc_44228_n2983_bF_buf99), .B(u2__abc_44228_n5923), .Y(u2__abc_44228_n13268) );
  AND2X2 AND2X2_5702 ( .A(u2__abc_44228_n13269), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n13270_1) );
  AND2X2 AND2X2_5703 ( .A(u2__abc_44228_n13267), .B(u2__abc_44228_n13270_1), .Y(u2__abc_44228_n13271) );
  AND2X2 AND2X2_5704 ( .A(u2__abc_44228_n13272), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_remHi_334__FF_INPUT) );
  AND2X2 AND2X2_5705 ( .A(u2__abc_44228_n3062_bF_buf36), .B(u2_remHi_335_), .Y(u2__abc_44228_n13274) );
  AND2X2 AND2X2_5706 ( .A(u2__abc_44228_n13279), .B(u2__abc_44228_n7547_bF_buf11), .Y(u2__abc_44228_n13280_1) );
  AND2X2 AND2X2_5707 ( .A(u2__abc_44228_n13280_1), .B(u2__abc_44228_n13278), .Y(u2__abc_44228_n13281) );
  AND2X2 AND2X2_5708 ( .A(u2__abc_44228_n7548_1_bF_buf12), .B(u2_remHi_333_), .Y(u2__abc_44228_n13282) );
  AND2X2 AND2X2_5709 ( .A(u2__abc_44228_n2983_bF_buf97), .B(u2__abc_44228_n5917), .Y(u2__abc_44228_n13285) );
  AND2X2 AND2X2_571 ( .A(u2__abc_44228_n3056), .B(u2__abc_44228_n3047), .Y(u2_cnt_7__FF_INPUT) );
  AND2X2 AND2X2_5710 ( .A(u2__abc_44228_n13286), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n13287_1) );
  AND2X2 AND2X2_5711 ( .A(u2__abc_44228_n13284), .B(u2__abc_44228_n13287_1), .Y(u2__abc_44228_n13288) );
  AND2X2 AND2X2_5712 ( .A(u2__abc_44228_n13289), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_remHi_335__FF_INPUT) );
  AND2X2 AND2X2_5713 ( .A(u2__abc_44228_n3062_bF_buf35), .B(u2_remHi_336_), .Y(u2__abc_44228_n13291) );
  AND2X2 AND2X2_5714 ( .A(u2__abc_44228_n13017), .B(u2__abc_44228_n6049_1), .Y(u2__abc_44228_n13292) );
  AND2X2 AND2X2_5715 ( .A(u2__abc_44228_n13293), .B(u2__abc_44228_n5926), .Y(u2__abc_44228_n13295_1) );
  AND2X2 AND2X2_5716 ( .A(u2__abc_44228_n13296), .B(u2__abc_44228_n13294), .Y(u2__abc_44228_n13297) );
  AND2X2 AND2X2_5717 ( .A(u2__abc_44228_n13298), .B(u2__abc_44228_n13299), .Y(u2__abc_44228_n13300) );
  AND2X2 AND2X2_5718 ( .A(u2__abc_44228_n2983_bF_buf95), .B(u2__abc_44228_n5909), .Y(u2__abc_44228_n13302_1) );
  AND2X2 AND2X2_5719 ( .A(u2__abc_44228_n13303), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n13304) );
  AND2X2 AND2X2_572 ( .A(ce), .B(u2_state_0_), .Y(u2__abc_44228_n3059) );
  AND2X2 AND2X2_5720 ( .A(u2__abc_44228_n13301), .B(u2__abc_44228_n13304), .Y(u2__abc_44228_n13305) );
  AND2X2 AND2X2_5721 ( .A(u2__abc_44228_n13306), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_remHi_336__FF_INPUT) );
  AND2X2 AND2X2_5722 ( .A(u2__abc_44228_n3062_bF_buf34), .B(u2_remHi_337_), .Y(u2__abc_44228_n13308) );
  AND2X2 AND2X2_5723 ( .A(u2__abc_44228_n13296), .B(u2__abc_44228_n6737), .Y(u2__abc_44228_n13310) );
  AND2X2 AND2X2_5724 ( .A(u2__abc_44228_n13313), .B(u2__abc_44228_n13311_1), .Y(u2__abc_44228_n13314) );
  AND2X2 AND2X2_5725 ( .A(u2__abc_44228_n13314), .B(u2__abc_44228_n7547_bF_buf9), .Y(u2__abc_44228_n13315) );
  AND2X2 AND2X2_5726 ( .A(u2__abc_44228_n7548_1_bF_buf10), .B(u2_remHi_335_), .Y(u2__abc_44228_n13316) );
  AND2X2 AND2X2_5727 ( .A(u2__abc_44228_n2983_bF_buf93), .B(u2__abc_44228_n5903), .Y(u2__abc_44228_n13319) );
  AND2X2 AND2X2_5728 ( .A(u2__abc_44228_n13320), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n13321) );
  AND2X2 AND2X2_5729 ( .A(u2__abc_44228_n13318_1), .B(u2__abc_44228_n13321), .Y(u2__abc_44228_n13322) );
  AND2X2 AND2X2_573 ( .A(u2__abc_44228_n3058), .B(u2__abc_44228_n3060), .Y(u2__abc_44228_n3061) );
  AND2X2 AND2X2_5730 ( .A(u2__abc_44228_n13323), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_remHi_337__FF_INPUT) );
  AND2X2 AND2X2_5731 ( .A(u2__abc_44228_n3062_bF_buf33), .B(u2_remHi_338_), .Y(u2__abc_44228_n13325) );
  AND2X2 AND2X2_5732 ( .A(u2__abc_44228_n13293), .B(u2__abc_44228_n5927), .Y(u2__abc_44228_n13326_1) );
  AND2X2 AND2X2_5733 ( .A(u2__abc_44228_n13327), .B(u2__abc_44228_n5912), .Y(u2__abc_44228_n13328) );
  AND2X2 AND2X2_5734 ( .A(u2__abc_44228_n13329), .B(u2__abc_44228_n13330), .Y(u2__abc_44228_n13331) );
  AND2X2 AND2X2_5735 ( .A(u2__abc_44228_n13331), .B(u2__abc_44228_n7547_bF_buf8), .Y(u2__abc_44228_n13332) );
  AND2X2 AND2X2_5736 ( .A(u2__abc_44228_n7548_1_bF_buf9), .B(u2_remHi_336_), .Y(u2__abc_44228_n13333_1) );
  AND2X2 AND2X2_5737 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n5887), .Y(u2__abc_44228_n13336) );
  AND2X2 AND2X2_5738 ( .A(u2__abc_44228_n13337), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n13338) );
  AND2X2 AND2X2_5739 ( .A(u2__abc_44228_n13335), .B(u2__abc_44228_n13338), .Y(u2__abc_44228_n13339) );
  AND2X2 AND2X2_574 ( .A(u2__abc_44228_n3062_bF_buf92), .B(u2_remHi_0_), .Y(u2__abc_44228_n3063) );
  AND2X2 AND2X2_5740 ( .A(u2__abc_44228_n13340), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_remHi_338__FF_INPUT) );
  AND2X2 AND2X2_5741 ( .A(u2__abc_44228_n3062_bF_buf32), .B(u2_remHi_339_), .Y(u2__abc_44228_n13342) );
  AND2X2 AND2X2_5742 ( .A(u2__abc_44228_n13347), .B(u2__abc_44228_n7547_bF_buf7), .Y(u2__abc_44228_n13348) );
  AND2X2 AND2X2_5743 ( .A(u2__abc_44228_n13348), .B(u2__abc_44228_n13346), .Y(u2__abc_44228_n13349) );
  AND2X2 AND2X2_5744 ( .A(u2__abc_44228_n7548_1_bF_buf8), .B(u2_remHi_337_), .Y(u2__abc_44228_n13350) );
  AND2X2 AND2X2_5745 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n5894), .Y(u2__abc_44228_n13353) );
  AND2X2 AND2X2_5746 ( .A(u2__abc_44228_n13354), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n13355) );
  AND2X2 AND2X2_5747 ( .A(u2__abc_44228_n13352), .B(u2__abc_44228_n13355), .Y(u2__abc_44228_n13356) );
  AND2X2 AND2X2_5748 ( .A(u2__abc_44228_n13357), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_remHi_339__FF_INPUT) );
  AND2X2 AND2X2_5749 ( .A(u2__abc_44228_n3062_bF_buf31), .B(u2_remHi_340_), .Y(u2__abc_44228_n13359_1) );
  AND2X2 AND2X2_575 ( .A(u2__abc_44228_n3065), .B(u2__abc_44228_n3068), .Y(u2__abc_44228_n3069) );
  AND2X2 AND2X2_5750 ( .A(u2__abc_44228_n13293), .B(u2__abc_44228_n5928), .Y(u2__abc_44228_n13360) );
  AND2X2 AND2X2_5751 ( .A(u2__abc_44228_n13361), .B(u2__abc_44228_n5890), .Y(u2__abc_44228_n13363) );
  AND2X2 AND2X2_5752 ( .A(u2__abc_44228_n13364), .B(u2__abc_44228_n13362), .Y(u2__abc_44228_n13365) );
  AND2X2 AND2X2_5753 ( .A(u2__abc_44228_n13365), .B(u2__abc_44228_n7547_bF_buf6), .Y(u2__abc_44228_n13366_1) );
  AND2X2 AND2X2_5754 ( .A(u2__abc_44228_n7548_1_bF_buf7), .B(u2_remHi_338_), .Y(u2__abc_44228_n13367) );
  AND2X2 AND2X2_5755 ( .A(u2__abc_44228_n2983_bF_buf89), .B(u2__abc_44228_n5880), .Y(u2__abc_44228_n13370) );
  AND2X2 AND2X2_5756 ( .A(u2__abc_44228_n13371), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n13372) );
  AND2X2 AND2X2_5757 ( .A(u2__abc_44228_n13369), .B(u2__abc_44228_n13372), .Y(u2__abc_44228_n13373) );
  AND2X2 AND2X2_5758 ( .A(u2__abc_44228_n13374), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_remHi_340__FF_INPUT) );
  AND2X2 AND2X2_5759 ( .A(u2__abc_44228_n3062_bF_buf30), .B(u2_remHi_341_), .Y(u2__abc_44228_n13376) );
  AND2X2 AND2X2_576 ( .A(u2__abc_44228_n3069), .B(u2_remHiShift_0_), .Y(u2__abc_44228_n3070) );
  AND2X2 AND2X2_5760 ( .A(u2__abc_44228_n13364), .B(u2__abc_44228_n6746), .Y(u2__abc_44228_n13377) );
  AND2X2 AND2X2_5761 ( .A(u2__abc_44228_n13377), .B(u2__abc_44228_n5897), .Y(u2__abc_44228_n13378) );
  AND2X2 AND2X2_5762 ( .A(u2__abc_44228_n13380), .B(u2__abc_44228_n13379), .Y(u2__abc_44228_n13381) );
  AND2X2 AND2X2_5763 ( .A(u2__abc_44228_n13382_1), .B(u2__abc_44228_n7547_bF_buf5), .Y(u2__abc_44228_n13383) );
  AND2X2 AND2X2_5764 ( .A(u2__abc_44228_n7548_1_bF_buf6), .B(u2_remHi_339_), .Y(u2__abc_44228_n13384) );
  AND2X2 AND2X2_5765 ( .A(u2__abc_44228_n2983_bF_buf87), .B(u2__abc_44228_n5874), .Y(u2__abc_44228_n13387) );
  AND2X2 AND2X2_5766 ( .A(u2__abc_44228_n13388), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n13389) );
  AND2X2 AND2X2_5767 ( .A(u2__abc_44228_n13386), .B(u2__abc_44228_n13389), .Y(u2__abc_44228_n13390_1) );
  AND2X2 AND2X2_5768 ( .A(u2__abc_44228_n13391), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_remHi_341__FF_INPUT) );
  AND2X2 AND2X2_5769 ( .A(u2__abc_44228_n3062_bF_buf29), .B(u2_remHi_342_), .Y(u2__abc_44228_n13393) );
  AND2X2 AND2X2_577 ( .A(u2__abc_44228_n3073), .B(u2__abc_44228_n3075), .Y(u2__abc_44228_n3076) );
  AND2X2 AND2X2_5770 ( .A(u2__abc_44228_n13364), .B(u2__abc_44228_n6747), .Y(u2__abc_44228_n13394) );
  AND2X2 AND2X2_5771 ( .A(u2__abc_44228_n13396), .B(u2__abc_44228_n5883_1), .Y(u2__abc_44228_n13397_1) );
  AND2X2 AND2X2_5772 ( .A(u2__abc_44228_n13398), .B(u2__abc_44228_n13399), .Y(u2__abc_44228_n13400) );
  AND2X2 AND2X2_5773 ( .A(u2__abc_44228_n13400), .B(u2__abc_44228_n7547_bF_buf4), .Y(u2__abc_44228_n13401) );
  AND2X2 AND2X2_5774 ( .A(u2__abc_44228_n7548_1_bF_buf5), .B(u2_remHi_340_), .Y(u2__abc_44228_n13402) );
  AND2X2 AND2X2_5775 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n5850), .Y(u2__abc_44228_n13405) );
  AND2X2 AND2X2_5776 ( .A(u2__abc_44228_n13406), .B(u2__abc_44228_n2972_bF_buf87), .Y(u2__abc_44228_n13407_1) );
  AND2X2 AND2X2_5777 ( .A(u2__abc_44228_n13404), .B(u2__abc_44228_n13407_1), .Y(u2__abc_44228_n13408) );
  AND2X2 AND2X2_5778 ( .A(u2__abc_44228_n13409), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_remHi_342__FF_INPUT) );
  AND2X2 AND2X2_5779 ( .A(u2__abc_44228_n3062_bF_buf28), .B(u2_remHi_343_), .Y(u2__abc_44228_n13411) );
  AND2X2 AND2X2_578 ( .A(u2__abc_44228_n3077), .B(u2_remHi_0_), .Y(u2__abc_44228_n3078) );
  AND2X2 AND2X2_5780 ( .A(u2__abc_44228_n13416), .B(u2__abc_44228_n7547_bF_buf3), .Y(u2__abc_44228_n13417) );
  AND2X2 AND2X2_5781 ( .A(u2__abc_44228_n13417), .B(u2__abc_44228_n13415), .Y(u2__abc_44228_n13418) );
  AND2X2 AND2X2_5782 ( .A(u2__abc_44228_n7548_1_bF_buf4), .B(u2_remHi_341_), .Y(u2__abc_44228_n13419) );
  AND2X2 AND2X2_5783 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n5844), .Y(u2__abc_44228_n13422_1) );
  AND2X2 AND2X2_5784 ( .A(u2__abc_44228_n13423), .B(u2__abc_44228_n2972_bF_buf86), .Y(u2__abc_44228_n13424) );
  AND2X2 AND2X2_5785 ( .A(u2__abc_44228_n13421), .B(u2__abc_44228_n13424), .Y(u2__abc_44228_n13425) );
  AND2X2 AND2X2_5786 ( .A(u2__abc_44228_n13426), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_remHi_343__FF_INPUT) );
  AND2X2 AND2X2_5787 ( .A(u2__abc_44228_n3062_bF_buf27), .B(u2_remHi_344_), .Y(u2__abc_44228_n13428) );
  AND2X2 AND2X2_5788 ( .A(u2__abc_44228_n13293), .B(u2__abc_44228_n5929), .Y(u2__abc_44228_n13429_1) );
  AND2X2 AND2X2_5789 ( .A(u2__abc_44228_n13430), .B(u2__abc_44228_n5853), .Y(u2__abc_44228_n13431) );
  AND2X2 AND2X2_579 ( .A(u2__abc_44228_n3079), .B(u2__abc_44228_n3080), .Y(u2__abc_44228_n3081) );
  AND2X2 AND2X2_5790 ( .A(u2__abc_44228_n13432), .B(u2__abc_44228_n13433), .Y(u2__abc_44228_n13434) );
  AND2X2 AND2X2_5791 ( .A(u2__abc_44228_n13434), .B(u2__abc_44228_n7547_bF_buf2), .Y(u2__abc_44228_n13435) );
  AND2X2 AND2X2_5792 ( .A(u2__abc_44228_n7548_1_bF_buf3), .B(u2_remHi_342_), .Y(u2__abc_44228_n13436) );
  AND2X2 AND2X2_5793 ( .A(u2__abc_44228_n2983_bF_buf83), .B(u2__abc_44228_n5864), .Y(u2__abc_44228_n13439) );
  AND2X2 AND2X2_5794 ( .A(u2__abc_44228_n13440), .B(u2__abc_44228_n2972_bF_buf85), .Y(u2__abc_44228_n13441) );
  AND2X2 AND2X2_5795 ( .A(u2__abc_44228_n13438_1), .B(u2__abc_44228_n13441), .Y(u2__abc_44228_n13442) );
  AND2X2 AND2X2_5796 ( .A(u2__abc_44228_n13443), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_remHi_344__FF_INPUT) );
  AND2X2 AND2X2_5797 ( .A(u2__abc_44228_n3062_bF_buf26), .B(u2_remHi_345_), .Y(u2__abc_44228_n13445_1) );
  AND2X2 AND2X2_5798 ( .A(u2__abc_44228_n13432), .B(u2__abc_44228_n6756), .Y(u2__abc_44228_n13447) );
  AND2X2 AND2X2_5799 ( .A(u2__abc_44228_n13450), .B(u2__abc_44228_n13448), .Y(u2__abc_44228_n13451) );
  AND2X2 AND2X2_58 ( .A(_abc_64468_n753_bF_buf12), .B(sqrto_57_), .Y(_auto_iopadmap_cc_313_execute_65414_93_) );
  AND2X2 AND2X2_580 ( .A(u2__abc_44228_n3081), .B(u2__abc_44228_n3076), .Y(u2__abc_44228_n3082) );
  AND2X2 AND2X2_5800 ( .A(u2__abc_44228_n13451), .B(u2__abc_44228_n7547_bF_buf1), .Y(u2__abc_44228_n13452) );
  AND2X2 AND2X2_5801 ( .A(u2__abc_44228_n7548_1_bF_buf2), .B(u2_remHi_343_), .Y(u2__abc_44228_n13453_1) );
  AND2X2 AND2X2_5802 ( .A(u2__abc_44228_n2983_bF_buf81), .B(u2__abc_44228_n5858), .Y(u2__abc_44228_n13456) );
  AND2X2 AND2X2_5803 ( .A(u2__abc_44228_n13457), .B(u2__abc_44228_n2972_bF_buf84), .Y(u2__abc_44228_n13458) );
  AND2X2 AND2X2_5804 ( .A(u2__abc_44228_n13455), .B(u2__abc_44228_n13458), .Y(u2__abc_44228_n13459) );
  AND2X2 AND2X2_5805 ( .A(u2__abc_44228_n13460_1), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_remHi_345__FF_INPUT) );
  AND2X2 AND2X2_5806 ( .A(u2__abc_44228_n3062_bF_buf25), .B(u2_remHi_346_), .Y(u2__abc_44228_n13462) );
  AND2X2 AND2X2_5807 ( .A(u2__abc_44228_n13430), .B(u2__abc_44228_n5854_1), .Y(u2__abc_44228_n13463) );
  AND2X2 AND2X2_5808 ( .A(u2__abc_44228_n13464), .B(u2__abc_44228_n5867), .Y(u2__abc_44228_n13465) );
  AND2X2 AND2X2_5809 ( .A(u2__abc_44228_n13466), .B(u2__abc_44228_n13467), .Y(u2__abc_44228_n13468) );
  AND2X2 AND2X2_581 ( .A(u2__abc_44228_n3071), .B(u2__abc_44228_n3082), .Y(u2__abc_44228_n3083) );
  AND2X2 AND2X2_5810 ( .A(u2__abc_44228_n13468), .B(u2__abc_44228_n7547_bF_buf0), .Y(u2__abc_44228_n13469) );
  AND2X2 AND2X2_5811 ( .A(u2__abc_44228_n7548_1_bF_buf1), .B(u2_remHi_344_), .Y(u2__abc_44228_n13470) );
  AND2X2 AND2X2_5812 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n5828), .Y(u2__abc_44228_n13473) );
  AND2X2 AND2X2_5813 ( .A(u2__abc_44228_n13474), .B(u2__abc_44228_n2972_bF_buf83), .Y(u2__abc_44228_n13475) );
  AND2X2 AND2X2_5814 ( .A(u2__abc_44228_n13472_1), .B(u2__abc_44228_n13475), .Y(u2__abc_44228_n13476) );
  AND2X2 AND2X2_5815 ( .A(u2__abc_44228_n13477), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_remHi_346__FF_INPUT) );
  AND2X2 AND2X2_5816 ( .A(u2__abc_44228_n3062_bF_buf24), .B(u2_remHi_347_), .Y(u2__abc_44228_n13479_1) );
  AND2X2 AND2X2_5817 ( .A(u2__abc_44228_n13466), .B(u2__abc_44228_n6761_1), .Y(u2__abc_44228_n13481) );
  AND2X2 AND2X2_5818 ( .A(u2__abc_44228_n13484), .B(u2__abc_44228_n13482), .Y(u2__abc_44228_n13485) );
  AND2X2 AND2X2_5819 ( .A(u2__abc_44228_n13485), .B(u2__abc_44228_n7547_bF_buf57), .Y(u2__abc_44228_n13486) );
  AND2X2 AND2X2_582 ( .A(u2__abc_44228_n3075), .B(u2__abc_44228_n3078), .Y(u2__abc_44228_n3085) );
  AND2X2 AND2X2_5820 ( .A(u2__abc_44228_n7548_1_bF_buf0), .B(u2_remHi_345_), .Y(u2__abc_44228_n13487_1) );
  AND2X2 AND2X2_5821 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n5835), .Y(u2__abc_44228_n13490) );
  AND2X2 AND2X2_5822 ( .A(u2__abc_44228_n13491), .B(u2__abc_44228_n2972_bF_buf82), .Y(u2__abc_44228_n13492) );
  AND2X2 AND2X2_5823 ( .A(u2__abc_44228_n13489), .B(u2__abc_44228_n13492), .Y(u2__abc_44228_n13493) );
  AND2X2 AND2X2_5824 ( .A(u2__abc_44228_n13494_1), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_remHi_347__FF_INPUT) );
  AND2X2 AND2X2_5825 ( .A(u2__abc_44228_n3062_bF_buf23), .B(u2_remHi_348_), .Y(u2__abc_44228_n13496) );
  AND2X2 AND2X2_5826 ( .A(u2__abc_44228_n13466), .B(u2__abc_44228_n6762), .Y(u2__abc_44228_n13497) );
  AND2X2 AND2X2_5827 ( .A(u2__abc_44228_n13499), .B(u2__abc_44228_n5831), .Y(u2__abc_44228_n13501) );
  AND2X2 AND2X2_5828 ( .A(u2__abc_44228_n13502), .B(u2__abc_44228_n13500), .Y(u2__abc_44228_n13503_1) );
  AND2X2 AND2X2_5829 ( .A(u2__abc_44228_n13503_1), .B(u2__abc_44228_n7547_bF_buf56), .Y(u2__abc_44228_n13504) );
  AND2X2 AND2X2_583 ( .A(u2__abc_44228_n3089), .B(u2__abc_44228_n3091), .Y(u2__abc_44228_n3092) );
  AND2X2 AND2X2_5830 ( .A(u2__abc_44228_n7548_1_bF_buf57), .B(u2_remHi_346_), .Y(u2__abc_44228_n13505) );
  AND2X2 AND2X2_5831 ( .A(u2__abc_44228_n2983_bF_buf77), .B(u2__abc_44228_n5821), .Y(u2__abc_44228_n13508) );
  AND2X2 AND2X2_5832 ( .A(u2__abc_44228_n13509), .B(u2__abc_44228_n2972_bF_buf81), .Y(u2__abc_44228_n13510_1) );
  AND2X2 AND2X2_5833 ( .A(u2__abc_44228_n13507), .B(u2__abc_44228_n13510_1), .Y(u2__abc_44228_n13511) );
  AND2X2 AND2X2_5834 ( .A(u2__abc_44228_n13512), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_remHi_348__FF_INPUT) );
  AND2X2 AND2X2_5835 ( .A(u2__abc_44228_n3062_bF_buf22), .B(u2_remHi_349_), .Y(u2__abc_44228_n13514) );
  AND2X2 AND2X2_5836 ( .A(u2__abc_44228_n13502), .B(u2__abc_44228_n6769), .Y(u2__abc_44228_n13515) );
  AND2X2 AND2X2_5837 ( .A(u2__abc_44228_n13519), .B(u2__abc_44228_n7547_bF_buf55), .Y(u2__abc_44228_n13520) );
  AND2X2 AND2X2_5838 ( .A(u2__abc_44228_n13520), .B(u2__abc_44228_n13517), .Y(u2__abc_44228_n13521) );
  AND2X2 AND2X2_5839 ( .A(u2__abc_44228_n7548_1_bF_buf56), .B(u2_remHi_347_), .Y(u2__abc_44228_n13522) );
  AND2X2 AND2X2_584 ( .A(u2__abc_44228_n3094), .B(u2__abc_44228_n3096), .Y(u2__abc_44228_n3097) );
  AND2X2 AND2X2_5840 ( .A(u2__abc_44228_n2983_bF_buf75), .B(u2__abc_44228_n5815), .Y(u2__abc_44228_n13525_1) );
  AND2X2 AND2X2_5841 ( .A(u2__abc_44228_n13526), .B(u2__abc_44228_n2972_bF_buf80), .Y(u2__abc_44228_n13527) );
  AND2X2 AND2X2_5842 ( .A(u2__abc_44228_n13524), .B(u2__abc_44228_n13527), .Y(u2__abc_44228_n13528) );
  AND2X2 AND2X2_5843 ( .A(u2__abc_44228_n13529), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_remHi_349__FF_INPUT) );
  AND2X2 AND2X2_5844 ( .A(u2__abc_44228_n3062_bF_buf21), .B(u2_remHi_350_), .Y(u2__abc_44228_n13531) );
  AND2X2 AND2X2_5845 ( .A(u2__abc_44228_n13502), .B(u2__abc_44228_n6770_1), .Y(u2__abc_44228_n13532) );
  AND2X2 AND2X2_5846 ( .A(u2__abc_44228_n13534), .B(u2__abc_44228_n5824), .Y(u2__abc_44228_n13535_1) );
  AND2X2 AND2X2_5847 ( .A(u2__abc_44228_n13537), .B(u2__abc_44228_n7547_bF_buf54), .Y(u2__abc_44228_n13538) );
  AND2X2 AND2X2_5848 ( .A(u2__abc_44228_n13538), .B(u2__abc_44228_n13536), .Y(u2__abc_44228_n13539) );
  AND2X2 AND2X2_5849 ( .A(u2__abc_44228_n7548_1_bF_buf55), .B(u2_remHi_348_), .Y(u2__abc_44228_n13540) );
  AND2X2 AND2X2_585 ( .A(u2__abc_44228_n3092), .B(u2__abc_44228_n3097), .Y(u2__abc_44228_n3098) );
  AND2X2 AND2X2_5850 ( .A(u2__abc_44228_n2983_bF_buf73), .B(u2__abc_44228_n5803), .Y(u2__abc_44228_n13543) );
  AND2X2 AND2X2_5851 ( .A(u2__abc_44228_n13544), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n13545) );
  AND2X2 AND2X2_5852 ( .A(u2__abc_44228_n13542_1), .B(u2__abc_44228_n13545), .Y(u2__abc_44228_n13546) );
  AND2X2 AND2X2_5853 ( .A(u2__abc_44228_n13547), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_remHi_350__FF_INPUT) );
  AND2X2 AND2X2_5854 ( .A(u2__abc_44228_n3062_bF_buf20), .B(u2_remHi_351_), .Y(u2__abc_44228_n13549) );
  AND2X2 AND2X2_5855 ( .A(u2__abc_44228_n13554), .B(u2__abc_44228_n7547_bF_buf53), .Y(u2__abc_44228_n13555) );
  AND2X2 AND2X2_5856 ( .A(u2__abc_44228_n13555), .B(u2__abc_44228_n13553), .Y(u2__abc_44228_n13556) );
  AND2X2 AND2X2_5857 ( .A(u2__abc_44228_n7548_1_bF_buf54), .B(u2_remHi_349_), .Y(u2__abc_44228_n13557_1) );
  AND2X2 AND2X2_5858 ( .A(u2__abc_44228_n2983_bF_buf71), .B(u2__abc_44228_n5797), .Y(u2__abc_44228_n13560) );
  AND2X2 AND2X2_5859 ( .A(u2__abc_44228_n13561), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n13562) );
  AND2X2 AND2X2_586 ( .A(u2__abc_44228_n3099), .B(u2_remHi_3_), .Y(u2__abc_44228_n3100) );
  AND2X2 AND2X2_5860 ( .A(u2__abc_44228_n13559), .B(u2__abc_44228_n13562), .Y(u2__abc_44228_n13563) );
  AND2X2 AND2X2_5861 ( .A(u2__abc_44228_n13564), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_remHi_351__FF_INPUT) );
  AND2X2 AND2X2_5862 ( .A(u2__abc_44228_n3062_bF_buf19), .B(u2_remHi_352_), .Y(u2__abc_44228_n13566_1) );
  AND2X2 AND2X2_5863 ( .A(u2__abc_44228_n13017), .B(u2__abc_44228_n6050), .Y(u2__abc_44228_n13567) );
  AND2X2 AND2X2_5864 ( .A(u2__abc_44228_n13568), .B(u2__abc_44228_n5806), .Y(u2__abc_44228_n13569) );
  AND2X2 AND2X2_5865 ( .A(u2__abc_44228_n13570), .B(u2__abc_44228_n13571), .Y(u2__abc_44228_n13572) );
  AND2X2 AND2X2_5866 ( .A(u2__abc_44228_n13573_1), .B(u2__abc_44228_n13574), .Y(u2__abc_44228_n13575) );
  AND2X2 AND2X2_5867 ( .A(u2__abc_44228_n2983_bF_buf69), .B(u2__abc_44228_n5789), .Y(u2__abc_44228_n13577) );
  AND2X2 AND2X2_5868 ( .A(u2__abc_44228_n13578), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n13579) );
  AND2X2 AND2X2_5869 ( .A(u2__abc_44228_n13576), .B(u2__abc_44228_n13579), .Y(u2__abc_44228_n13580) );
  AND2X2 AND2X2_587 ( .A(u2__abc_44228_n3101), .B(u2__abc_44228_n3102), .Y(u2__abc_44228_n3103) );
  AND2X2 AND2X2_5870 ( .A(u2__abc_44228_n13581_1), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_remHi_352__FF_INPUT) );
  AND2X2 AND2X2_5871 ( .A(u2__abc_44228_n3062_bF_buf18), .B(u2_remHi_353_), .Y(u2__abc_44228_n13583) );
  AND2X2 AND2X2_5872 ( .A(u2__abc_44228_n13570), .B(u2__abc_44228_n6779_1), .Y(u2__abc_44228_n13585) );
  AND2X2 AND2X2_5873 ( .A(u2__abc_44228_n13588_1), .B(u2__abc_44228_n13586), .Y(u2__abc_44228_n13589) );
  AND2X2 AND2X2_5874 ( .A(u2__abc_44228_n13589), .B(u2__abc_44228_n7547_bF_buf51), .Y(u2__abc_44228_n13590) );
  AND2X2 AND2X2_5875 ( .A(u2__abc_44228_n7548_1_bF_buf52), .B(u2_remHi_351_), .Y(u2__abc_44228_n13591) );
  AND2X2 AND2X2_5876 ( .A(u2__abc_44228_n2983_bF_buf67), .B(u2__abc_44228_n5783_1), .Y(u2__abc_44228_n13594) );
  AND2X2 AND2X2_5877 ( .A(u2__abc_44228_n13595), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n13596) );
  AND2X2 AND2X2_5878 ( .A(u2__abc_44228_n13593), .B(u2__abc_44228_n13596), .Y(u2__abc_44228_n13597) );
  AND2X2 AND2X2_5879 ( .A(u2__abc_44228_n13598), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_remHi_353__FF_INPUT) );
  AND2X2 AND2X2_588 ( .A(u2__abc_44228_n3104), .B(u2_remHi_2_), .Y(u2__abc_44228_n3105) );
  AND2X2 AND2X2_5880 ( .A(u2__abc_44228_n3062_bF_buf17), .B(u2_remHi_354_), .Y(u2__abc_44228_n13600) );
  AND2X2 AND2X2_5881 ( .A(u2__abc_44228_n13568), .B(u2__abc_44228_n5807), .Y(u2__abc_44228_n13601) );
  AND2X2 AND2X2_5882 ( .A(u2__abc_44228_n13602), .B(u2__abc_44228_n5792), .Y(u2__abc_44228_n13603) );
  AND2X2 AND2X2_5883 ( .A(u2__abc_44228_n13604), .B(u2__abc_44228_n13605), .Y(u2__abc_44228_n13606_1) );
  AND2X2 AND2X2_5884 ( .A(u2__abc_44228_n13606_1), .B(u2__abc_44228_n7547_bF_buf50), .Y(u2__abc_44228_n13607) );
  AND2X2 AND2X2_5885 ( .A(u2__abc_44228_n7548_1_bF_buf51), .B(u2_remHi_352_), .Y(u2__abc_44228_n13608) );
  AND2X2 AND2X2_5886 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n5767), .Y(u2__abc_44228_n13611) );
  AND2X2 AND2X2_5887 ( .A(u2__abc_44228_n13612), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n13613) );
  AND2X2 AND2X2_5888 ( .A(u2__abc_44228_n13610), .B(u2__abc_44228_n13613), .Y(u2__abc_44228_n13614_1) );
  AND2X2 AND2X2_5889 ( .A(u2__abc_44228_n13615), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_remHi_354__FF_INPUT) );
  AND2X2 AND2X2_589 ( .A(u2__abc_44228_n3106), .B(u2__abc_44228_n3107), .Y(u2__abc_44228_n3108) );
  AND2X2 AND2X2_5890 ( .A(u2__abc_44228_n3062_bF_buf16), .B(u2_remHi_355_), .Y(u2__abc_44228_n13617) );
  AND2X2 AND2X2_5891 ( .A(u2__abc_44228_n13622), .B(u2__abc_44228_n7547_bF_buf49), .Y(u2__abc_44228_n13623) );
  AND2X2 AND2X2_5892 ( .A(u2__abc_44228_n13623), .B(u2__abc_44228_n13621_1), .Y(u2__abc_44228_n13624) );
  AND2X2 AND2X2_5893 ( .A(u2__abc_44228_n7548_1_bF_buf50), .B(u2_remHi_353_), .Y(u2__abc_44228_n13625) );
  AND2X2 AND2X2_5894 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n5774_1), .Y(u2__abc_44228_n13628) );
  AND2X2 AND2X2_5895 ( .A(u2__abc_44228_n13629), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n13630_1) );
  AND2X2 AND2X2_5896 ( .A(u2__abc_44228_n13627), .B(u2__abc_44228_n13630_1), .Y(u2__abc_44228_n13631) );
  AND2X2 AND2X2_5897 ( .A(u2__abc_44228_n13632), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_remHi_355__FF_INPUT) );
  AND2X2 AND2X2_5898 ( .A(u2__abc_44228_n3062_bF_buf15), .B(u2_remHi_356_), .Y(u2__abc_44228_n13634) );
  AND2X2 AND2X2_5899 ( .A(u2__abc_44228_n13568), .B(u2__abc_44228_n5808), .Y(u2__abc_44228_n13635) );
  AND2X2 AND2X2_59 ( .A(_abc_64468_n753_bF_buf11), .B(sqrto_58_), .Y(_auto_iopadmap_cc_313_execute_65414_94_) );
  AND2X2 AND2X2_590 ( .A(u2__abc_44228_n3103), .B(u2__abc_44228_n3108), .Y(u2__abc_44228_n3109) );
  AND2X2 AND2X2_5900 ( .A(u2__abc_44228_n13636), .B(u2__abc_44228_n5770), .Y(u2__abc_44228_n13638) );
  AND2X2 AND2X2_5901 ( .A(u2__abc_44228_n13639), .B(u2__abc_44228_n13637_1), .Y(u2__abc_44228_n13640) );
  AND2X2 AND2X2_5902 ( .A(u2__abc_44228_n13640), .B(u2__abc_44228_n7547_bF_buf48), .Y(u2__abc_44228_n13641) );
  AND2X2 AND2X2_5903 ( .A(u2__abc_44228_n7548_1_bF_buf49), .B(u2_remHi_354_), .Y(u2__abc_44228_n13642) );
  AND2X2 AND2X2_5904 ( .A(u2__abc_44228_n2983_bF_buf63), .B(u2__abc_44228_n5760), .Y(u2__abc_44228_n13645_1) );
  AND2X2 AND2X2_5905 ( .A(u2__abc_44228_n13646), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n13647) );
  AND2X2 AND2X2_5906 ( .A(u2__abc_44228_n13644), .B(u2__abc_44228_n13647), .Y(u2__abc_44228_n13648) );
  AND2X2 AND2X2_5907 ( .A(u2__abc_44228_n13649), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_remHi_356__FF_INPUT) );
  AND2X2 AND2X2_5908 ( .A(u2__abc_44228_n3062_bF_buf14), .B(u2_remHi_357_), .Y(u2__abc_44228_n13651) );
  AND2X2 AND2X2_5909 ( .A(u2__abc_44228_n13639), .B(u2__abc_44228_n6788), .Y(u2__abc_44228_n13652_1) );
  AND2X2 AND2X2_591 ( .A(u2__abc_44228_n3109), .B(u2__abc_44228_n3098), .Y(u2__abc_44228_n3110) );
  AND2X2 AND2X2_5910 ( .A(u2__abc_44228_n13652_1), .B(u2__abc_44228_n5777), .Y(u2__abc_44228_n13653) );
  AND2X2 AND2X2_5911 ( .A(u2__abc_44228_n13655), .B(u2__abc_44228_n13654), .Y(u2__abc_44228_n13656) );
  AND2X2 AND2X2_5912 ( .A(u2__abc_44228_n13657), .B(u2__abc_44228_n7547_bF_buf47), .Y(u2__abc_44228_n13658) );
  AND2X2 AND2X2_5913 ( .A(u2__abc_44228_n7548_1_bF_buf48), .B(u2_remHi_355_), .Y(u2__abc_44228_n13659) );
  AND2X2 AND2X2_5914 ( .A(u2__abc_44228_n2983_bF_buf61), .B(u2__abc_44228_n5754), .Y(u2__abc_44228_n13662_1) );
  AND2X2 AND2X2_5915 ( .A(u2__abc_44228_n13663), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n13664) );
  AND2X2 AND2X2_5916 ( .A(u2__abc_44228_n13661), .B(u2__abc_44228_n13664), .Y(u2__abc_44228_n13665) );
  AND2X2 AND2X2_5917 ( .A(u2__abc_44228_n13666), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_remHi_357__FF_INPUT) );
  AND2X2 AND2X2_5918 ( .A(u2__abc_44228_n3062_bF_buf13), .B(u2_remHi_358_), .Y(u2__abc_44228_n13668) );
  AND2X2 AND2X2_5919 ( .A(u2__abc_44228_n13639), .B(u2__abc_44228_n6789_1), .Y(u2__abc_44228_n13669_1) );
  AND2X2 AND2X2_592 ( .A(u2__abc_44228_n3087), .B(u2__abc_44228_n3110), .Y(u2__abc_44228_n3111) );
  AND2X2 AND2X2_5920 ( .A(u2__abc_44228_n13671), .B(u2__abc_44228_n5763), .Y(u2__abc_44228_n13672) );
  AND2X2 AND2X2_5921 ( .A(u2__abc_44228_n13673), .B(u2__abc_44228_n13674), .Y(u2__abc_44228_n13675) );
  AND2X2 AND2X2_5922 ( .A(u2__abc_44228_n13675), .B(u2__abc_44228_n7547_bF_buf46), .Y(u2__abc_44228_n13676) );
  AND2X2 AND2X2_5923 ( .A(u2__abc_44228_n7548_1_bF_buf47), .B(u2_remHi_356_), .Y(u2__abc_44228_n13677_1) );
  AND2X2 AND2X2_5924 ( .A(u2__abc_44228_n2983_bF_buf60), .B(u2__abc_44228_n5730), .Y(u2__abc_44228_n13680) );
  AND2X2 AND2X2_5925 ( .A(u2__abc_44228_n13681), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n13682) );
  AND2X2 AND2X2_5926 ( .A(u2__abc_44228_n13679), .B(u2__abc_44228_n13682), .Y(u2__abc_44228_n13683) );
  AND2X2 AND2X2_5927 ( .A(u2__abc_44228_n13684_1), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_remHi_358__FF_INPUT) );
  AND2X2 AND2X2_5928 ( .A(u2__abc_44228_n3062_bF_buf12), .B(u2_remHi_359_), .Y(u2__abc_44228_n13686) );
  AND2X2 AND2X2_5929 ( .A(u2__abc_44228_n13691), .B(u2__abc_44228_n7547_bF_buf45), .Y(u2__abc_44228_n13692) );
  AND2X2 AND2X2_593 ( .A(u2__abc_44228_n3112), .B(u2__abc_44228_n3102), .Y(u2__abc_44228_n3113) );
  AND2X2 AND2X2_5930 ( .A(u2__abc_44228_n13692), .B(u2__abc_44228_n13690), .Y(u2__abc_44228_n13693_1) );
  AND2X2 AND2X2_5931 ( .A(u2__abc_44228_n7548_1_bF_buf46), .B(u2_remHi_357_), .Y(u2__abc_44228_n13694) );
  AND2X2 AND2X2_5932 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n5724), .Y(u2__abc_44228_n13697) );
  AND2X2 AND2X2_5933 ( .A(u2__abc_44228_n13698), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n13699) );
  AND2X2 AND2X2_5934 ( .A(u2__abc_44228_n13696), .B(u2__abc_44228_n13699), .Y(u2__abc_44228_n13700_1) );
  AND2X2 AND2X2_5935 ( .A(u2__abc_44228_n13701), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_remHi_359__FF_INPUT) );
  AND2X2 AND2X2_5936 ( .A(u2__abc_44228_n3062_bF_buf11), .B(u2_remHi_360_), .Y(u2__abc_44228_n13703) );
  AND2X2 AND2X2_5937 ( .A(u2__abc_44228_n13568), .B(u2__abc_44228_n5809), .Y(u2__abc_44228_n13704) );
  AND2X2 AND2X2_5938 ( .A(u2__abc_44228_n13705), .B(u2__abc_44228_n5733), .Y(u2__abc_44228_n13706) );
  AND2X2 AND2X2_5939 ( .A(u2__abc_44228_n13707), .B(u2__abc_44228_n13708), .Y(u2__abc_44228_n13709_1) );
  AND2X2 AND2X2_594 ( .A(u2__abc_44228_n3113), .B(u2__abc_44228_n3098), .Y(u2__abc_44228_n3114) );
  AND2X2 AND2X2_5940 ( .A(u2__abc_44228_n13709_1), .B(u2__abc_44228_n7547_bF_buf44), .Y(u2__abc_44228_n13710) );
  AND2X2 AND2X2_5941 ( .A(u2__abc_44228_n7548_1_bF_buf45), .B(u2_remHi_358_), .Y(u2__abc_44228_n13711) );
  AND2X2 AND2X2_5942 ( .A(u2__abc_44228_n2983_bF_buf57), .B(u2__abc_44228_n5744), .Y(u2__abc_44228_n13714) );
  AND2X2 AND2X2_5943 ( .A(u2__abc_44228_n13715), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n13716) );
  AND2X2 AND2X2_5944 ( .A(u2__abc_44228_n13713), .B(u2__abc_44228_n13716), .Y(u2__abc_44228_n13717_1) );
  AND2X2 AND2X2_5945 ( .A(u2__abc_44228_n13718), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_remHi_360__FF_INPUT) );
  AND2X2 AND2X2_5946 ( .A(u2__abc_44228_n3062_bF_buf10), .B(u2_remHi_361_), .Y(u2__abc_44228_n13720) );
  AND2X2 AND2X2_5947 ( .A(u2__abc_44228_n13707), .B(u2__abc_44228_n6798), .Y(u2__abc_44228_n13722) );
  AND2X2 AND2X2_5948 ( .A(u2__abc_44228_n13725), .B(u2__abc_44228_n13723), .Y(u2__abc_44228_n13726) );
  AND2X2 AND2X2_5949 ( .A(u2__abc_44228_n13726), .B(u2__abc_44228_n7547_bF_buf43), .Y(u2__abc_44228_n13727) );
  AND2X2 AND2X2_595 ( .A(u2__abc_44228_n3116), .B(u2__abc_44228_n3091), .Y(u2__abc_44228_n3117) );
  AND2X2 AND2X2_5950 ( .A(u2__abc_44228_n7548_1_bF_buf44), .B(u2_remHi_359_), .Y(u2__abc_44228_n13728) );
  AND2X2 AND2X2_5951 ( .A(u2__abc_44228_n2983_bF_buf55), .B(u2__abc_44228_n5738), .Y(u2__abc_44228_n13731) );
  AND2X2 AND2X2_5952 ( .A(u2__abc_44228_n13732_1), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n13733) );
  AND2X2 AND2X2_5953 ( .A(u2__abc_44228_n13730), .B(u2__abc_44228_n13733), .Y(u2__abc_44228_n13734) );
  AND2X2 AND2X2_5954 ( .A(u2__abc_44228_n13735), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_remHi_361__FF_INPUT) );
  AND2X2 AND2X2_5955 ( .A(u2__abc_44228_n3062_bF_buf9), .B(u2_remHi_362_), .Y(u2__abc_44228_n13737) );
  AND2X2 AND2X2_5956 ( .A(u2__abc_44228_n13705), .B(u2__abc_44228_n5734), .Y(u2__abc_44228_n13738) );
  AND2X2 AND2X2_5957 ( .A(u2__abc_44228_n13739), .B(u2__abc_44228_n5747_1), .Y(u2__abc_44228_n13740_1) );
  AND2X2 AND2X2_5958 ( .A(u2__abc_44228_n13741), .B(u2__abc_44228_n13742), .Y(u2__abc_44228_n13743) );
  AND2X2 AND2X2_5959 ( .A(u2__abc_44228_n13743), .B(u2__abc_44228_n7547_bF_buf42), .Y(u2__abc_44228_n13744) );
  AND2X2 AND2X2_596 ( .A(u2__abc_44228_n3121), .B(u2_remHi_13_), .Y(u2__abc_44228_n3122) );
  AND2X2 AND2X2_5960 ( .A(u2__abc_44228_n7548_1_bF_buf43), .B(u2_remHi_360_), .Y(u2__abc_44228_n13745) );
  AND2X2 AND2X2_5961 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n5715), .Y(u2__abc_44228_n13748) );
  AND2X2 AND2X2_5962 ( .A(u2__abc_44228_n13749_1), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n13750) );
  AND2X2 AND2X2_5963 ( .A(u2__abc_44228_n13747), .B(u2__abc_44228_n13750), .Y(u2__abc_44228_n13751) );
  AND2X2 AND2X2_5964 ( .A(u2__abc_44228_n13752), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_remHi_362__FF_INPUT) );
  AND2X2 AND2X2_5965 ( .A(u2__abc_44228_n3062_bF_buf8), .B(u2_remHi_363_), .Y(u2__abc_44228_n13754) );
  AND2X2 AND2X2_5966 ( .A(u2__abc_44228_n13741), .B(u2__abc_44228_n6803), .Y(u2__abc_44228_n13756) );
  AND2X2 AND2X2_5967 ( .A(u2__abc_44228_n13759), .B(u2__abc_44228_n13757_1), .Y(u2__abc_44228_n13760) );
  AND2X2 AND2X2_5968 ( .A(u2__abc_44228_n13760), .B(u2__abc_44228_n7547_bF_buf41), .Y(u2__abc_44228_n13761) );
  AND2X2 AND2X2_5969 ( .A(u2__abc_44228_n7548_1_bF_buf42), .B(u2_remHi_361_), .Y(u2__abc_44228_n13762) );
  AND2X2 AND2X2_597 ( .A(u2__abc_44228_n3124), .B(sqrto_13_), .Y(u2__abc_44228_n3125) );
  AND2X2 AND2X2_5970 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n5709), .Y(u2__abc_44228_n13765) );
  AND2X2 AND2X2_5971 ( .A(u2__abc_44228_n13766), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n13767_1) );
  AND2X2 AND2X2_5972 ( .A(u2__abc_44228_n13764), .B(u2__abc_44228_n13767_1), .Y(u2__abc_44228_n13768) );
  AND2X2 AND2X2_5973 ( .A(u2__abc_44228_n13769), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_remHi_363__FF_INPUT) );
  AND2X2 AND2X2_5974 ( .A(u2__abc_44228_n3062_bF_buf7), .B(u2_remHi_364_), .Y(u2__abc_44228_n13771) );
  AND2X2 AND2X2_5975 ( .A(u2__abc_44228_n13741), .B(u2__abc_44228_n6804), .Y(u2__abc_44228_n13772) );
  AND2X2 AND2X2_5976 ( .A(u2__abc_44228_n13774), .B(u2__abc_44228_n5718), .Y(u2__abc_44228_n13776) );
  AND2X2 AND2X2_5977 ( .A(u2__abc_44228_n13777), .B(u2__abc_44228_n13775_1), .Y(u2__abc_44228_n13778) );
  AND2X2 AND2X2_5978 ( .A(u2__abc_44228_n13778), .B(u2__abc_44228_n7547_bF_buf40), .Y(u2__abc_44228_n13779) );
  AND2X2 AND2X2_5979 ( .A(u2__abc_44228_n7548_1_bF_buf41), .B(u2_remHi_362_), .Y(u2__abc_44228_n13780) );
  AND2X2 AND2X2_598 ( .A(u2__abc_44228_n3123), .B(u2__abc_44228_n3126), .Y(u2__abc_44228_n3127) );
  AND2X2 AND2X2_5980 ( .A(u2__abc_44228_n2983_bF_buf51), .B(u2__abc_44228_n5701), .Y(u2__abc_44228_n13783) );
  AND2X2 AND2X2_5981 ( .A(u2__abc_44228_n13784_1), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n13785) );
  AND2X2 AND2X2_5982 ( .A(u2__abc_44228_n13782), .B(u2__abc_44228_n13785), .Y(u2__abc_44228_n13786) );
  AND2X2 AND2X2_5983 ( .A(u2__abc_44228_n13787), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_remHi_364__FF_INPUT) );
  AND2X2 AND2X2_5984 ( .A(u2__abc_44228_n3062_bF_buf6), .B(u2_remHi_365_), .Y(u2__abc_44228_n13789) );
  AND2X2 AND2X2_5985 ( .A(u2__abc_44228_n13777), .B(u2__abc_44228_n6811), .Y(u2__abc_44228_n13791) );
  AND2X2 AND2X2_5986 ( .A(u2__abc_44228_n13794), .B(u2__abc_44228_n13792_1), .Y(u2__abc_44228_n13795) );
  AND2X2 AND2X2_5987 ( .A(u2__abc_44228_n13795), .B(u2__abc_44228_n7547_bF_buf39), .Y(u2__abc_44228_n13796) );
  AND2X2 AND2X2_5988 ( .A(u2__abc_44228_n7548_1_bF_buf40), .B(u2_remHi_363_), .Y(u2__abc_44228_n13797) );
  AND2X2 AND2X2_5989 ( .A(u2__abc_44228_n2983_bF_buf49), .B(u2__abc_44228_n5695), .Y(u2__abc_44228_n13800) );
  AND2X2 AND2X2_599 ( .A(u2__abc_44228_n3128), .B(u2_remHi_12_), .Y(u2__abc_44228_n3129) );
  AND2X2 AND2X2_5990 ( .A(u2__abc_44228_n13801), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n13802) );
  AND2X2 AND2X2_5991 ( .A(u2__abc_44228_n13799), .B(u2__abc_44228_n13802), .Y(u2__abc_44228_n13803_1) );
  AND2X2 AND2X2_5992 ( .A(u2__abc_44228_n13804), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_remHi_365__FF_INPUT) );
  AND2X2 AND2X2_5993 ( .A(u2__abc_44228_n3062_bF_buf5), .B(u2_remHi_366_), .Y(u2__abc_44228_n13806) );
  AND2X2 AND2X2_5994 ( .A(u2__abc_44228_n13774), .B(u2__abc_44228_n5719_1), .Y(u2__abc_44228_n13807) );
  AND2X2 AND2X2_5995 ( .A(u2__abc_44228_n13808), .B(u2__abc_44228_n5704), .Y(u2__abc_44228_n13809) );
  AND2X2 AND2X2_5996 ( .A(u2__abc_44228_n13811_1), .B(u2__abc_44228_n7547_bF_buf38), .Y(u2__abc_44228_n13812) );
  AND2X2 AND2X2_5997 ( .A(u2__abc_44228_n13812), .B(u2__abc_44228_n13810), .Y(u2__abc_44228_n13813) );
  AND2X2 AND2X2_5998 ( .A(u2__abc_44228_n7548_1_bF_buf39), .B(u2_remHi_364_), .Y(u2__abc_44228_n13814) );
  AND2X2 AND2X2_5999 ( .A(u2__abc_44228_n2983_bF_buf47), .B(u2__abc_44228_n5670), .Y(u2__abc_44228_n13817) );
  AND2X2 AND2X2_6 ( .A(_abc_64468_n753_bF_buf8), .B(sqrto_5_), .Y(_auto_iopadmap_cc_313_execute_65414_41_) );
  AND2X2 AND2X2_60 ( .A(_abc_64468_n753_bF_buf10), .B(sqrto_59_), .Y(_auto_iopadmap_cc_313_execute_65414_95_) );
  AND2X2 AND2X2_600 ( .A(u2__abc_44228_n3130), .B(sqrto_12_), .Y(u2__abc_44228_n3131) );
  AND2X2 AND2X2_6000 ( .A(u2__abc_44228_n13818), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n13819) );
  AND2X2 AND2X2_6001 ( .A(u2__abc_44228_n13816), .B(u2__abc_44228_n13819), .Y(u2__abc_44228_n13820_1) );
  AND2X2 AND2X2_6002 ( .A(u2__abc_44228_n13821), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_remHi_366__FF_INPUT) );
  AND2X2 AND2X2_6003 ( .A(u2__abc_44228_n3062_bF_buf4), .B(u2_remHi_367_), .Y(u2__abc_44228_n13823) );
  AND2X2 AND2X2_6004 ( .A(u2__abc_44228_n13828_1), .B(u2__abc_44228_n7547_bF_buf37), .Y(u2__abc_44228_n13829) );
  AND2X2 AND2X2_6005 ( .A(u2__abc_44228_n13829), .B(u2__abc_44228_n13827), .Y(u2__abc_44228_n13830) );
  AND2X2 AND2X2_6006 ( .A(u2__abc_44228_n7548_1_bF_buf38), .B(u2_remHi_365_), .Y(u2__abc_44228_n13831) );
  AND2X2 AND2X2_6007 ( .A(u2__abc_44228_n2983_bF_buf45), .B(u2__abc_44228_n5664), .Y(u2__abc_44228_n13834) );
  AND2X2 AND2X2_6008 ( .A(u2__abc_44228_n13835), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n13836) );
  AND2X2 AND2X2_6009 ( .A(u2__abc_44228_n13833), .B(u2__abc_44228_n13836), .Y(u2__abc_44228_n13837) );
  AND2X2 AND2X2_601 ( .A(u2__abc_44228_n3133), .B(u2__abc_44228_n3127), .Y(u2__abc_44228_n3134) );
  AND2X2 AND2X2_6010 ( .A(u2__abc_44228_n13838_1), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_remHi_367__FF_INPUT) );
  AND2X2 AND2X2_6011 ( .A(u2__abc_44228_n3062_bF_buf3), .B(u2_remHi_368_), .Y(u2__abc_44228_n13840) );
  AND2X2 AND2X2_6012 ( .A(u2__abc_44228_n13568), .B(u2__abc_44228_n5810), .Y(u2__abc_44228_n13841) );
  AND2X2 AND2X2_6013 ( .A(u2__abc_44228_n13842), .B(u2__abc_44228_n5673), .Y(u2__abc_44228_n13844) );
  AND2X2 AND2X2_6014 ( .A(u2__abc_44228_n13845), .B(u2__abc_44228_n13843), .Y(u2__abc_44228_n13846_1) );
  AND2X2 AND2X2_6015 ( .A(u2__abc_44228_n13846_1), .B(u2__abc_44228_n7547_bF_buf36), .Y(u2__abc_44228_n13847) );
  AND2X2 AND2X2_6016 ( .A(u2__abc_44228_n7548_1_bF_buf37), .B(u2_remHi_366_), .Y(u2__abc_44228_n13848) );
  AND2X2 AND2X2_6017 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n5684), .Y(u2__abc_44228_n13851) );
  AND2X2 AND2X2_6018 ( .A(u2__abc_44228_n13852), .B(u2__abc_44228_n2972_bF_buf61), .Y(u2__abc_44228_n13853) );
  AND2X2 AND2X2_6019 ( .A(u2__abc_44228_n13850), .B(u2__abc_44228_n13853), .Y(u2__abc_44228_n13854) );
  AND2X2 AND2X2_602 ( .A(u2__abc_44228_n3135), .B(u2_remHi_11_), .Y(u2__abc_44228_n3136) );
  AND2X2 AND2X2_6020 ( .A(u2__abc_44228_n13855_1), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_remHi_368__FF_INPUT) );
  AND2X2 AND2X2_6021 ( .A(u2__abc_44228_n3062_bF_buf2), .B(u2_remHi_369_), .Y(u2__abc_44228_n13857) );
  AND2X2 AND2X2_6022 ( .A(u2__abc_44228_n7548_1_bF_buf36), .B(u2_remHi_367_), .Y(u2__abc_44228_n13858) );
  AND2X2 AND2X2_6023 ( .A(u2__abc_44228_n13845), .B(u2__abc_44228_n6820), .Y(u2__abc_44228_n13861) );
  AND2X2 AND2X2_6024 ( .A(u2__abc_44228_n13864), .B(u2__abc_44228_n13862), .Y(u2__abc_44228_n13865) );
  AND2X2 AND2X2_6025 ( .A(u2__abc_44228_n13865), .B(u2__abc_44228_n7547_bF_buf35), .Y(u2__abc_44228_n13866) );
  AND2X2 AND2X2_6026 ( .A(u2__abc_44228_n2983_bF_buf43), .B(u2__abc_44228_n5678), .Y(u2__abc_44228_n13868) );
  AND2X2 AND2X2_6027 ( .A(u2__abc_44228_n13869), .B(u2__abc_44228_n2972_bF_buf60), .Y(u2__abc_44228_n13870) );
  AND2X2 AND2X2_6028 ( .A(u2__abc_44228_n13867), .B(u2__abc_44228_n13870), .Y(u2__abc_44228_n13871) );
  AND2X2 AND2X2_6029 ( .A(u2__abc_44228_n13872), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_remHi_369__FF_INPUT) );
  AND2X2 AND2X2_603 ( .A(u2__abc_44228_n3138), .B(sqrto_11_), .Y(u2__abc_44228_n3139) );
  AND2X2 AND2X2_6030 ( .A(u2__abc_44228_n3062_bF_buf1), .B(u2_remHi_370_), .Y(u2__abc_44228_n13874) );
  AND2X2 AND2X2_6031 ( .A(u2__abc_44228_n13842), .B(u2__abc_44228_n5674), .Y(u2__abc_44228_n13875_1) );
  AND2X2 AND2X2_6032 ( .A(u2__abc_44228_n13876), .B(u2__abc_44228_n5687), .Y(u2__abc_44228_n13877) );
  AND2X2 AND2X2_6033 ( .A(u2__abc_44228_n13878), .B(u2__abc_44228_n13879), .Y(u2__abc_44228_n13880) );
  AND2X2 AND2X2_6034 ( .A(u2__abc_44228_n13880), .B(u2__abc_44228_n7547_bF_buf34), .Y(u2__abc_44228_n13881) );
  AND2X2 AND2X2_6035 ( .A(u2__abc_44228_n7548_1_bF_buf35), .B(u2_remHi_368_), .Y(u2__abc_44228_n13882) );
  AND2X2 AND2X2_6036 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n5648), .Y(u2__abc_44228_n13885) );
  AND2X2 AND2X2_6037 ( .A(u2__abc_44228_n13886), .B(u2__abc_44228_n2972_bF_buf59), .Y(u2__abc_44228_n13887) );
  AND2X2 AND2X2_6038 ( .A(u2__abc_44228_n13884), .B(u2__abc_44228_n13887), .Y(u2__abc_44228_n13888) );
  AND2X2 AND2X2_6039 ( .A(u2__abc_44228_n13889), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_remHi_370__FF_INPUT) );
  AND2X2 AND2X2_604 ( .A(u2__abc_44228_n3137), .B(u2__abc_44228_n3140), .Y(u2__abc_44228_n3141) );
  AND2X2 AND2X2_6040 ( .A(u2__abc_44228_n3062_bF_buf0), .B(u2_remHi_371_), .Y(u2__abc_44228_n13891) );
  AND2X2 AND2X2_6041 ( .A(u2__abc_44228_n13878), .B(u2__abc_44228_n6825_1), .Y(u2__abc_44228_n13893) );
  AND2X2 AND2X2_6042 ( .A(u2__abc_44228_n13896), .B(u2__abc_44228_n13894), .Y(u2__abc_44228_n13897) );
  AND2X2 AND2X2_6043 ( .A(u2__abc_44228_n13897), .B(u2__abc_44228_n7547_bF_buf33), .Y(u2__abc_44228_n13898) );
  AND2X2 AND2X2_6044 ( .A(u2__abc_44228_n7548_1_bF_buf34), .B(u2_remHi_369_), .Y(u2__abc_44228_n13899) );
  AND2X2 AND2X2_6045 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n5655), .Y(u2__abc_44228_n13902) );
  AND2X2 AND2X2_6046 ( .A(u2__abc_44228_n13903), .B(u2__abc_44228_n2972_bF_buf58), .Y(u2__abc_44228_n13904) );
  AND2X2 AND2X2_6047 ( .A(u2__abc_44228_n13901), .B(u2__abc_44228_n13904), .Y(u2__abc_44228_n13905) );
  AND2X2 AND2X2_6048 ( .A(u2__abc_44228_n13906), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_remHi_371__FF_INPUT) );
  AND2X2 AND2X2_6049 ( .A(u2__abc_44228_n3062_bF_buf92), .B(u2_remHi_372_), .Y(u2__abc_44228_n13908) );
  AND2X2 AND2X2_605 ( .A(u2__abc_44228_n3142), .B(u2_remHi_10_), .Y(u2__abc_44228_n3143) );
  AND2X2 AND2X2_6050 ( .A(u2__abc_44228_n13878), .B(u2__abc_44228_n6826), .Y(u2__abc_44228_n13909) );
  AND2X2 AND2X2_6051 ( .A(u2__abc_44228_n13911), .B(u2__abc_44228_n5651), .Y(u2__abc_44228_n13912) );
  AND2X2 AND2X2_6052 ( .A(u2__abc_44228_n13914), .B(u2__abc_44228_n7547_bF_buf32), .Y(u2__abc_44228_n13915) );
  AND2X2 AND2X2_6053 ( .A(u2__abc_44228_n13915), .B(u2__abc_44228_n13913), .Y(u2__abc_44228_n13916) );
  AND2X2 AND2X2_6054 ( .A(u2__abc_44228_n7548_1_bF_buf33), .B(u2_remHi_370_), .Y(u2__abc_44228_n13917) );
  AND2X2 AND2X2_6055 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n5641), .Y(u2__abc_44228_n13920) );
  AND2X2 AND2X2_6056 ( .A(u2__abc_44228_n13921), .B(u2__abc_44228_n2972_bF_buf57), .Y(u2__abc_44228_n13922) );
  AND2X2 AND2X2_6057 ( .A(u2__abc_44228_n13919), .B(u2__abc_44228_n13922), .Y(u2__abc_44228_n13923) );
  AND2X2 AND2X2_6058 ( .A(u2__abc_44228_n13924), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_remHi_372__FF_INPUT) );
  AND2X2 AND2X2_6059 ( .A(u2__abc_44228_n3062_bF_buf91), .B(u2_remHi_373_), .Y(u2__abc_44228_n13926) );
  AND2X2 AND2X2_606 ( .A(u2__abc_44228_n3144), .B(sqrto_10_), .Y(u2__abc_44228_n3145) );
  AND2X2 AND2X2_6060 ( .A(u2__abc_44228_n13913), .B(u2__abc_44228_n6831), .Y(u2__abc_44228_n13927_1) );
  AND2X2 AND2X2_6061 ( .A(u2__abc_44228_n13927_1), .B(u2__abc_44228_n5658), .Y(u2__abc_44228_n13928) );
  AND2X2 AND2X2_6062 ( .A(u2__abc_44228_n13930), .B(u2__abc_44228_n13929), .Y(u2__abc_44228_n13931) );
  AND2X2 AND2X2_6063 ( .A(u2__abc_44228_n13932), .B(u2__abc_44228_n7547_bF_buf31), .Y(u2__abc_44228_n13933) );
  AND2X2 AND2X2_6064 ( .A(u2__abc_44228_n7548_1_bF_buf32), .B(u2_remHi_371_), .Y(u2__abc_44228_n13934) );
  AND2X2 AND2X2_6065 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n5635), .Y(u2__abc_44228_n13937) );
  AND2X2 AND2X2_6066 ( .A(u2__abc_44228_n13938), .B(u2__abc_44228_n2972_bF_buf56), .Y(u2__abc_44228_n13939) );
  AND2X2 AND2X2_6067 ( .A(u2__abc_44228_n13936), .B(u2__abc_44228_n13939), .Y(u2__abc_44228_n13940) );
  AND2X2 AND2X2_6068 ( .A(u2__abc_44228_n13941), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_remHi_373__FF_INPUT) );
  AND2X2 AND2X2_6069 ( .A(u2__abc_44228_n3062_bF_buf90), .B(u2_remHi_374_), .Y(u2__abc_44228_n13943) );
  AND2X2 AND2X2_607 ( .A(u2__abc_44228_n3147), .B(u2__abc_44228_n3141), .Y(u2__abc_44228_n3148) );
  AND2X2 AND2X2_6070 ( .A(u2__abc_44228_n13913), .B(u2__abc_44228_n6832), .Y(u2__abc_44228_n13944) );
  AND2X2 AND2X2_6071 ( .A(u2__abc_44228_n13946_1), .B(u2__abc_44228_n5644), .Y(u2__abc_44228_n13947) );
  AND2X2 AND2X2_6072 ( .A(u2__abc_44228_n13949), .B(u2__abc_44228_n7547_bF_buf30), .Y(u2__abc_44228_n13950) );
  AND2X2 AND2X2_6073 ( .A(u2__abc_44228_n13950), .B(u2__abc_44228_n13948), .Y(u2__abc_44228_n13951) );
  AND2X2 AND2X2_6074 ( .A(u2__abc_44228_n7548_1_bF_buf31), .B(u2_remHi_372_), .Y(u2__abc_44228_n13952) );
  AND2X2 AND2X2_6075 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n5611), .Y(u2__abc_44228_n13955) );
  AND2X2 AND2X2_6076 ( .A(u2__abc_44228_n13956), .B(u2__abc_44228_n2972_bF_buf55), .Y(u2__abc_44228_n13957) );
  AND2X2 AND2X2_6077 ( .A(u2__abc_44228_n13954_1), .B(u2__abc_44228_n13957), .Y(u2__abc_44228_n13958) );
  AND2X2 AND2X2_6078 ( .A(u2__abc_44228_n13959), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_remHi_374__FF_INPUT) );
  AND2X2 AND2X2_6079 ( .A(u2__abc_44228_n3062_bF_buf89), .B(u2_remHi_375_), .Y(u2__abc_44228_n13961) );
  AND2X2 AND2X2_608 ( .A(u2__abc_44228_n3134), .B(u2__abc_44228_n3148), .Y(u2__abc_44228_n3149) );
  AND2X2 AND2X2_6080 ( .A(u2__abc_44228_n13966), .B(u2__abc_44228_n7547_bF_buf29), .Y(u2__abc_44228_n13967) );
  AND2X2 AND2X2_6081 ( .A(u2__abc_44228_n13967), .B(u2__abc_44228_n13965), .Y(u2__abc_44228_n13968) );
  AND2X2 AND2X2_6082 ( .A(u2__abc_44228_n7548_1_bF_buf30), .B(u2_remHi_373_), .Y(u2__abc_44228_n13969) );
  AND2X2 AND2X2_6083 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n5605), .Y(u2__abc_44228_n13972) );
  AND2X2 AND2X2_6084 ( .A(u2__abc_44228_n13973), .B(u2__abc_44228_n2972_bF_buf54), .Y(u2__abc_44228_n13974) );
  AND2X2 AND2X2_6085 ( .A(u2__abc_44228_n13971_1), .B(u2__abc_44228_n13974), .Y(u2__abc_44228_n13975) );
  AND2X2 AND2X2_6086 ( .A(u2__abc_44228_n13976), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_remHi_375__FF_INPUT) );
  AND2X2 AND2X2_6087 ( .A(u2__abc_44228_n3062_bF_buf88), .B(u2_remHi_376_), .Y(u2__abc_44228_n13978) );
  AND2X2 AND2X2_6088 ( .A(u2__abc_44228_n13842), .B(u2__abc_44228_n5690_1), .Y(u2__abc_44228_n13979) );
  AND2X2 AND2X2_6089 ( .A(u2__abc_44228_n13980), .B(u2__abc_44228_n5614), .Y(u2__abc_44228_n13981_1) );
  AND2X2 AND2X2_609 ( .A(u2__abc_44228_n3151), .B(u2__abc_44228_n3153), .Y(u2__abc_44228_n3154) );
  AND2X2 AND2X2_6090 ( .A(u2__abc_44228_n13982), .B(u2__abc_44228_n13983), .Y(u2__abc_44228_n13984) );
  AND2X2 AND2X2_6091 ( .A(u2__abc_44228_n13984), .B(u2__abc_44228_n7547_bF_buf28), .Y(u2__abc_44228_n13985) );
  AND2X2 AND2X2_6092 ( .A(u2__abc_44228_n7548_1_bF_buf29), .B(u2_remHi_374_), .Y(u2__abc_44228_n13986) );
  AND2X2 AND2X2_6093 ( .A(u2__abc_44228_n2983_bF_buf31), .B(u2__abc_44228_n5625), .Y(u2__abc_44228_n13989_1) );
  AND2X2 AND2X2_6094 ( .A(u2__abc_44228_n13990), .B(u2__abc_44228_n2972_bF_buf53), .Y(u2__abc_44228_n13991) );
  AND2X2 AND2X2_6095 ( .A(u2__abc_44228_n13988), .B(u2__abc_44228_n13991), .Y(u2__abc_44228_n13992) );
  AND2X2 AND2X2_6096 ( .A(u2__abc_44228_n13993), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_remHi_376__FF_INPUT) );
  AND2X2 AND2X2_6097 ( .A(u2__abc_44228_n3062_bF_buf87), .B(u2_remHi_377_), .Y(u2__abc_44228_n13995) );
  AND2X2 AND2X2_6098 ( .A(u2__abc_44228_n13982), .B(u2__abc_44228_n6841), .Y(u2__abc_44228_n13997) );
  AND2X2 AND2X2_6099 ( .A(u2__abc_44228_n14000), .B(u2__abc_44228_n13998_1), .Y(u2__abc_44228_n14001) );
  AND2X2 AND2X2_61 ( .A(_abc_64468_n753_bF_buf9), .B(sqrto_60_), .Y(_auto_iopadmap_cc_313_execute_65414_96_) );
  AND2X2 AND2X2_610 ( .A(u2__abc_44228_n3156), .B(u2__abc_44228_n3158), .Y(u2__abc_44228_n3159) );
  AND2X2 AND2X2_6100 ( .A(u2__abc_44228_n14001), .B(u2__abc_44228_n7547_bF_buf27), .Y(u2__abc_44228_n14002) );
  AND2X2 AND2X2_6101 ( .A(u2__abc_44228_n7548_1_bF_buf28), .B(u2_remHi_375_), .Y(u2__abc_44228_n14003) );
  AND2X2 AND2X2_6102 ( .A(u2__abc_44228_n2983_bF_buf29), .B(u2__abc_44228_n5619), .Y(u2__abc_44228_n14006_1) );
  AND2X2 AND2X2_6103 ( .A(u2__abc_44228_n14007), .B(u2__abc_44228_n2972_bF_buf52), .Y(u2__abc_44228_n14008) );
  AND2X2 AND2X2_6104 ( .A(u2__abc_44228_n14005), .B(u2__abc_44228_n14008), .Y(u2__abc_44228_n14009) );
  AND2X2 AND2X2_6105 ( .A(u2__abc_44228_n14010), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_remHi_377__FF_INPUT) );
  AND2X2 AND2X2_6106 ( .A(u2__abc_44228_n3062_bF_buf86), .B(u2_remHi_378_), .Y(u2__abc_44228_n14012) );
  AND2X2 AND2X2_6107 ( .A(u2__abc_44228_n13980), .B(u2__abc_44228_n5615_1), .Y(u2__abc_44228_n14013) );
  AND2X2 AND2X2_6108 ( .A(u2__abc_44228_n14014), .B(u2__abc_44228_n5628), .Y(u2__abc_44228_n14015) );
  AND2X2 AND2X2_6109 ( .A(u2__abc_44228_n14016), .B(u2__abc_44228_n14017), .Y(u2__abc_44228_n14018) );
  AND2X2 AND2X2_611 ( .A(u2__abc_44228_n3154), .B(u2__abc_44228_n3159), .Y(u2__abc_44228_n3160) );
  AND2X2 AND2X2_6110 ( .A(u2__abc_44228_n14018), .B(u2__abc_44228_n7547_bF_buf26), .Y(u2__abc_44228_n14019_1) );
  AND2X2 AND2X2_6111 ( .A(u2__abc_44228_n7548_1_bF_buf27), .B(u2_remHi_376_), .Y(u2__abc_44228_n14020) );
  AND2X2 AND2X2_6112 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n5596), .Y(u2__abc_44228_n14023) );
  AND2X2 AND2X2_6113 ( .A(u2__abc_44228_n14024), .B(u2__abc_44228_n2972_bF_buf51), .Y(u2__abc_44228_n14025) );
  AND2X2 AND2X2_6114 ( .A(u2__abc_44228_n14022), .B(u2__abc_44228_n14025), .Y(u2__abc_44228_n14026) );
  AND2X2 AND2X2_6115 ( .A(u2__abc_44228_n14027_1), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_remHi_378__FF_INPUT) );
  AND2X2 AND2X2_6116 ( .A(u2__abc_44228_n3062_bF_buf85), .B(u2_remHi_379_), .Y(u2__abc_44228_n14029) );
  AND2X2 AND2X2_6117 ( .A(u2__abc_44228_n14016), .B(u2__abc_44228_n6846), .Y(u2__abc_44228_n14031) );
  AND2X2 AND2X2_6118 ( .A(u2__abc_44228_n14034), .B(u2__abc_44228_n14032), .Y(u2__abc_44228_n14035) );
  AND2X2 AND2X2_6119 ( .A(u2__abc_44228_n14035), .B(u2__abc_44228_n7547_bF_buf25), .Y(u2__abc_44228_n14036_1) );
  AND2X2 AND2X2_612 ( .A(u2__abc_44228_n3161), .B(u2_remHi_6_), .Y(u2__abc_44228_n3162) );
  AND2X2 AND2X2_6120 ( .A(u2__abc_44228_n7548_1_bF_buf26), .B(u2_remHi_377_), .Y(u2__abc_44228_n14037) );
  AND2X2 AND2X2_6121 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n5590), .Y(u2__abc_44228_n14040) );
  AND2X2 AND2X2_6122 ( .A(u2__abc_44228_n14041), .B(u2__abc_44228_n2972_bF_buf50), .Y(u2__abc_44228_n14042) );
  AND2X2 AND2X2_6123 ( .A(u2__abc_44228_n14039), .B(u2__abc_44228_n14042), .Y(u2__abc_44228_n14043) );
  AND2X2 AND2X2_6124 ( .A(u2__abc_44228_n14044_1), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_remHi_379__FF_INPUT) );
  AND2X2 AND2X2_6125 ( .A(u2__abc_44228_n3062_bF_buf84), .B(u2_remHi_380_), .Y(u2__abc_44228_n14046) );
  AND2X2 AND2X2_6126 ( .A(u2__abc_44228_n14016), .B(u2__abc_44228_n6847), .Y(u2__abc_44228_n14047) );
  AND2X2 AND2X2_6127 ( .A(u2__abc_44228_n14049), .B(u2__abc_44228_n5599), .Y(u2__abc_44228_n14050) );
  AND2X2 AND2X2_6128 ( .A(u2__abc_44228_n14052), .B(u2__abc_44228_n7547_bF_buf24), .Y(u2__abc_44228_n14053) );
  AND2X2 AND2X2_6129 ( .A(u2__abc_44228_n14053), .B(u2__abc_44228_n14051), .Y(u2__abc_44228_n14054_1) );
  AND2X2 AND2X2_613 ( .A(u2__abc_44228_n3163), .B(sqrto_6_), .Y(u2__abc_44228_n3164) );
  AND2X2 AND2X2_6130 ( .A(u2__abc_44228_n7548_1_bF_buf25), .B(u2_remHi_378_), .Y(u2__abc_44228_n14055) );
  AND2X2 AND2X2_6131 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n5582), .Y(u2__abc_44228_n14058) );
  AND2X2 AND2X2_6132 ( .A(u2__abc_44228_n14059), .B(u2__abc_44228_n2972_bF_buf49), .Y(u2__abc_44228_n14060) );
  AND2X2 AND2X2_6133 ( .A(u2__abc_44228_n14057), .B(u2__abc_44228_n14060), .Y(u2__abc_44228_n14061) );
  AND2X2 AND2X2_6134 ( .A(u2__abc_44228_n14062_1), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_remHi_380__FF_INPUT) );
  AND2X2 AND2X2_6135 ( .A(u2__abc_44228_n3062_bF_buf83), .B(u2_remHi_381_), .Y(u2__abc_44228_n14064) );
  AND2X2 AND2X2_6136 ( .A(u2__abc_44228_n14051), .B(u2__abc_44228_n6854), .Y(u2__abc_44228_n14065) );
  AND2X2 AND2X2_6137 ( .A(u2__abc_44228_n14065), .B(u2__abc_44228_n5593), .Y(u2__abc_44228_n14066) );
  AND2X2 AND2X2_6138 ( .A(u2__abc_44228_n14068), .B(u2__abc_44228_n14067), .Y(u2__abc_44228_n14069) );
  AND2X2 AND2X2_6139 ( .A(u2__abc_44228_n14070), .B(u2__abc_44228_n7547_bF_buf23), .Y(u2__abc_44228_n14071_1) );
  AND2X2 AND2X2_614 ( .A(u2__abc_44228_n3167), .B(u2_remHi_7_), .Y(u2__abc_44228_n3168) );
  AND2X2 AND2X2_6140 ( .A(u2__abc_44228_n7548_1_bF_buf24), .B(u2_remHi_379_), .Y(u2__abc_44228_n14072) );
  AND2X2 AND2X2_6141 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n5576), .Y(u2__abc_44228_n14075) );
  AND2X2 AND2X2_6142 ( .A(u2__abc_44228_n14076), .B(u2__abc_44228_n2972_bF_buf48), .Y(u2__abc_44228_n14077) );
  AND2X2 AND2X2_6143 ( .A(u2__abc_44228_n14074), .B(u2__abc_44228_n14077), .Y(u2__abc_44228_n14078) );
  AND2X2 AND2X2_6144 ( .A(u2__abc_44228_n14079_1), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_remHi_381__FF_INPUT) );
  AND2X2 AND2X2_6145 ( .A(u2__abc_44228_n3062_bF_buf82), .B(u2_remHi_382_), .Y(u2__abc_44228_n14081) );
  AND2X2 AND2X2_6146 ( .A(u2__abc_44228_n14051), .B(u2__abc_44228_n6855), .Y(u2__abc_44228_n14082) );
  AND2X2 AND2X2_6147 ( .A(u2__abc_44228_n14084), .B(u2__abc_44228_n5585), .Y(u2__abc_44228_n14085) );
  AND2X2 AND2X2_6148 ( .A(u2__abc_44228_n14087), .B(u2__abc_44228_n7547_bF_buf22), .Y(u2__abc_44228_n14088) );
  AND2X2 AND2X2_6149 ( .A(u2__abc_44228_n14088), .B(u2__abc_44228_n14086), .Y(u2__abc_44228_n14089) );
  AND2X2 AND2X2_615 ( .A(u2__abc_44228_n3170), .B(sqrto_7_), .Y(u2__abc_44228_n3171) );
  AND2X2 AND2X2_6150 ( .A(u2__abc_44228_n7548_1_bF_buf23), .B(u2_remHi_380_), .Y(u2__abc_44228_n14090_1) );
  AND2X2 AND2X2_6151 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n7335), .Y(u2__abc_44228_n14093) );
  AND2X2 AND2X2_6152 ( .A(u2__abc_44228_n14094), .B(u2__abc_44228_n2972_bF_buf47), .Y(u2__abc_44228_n14095) );
  AND2X2 AND2X2_6153 ( .A(u2__abc_44228_n14092), .B(u2__abc_44228_n14095), .Y(u2__abc_44228_n14096) );
  AND2X2 AND2X2_6154 ( .A(u2__abc_44228_n14097), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_remHi_382__FF_INPUT) );
  AND2X2 AND2X2_6155 ( .A(u2__abc_44228_n3062_bF_buf81), .B(u2_remHi_383_), .Y(u2__abc_44228_n14099) );
  AND2X2 AND2X2_6156 ( .A(u2__abc_44228_n14104), .B(u2__abc_44228_n7547_bF_buf21), .Y(u2__abc_44228_n14105) );
  AND2X2 AND2X2_6157 ( .A(u2__abc_44228_n14105), .B(u2__abc_44228_n14103), .Y(u2__abc_44228_n14106) );
  AND2X2 AND2X2_6158 ( .A(u2__abc_44228_n7548_1_bF_buf22), .B(u2_remHi_381_), .Y(u2__abc_44228_n14107_1) );
  AND2X2 AND2X2_6159 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n7329), .Y(u2__abc_44228_n14110) );
  AND2X2 AND2X2_616 ( .A(u2__abc_44228_n3169), .B(u2__abc_44228_n3172), .Y(u2__abc_44228_n3173) );
  AND2X2 AND2X2_6160 ( .A(u2__abc_44228_n14111), .B(u2__abc_44228_n2972_bF_buf46), .Y(u2__abc_44228_n14112) );
  AND2X2 AND2X2_6161 ( .A(u2__abc_44228_n14109), .B(u2__abc_44228_n14112), .Y(u2__abc_44228_n14113) );
  AND2X2 AND2X2_6162 ( .A(u2__abc_44228_n14114), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_remHi_383__FF_INPUT) );
  AND2X2 AND2X2_6163 ( .A(u2__abc_44228_n3062_bF_buf80), .B(u2_remHi_384_), .Y(u2__abc_44228_n14116) );
  AND2X2 AND2X2_6164 ( .A(u2__abc_44228_n6865), .B(u2__abc_44228_n7338), .Y(u2__abc_44228_n14117) );
  AND2X2 AND2X2_6165 ( .A(u2__abc_44228_n14118), .B(u2__abc_44228_n14119), .Y(u2__abc_44228_n14120) );
  AND2X2 AND2X2_6166 ( .A(u2__abc_44228_n14121), .B(u2__abc_44228_n14122), .Y(u2__abc_44228_n14123) );
  AND2X2 AND2X2_6167 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n7321), .Y(u2__abc_44228_n14125_1) );
  AND2X2 AND2X2_6168 ( .A(u2__abc_44228_n14126), .B(u2__abc_44228_n2972_bF_buf45), .Y(u2__abc_44228_n14127) );
  AND2X2 AND2X2_6169 ( .A(u2__abc_44228_n14124), .B(u2__abc_44228_n14127), .Y(u2__abc_44228_n14128) );
  AND2X2 AND2X2_617 ( .A(u2__abc_44228_n3166), .B(u2__abc_44228_n3173), .Y(u2__abc_44228_n3174) );
  AND2X2 AND2X2_6170 ( .A(u2__abc_44228_n14129), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_remHi_384__FF_INPUT) );
  AND2X2 AND2X2_6171 ( .A(u2__abc_44228_n3062_bF_buf79), .B(u2_remHi_385_), .Y(u2__abc_44228_n14131) );
  AND2X2 AND2X2_6172 ( .A(u2__abc_44228_n14118), .B(u2__abc_44228_n7346_1), .Y(u2__abc_44228_n14133_1) );
  AND2X2 AND2X2_6173 ( .A(u2__abc_44228_n14136), .B(u2__abc_44228_n14134), .Y(u2__abc_44228_n14137) );
  AND2X2 AND2X2_6174 ( .A(u2__abc_44228_n14137), .B(u2__abc_44228_n7547_bF_buf19), .Y(u2__abc_44228_n14138) );
  AND2X2 AND2X2_6175 ( .A(u2__abc_44228_n7548_1_bF_buf20), .B(u2_remHi_383_), .Y(u2__abc_44228_n14139) );
  AND2X2 AND2X2_6176 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n7315), .Y(u2__abc_44228_n14142_1) );
  AND2X2 AND2X2_6177 ( .A(u2__abc_44228_n14143), .B(u2__abc_44228_n2972_bF_buf44), .Y(u2__abc_44228_n14144) );
  AND2X2 AND2X2_6178 ( .A(u2__abc_44228_n14141), .B(u2__abc_44228_n14144), .Y(u2__abc_44228_n14145) );
  AND2X2 AND2X2_6179 ( .A(u2__abc_44228_n14146), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_remHi_385__FF_INPUT) );
  AND2X2 AND2X2_618 ( .A(u2__abc_44228_n3174), .B(u2__abc_44228_n3160), .Y(u2__abc_44228_n3175) );
  AND2X2 AND2X2_6180 ( .A(u2__abc_44228_n3062_bF_buf78), .B(u2_remHi_386_), .Y(u2__abc_44228_n14148) );
  AND2X2 AND2X2_6181 ( .A(u2__abc_44228_n6865), .B(u2__abc_44228_n7339), .Y(u2__abc_44228_n14149) );
  AND2X2 AND2X2_6182 ( .A(u2__abc_44228_n14150_1), .B(u2__abc_44228_n7324), .Y(u2__abc_44228_n14151) );
  AND2X2 AND2X2_6183 ( .A(u2__abc_44228_n14152), .B(u2__abc_44228_n14153), .Y(u2__abc_44228_n14154) );
  AND2X2 AND2X2_6184 ( .A(u2__abc_44228_n14155), .B(u2__abc_44228_n14156), .Y(u2__abc_44228_n14157) );
  AND2X2 AND2X2_6185 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n7299_1), .Y(u2__abc_44228_n14159) );
  AND2X2 AND2X2_6186 ( .A(u2__abc_44228_n14160), .B(u2__abc_44228_n2972_bF_buf43), .Y(u2__abc_44228_n14161) );
  AND2X2 AND2X2_6187 ( .A(u2__abc_44228_n14158), .B(u2__abc_44228_n14161), .Y(u2__abc_44228_n14162_1) );
  AND2X2 AND2X2_6188 ( .A(u2__abc_44228_n14163), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_remHi_386__FF_INPUT) );
  AND2X2 AND2X2_6189 ( .A(u2__abc_44228_n3062_bF_buf77), .B(u2_remHi_387_), .Y(u2__abc_44228_n14165) );
  AND2X2 AND2X2_619 ( .A(u2__abc_44228_n3149), .B(u2__abc_44228_n3175), .Y(u2__abc_44228_n3176) );
  AND2X2 AND2X2_6190 ( .A(u2__abc_44228_n14170_1), .B(u2__abc_44228_n7547_bF_buf17), .Y(u2__abc_44228_n14171) );
  AND2X2 AND2X2_6191 ( .A(u2__abc_44228_n14171), .B(u2__abc_44228_n14169), .Y(u2__abc_44228_n14172) );
  AND2X2 AND2X2_6192 ( .A(u2__abc_44228_n7548_1_bF_buf18), .B(u2_remHi_385_), .Y(u2__abc_44228_n14173) );
  AND2X2 AND2X2_6193 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n7306), .Y(u2__abc_44228_n14176) );
  AND2X2 AND2X2_6194 ( .A(u2__abc_44228_n14177), .B(u2__abc_44228_n2972_bF_buf42), .Y(u2__abc_44228_n14178) );
  AND2X2 AND2X2_6195 ( .A(u2__abc_44228_n14175), .B(u2__abc_44228_n14178), .Y(u2__abc_44228_n14179_1) );
  AND2X2 AND2X2_6196 ( .A(u2__abc_44228_n14180), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_remHi_387__FF_INPUT) );
  AND2X2 AND2X2_6197 ( .A(u2__abc_44228_n3062_bF_buf76), .B(u2_remHi_388_), .Y(u2__abc_44228_n14182) );
  AND2X2 AND2X2_6198 ( .A(u2__abc_44228_n6865), .B(u2__abc_44228_n7340), .Y(u2__abc_44228_n14183) );
  AND2X2 AND2X2_6199 ( .A(u2__abc_44228_n14184), .B(u2__abc_44228_n7302), .Y(u2__abc_44228_n14186) );
  AND2X2 AND2X2_62 ( .A(_abc_64468_n753_bF_buf8), .B(sqrto_61_), .Y(_auto_iopadmap_cc_313_execute_65414_97_) );
  AND2X2 AND2X2_620 ( .A(u2__abc_44228_n3120), .B(u2__abc_44228_n3176), .Y(u2__abc_44228_n3177) );
  AND2X2 AND2X2_6200 ( .A(u2__abc_44228_n14187_1), .B(u2__abc_44228_n14185), .Y(u2__abc_44228_n14188) );
  AND2X2 AND2X2_6201 ( .A(u2__abc_44228_n14189), .B(u2__abc_44228_n14190), .Y(u2__abc_44228_n14191) );
  AND2X2 AND2X2_6202 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n7292), .Y(u2__abc_44228_n14193) );
  AND2X2 AND2X2_6203 ( .A(u2__abc_44228_n14194), .B(u2__abc_44228_n2972_bF_buf41), .Y(u2__abc_44228_n14195) );
  AND2X2 AND2X2_6204 ( .A(u2__abc_44228_n14192), .B(u2__abc_44228_n14195), .Y(u2__abc_44228_n14196) );
  AND2X2 AND2X2_6205 ( .A(u2__abc_44228_n14197_1), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_remHi_388__FF_INPUT) );
  AND2X2 AND2X2_6206 ( .A(u2__abc_44228_n3062_bF_buf75), .B(u2_remHi_389_), .Y(u2__abc_44228_n14199) );
  AND2X2 AND2X2_6207 ( .A(u2__abc_44228_n14187_1), .B(u2__abc_44228_n7355_1), .Y(u2__abc_44228_n14200) );
  AND2X2 AND2X2_6208 ( .A(u2__abc_44228_n14204), .B(u2__abc_44228_n7547_bF_buf15), .Y(u2__abc_44228_n14205_1) );
  AND2X2 AND2X2_6209 ( .A(u2__abc_44228_n14205_1), .B(u2__abc_44228_n14202), .Y(u2__abc_44228_n14206) );
  AND2X2 AND2X2_621 ( .A(u2__abc_44228_n3178), .B(u2__abc_44228_n3172), .Y(u2__abc_44228_n3179) );
  AND2X2 AND2X2_6210 ( .A(u2__abc_44228_n7548_1_bF_buf16), .B(u2_remHi_387_), .Y(u2__abc_44228_n14207) );
  AND2X2 AND2X2_6211 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n7286), .Y(u2__abc_44228_n14210) );
  AND2X2 AND2X2_6212 ( .A(u2__abc_44228_n14211), .B(u2__abc_44228_n2972_bF_buf40), .Y(u2__abc_44228_n14212) );
  AND2X2 AND2X2_6213 ( .A(u2__abc_44228_n14209), .B(u2__abc_44228_n14212), .Y(u2__abc_44228_n14213) );
  AND2X2 AND2X2_6214 ( .A(u2__abc_44228_n14214_1), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_remHi_389__FF_INPUT) );
  AND2X2 AND2X2_6215 ( .A(u2__abc_44228_n3062_bF_buf74), .B(u2_remHi_390_), .Y(u2__abc_44228_n14216) );
  AND2X2 AND2X2_6216 ( .A(u2__abc_44228_n14187_1), .B(u2__abc_44228_n7356), .Y(u2__abc_44228_n14217) );
  AND2X2 AND2X2_6217 ( .A(u2__abc_44228_n14219), .B(u2__abc_44228_n7295), .Y(u2__abc_44228_n14220) );
  AND2X2 AND2X2_6218 ( .A(u2__abc_44228_n14221), .B(u2__abc_44228_n14222_1), .Y(u2__abc_44228_n14223) );
  AND2X2 AND2X2_6219 ( .A(u2__abc_44228_n14223), .B(u2__abc_44228_n7547_bF_buf14), .Y(u2__abc_44228_n14224) );
  AND2X2 AND2X2_622 ( .A(u2__abc_44228_n3179), .B(u2__abc_44228_n3160), .Y(u2__abc_44228_n3180) );
  AND2X2 AND2X2_6220 ( .A(u2__abc_44228_n7548_1_bF_buf15), .B(u2_remHi_388_), .Y(u2__abc_44228_n14225) );
  AND2X2 AND2X2_6221 ( .A(u2__abc_44228_n2983_bF_buf5), .B(u2__abc_44228_n7269), .Y(u2__abc_44228_n14228) );
  AND2X2 AND2X2_6222 ( .A(u2__abc_44228_n14229), .B(u2__abc_44228_n2972_bF_buf39), .Y(u2__abc_44228_n14230) );
  AND2X2 AND2X2_6223 ( .A(u2__abc_44228_n14227), .B(u2__abc_44228_n14230), .Y(u2__abc_44228_n14231) );
  AND2X2 AND2X2_6224 ( .A(u2__abc_44228_n14232), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_remHi_390__FF_INPUT) );
  AND2X2 AND2X2_6225 ( .A(u2__abc_44228_n3062_bF_buf73), .B(u2_remHi_391_), .Y(u2__abc_44228_n14234) );
  AND2X2 AND2X2_6226 ( .A(u2__abc_44228_n14239), .B(u2__abc_44228_n7547_bF_buf13), .Y(u2__abc_44228_n14240) );
  AND2X2 AND2X2_6227 ( .A(u2__abc_44228_n14240), .B(u2__abc_44228_n14238), .Y(u2__abc_44228_n14241_1) );
  AND2X2 AND2X2_6228 ( .A(u2__abc_44228_n7548_1_bF_buf14), .B(u2_remHi_389_), .Y(u2__abc_44228_n14242) );
  AND2X2 AND2X2_6229 ( .A(u2__abc_44228_n2983_bF_buf3), .B(u2__abc_44228_n7276), .Y(u2__abc_44228_n14245) );
  AND2X2 AND2X2_623 ( .A(u2__abc_44228_n3182), .B(u2__abc_44228_n3153), .Y(u2__abc_44228_n3183) );
  AND2X2 AND2X2_6230 ( .A(u2__abc_44228_n14246), .B(u2__abc_44228_n2972_bF_buf38), .Y(u2__abc_44228_n14247) );
  AND2X2 AND2X2_6231 ( .A(u2__abc_44228_n14244), .B(u2__abc_44228_n14247), .Y(u2__abc_44228_n14248) );
  AND2X2 AND2X2_6232 ( .A(u2__abc_44228_n14249), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_remHi_391__FF_INPUT) );
  AND2X2 AND2X2_6233 ( .A(u2__abc_44228_n3062_bF_buf72), .B(u2_remHi_392_), .Y(u2__abc_44228_n14251) );
  AND2X2 AND2X2_6234 ( .A(u2__abc_44228_n6865), .B(u2__abc_44228_n7341), .Y(u2__abc_44228_n14252) );
  AND2X2 AND2X2_6235 ( .A(u2__abc_44228_n14253), .B(u2__abc_44228_n7272), .Y(u2__abc_44228_n14254) );
  AND2X2 AND2X2_6236 ( .A(u2__abc_44228_n14255), .B(u2__abc_44228_n14256), .Y(u2__abc_44228_n14257) );
  AND2X2 AND2X2_6237 ( .A(u2__abc_44228_n14258_1), .B(u2__abc_44228_n14259), .Y(u2__abc_44228_n14260) );
  AND2X2 AND2X2_6238 ( .A(u2__abc_44228_n2983_bF_buf1), .B(u2__abc_44228_n7262_1), .Y(u2__abc_44228_n14262) );
  AND2X2 AND2X2_6239 ( .A(u2__abc_44228_n14263), .B(u2__abc_44228_n2972_bF_buf37), .Y(u2__abc_44228_n14264) );
  AND2X2 AND2X2_624 ( .A(u2__abc_44228_n3185), .B(u2__abc_44228_n3149), .Y(u2__abc_44228_n3186) );
  AND2X2 AND2X2_6240 ( .A(u2__abc_44228_n14261), .B(u2__abc_44228_n14264), .Y(u2__abc_44228_n14265) );
  AND2X2 AND2X2_6241 ( .A(u2__abc_44228_n14266), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_remHi_392__FF_INPUT) );
  AND2X2 AND2X2_6242 ( .A(u2__abc_44228_n3062_bF_buf71), .B(u2_remHi_393_), .Y(u2__abc_44228_n14268_1) );
  AND2X2 AND2X2_6243 ( .A(u2__abc_44228_n14255), .B(u2__abc_44228_n7365), .Y(u2__abc_44228_n14270) );
  AND2X2 AND2X2_6244 ( .A(u2__abc_44228_n14273), .B(u2__abc_44228_n14271), .Y(u2__abc_44228_n14274) );
  AND2X2 AND2X2_6245 ( .A(u2__abc_44228_n14274), .B(u2__abc_44228_n7547_bF_buf11), .Y(u2__abc_44228_n14275) );
  AND2X2 AND2X2_6246 ( .A(u2__abc_44228_n7548_1_bF_buf12), .B(u2_remHi_391_), .Y(u2__abc_44228_n14276_1) );
  AND2X2 AND2X2_6247 ( .A(u2__abc_44228_n2983_bF_buf141), .B(u2__abc_44228_n7256), .Y(u2__abc_44228_n14279) );
  AND2X2 AND2X2_6248 ( .A(u2__abc_44228_n14280), .B(u2__abc_44228_n2972_bF_buf36), .Y(u2__abc_44228_n14281) );
  AND2X2 AND2X2_6249 ( .A(u2__abc_44228_n14278), .B(u2__abc_44228_n14281), .Y(u2__abc_44228_n14282) );
  AND2X2 AND2X2_625 ( .A(u2__abc_44228_n3187), .B(u2__abc_44228_n3140), .Y(u2__abc_44228_n3188) );
  AND2X2 AND2X2_6250 ( .A(u2__abc_44228_n14283), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_remHi_393__FF_INPUT) );
  AND2X2 AND2X2_6251 ( .A(u2__abc_44228_n3062_bF_buf70), .B(u2_remHi_394_), .Y(u2__abc_44228_n14285_1) );
  AND2X2 AND2X2_6252 ( .A(u2__abc_44228_n14255), .B(u2__abc_44228_n7366), .Y(u2__abc_44228_n14286) );
  AND2X2 AND2X2_6253 ( .A(u2__abc_44228_n14288), .B(u2__abc_44228_n7265), .Y(u2__abc_44228_n14289) );
  AND2X2 AND2X2_6254 ( .A(u2__abc_44228_n14290), .B(u2__abc_44228_n14291), .Y(u2__abc_44228_n14292) );
  AND2X2 AND2X2_6255 ( .A(u2__abc_44228_n14292), .B(u2__abc_44228_n7547_bF_buf10), .Y(u2__abc_44228_n14293_1) );
  AND2X2 AND2X2_6256 ( .A(u2__abc_44228_n7548_1_bF_buf11), .B(u2_remHi_392_), .Y(u2__abc_44228_n14294) );
  AND2X2 AND2X2_6257 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n7240), .Y(u2__abc_44228_n14297) );
  AND2X2 AND2X2_6258 ( .A(u2__abc_44228_n14298), .B(u2__abc_44228_n2972_bF_buf35), .Y(u2__abc_44228_n14299) );
  AND2X2 AND2X2_6259 ( .A(u2__abc_44228_n14296), .B(u2__abc_44228_n14299), .Y(u2__abc_44228_n14300) );
  AND2X2 AND2X2_626 ( .A(u2__abc_44228_n3134), .B(u2__abc_44228_n3188), .Y(u2__abc_44228_n3189) );
  AND2X2 AND2X2_6260 ( .A(u2__abc_44228_n14301), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_remHi_394__FF_INPUT) );
  AND2X2 AND2X2_6261 ( .A(u2__abc_44228_n3062_bF_buf69), .B(u2_remHi_395_), .Y(u2__abc_44228_n14303) );
  AND2X2 AND2X2_6262 ( .A(u2__abc_44228_n14308), .B(u2__abc_44228_n7547_bF_buf9), .Y(u2__abc_44228_n14309) );
  AND2X2 AND2X2_6263 ( .A(u2__abc_44228_n14309), .B(u2__abc_44228_n14307_1), .Y(u2__abc_44228_n14310) );
  AND2X2 AND2X2_6264 ( .A(u2__abc_44228_n7548_1_bF_buf10), .B(u2_remHi_393_), .Y(u2__abc_44228_n14311) );
  AND2X2 AND2X2_6265 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n7247), .Y(u2__abc_44228_n14314) );
  AND2X2 AND2X2_6266 ( .A(u2__abc_44228_n14315_1), .B(u2__abc_44228_n2972_bF_buf34), .Y(u2__abc_44228_n14316) );
  AND2X2 AND2X2_6267 ( .A(u2__abc_44228_n14313), .B(u2__abc_44228_n14316), .Y(u2__abc_44228_n14317) );
  AND2X2 AND2X2_6268 ( .A(u2__abc_44228_n14318), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_remHi_395__FF_INPUT) );
  AND2X2 AND2X2_6269 ( .A(u2__abc_44228_n3062_bF_buf68), .B(u2_remHi_396_), .Y(u2__abc_44228_n14320) );
  AND2X2 AND2X2_627 ( .A(u2__abc_44228_n3126), .B(u2__abc_44228_n3129), .Y(u2__abc_44228_n3190) );
  AND2X2 AND2X2_6270 ( .A(u2__abc_44228_n14253), .B(u2__abc_44228_n7281), .Y(u2__abc_44228_n14321) );
  AND2X2 AND2X2_6271 ( .A(u2__abc_44228_n14322), .B(u2__abc_44228_n7243), .Y(u2__abc_44228_n14324_1) );
  AND2X2 AND2X2_6272 ( .A(u2__abc_44228_n14325), .B(u2__abc_44228_n14323), .Y(u2__abc_44228_n14326) );
  AND2X2 AND2X2_6273 ( .A(u2__abc_44228_n14326), .B(u2__abc_44228_n7547_bF_buf8), .Y(u2__abc_44228_n14327) );
  AND2X2 AND2X2_6274 ( .A(u2__abc_44228_n7548_1_bF_buf9), .B(u2_remHi_394_), .Y(u2__abc_44228_n14328) );
  AND2X2 AND2X2_6275 ( .A(u2__abc_44228_n2983_bF_buf137), .B(u2__abc_44228_n7233), .Y(u2__abc_44228_n14331) );
  AND2X2 AND2X2_6276 ( .A(u2__abc_44228_n14332_1), .B(u2__abc_44228_n2972_bF_buf33), .Y(u2__abc_44228_n14333) );
  AND2X2 AND2X2_6277 ( .A(u2__abc_44228_n14330), .B(u2__abc_44228_n14333), .Y(u2__abc_44228_n14334) );
  AND2X2 AND2X2_6278 ( .A(u2__abc_44228_n14335), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_remHi_396__FF_INPUT) );
  AND2X2 AND2X2_6279 ( .A(u2__abc_44228_n3062_bF_buf67), .B(u2_remHi_397_), .Y(u2__abc_44228_n14337) );
  AND2X2 AND2X2_628 ( .A(u2__abc_44228_n3195), .B(u2_remHi_29_), .Y(u2__abc_44228_n3196) );
  AND2X2 AND2X2_6280 ( .A(u2__abc_44228_n14325), .B(u2__abc_44228_n7376), .Y(u2__abc_44228_n14338) );
  AND2X2 AND2X2_6281 ( .A(u2__abc_44228_n14338), .B(u2__abc_44228_n7250), .Y(u2__abc_44228_n14339) );
  AND2X2 AND2X2_6282 ( .A(u2__abc_44228_n14341), .B(u2__abc_44228_n14340), .Y(u2__abc_44228_n14342_1) );
  AND2X2 AND2X2_6283 ( .A(u2__abc_44228_n14343), .B(u2__abc_44228_n7547_bF_buf7), .Y(u2__abc_44228_n14344) );
  AND2X2 AND2X2_6284 ( .A(u2__abc_44228_n7548_1_bF_buf8), .B(u2_remHi_395_), .Y(u2__abc_44228_n14345) );
  AND2X2 AND2X2_6285 ( .A(u2__abc_44228_n2983_bF_buf135), .B(u2__abc_44228_n7227), .Y(u2__abc_44228_n14348) );
  AND2X2 AND2X2_6286 ( .A(u2__abc_44228_n14349), .B(u2__abc_44228_n2972_bF_buf32), .Y(u2__abc_44228_n14350_1) );
  AND2X2 AND2X2_6287 ( .A(u2__abc_44228_n14347), .B(u2__abc_44228_n14350_1), .Y(u2__abc_44228_n14351) );
  AND2X2 AND2X2_6288 ( .A(u2__abc_44228_n14352), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_remHi_397__FF_INPUT) );
  AND2X2 AND2X2_6289 ( .A(u2__abc_44228_n3062_bF_buf66), .B(u2_remHi_398_), .Y(u2__abc_44228_n14354) );
  AND2X2 AND2X2_629 ( .A(u2__abc_44228_n3198), .B(sqrto_29_), .Y(u2__abc_44228_n3199) );
  AND2X2 AND2X2_6290 ( .A(u2__abc_44228_n14325), .B(u2__abc_44228_n7377), .Y(u2__abc_44228_n14355) );
  AND2X2 AND2X2_6291 ( .A(u2__abc_44228_n14357), .B(u2__abc_44228_n7236), .Y(u2__abc_44228_n14358) );
  AND2X2 AND2X2_6292 ( .A(u2__abc_44228_n14359_1), .B(u2__abc_44228_n14360), .Y(u2__abc_44228_n14361) );
  AND2X2 AND2X2_6293 ( .A(u2__abc_44228_n14361), .B(u2__abc_44228_n7547_bF_buf6), .Y(u2__abc_44228_n14362) );
  AND2X2 AND2X2_6294 ( .A(u2__abc_44228_n7548_1_bF_buf7), .B(u2_remHi_396_), .Y(u2__abc_44228_n14363) );
  AND2X2 AND2X2_6295 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n7209), .Y(u2__abc_44228_n14366) );
  AND2X2 AND2X2_6296 ( .A(u2__abc_44228_n14367_1), .B(u2__abc_44228_n2972_bF_buf31), .Y(u2__abc_44228_n14368) );
  AND2X2 AND2X2_6297 ( .A(u2__abc_44228_n14365), .B(u2__abc_44228_n14368), .Y(u2__abc_44228_n14369) );
  AND2X2 AND2X2_6298 ( .A(u2__abc_44228_n14370), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_remHi_398__FF_INPUT) );
  AND2X2 AND2X2_6299 ( .A(u2__abc_44228_n3062_bF_buf65), .B(u2_remHi_399_), .Y(u2__abc_44228_n14372) );
  AND2X2 AND2X2_63 ( .A(_abc_64468_n753_bF_buf7), .B(sqrto_62_), .Y(_auto_iopadmap_cc_313_execute_65414_98_) );
  AND2X2 AND2X2_630 ( .A(u2__abc_44228_n3197), .B(u2__abc_44228_n3200), .Y(u2__abc_44228_n3201) );
  AND2X2 AND2X2_6300 ( .A(u2__abc_44228_n14377), .B(u2__abc_44228_n7547_bF_buf5), .Y(u2__abc_44228_n14378_1) );
  AND2X2 AND2X2_6301 ( .A(u2__abc_44228_n14378_1), .B(u2__abc_44228_n14376), .Y(u2__abc_44228_n14379) );
  AND2X2 AND2X2_6302 ( .A(u2__abc_44228_n7548_1_bF_buf6), .B(u2_remHi_397_), .Y(u2__abc_44228_n14380) );
  AND2X2 AND2X2_6303 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n7216), .Y(u2__abc_44228_n14383) );
  AND2X2 AND2X2_6304 ( .A(u2__abc_44228_n14384), .B(u2__abc_44228_n2972_bF_buf30), .Y(u2__abc_44228_n14385) );
  AND2X2 AND2X2_6305 ( .A(u2__abc_44228_n14382), .B(u2__abc_44228_n14385), .Y(u2__abc_44228_n14386_1) );
  AND2X2 AND2X2_6306 ( .A(u2__abc_44228_n14387), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_remHi_399__FF_INPUT) );
  AND2X2 AND2X2_6307 ( .A(u2__abc_44228_n3062_bF_buf64), .B(u2_remHi_400_), .Y(u2__abc_44228_n14389) );
  AND2X2 AND2X2_6308 ( .A(u2__abc_44228_n6865), .B(u2__abc_44228_n7342), .Y(u2__abc_44228_n14390) );
  AND2X2 AND2X2_6309 ( .A(u2__abc_44228_n14391), .B(u2__abc_44228_n7212), .Y(u2__abc_44228_n14393) );
  AND2X2 AND2X2_631 ( .A(u2__abc_44228_n3202), .B(u2_remHi_28_), .Y(u2__abc_44228_n3203) );
  AND2X2 AND2X2_6310 ( .A(u2__abc_44228_n14394), .B(u2__abc_44228_n14392), .Y(u2__abc_44228_n14395_1) );
  AND2X2 AND2X2_6311 ( .A(u2__abc_44228_n14396), .B(u2__abc_44228_n14397), .Y(u2__abc_44228_n14398) );
  AND2X2 AND2X2_6312 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n7202), .Y(u2__abc_44228_n14400) );
  AND2X2 AND2X2_6313 ( .A(u2__abc_44228_n14401), .B(u2__abc_44228_n2972_bF_buf29), .Y(u2__abc_44228_n14402) );
  AND2X2 AND2X2_6314 ( .A(u2__abc_44228_n14399), .B(u2__abc_44228_n14402), .Y(u2__abc_44228_n14403_1) );
  AND2X2 AND2X2_6315 ( .A(u2__abc_44228_n14404), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_remHi_400__FF_INPUT) );
  AND2X2 AND2X2_6316 ( .A(u2__abc_44228_n3062_bF_buf63), .B(u2_remHi_401_), .Y(u2__abc_44228_n14406) );
  AND2X2 AND2X2_6317 ( .A(u2__abc_44228_n14394), .B(u2__abc_44228_n7385), .Y(u2__abc_44228_n14407) );
  AND2X2 AND2X2_6318 ( .A(u2__abc_44228_n14407), .B(u2__abc_44228_n7219), .Y(u2__abc_44228_n14408) );
  AND2X2 AND2X2_6319 ( .A(u2__abc_44228_n14410), .B(u2__abc_44228_n14409), .Y(u2__abc_44228_n14411) );
  AND2X2 AND2X2_632 ( .A(u2__abc_44228_n3204), .B(sqrto_28_), .Y(u2__abc_44228_n3205) );
  AND2X2 AND2X2_6320 ( .A(u2__abc_44228_n14412), .B(u2__abc_44228_n7547_bF_buf3), .Y(u2__abc_44228_n14413_1) );
  AND2X2 AND2X2_6321 ( .A(u2__abc_44228_n7548_1_bF_buf4), .B(u2_remHi_399_), .Y(u2__abc_44228_n14414) );
  AND2X2 AND2X2_6322 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n7196), .Y(u2__abc_44228_n14417) );
  AND2X2 AND2X2_6323 ( .A(u2__abc_44228_n14418), .B(u2__abc_44228_n2972_bF_buf28), .Y(u2__abc_44228_n14419) );
  AND2X2 AND2X2_6324 ( .A(u2__abc_44228_n14416), .B(u2__abc_44228_n14419), .Y(u2__abc_44228_n14420) );
  AND2X2 AND2X2_6325 ( .A(u2__abc_44228_n14421_1), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_remHi_401__FF_INPUT) );
  AND2X2 AND2X2_6326 ( .A(u2__abc_44228_n3062_bF_buf62), .B(u2_remHi_402_), .Y(u2__abc_44228_n14423) );
  AND2X2 AND2X2_6327 ( .A(u2__abc_44228_n14394), .B(u2__abc_44228_n7386), .Y(u2__abc_44228_n14424) );
  AND2X2 AND2X2_6328 ( .A(u2__abc_44228_n14426), .B(u2__abc_44228_n7205), .Y(u2__abc_44228_n14427) );
  AND2X2 AND2X2_6329 ( .A(u2__abc_44228_n14428), .B(u2__abc_44228_n14429), .Y(u2__abc_44228_n14430_1) );
  AND2X2 AND2X2_633 ( .A(u2__abc_44228_n3207), .B(u2__abc_44228_n3201), .Y(u2__abc_44228_n3208) );
  AND2X2 AND2X2_6330 ( .A(u2__abc_44228_n14430_1), .B(u2__abc_44228_n7547_bF_buf2), .Y(u2__abc_44228_n14431) );
  AND2X2 AND2X2_6331 ( .A(u2__abc_44228_n7548_1_bF_buf3), .B(u2_remHi_400_), .Y(u2__abc_44228_n14432) );
  AND2X2 AND2X2_6332 ( .A(u2__abc_44228_n2983_bF_buf127), .B(u2__abc_44228_n7187), .Y(u2__abc_44228_n14435) );
  AND2X2 AND2X2_6333 ( .A(u2__abc_44228_n14436), .B(u2__abc_44228_n2972_bF_buf27), .Y(u2__abc_44228_n14437) );
  AND2X2 AND2X2_6334 ( .A(u2__abc_44228_n14434), .B(u2__abc_44228_n14437), .Y(u2__abc_44228_n14438_1) );
  AND2X2 AND2X2_6335 ( .A(u2__abc_44228_n14439), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_remHi_402__FF_INPUT) );
  AND2X2 AND2X2_6336 ( .A(u2__abc_44228_n3062_bF_buf61), .B(u2_remHi_403_), .Y(u2__abc_44228_n14441) );
  AND2X2 AND2X2_6337 ( .A(u2__abc_44228_n14446), .B(u2__abc_44228_n7547_bF_buf1), .Y(u2__abc_44228_n14447) );
  AND2X2 AND2X2_6338 ( .A(u2__abc_44228_n14447), .B(u2__abc_44228_n14445), .Y(u2__abc_44228_n14448) );
  AND2X2 AND2X2_6339 ( .A(u2__abc_44228_n7548_1_bF_buf2), .B(u2_remHi_401_), .Y(u2__abc_44228_n14449) );
  AND2X2 AND2X2_634 ( .A(u2__abc_44228_n3209), .B(u2_remHi_26_), .Y(u2__abc_44228_n3210) );
  AND2X2 AND2X2_6340 ( .A(u2__abc_44228_n2983_bF_buf125), .B(u2__abc_44228_n7181), .Y(u2__abc_44228_n14452) );
  AND2X2 AND2X2_6341 ( .A(u2__abc_44228_n14453), .B(u2__abc_44228_n2972_bF_buf26), .Y(u2__abc_44228_n14454) );
  AND2X2 AND2X2_6342 ( .A(u2__abc_44228_n14451), .B(u2__abc_44228_n14454), .Y(u2__abc_44228_n14455) );
  AND2X2 AND2X2_6343 ( .A(u2__abc_44228_n14456), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_remHi_403__FF_INPUT) );
  AND2X2 AND2X2_6344 ( .A(u2__abc_44228_n3062_bF_buf60), .B(u2_remHi_404_), .Y(u2__abc_44228_n14458_1) );
  AND2X2 AND2X2_6345 ( .A(u2__abc_44228_n14391), .B(u2__abc_44228_n7221), .Y(u2__abc_44228_n14459) );
  AND2X2 AND2X2_6346 ( .A(u2__abc_44228_n14460), .B(u2__abc_44228_n7190), .Y(u2__abc_44228_n14462) );
  AND2X2 AND2X2_6347 ( .A(u2__abc_44228_n14463), .B(u2__abc_44228_n14461), .Y(u2__abc_44228_n14464) );
  AND2X2 AND2X2_6348 ( .A(u2__abc_44228_n14464), .B(u2__abc_44228_n7547_bF_buf0), .Y(u2__abc_44228_n14465) );
  AND2X2 AND2X2_6349 ( .A(u2__abc_44228_n7548_1_bF_buf1), .B(u2_remHi_402_), .Y(u2__abc_44228_n14466) );
  AND2X2 AND2X2_635 ( .A(u2__abc_44228_n3211), .B(sqrto_26_), .Y(u2__abc_44228_n3212) );
  AND2X2 AND2X2_6350 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n7173), .Y(u2__abc_44228_n14469) );
  AND2X2 AND2X2_6351 ( .A(u2__abc_44228_n14470), .B(u2__abc_44228_n2972_bF_buf25), .Y(u2__abc_44228_n14471) );
  AND2X2 AND2X2_6352 ( .A(u2__abc_44228_n14468), .B(u2__abc_44228_n14471), .Y(u2__abc_44228_n14472) );
  AND2X2 AND2X2_6353 ( .A(u2__abc_44228_n14473), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_remHi_404__FF_INPUT) );
  AND2X2 AND2X2_6354 ( .A(u2__abc_44228_n3062_bF_buf59), .B(u2_remHi_405_), .Y(u2__abc_44228_n14475_1) );
  AND2X2 AND2X2_6355 ( .A(u2__abc_44228_n14463), .B(u2__abc_44228_n7394), .Y(u2__abc_44228_n14477) );
  AND2X2 AND2X2_6356 ( .A(u2__abc_44228_n14480), .B(u2__abc_44228_n14478), .Y(u2__abc_44228_n14481) );
  AND2X2 AND2X2_6357 ( .A(u2__abc_44228_n14481), .B(u2__abc_44228_n7547_bF_buf57), .Y(u2__abc_44228_n14482) );
  AND2X2 AND2X2_6358 ( .A(u2__abc_44228_n7548_1_bF_buf0), .B(u2_remHi_403_), .Y(u2__abc_44228_n14483) );
  AND2X2 AND2X2_6359 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n7167), .Y(u2__abc_44228_n14486) );
  AND2X2 AND2X2_636 ( .A(u2__abc_44228_n3215), .B(u2_remHi_27_), .Y(u2__abc_44228_n3216) );
  AND2X2 AND2X2_6360 ( .A(u2__abc_44228_n14487), .B(u2__abc_44228_n2972_bF_buf24), .Y(u2__abc_44228_n14488) );
  AND2X2 AND2X2_6361 ( .A(u2__abc_44228_n14485_1), .B(u2__abc_44228_n14488), .Y(u2__abc_44228_n14489) );
  AND2X2 AND2X2_6362 ( .A(u2__abc_44228_n14490), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_remHi_405__FF_INPUT) );
  AND2X2 AND2X2_6363 ( .A(u2__abc_44228_n3062_bF_buf58), .B(u2_remHi_406_), .Y(u2__abc_44228_n14492) );
  AND2X2 AND2X2_6364 ( .A(u2__abc_44228_n14460), .B(u2__abc_44228_n7191), .Y(u2__abc_44228_n14493_1) );
  AND2X2 AND2X2_6365 ( .A(u2__abc_44228_n14494), .B(u2__abc_44228_n7176), .Y(u2__abc_44228_n14495) );
  AND2X2 AND2X2_6366 ( .A(u2__abc_44228_n14496), .B(u2__abc_44228_n14497), .Y(u2__abc_44228_n14498) );
  AND2X2 AND2X2_6367 ( .A(u2__abc_44228_n14498), .B(u2__abc_44228_n7547_bF_buf56), .Y(u2__abc_44228_n14499) );
  AND2X2 AND2X2_6368 ( .A(u2__abc_44228_n7548_1_bF_buf57), .B(u2_remHi_404_), .Y(u2__abc_44228_n14500) );
  AND2X2 AND2X2_6369 ( .A(u2__abc_44228_n2983_bF_buf121), .B(u2__abc_44228_n7157), .Y(u2__abc_44228_n14503) );
  AND2X2 AND2X2_637 ( .A(u2__abc_44228_n3218), .B(sqrto_27_), .Y(u2__abc_44228_n3219) );
  AND2X2 AND2X2_6370 ( .A(u2__abc_44228_n14504), .B(u2__abc_44228_n2972_bF_buf23), .Y(u2__abc_44228_n14505) );
  AND2X2 AND2X2_6371 ( .A(u2__abc_44228_n14502_1), .B(u2__abc_44228_n14505), .Y(u2__abc_44228_n14506) );
  AND2X2 AND2X2_6372 ( .A(u2__abc_44228_n14507), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_remHi_406__FF_INPUT) );
  AND2X2 AND2X2_6373 ( .A(u2__abc_44228_n3062_bF_buf57), .B(u2_remHi_407_), .Y(u2__abc_44228_n14509) );
  AND2X2 AND2X2_6374 ( .A(u2__abc_44228_n14514), .B(u2__abc_44228_n7547_bF_buf55), .Y(u2__abc_44228_n14515) );
  AND2X2 AND2X2_6375 ( .A(u2__abc_44228_n14515), .B(u2__abc_44228_n14513), .Y(u2__abc_44228_n14516) );
  AND2X2 AND2X2_6376 ( .A(u2__abc_44228_n7548_1_bF_buf56), .B(u2_remHi_405_), .Y(u2__abc_44228_n14517) );
  AND2X2 AND2X2_6377 ( .A(u2__abc_44228_n2983_bF_buf119), .B(u2__abc_44228_n7151), .Y(u2__abc_44228_n14520) );
  AND2X2 AND2X2_6378 ( .A(u2__abc_44228_n14521_1), .B(u2__abc_44228_n2972_bF_buf22), .Y(u2__abc_44228_n14522) );
  AND2X2 AND2X2_6379 ( .A(u2__abc_44228_n14519), .B(u2__abc_44228_n14522), .Y(u2__abc_44228_n14523) );
  AND2X2 AND2X2_638 ( .A(u2__abc_44228_n3217), .B(u2__abc_44228_n3220), .Y(u2__abc_44228_n3221) );
  AND2X2 AND2X2_6380 ( .A(u2__abc_44228_n14524), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_remHi_407__FF_INPUT) );
  AND2X2 AND2X2_6381 ( .A(u2__abc_44228_n3062_bF_buf56), .B(u2_remHi_408_), .Y(u2__abc_44228_n14526) );
  AND2X2 AND2X2_6382 ( .A(u2__abc_44228_n14391), .B(u2__abc_44228_n7222), .Y(u2__abc_44228_n14527) );
  AND2X2 AND2X2_6383 ( .A(u2__abc_44228_n14528), .B(u2__abc_44228_n7160), .Y(u2__abc_44228_n14529_1) );
  AND2X2 AND2X2_6384 ( .A(u2__abc_44228_n14530), .B(u2__abc_44228_n14531), .Y(u2__abc_44228_n14532) );
  AND2X2 AND2X2_6385 ( .A(u2__abc_44228_n14532), .B(u2__abc_44228_n7547_bF_buf54), .Y(u2__abc_44228_n14533) );
  AND2X2 AND2X2_6386 ( .A(u2__abc_44228_n7548_1_bF_buf55), .B(u2_remHi_406_), .Y(u2__abc_44228_n14534) );
  AND2X2 AND2X2_6387 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n7143_1), .Y(u2__abc_44228_n14537) );
  AND2X2 AND2X2_6388 ( .A(u2__abc_44228_n14538_1), .B(u2__abc_44228_n2972_bF_buf21), .Y(u2__abc_44228_n14539) );
  AND2X2 AND2X2_6389 ( .A(u2__abc_44228_n14536), .B(u2__abc_44228_n14539), .Y(u2__abc_44228_n14540) );
  AND2X2 AND2X2_639 ( .A(u2__abc_44228_n3214), .B(u2__abc_44228_n3221), .Y(u2__abc_44228_n3222) );
  AND2X2 AND2X2_6390 ( .A(u2__abc_44228_n14541), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_remHi_408__FF_INPUT) );
  AND2X2 AND2X2_6391 ( .A(u2__abc_44228_n3062_bF_buf55), .B(u2_remHi_409_), .Y(u2__abc_44228_n14543) );
  AND2X2 AND2X2_6392 ( .A(u2__abc_44228_n14530), .B(u2__abc_44228_n7406), .Y(u2__abc_44228_n14545) );
  AND2X2 AND2X2_6393 ( .A(u2__abc_44228_n14548), .B(u2__abc_44228_n14546_1), .Y(u2__abc_44228_n14549) );
  AND2X2 AND2X2_6394 ( .A(u2__abc_44228_n14549), .B(u2__abc_44228_n7547_bF_buf53), .Y(u2__abc_44228_n14550) );
  AND2X2 AND2X2_6395 ( .A(u2__abc_44228_n7548_1_bF_buf54), .B(u2_remHi_407_), .Y(u2__abc_44228_n14551) );
  AND2X2 AND2X2_6396 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n7137), .Y(u2__abc_44228_n14554) );
  AND2X2 AND2X2_6397 ( .A(u2__abc_44228_n14555), .B(u2__abc_44228_n2972_bF_buf20), .Y(u2__abc_44228_n14556_1) );
  AND2X2 AND2X2_6398 ( .A(u2__abc_44228_n14553), .B(u2__abc_44228_n14556_1), .Y(u2__abc_44228_n14557) );
  AND2X2 AND2X2_6399 ( .A(u2__abc_44228_n14558), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_remHi_409__FF_INPUT) );
  AND2X2 AND2X2_64 ( .A(_abc_64468_n753_bF_buf6), .B(sqrto_63_), .Y(_auto_iopadmap_cc_313_execute_65414_99_) );
  AND2X2 AND2X2_640 ( .A(u2__abc_44228_n3208), .B(u2__abc_44228_n3222), .Y(u2__abc_44228_n3223) );
  AND2X2 AND2X2_6400 ( .A(u2__abc_44228_n3062_bF_buf54), .B(u2_remHi_410_), .Y(u2__abc_44228_n14560) );
  AND2X2 AND2X2_6401 ( .A(u2__abc_44228_n14530), .B(u2__abc_44228_n7407), .Y(u2__abc_44228_n14561) );
  AND2X2 AND2X2_6402 ( .A(u2__abc_44228_n14563), .B(u2__abc_44228_n7146), .Y(u2__abc_44228_n14564_1) );
  AND2X2 AND2X2_6403 ( .A(u2__abc_44228_n14565), .B(u2__abc_44228_n14566), .Y(u2__abc_44228_n14567) );
  AND2X2 AND2X2_6404 ( .A(u2__abc_44228_n14567), .B(u2__abc_44228_n7547_bF_buf52), .Y(u2__abc_44228_n14568) );
  AND2X2 AND2X2_6405 ( .A(u2__abc_44228_n7548_1_bF_buf53), .B(u2_remHi_408_), .Y(u2__abc_44228_n14569) );
  AND2X2 AND2X2_6406 ( .A(u2__abc_44228_n2983_bF_buf115), .B(u2__abc_44228_n7128), .Y(u2__abc_44228_n14572) );
  AND2X2 AND2X2_6407 ( .A(u2__abc_44228_n14573_1), .B(u2__abc_44228_n2972_bF_buf19), .Y(u2__abc_44228_n14574) );
  AND2X2 AND2X2_6408 ( .A(u2__abc_44228_n14571), .B(u2__abc_44228_n14574), .Y(u2__abc_44228_n14575) );
  AND2X2 AND2X2_6409 ( .A(u2__abc_44228_n14576), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_remHi_410__FF_INPUT) );
  AND2X2 AND2X2_641 ( .A(u2__abc_44228_n3224), .B(u2_remHi_23_), .Y(u2__abc_44228_n3225) );
  AND2X2 AND2X2_6410 ( .A(u2__abc_44228_n3062_bF_buf53), .B(u2_remHi_411_), .Y(u2__abc_44228_n14578) );
  AND2X2 AND2X2_6411 ( .A(u2__abc_44228_n14583), .B(u2__abc_44228_n7547_bF_buf51), .Y(u2__abc_44228_n14584) );
  AND2X2 AND2X2_6412 ( .A(u2__abc_44228_n14584), .B(u2__abc_44228_n14582), .Y(u2__abc_44228_n14585) );
  AND2X2 AND2X2_6413 ( .A(u2__abc_44228_n7548_1_bF_buf52), .B(u2_remHi_409_), .Y(u2__abc_44228_n14586) );
  AND2X2 AND2X2_6414 ( .A(u2__abc_44228_n2983_bF_buf113), .B(u2__abc_44228_n7122), .Y(u2__abc_44228_n14589) );
  AND2X2 AND2X2_6415 ( .A(u2__abc_44228_n14590), .B(u2__abc_44228_n2972_bF_buf18), .Y(u2__abc_44228_n14591) );
  AND2X2 AND2X2_6416 ( .A(u2__abc_44228_n14588), .B(u2__abc_44228_n14591), .Y(u2__abc_44228_n14592) );
  AND2X2 AND2X2_6417 ( .A(u2__abc_44228_n14593), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_remHi_411__FF_INPUT) );
  AND2X2 AND2X2_6418 ( .A(u2__abc_44228_n3062_bF_buf52), .B(u2_remHi_412_), .Y(u2__abc_44228_n14595) );
  AND2X2 AND2X2_6419 ( .A(u2__abc_44228_n14528), .B(u2__abc_44228_n7162), .Y(u2__abc_44228_n14596) );
  AND2X2 AND2X2_642 ( .A(u2__abc_44228_n3227), .B(sqrto_23_), .Y(u2__abc_44228_n3228) );
  AND2X2 AND2X2_6420 ( .A(u2__abc_44228_n14597), .B(u2__abc_44228_n7131), .Y(u2__abc_44228_n14599) );
  AND2X2 AND2X2_6421 ( .A(u2__abc_44228_n14600), .B(u2__abc_44228_n14598), .Y(u2__abc_44228_n14601) );
  AND2X2 AND2X2_6422 ( .A(u2__abc_44228_n14601), .B(u2__abc_44228_n7547_bF_buf50), .Y(u2__abc_44228_n14602_1) );
  AND2X2 AND2X2_6423 ( .A(u2__abc_44228_n7548_1_bF_buf51), .B(u2_remHi_410_), .Y(u2__abc_44228_n14603) );
  AND2X2 AND2X2_6424 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n7114), .Y(u2__abc_44228_n14606) );
  AND2X2 AND2X2_6425 ( .A(u2__abc_44228_n14607), .B(u2__abc_44228_n2972_bF_buf17), .Y(u2__abc_44228_n14608) );
  AND2X2 AND2X2_6426 ( .A(u2__abc_44228_n14605), .B(u2__abc_44228_n14608), .Y(u2__abc_44228_n14609) );
  AND2X2 AND2X2_6427 ( .A(u2__abc_44228_n14610), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_remHi_412__FF_INPUT) );
  AND2X2 AND2X2_6428 ( .A(u2__abc_44228_n3062_bF_buf51), .B(u2_remHi_413_), .Y(u2__abc_44228_n14612) );
  AND2X2 AND2X2_6429 ( .A(u2__abc_44228_n14600), .B(u2__abc_44228_n7413), .Y(u2__abc_44228_n14613) );
  AND2X2 AND2X2_643 ( .A(u2__abc_44228_n3226), .B(u2__abc_44228_n3229), .Y(u2__abc_44228_n3230) );
  AND2X2 AND2X2_6430 ( .A(u2__abc_44228_n14617), .B(u2__abc_44228_n7547_bF_buf49), .Y(u2__abc_44228_n14618) );
  AND2X2 AND2X2_6431 ( .A(u2__abc_44228_n14618), .B(u2__abc_44228_n14615), .Y(u2__abc_44228_n14619_1) );
  AND2X2 AND2X2_6432 ( .A(u2__abc_44228_n7548_1_bF_buf50), .B(u2_remHi_411_), .Y(u2__abc_44228_n14620) );
  AND2X2 AND2X2_6433 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n7108), .Y(u2__abc_44228_n14623) );
  AND2X2 AND2X2_6434 ( .A(u2__abc_44228_n14624), .B(u2__abc_44228_n2972_bF_buf16), .Y(u2__abc_44228_n14625) );
  AND2X2 AND2X2_6435 ( .A(u2__abc_44228_n14622), .B(u2__abc_44228_n14625), .Y(u2__abc_44228_n14626) );
  AND2X2 AND2X2_6436 ( .A(u2__abc_44228_n14627), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_remHi_413__FF_INPUT) );
  AND2X2 AND2X2_6437 ( .A(u2__abc_44228_n3062_bF_buf50), .B(u2_remHi_414_), .Y(u2__abc_44228_n14629_1) );
  AND2X2 AND2X2_6438 ( .A(u2__abc_44228_n14600), .B(u2__abc_44228_n7414), .Y(u2__abc_44228_n14630) );
  AND2X2 AND2X2_6439 ( .A(u2__abc_44228_n14632), .B(u2__abc_44228_n7117), .Y(u2__abc_44228_n14633) );
  AND2X2 AND2X2_644 ( .A(u2__abc_44228_n3231), .B(u2_remHi_22_), .Y(u2__abc_44228_n3232) );
  AND2X2 AND2X2_6440 ( .A(u2__abc_44228_n14634), .B(u2__abc_44228_n14635), .Y(u2__abc_44228_n14636) );
  AND2X2 AND2X2_6441 ( .A(u2__abc_44228_n14636), .B(u2__abc_44228_n7547_bF_buf48), .Y(u2__abc_44228_n14637_1) );
  AND2X2 AND2X2_6442 ( .A(u2__abc_44228_n7548_1_bF_buf49), .B(u2_remHi_412_), .Y(u2__abc_44228_n14638) );
  AND2X2 AND2X2_6443 ( .A(u2__abc_44228_n2983_bF_buf109), .B(u2__abc_44228_n7089), .Y(u2__abc_44228_n14641) );
  AND2X2 AND2X2_6444 ( .A(u2__abc_44228_n14642), .B(u2__abc_44228_n2972_bF_buf15), .Y(u2__abc_44228_n14643) );
  AND2X2 AND2X2_6445 ( .A(u2__abc_44228_n14640), .B(u2__abc_44228_n14643), .Y(u2__abc_44228_n14644) );
  AND2X2 AND2X2_6446 ( .A(u2__abc_44228_n14645), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_remHi_414__FF_INPUT) );
  AND2X2 AND2X2_6447 ( .A(u2__abc_44228_n3062_bF_buf49), .B(u2_remHi_415_), .Y(u2__abc_44228_n14647) );
  AND2X2 AND2X2_6448 ( .A(u2__abc_44228_n14652), .B(u2__abc_44228_n7547_bF_buf47), .Y(u2__abc_44228_n14653) );
  AND2X2 AND2X2_6449 ( .A(u2__abc_44228_n14653), .B(u2__abc_44228_n14651), .Y(u2__abc_44228_n14654_1) );
  AND2X2 AND2X2_645 ( .A(u2__abc_44228_n3233), .B(sqrto_22_), .Y(u2__abc_44228_n3234) );
  AND2X2 AND2X2_6450 ( .A(u2__abc_44228_n7548_1_bF_buf48), .B(u2_remHi_413_), .Y(u2__abc_44228_n14655) );
  AND2X2 AND2X2_6451 ( .A(u2__abc_44228_n2983_bF_buf107), .B(u2__abc_44228_n7096), .Y(u2__abc_44228_n14658) );
  AND2X2 AND2X2_6452 ( .A(u2__abc_44228_n14659), .B(u2__abc_44228_n2972_bF_buf14), .Y(u2__abc_44228_n14660) );
  AND2X2 AND2X2_6453 ( .A(u2__abc_44228_n14657), .B(u2__abc_44228_n14660), .Y(u2__abc_44228_n14661) );
  AND2X2 AND2X2_6454 ( .A(u2__abc_44228_n14662), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_remHi_415__FF_INPUT) );
  AND2X2 AND2X2_6455 ( .A(u2__abc_44228_n3062_bF_buf48), .B(u2_remHi_416_), .Y(u2__abc_44228_n14664) );
  AND2X2 AND2X2_6456 ( .A(u2__abc_44228_n6865), .B(u2__abc_44228_n7343), .Y(u2__abc_44228_n14665_1) );
  AND2X2 AND2X2_6457 ( .A(u2__abc_44228_n14666), .B(u2__abc_44228_n7092), .Y(u2__abc_44228_n14667) );
  AND2X2 AND2X2_6458 ( .A(u2__abc_44228_n14668), .B(u2__abc_44228_n14669), .Y(u2__abc_44228_n14670) );
  AND2X2 AND2X2_6459 ( .A(u2__abc_44228_n14671), .B(u2__abc_44228_n14672), .Y(u2__abc_44228_n14673_1) );
  AND2X2 AND2X2_646 ( .A(u2__abc_44228_n3236), .B(u2__abc_44228_n3230), .Y(u2__abc_44228_n3237) );
  AND2X2 AND2X2_6460 ( .A(u2__abc_44228_n2983_bF_buf105), .B(u2__abc_44228_n7082), .Y(u2__abc_44228_n14675) );
  AND2X2 AND2X2_6461 ( .A(u2__abc_44228_n14676), .B(u2__abc_44228_n2972_bF_buf13), .Y(u2__abc_44228_n14677) );
  AND2X2 AND2X2_6462 ( .A(u2__abc_44228_n14674), .B(u2__abc_44228_n14677), .Y(u2__abc_44228_n14678) );
  AND2X2 AND2X2_6463 ( .A(u2__abc_44228_n14679), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_remHi_416__FF_INPUT) );
  AND2X2 AND2X2_6464 ( .A(u2__abc_44228_n3062_bF_buf47), .B(u2_remHi_417_), .Y(u2__abc_44228_n14681) );
  AND2X2 AND2X2_6465 ( .A(u2__abc_44228_n14668), .B(u2__abc_44228_n7425), .Y(u2__abc_44228_n14682_1) );
  AND2X2 AND2X2_6466 ( .A(u2__abc_44228_n14682_1), .B(u2__abc_44228_n7099), .Y(u2__abc_44228_n14683) );
  AND2X2 AND2X2_6467 ( .A(u2__abc_44228_n14685), .B(u2__abc_44228_n14684), .Y(u2__abc_44228_n14686) );
  AND2X2 AND2X2_6468 ( .A(u2__abc_44228_n14687), .B(u2__abc_44228_n7547_bF_buf45), .Y(u2__abc_44228_n14688) );
  AND2X2 AND2X2_6469 ( .A(u2__abc_44228_n7548_1_bF_buf46), .B(u2_remHi_415_), .Y(u2__abc_44228_n14689) );
  AND2X2 AND2X2_647 ( .A(u2__abc_44228_n3238), .B(u2_remHi_25_), .Y(u2__abc_44228_n3239) );
  AND2X2 AND2X2_6470 ( .A(u2__abc_44228_n2983_bF_buf103), .B(u2__abc_44228_n7076), .Y(u2__abc_44228_n14692) );
  AND2X2 AND2X2_6471 ( .A(u2__abc_44228_n14693), .B(u2__abc_44228_n2972_bF_buf12), .Y(u2__abc_44228_n14694) );
  AND2X2 AND2X2_6472 ( .A(u2__abc_44228_n14691), .B(u2__abc_44228_n14694), .Y(u2__abc_44228_n14695) );
  AND2X2 AND2X2_6473 ( .A(u2__abc_44228_n14696), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_remHi_417__FF_INPUT) );
  AND2X2 AND2X2_6474 ( .A(u2__abc_44228_n3062_bF_buf46), .B(u2_remHi_418_), .Y(u2__abc_44228_n14698) );
  AND2X2 AND2X2_6475 ( .A(u2__abc_44228_n14668), .B(u2__abc_44228_n7426), .Y(u2__abc_44228_n14699) );
  AND2X2 AND2X2_6476 ( .A(u2__abc_44228_n14701), .B(u2__abc_44228_n7085), .Y(u2__abc_44228_n14702) );
  AND2X2 AND2X2_6477 ( .A(u2__abc_44228_n14703), .B(u2__abc_44228_n14704), .Y(u2__abc_44228_n14705) );
  AND2X2 AND2X2_6478 ( .A(u2__abc_44228_n14705), .B(u2__abc_44228_n7547_bF_buf44), .Y(u2__abc_44228_n14706) );
  AND2X2 AND2X2_6479 ( .A(u2__abc_44228_n7548_1_bF_buf45), .B(u2_remHi_416_), .Y(u2__abc_44228_n14707) );
  AND2X2 AND2X2_648 ( .A(u2__abc_44228_n3241), .B(sqrto_25_), .Y(u2__abc_44228_n3242) );
  AND2X2 AND2X2_6480 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n7067), .Y(u2__abc_44228_n14710) );
  AND2X2 AND2X2_6481 ( .A(u2__abc_44228_n14711), .B(u2__abc_44228_n2972_bF_buf11), .Y(u2__abc_44228_n14712) );
  AND2X2 AND2X2_6482 ( .A(u2__abc_44228_n14709), .B(u2__abc_44228_n14712), .Y(u2__abc_44228_n14713) );
  AND2X2 AND2X2_6483 ( .A(u2__abc_44228_n14714), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_remHi_418__FF_INPUT) );
  AND2X2 AND2X2_6484 ( .A(u2__abc_44228_n3062_bF_buf45), .B(u2_remHi_419_), .Y(u2__abc_44228_n14716) );
  AND2X2 AND2X2_6485 ( .A(u2__abc_44228_n14721), .B(u2__abc_44228_n7547_bF_buf43), .Y(u2__abc_44228_n14722) );
  AND2X2 AND2X2_6486 ( .A(u2__abc_44228_n14722), .B(u2__abc_44228_n14720), .Y(u2__abc_44228_n14723) );
  AND2X2 AND2X2_6487 ( .A(u2__abc_44228_n7548_1_bF_buf44), .B(u2_remHi_417_), .Y(u2__abc_44228_n14724) );
  AND2X2 AND2X2_6488 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n7061), .Y(u2__abc_44228_n14727) );
  AND2X2 AND2X2_6489 ( .A(u2__abc_44228_n14728), .B(u2__abc_44228_n2972_bF_buf10), .Y(u2__abc_44228_n14729) );
  AND2X2 AND2X2_649 ( .A(u2__abc_44228_n3240), .B(u2__abc_44228_n3243), .Y(u2__abc_44228_n3244) );
  AND2X2 AND2X2_6490 ( .A(u2__abc_44228_n14726), .B(u2__abc_44228_n14729), .Y(u2__abc_44228_n14730) );
  AND2X2 AND2X2_6491 ( .A(u2__abc_44228_n14731), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_remHi_419__FF_INPUT) );
  AND2X2 AND2X2_6492 ( .A(u2__abc_44228_n3062_bF_buf44), .B(u2_remHi_420_), .Y(u2__abc_44228_n14733) );
  AND2X2 AND2X2_6493 ( .A(u2__abc_44228_n14666), .B(u2__abc_44228_n7101), .Y(u2__abc_44228_n14734) );
  AND2X2 AND2X2_6494 ( .A(u2__abc_44228_n14735), .B(u2__abc_44228_n7070), .Y(u2__abc_44228_n14737_1) );
  AND2X2 AND2X2_6495 ( .A(u2__abc_44228_n14738), .B(u2__abc_44228_n14736), .Y(u2__abc_44228_n14739) );
  AND2X2 AND2X2_6496 ( .A(u2__abc_44228_n14739), .B(u2__abc_44228_n7547_bF_buf42), .Y(u2__abc_44228_n14740) );
  AND2X2 AND2X2_6497 ( .A(u2__abc_44228_n7548_1_bF_buf43), .B(u2_remHi_418_), .Y(u2__abc_44228_n14741) );
  AND2X2 AND2X2_6498 ( .A(u2__abc_44228_n2983_bF_buf99), .B(u2__abc_44228_n7053), .Y(u2__abc_44228_n14744) );
  AND2X2 AND2X2_6499 ( .A(u2__abc_44228_n14745_1), .B(u2__abc_44228_n2972_bF_buf9), .Y(u2__abc_44228_n14746) );
  AND2X2 AND2X2_65 ( .A(_abc_64468_n753_bF_buf5), .B(sqrto_64_), .Y(_auto_iopadmap_cc_313_execute_65414_100_) );
  AND2X2 AND2X2_650 ( .A(u2__abc_44228_n3245), .B(u2_remHi_24_), .Y(u2__abc_44228_n3246) );
  AND2X2 AND2X2_6500 ( .A(u2__abc_44228_n14743), .B(u2__abc_44228_n14746), .Y(u2__abc_44228_n14747) );
  AND2X2 AND2X2_6501 ( .A(u2__abc_44228_n14748), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_remHi_420__FF_INPUT) );
  AND2X2 AND2X2_6502 ( .A(u2__abc_44228_n3062_bF_buf43), .B(u2_remHi_421_), .Y(u2__abc_44228_n14750) );
  AND2X2 AND2X2_6503 ( .A(u2__abc_44228_n14738), .B(u2__abc_44228_n7434), .Y(u2__abc_44228_n14752) );
  AND2X2 AND2X2_6504 ( .A(u2__abc_44228_n14755), .B(u2__abc_44228_n14753), .Y(u2__abc_44228_n14756) );
  AND2X2 AND2X2_6505 ( .A(u2__abc_44228_n14756), .B(u2__abc_44228_n7547_bF_buf41), .Y(u2__abc_44228_n14757) );
  AND2X2 AND2X2_6506 ( .A(u2__abc_44228_n7548_1_bF_buf42), .B(u2_remHi_419_), .Y(u2__abc_44228_n14758) );
  AND2X2 AND2X2_6507 ( .A(u2__abc_44228_n2983_bF_buf97), .B(u2__abc_44228_n7047), .Y(u2__abc_44228_n14761) );
  AND2X2 AND2X2_6508 ( .A(u2__abc_44228_n14762_1), .B(u2__abc_44228_n2972_bF_buf8), .Y(u2__abc_44228_n14763) );
  AND2X2 AND2X2_6509 ( .A(u2__abc_44228_n14760), .B(u2__abc_44228_n14763), .Y(u2__abc_44228_n14764) );
  AND2X2 AND2X2_651 ( .A(u2__abc_44228_n3247), .B(sqrto_24_), .Y(u2__abc_44228_n3248) );
  AND2X2 AND2X2_6510 ( .A(u2__abc_44228_n14765), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_remHi_421__FF_INPUT) );
  AND2X2 AND2X2_6511 ( .A(u2__abc_44228_n3062_bF_buf42), .B(u2_remHi_422_), .Y(u2__abc_44228_n14767) );
  AND2X2 AND2X2_6512 ( .A(u2__abc_44228_n14735), .B(u2__abc_44228_n7071), .Y(u2__abc_44228_n14768) );
  AND2X2 AND2X2_6513 ( .A(u2__abc_44228_n14769), .B(u2__abc_44228_n7056), .Y(u2__abc_44228_n14770) );
  AND2X2 AND2X2_6514 ( .A(u2__abc_44228_n14771), .B(u2__abc_44228_n14772_1), .Y(u2__abc_44228_n14773) );
  AND2X2 AND2X2_6515 ( .A(u2__abc_44228_n14773), .B(u2__abc_44228_n7547_bF_buf40), .Y(u2__abc_44228_n14774) );
  AND2X2 AND2X2_6516 ( .A(u2__abc_44228_n7548_1_bF_buf41), .B(u2_remHi_420_), .Y(u2__abc_44228_n14775) );
  AND2X2 AND2X2_6517 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n7037), .Y(u2__abc_44228_n14778) );
  AND2X2 AND2X2_6518 ( .A(u2__abc_44228_n14779), .B(u2__abc_44228_n2972_bF_buf7), .Y(u2__abc_44228_n14780_1) );
  AND2X2 AND2X2_6519 ( .A(u2__abc_44228_n14777), .B(u2__abc_44228_n14780_1), .Y(u2__abc_44228_n14781) );
  AND2X2 AND2X2_652 ( .A(u2__abc_44228_n3250), .B(u2__abc_44228_n3244), .Y(u2__abc_44228_n3251) );
  AND2X2 AND2X2_6520 ( .A(u2__abc_44228_n14782), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_remHi_422__FF_INPUT) );
  AND2X2 AND2X2_6521 ( .A(u2__abc_44228_n3062_bF_buf41), .B(u2_remHi_423_), .Y(u2__abc_44228_n14784) );
  AND2X2 AND2X2_6522 ( .A(u2__abc_44228_n14789_1), .B(u2__abc_44228_n7547_bF_buf39), .Y(u2__abc_44228_n14790) );
  AND2X2 AND2X2_6523 ( .A(u2__abc_44228_n14790), .B(u2__abc_44228_n14788), .Y(u2__abc_44228_n14791) );
  AND2X2 AND2X2_6524 ( .A(u2__abc_44228_n7548_1_bF_buf40), .B(u2_remHi_421_), .Y(u2__abc_44228_n14792) );
  AND2X2 AND2X2_6525 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n7031), .Y(u2__abc_44228_n14795) );
  AND2X2 AND2X2_6526 ( .A(u2__abc_44228_n14796), .B(u2__abc_44228_n2972_bF_buf6), .Y(u2__abc_44228_n14797_1) );
  AND2X2 AND2X2_6527 ( .A(u2__abc_44228_n14794), .B(u2__abc_44228_n14797_1), .Y(u2__abc_44228_n14798) );
  AND2X2 AND2X2_6528 ( .A(u2__abc_44228_n14799), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_remHi_423__FF_INPUT) );
  AND2X2 AND2X2_6529 ( .A(u2__abc_44228_n3062_bF_buf40), .B(u2_remHi_424_), .Y(u2__abc_44228_n14801) );
  AND2X2 AND2X2_653 ( .A(u2__abc_44228_n3237), .B(u2__abc_44228_n3251), .Y(u2__abc_44228_n3252) );
  AND2X2 AND2X2_6530 ( .A(u2__abc_44228_n14666), .B(u2__abc_44228_n7102), .Y(u2__abc_44228_n14802) );
  AND2X2 AND2X2_6531 ( .A(u2__abc_44228_n14803), .B(u2__abc_44228_n7040), .Y(u2__abc_44228_n14804) );
  AND2X2 AND2X2_6532 ( .A(u2__abc_44228_n14805), .B(u2__abc_44228_n14806), .Y(u2__abc_44228_n14807) );
  AND2X2 AND2X2_6533 ( .A(u2__abc_44228_n14807), .B(u2__abc_44228_n7547_bF_buf38), .Y(u2__abc_44228_n14808_1) );
  AND2X2 AND2X2_6534 ( .A(u2__abc_44228_n7548_1_bF_buf39), .B(u2_remHi_422_), .Y(u2__abc_44228_n14809) );
  AND2X2 AND2X2_6535 ( .A(u2__abc_44228_n2983_bF_buf93), .B(u2__abc_44228_n7023), .Y(u2__abc_44228_n14812) );
  AND2X2 AND2X2_6536 ( .A(u2__abc_44228_n14813), .B(u2__abc_44228_n2972_bF_buf5), .Y(u2__abc_44228_n14814) );
  AND2X2 AND2X2_6537 ( .A(u2__abc_44228_n14811), .B(u2__abc_44228_n14814), .Y(u2__abc_44228_n14815) );
  AND2X2 AND2X2_6538 ( .A(u2__abc_44228_n14816_1), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_remHi_424__FF_INPUT) );
  AND2X2 AND2X2_6539 ( .A(u2__abc_44228_n3062_bF_buf39), .B(u2_remHi_425_), .Y(u2__abc_44228_n14818) );
  AND2X2 AND2X2_654 ( .A(u2__abc_44228_n3223), .B(u2__abc_44228_n3252), .Y(u2__abc_44228_n3253) );
  AND2X2 AND2X2_6540 ( .A(u2__abc_44228_n7548_1_bF_buf38), .B(u2_remHi_423_), .Y(u2__abc_44228_n14819) );
  AND2X2 AND2X2_6541 ( .A(u2__abc_44228_n14805), .B(u2__abc_44228_n7444), .Y(u2__abc_44228_n14822) );
  AND2X2 AND2X2_6542 ( .A(u2__abc_44228_n14825_1), .B(u2__abc_44228_n14823), .Y(u2__abc_44228_n14826) );
  AND2X2 AND2X2_6543 ( .A(u2__abc_44228_n14826), .B(u2__abc_44228_n7547_bF_buf37), .Y(u2__abc_44228_n14827) );
  AND2X2 AND2X2_6544 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n7017), .Y(u2__abc_44228_n14829) );
  AND2X2 AND2X2_6545 ( .A(u2__abc_44228_n14830), .B(u2__abc_44228_n2972_bF_buf4), .Y(u2__abc_44228_n14831) );
  AND2X2 AND2X2_6546 ( .A(u2__abc_44228_n14828), .B(u2__abc_44228_n14831), .Y(u2__abc_44228_n14832) );
  AND2X2 AND2X2_6547 ( .A(u2__abc_44228_n14833_1), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_remHi_425__FF_INPUT) );
  AND2X2 AND2X2_6548 ( .A(u2__abc_44228_n3062_bF_buf38), .B(u2_remHi_426_), .Y(u2__abc_44228_n14835) );
  AND2X2 AND2X2_6549 ( .A(u2__abc_44228_n14803), .B(u2__abc_44228_n7041), .Y(u2__abc_44228_n14836) );
  AND2X2 AND2X2_655 ( .A(u2__abc_44228_n3254), .B(u2_remHi_21_), .Y(u2__abc_44228_n3255) );
  AND2X2 AND2X2_6550 ( .A(u2__abc_44228_n14837), .B(u2__abc_44228_n7026), .Y(u2__abc_44228_n14838) );
  AND2X2 AND2X2_6551 ( .A(u2__abc_44228_n14839), .B(u2__abc_44228_n14840), .Y(u2__abc_44228_n14841) );
  AND2X2 AND2X2_6552 ( .A(u2__abc_44228_n14841), .B(u2__abc_44228_n7547_bF_buf36), .Y(u2__abc_44228_n14842) );
  AND2X2 AND2X2_6553 ( .A(u2__abc_44228_n7548_1_bF_buf37), .B(u2_remHi_424_), .Y(u2__abc_44228_n14843_1) );
  AND2X2 AND2X2_6554 ( .A(u2__abc_44228_n2983_bF_buf91), .B(u2__abc_44228_n7008), .Y(u2__abc_44228_n14846) );
  AND2X2 AND2X2_6555 ( .A(u2__abc_44228_n14847), .B(u2__abc_44228_n2972_bF_buf3), .Y(u2__abc_44228_n14848) );
  AND2X2 AND2X2_6556 ( .A(u2__abc_44228_n14845), .B(u2__abc_44228_n14848), .Y(u2__abc_44228_n14849) );
  AND2X2 AND2X2_6557 ( .A(u2__abc_44228_n14850), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_remHi_426__FF_INPUT) );
  AND2X2 AND2X2_6558 ( .A(u2__abc_44228_n3062_bF_buf37), .B(u2_remHi_427_), .Y(u2__abc_44228_n14852) );
  AND2X2 AND2X2_6559 ( .A(u2__abc_44228_n14839), .B(u2__abc_44228_n7449), .Y(u2__abc_44228_n14854) );
  AND2X2 AND2X2_656 ( .A(u2__abc_44228_n3257), .B(sqrto_21_), .Y(u2__abc_44228_n3258) );
  AND2X2 AND2X2_6560 ( .A(u2__abc_44228_n14857), .B(u2__abc_44228_n14855), .Y(u2__abc_44228_n14858) );
  AND2X2 AND2X2_6561 ( .A(u2__abc_44228_n14858), .B(u2__abc_44228_n7547_bF_buf35), .Y(u2__abc_44228_n14859) );
  AND2X2 AND2X2_6562 ( .A(u2__abc_44228_n7548_1_bF_buf36), .B(u2_remHi_425_), .Y(u2__abc_44228_n14860_1) );
  AND2X2 AND2X2_6563 ( .A(u2__abc_44228_n2983_bF_buf89), .B(u2__abc_44228_n7002), .Y(u2__abc_44228_n14863) );
  AND2X2 AND2X2_6564 ( .A(u2__abc_44228_n14864), .B(u2__abc_44228_n2972_bF_buf2), .Y(u2__abc_44228_n14865) );
  AND2X2 AND2X2_6565 ( .A(u2__abc_44228_n14862), .B(u2__abc_44228_n14865), .Y(u2__abc_44228_n14866) );
  AND2X2 AND2X2_6566 ( .A(u2__abc_44228_n14867), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_remHi_427__FF_INPUT) );
  AND2X2 AND2X2_6567 ( .A(u2__abc_44228_n3062_bF_buf36), .B(u2_remHi_428_), .Y(u2__abc_44228_n14869) );
  AND2X2 AND2X2_6568 ( .A(u2__abc_44228_n14839), .B(u2__abc_44228_n7450), .Y(u2__abc_44228_n14870) );
  AND2X2 AND2X2_6569 ( .A(u2__abc_44228_n14872), .B(u2__abc_44228_n7011), .Y(u2__abc_44228_n14873) );
  AND2X2 AND2X2_657 ( .A(u2__abc_44228_n3256), .B(u2__abc_44228_n3259), .Y(u2__abc_44228_n3260) );
  AND2X2 AND2X2_6570 ( .A(u2__abc_44228_n14875), .B(u2__abc_44228_n7547_bF_buf34), .Y(u2__abc_44228_n14876) );
  AND2X2 AND2X2_6571 ( .A(u2__abc_44228_n14876), .B(u2__abc_44228_n14874), .Y(u2__abc_44228_n14877) );
  AND2X2 AND2X2_6572 ( .A(u2__abc_44228_n7548_1_bF_buf35), .B(u2_remHi_426_), .Y(u2__abc_44228_n14878) );
  AND2X2 AND2X2_6573 ( .A(u2__abc_44228_n2983_bF_buf87), .B(u2__abc_44228_n6994), .Y(u2__abc_44228_n14881) );
  AND2X2 AND2X2_6574 ( .A(u2__abc_44228_n14882), .B(u2__abc_44228_n2972_bF_buf1), .Y(u2__abc_44228_n14883_1) );
  AND2X2 AND2X2_6575 ( .A(u2__abc_44228_n14880), .B(u2__abc_44228_n14883_1), .Y(u2__abc_44228_n14884) );
  AND2X2 AND2X2_6576 ( .A(u2__abc_44228_n14885), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_remHi_428__FF_INPUT) );
  AND2X2 AND2X2_6577 ( .A(u2__abc_44228_n3062_bF_buf35), .B(u2_remHi_429_), .Y(u2__abc_44228_n14887) );
  AND2X2 AND2X2_6578 ( .A(u2__abc_44228_n14874), .B(u2__abc_44228_n7457), .Y(u2__abc_44228_n14888) );
  AND2X2 AND2X2_6579 ( .A(u2__abc_44228_n14888), .B(u2__abc_44228_n7005), .Y(u2__abc_44228_n14889) );
  AND2X2 AND2X2_658 ( .A(u2__abc_44228_n3261), .B(u2_remHi_20_), .Y(u2__abc_44228_n3262) );
  AND2X2 AND2X2_6580 ( .A(u2__abc_44228_n14891_1), .B(u2__abc_44228_n14890), .Y(u2__abc_44228_n14892) );
  AND2X2 AND2X2_6581 ( .A(u2__abc_44228_n14893), .B(u2__abc_44228_n7547_bF_buf33), .Y(u2__abc_44228_n14894) );
  AND2X2 AND2X2_6582 ( .A(u2__abc_44228_n7548_1_bF_buf34), .B(u2_remHi_427_), .Y(u2__abc_44228_n14895) );
  AND2X2 AND2X2_6583 ( .A(u2__abc_44228_n2983_bF_buf85), .B(u2__abc_44228_n6988_1), .Y(u2__abc_44228_n14898) );
  AND2X2 AND2X2_6584 ( .A(u2__abc_44228_n14899), .B(u2__abc_44228_n2972_bF_buf0), .Y(u2__abc_44228_n14900_1) );
  AND2X2 AND2X2_6585 ( .A(u2__abc_44228_n14897), .B(u2__abc_44228_n14900_1), .Y(u2__abc_44228_n14901) );
  AND2X2 AND2X2_6586 ( .A(u2__abc_44228_n14902), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_remHi_429__FF_INPUT) );
  AND2X2 AND2X2_6587 ( .A(u2__abc_44228_n3062_bF_buf34), .B(u2_remHi_430_), .Y(u2__abc_44228_n14904) );
  AND2X2 AND2X2_6588 ( .A(u2__abc_44228_n14874), .B(u2__abc_44228_n7458), .Y(u2__abc_44228_n14905) );
  AND2X2 AND2X2_6589 ( .A(u2__abc_44228_n14907), .B(u2__abc_44228_n6997_1), .Y(u2__abc_44228_n14908_1) );
  AND2X2 AND2X2_659 ( .A(u2__abc_44228_n3263), .B(sqrto_20_), .Y(u2__abc_44228_n3264) );
  AND2X2 AND2X2_6590 ( .A(u2__abc_44228_n14910), .B(u2__abc_44228_n7547_bF_buf32), .Y(u2__abc_44228_n14911) );
  AND2X2 AND2X2_6591 ( .A(u2__abc_44228_n14911), .B(u2__abc_44228_n14909), .Y(u2__abc_44228_n14912) );
  AND2X2 AND2X2_6592 ( .A(u2__abc_44228_n7548_1_bF_buf33), .B(u2_remHi_428_), .Y(u2__abc_44228_n14913) );
  AND2X2 AND2X2_6593 ( .A(u2__abc_44228_n2983_bF_buf83), .B(u2__abc_44228_n6963), .Y(u2__abc_44228_n14916) );
  AND2X2 AND2X2_6594 ( .A(u2__abc_44228_n14917), .B(u2__abc_44228_n2972_bF_buf107), .Y(u2__abc_44228_n14918_1) );
  AND2X2 AND2X2_6595 ( .A(u2__abc_44228_n14915), .B(u2__abc_44228_n14918_1), .Y(u2__abc_44228_n14919) );
  AND2X2 AND2X2_6596 ( .A(u2__abc_44228_n14920), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_remHi_430__FF_INPUT) );
  AND2X2 AND2X2_6597 ( .A(u2__abc_44228_n3062_bF_buf33), .B(u2_remHi_431_), .Y(u2__abc_44228_n14922) );
  AND2X2 AND2X2_6598 ( .A(u2__abc_44228_n14927), .B(u2__abc_44228_n7547_bF_buf31), .Y(u2__abc_44228_n14928) );
  AND2X2 AND2X2_6599 ( .A(u2__abc_44228_n14928), .B(u2__abc_44228_n14926_1), .Y(u2__abc_44228_n14929) );
  AND2X2 AND2X2_66 ( .A(_abc_64468_n753_bF_buf4), .B(sqrto_65_), .Y(_auto_iopadmap_cc_313_execute_65414_101_) );
  AND2X2 AND2X2_660 ( .A(u2__abc_44228_n3266), .B(u2__abc_44228_n3260), .Y(u2__abc_44228_n3267) );
  AND2X2 AND2X2_6600 ( .A(u2__abc_44228_n7548_1_bF_buf32), .B(u2_remHi_429_), .Y(u2__abc_44228_n14930) );
  AND2X2 AND2X2_6601 ( .A(u2__abc_44228_n2983_bF_buf81), .B(u2__abc_44228_n6957), .Y(u2__abc_44228_n14933) );
  AND2X2 AND2X2_6602 ( .A(u2__abc_44228_n14934), .B(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n14935_1) );
  AND2X2 AND2X2_6603 ( .A(u2__abc_44228_n14932), .B(u2__abc_44228_n14935_1), .Y(u2__abc_44228_n14936) );
  AND2X2 AND2X2_6604 ( .A(u2__abc_44228_n14937), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_remHi_431__FF_INPUT) );
  AND2X2 AND2X2_6605 ( .A(u2__abc_44228_n3062_bF_buf32), .B(u2_remHi_432_), .Y(u2__abc_44228_n14939) );
  AND2X2 AND2X2_6606 ( .A(u2__abc_44228_n14666), .B(u2__abc_44228_n7103), .Y(u2__abc_44228_n14940) );
  AND2X2 AND2X2_6607 ( .A(u2__abc_44228_n14941), .B(u2__abc_44228_n6966), .Y(u2__abc_44228_n14943_1) );
  AND2X2 AND2X2_6608 ( .A(u2__abc_44228_n14944), .B(u2__abc_44228_n14942), .Y(u2__abc_44228_n14945) );
  AND2X2 AND2X2_6609 ( .A(u2__abc_44228_n14945), .B(u2__abc_44228_n7547_bF_buf30), .Y(u2__abc_44228_n14946) );
  AND2X2 AND2X2_661 ( .A(u2__abc_44228_n3268), .B(u2_remHi_18_), .Y(u2__abc_44228_n3269) );
  AND2X2 AND2X2_6610 ( .A(u2__abc_44228_n7548_1_bF_buf31), .B(u2_remHi_430_), .Y(u2__abc_44228_n14947) );
  AND2X2 AND2X2_6611 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n6977), .Y(u2__abc_44228_n14950) );
  AND2X2 AND2X2_6612 ( .A(u2__abc_44228_n14951), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n14952) );
  AND2X2 AND2X2_6613 ( .A(u2__abc_44228_n14949), .B(u2__abc_44228_n14952), .Y(u2__abc_44228_n14953) );
  AND2X2 AND2X2_6614 ( .A(u2__abc_44228_n14954_1), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_remHi_432__FF_INPUT) );
  AND2X2 AND2X2_6615 ( .A(u2__abc_44228_n3062_bF_buf31), .B(u2_remHi_433_), .Y(u2__abc_44228_n14956) );
  AND2X2 AND2X2_6616 ( .A(u2__abc_44228_n14944), .B(u2__abc_44228_n7466), .Y(u2__abc_44228_n14958) );
  AND2X2 AND2X2_6617 ( .A(u2__abc_44228_n14961), .B(u2__abc_44228_n14959), .Y(u2__abc_44228_n14962_1) );
  AND2X2 AND2X2_6618 ( .A(u2__abc_44228_n14962_1), .B(u2__abc_44228_n7547_bF_buf29), .Y(u2__abc_44228_n14963) );
  AND2X2 AND2X2_6619 ( .A(u2__abc_44228_n7548_1_bF_buf30), .B(u2_remHi_431_), .Y(u2__abc_44228_n14964) );
  AND2X2 AND2X2_662 ( .A(u2__abc_44228_n3270), .B(sqrto_18_), .Y(u2__abc_44228_n3271) );
  AND2X2 AND2X2_6620 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n6971_1), .Y(u2__abc_44228_n14967) );
  AND2X2 AND2X2_6621 ( .A(u2__abc_44228_n14968), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n14969) );
  AND2X2 AND2X2_6622 ( .A(u2__abc_44228_n14966), .B(u2__abc_44228_n14969), .Y(u2__abc_44228_n14970) );
  AND2X2 AND2X2_6623 ( .A(u2__abc_44228_n14971_1), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_remHi_433__FF_INPUT) );
  AND2X2 AND2X2_6624 ( .A(u2__abc_44228_n3062_bF_buf30), .B(u2_remHi_434_), .Y(u2__abc_44228_n14973) );
  AND2X2 AND2X2_6625 ( .A(u2__abc_44228_n14941), .B(u2__abc_44228_n6967), .Y(u2__abc_44228_n14974) );
  AND2X2 AND2X2_6626 ( .A(u2__abc_44228_n14975), .B(u2__abc_44228_n6980), .Y(u2__abc_44228_n14976) );
  AND2X2 AND2X2_6627 ( .A(u2__abc_44228_n14977), .B(u2__abc_44228_n14978), .Y(u2__abc_44228_n14979_1) );
  AND2X2 AND2X2_6628 ( .A(u2__abc_44228_n14979_1), .B(u2__abc_44228_n7547_bF_buf28), .Y(u2__abc_44228_n14980) );
  AND2X2 AND2X2_6629 ( .A(u2__abc_44228_n7548_1_bF_buf29), .B(u2_remHi_432_), .Y(u2__abc_44228_n14981) );
  AND2X2 AND2X2_663 ( .A(u2__abc_44228_n3274), .B(u2_remHi_19_), .Y(u2__abc_44228_n3275) );
  AND2X2 AND2X2_6630 ( .A(u2__abc_44228_n2983_bF_buf77), .B(u2__abc_44228_n6941), .Y(u2__abc_44228_n14984) );
  AND2X2 AND2X2_6631 ( .A(u2__abc_44228_n14985), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n14986) );
  AND2X2 AND2X2_6632 ( .A(u2__abc_44228_n14983), .B(u2__abc_44228_n14986), .Y(u2__abc_44228_n14987) );
  AND2X2 AND2X2_6633 ( .A(u2__abc_44228_n14988), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_remHi_434__FF_INPUT) );
  AND2X2 AND2X2_6634 ( .A(u2__abc_44228_n3062_bF_buf29), .B(u2_remHi_435_), .Y(u2__abc_44228_n14990) );
  AND2X2 AND2X2_6635 ( .A(u2__abc_44228_n14977), .B(u2__abc_44228_n7471), .Y(u2__abc_44228_n14992) );
  AND2X2 AND2X2_6636 ( .A(u2__abc_44228_n14995), .B(u2__abc_44228_n14993), .Y(u2__abc_44228_n14996) );
  AND2X2 AND2X2_6637 ( .A(u2__abc_44228_n14996), .B(u2__abc_44228_n7547_bF_buf27), .Y(u2__abc_44228_n14997_1) );
  AND2X2 AND2X2_6638 ( .A(u2__abc_44228_n7548_1_bF_buf28), .B(u2_remHi_433_), .Y(u2__abc_44228_n14998) );
  AND2X2 AND2X2_6639 ( .A(u2__abc_44228_n2983_bF_buf75), .B(u2__abc_44228_n6948), .Y(u2__abc_44228_n15001) );
  AND2X2 AND2X2_664 ( .A(u2__abc_44228_n3277), .B(sqrto_19_), .Y(u2__abc_44228_n3278) );
  AND2X2 AND2X2_6640 ( .A(u2__abc_44228_n15002), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n15003) );
  AND2X2 AND2X2_6641 ( .A(u2__abc_44228_n15000), .B(u2__abc_44228_n15003), .Y(u2__abc_44228_n15004) );
  AND2X2 AND2X2_6642 ( .A(u2__abc_44228_n15005), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_remHi_435__FF_INPUT) );
  AND2X2 AND2X2_6643 ( .A(u2__abc_44228_n3062_bF_buf28), .B(u2_remHi_436_), .Y(u2__abc_44228_n15007) );
  AND2X2 AND2X2_6644 ( .A(u2__abc_44228_n14977), .B(u2__abc_44228_n7472), .Y(u2__abc_44228_n15008) );
  AND2X2 AND2X2_6645 ( .A(u2__abc_44228_n15010), .B(u2__abc_44228_n6944), .Y(u2__abc_44228_n15012) );
  AND2X2 AND2X2_6646 ( .A(u2__abc_44228_n15013), .B(u2__abc_44228_n15011), .Y(u2__abc_44228_n15014_1) );
  AND2X2 AND2X2_6647 ( .A(u2__abc_44228_n15014_1), .B(u2__abc_44228_n7547_bF_buf26), .Y(u2__abc_44228_n15015) );
  AND2X2 AND2X2_6648 ( .A(u2__abc_44228_n7548_1_bF_buf27), .B(u2_remHi_434_), .Y(u2__abc_44228_n15016) );
  AND2X2 AND2X2_6649 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n6934_1), .Y(u2__abc_44228_n15019) );
  AND2X2 AND2X2_665 ( .A(u2__abc_44228_n3276), .B(u2__abc_44228_n3279), .Y(u2__abc_44228_n3280) );
  AND2X2 AND2X2_6650 ( .A(u2__abc_44228_n15020), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n15021) );
  AND2X2 AND2X2_6651 ( .A(u2__abc_44228_n15018), .B(u2__abc_44228_n15021), .Y(u2__abc_44228_n15022) );
  AND2X2 AND2X2_6652 ( .A(u2__abc_44228_n15023), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_remHi_436__FF_INPUT) );
  AND2X2 AND2X2_6653 ( .A(u2__abc_44228_n3062_bF_buf27), .B(u2_remHi_437_), .Y(u2__abc_44228_n15025) );
  AND2X2 AND2X2_6654 ( .A(u2__abc_44228_n15013), .B(u2__abc_44228_n7477), .Y(u2__abc_44228_n15026_1) );
  AND2X2 AND2X2_6655 ( .A(u2__abc_44228_n15030), .B(u2__abc_44228_n7547_bF_buf25), .Y(u2__abc_44228_n15031) );
  AND2X2 AND2X2_6656 ( .A(u2__abc_44228_n15031), .B(u2__abc_44228_n15028), .Y(u2__abc_44228_n15032) );
  AND2X2 AND2X2_6657 ( .A(u2__abc_44228_n7548_1_bF_buf26), .B(u2_remHi_435_), .Y(u2__abc_44228_n15033) );
  AND2X2 AND2X2_6658 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n6928), .Y(u2__abc_44228_n15036) );
  AND2X2 AND2X2_6659 ( .A(u2__abc_44228_n15037), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n15038) );
  AND2X2 AND2X2_666 ( .A(u2__abc_44228_n3273), .B(u2__abc_44228_n3280), .Y(u2__abc_44228_n3281) );
  AND2X2 AND2X2_6660 ( .A(u2__abc_44228_n15035), .B(u2__abc_44228_n15038), .Y(u2__abc_44228_n15039) );
  AND2X2 AND2X2_6661 ( .A(u2__abc_44228_n15040), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_remHi_437__FF_INPUT) );
  AND2X2 AND2X2_6662 ( .A(u2__abc_44228_n3062_bF_buf26), .B(u2_remHi_438_), .Y(u2__abc_44228_n15042) );
  AND2X2 AND2X2_6663 ( .A(u2__abc_44228_n15013), .B(u2__abc_44228_n7478), .Y(u2__abc_44228_n15043_1) );
  AND2X2 AND2X2_6664 ( .A(u2__abc_44228_n15045), .B(u2__abc_44228_n6937), .Y(u2__abc_44228_n15046) );
  AND2X2 AND2X2_6665 ( .A(u2__abc_44228_n15048), .B(u2__abc_44228_n7547_bF_buf24), .Y(u2__abc_44228_n15049) );
  AND2X2 AND2X2_6666 ( .A(u2__abc_44228_n15049), .B(u2__abc_44228_n15047), .Y(u2__abc_44228_n15050) );
  AND2X2 AND2X2_6667 ( .A(u2__abc_44228_n7548_1_bF_buf25), .B(u2_remHi_436_), .Y(u2__abc_44228_n15051_1) );
  AND2X2 AND2X2_6668 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n6918), .Y(u2__abc_44228_n15054) );
  AND2X2 AND2X2_6669 ( .A(u2__abc_44228_n15055), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n15056) );
  AND2X2 AND2X2_667 ( .A(u2__abc_44228_n3267), .B(u2__abc_44228_n3281), .Y(u2__abc_44228_n3282) );
  AND2X2 AND2X2_6670 ( .A(u2__abc_44228_n15053), .B(u2__abc_44228_n15056), .Y(u2__abc_44228_n15057) );
  AND2X2 AND2X2_6671 ( .A(u2__abc_44228_n15058), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_remHi_438__FF_INPUT) );
  AND2X2 AND2X2_6672 ( .A(u2__abc_44228_n3062_bF_buf25), .B(u2_remHi_439_), .Y(u2__abc_44228_n15060) );
  AND2X2 AND2X2_6673 ( .A(u2__abc_44228_n15065), .B(u2__abc_44228_n7547_bF_buf23), .Y(u2__abc_44228_n15066) );
  AND2X2 AND2X2_6674 ( .A(u2__abc_44228_n15066), .B(u2__abc_44228_n15064), .Y(u2__abc_44228_n15067) );
  AND2X2 AND2X2_6675 ( .A(u2__abc_44228_n7548_1_bF_buf24), .B(u2_remHi_437_), .Y(u2__abc_44228_n15068) );
  AND2X2 AND2X2_6676 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n6912), .Y(u2__abc_44228_n15071) );
  AND2X2 AND2X2_6677 ( .A(u2__abc_44228_n15072), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n15073) );
  AND2X2 AND2X2_6678 ( .A(u2__abc_44228_n15070), .B(u2__abc_44228_n15073), .Y(u2__abc_44228_n15074) );
  AND2X2 AND2X2_6679 ( .A(u2__abc_44228_n15075), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_remHi_439__FF_INPUT) );
  AND2X2 AND2X2_668 ( .A(u2__abc_44228_n3284), .B(u2__abc_44228_n3286), .Y(u2__abc_44228_n3287) );
  AND2X2 AND2X2_6680 ( .A(u2__abc_44228_n3062_bF_buf24), .B(u2_remHi_440_), .Y(u2__abc_44228_n15077) );
  AND2X2 AND2X2_6681 ( .A(u2__abc_44228_n14941), .B(u2__abc_44228_n6983), .Y(u2__abc_44228_n15078_1) );
  AND2X2 AND2X2_6682 ( .A(u2__abc_44228_n15079), .B(u2__abc_44228_n6921), .Y(u2__abc_44228_n15080) );
  AND2X2 AND2X2_6683 ( .A(u2__abc_44228_n15081), .B(u2__abc_44228_n15082), .Y(u2__abc_44228_n15083) );
  AND2X2 AND2X2_6684 ( .A(u2__abc_44228_n15083), .B(u2__abc_44228_n7547_bF_buf22), .Y(u2__abc_44228_n15084) );
  AND2X2 AND2X2_6685 ( .A(u2__abc_44228_n7548_1_bF_buf23), .B(u2_remHi_438_), .Y(u2__abc_44228_n15085) );
  AND2X2 AND2X2_6686 ( .A(u2__abc_44228_n2983_bF_buf67), .B(u2__abc_44228_n6904), .Y(u2__abc_44228_n15088) );
  AND2X2 AND2X2_6687 ( .A(u2__abc_44228_n15089), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n15090) );
  AND2X2 AND2X2_6688 ( .A(u2__abc_44228_n15087), .B(u2__abc_44228_n15090), .Y(u2__abc_44228_n15091) );
  AND2X2 AND2X2_6689 ( .A(u2__abc_44228_n15092), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_remHi_440__FF_INPUT) );
  AND2X2 AND2X2_669 ( .A(u2__abc_44228_n3289), .B(u2__abc_44228_n3291), .Y(u2__abc_44228_n3292) );
  AND2X2 AND2X2_6690 ( .A(u2__abc_44228_n3062_bF_buf23), .B(u2_remHi_441_), .Y(u2__abc_44228_n15094) );
  AND2X2 AND2X2_6691 ( .A(u2__abc_44228_n15081), .B(u2__abc_44228_n7489), .Y(u2__abc_44228_n15095) );
  AND2X2 AND2X2_6692 ( .A(u2__abc_44228_n15095), .B(u2__abc_44228_n6915_1), .Y(u2__abc_44228_n15096) );
  AND2X2 AND2X2_6693 ( .A(u2__abc_44228_n15098), .B(u2__abc_44228_n15097_1), .Y(u2__abc_44228_n15099) );
  AND2X2 AND2X2_6694 ( .A(u2__abc_44228_n15100), .B(u2__abc_44228_n7547_bF_buf21), .Y(u2__abc_44228_n15101) );
  AND2X2 AND2X2_6695 ( .A(u2__abc_44228_n7548_1_bF_buf22), .B(u2_remHi_439_), .Y(u2__abc_44228_n15102) );
  AND2X2 AND2X2_6696 ( .A(u2__abc_44228_n2983_bF_buf65), .B(u2__abc_44228_n6898), .Y(u2__abc_44228_n15105_1) );
  AND2X2 AND2X2_6697 ( .A(u2__abc_44228_n15106), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n15107) );
  AND2X2 AND2X2_6698 ( .A(u2__abc_44228_n15104), .B(u2__abc_44228_n15107), .Y(u2__abc_44228_n15108) );
  AND2X2 AND2X2_6699 ( .A(u2__abc_44228_n15109), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_remHi_441__FF_INPUT) );
  AND2X2 AND2X2_67 ( .A(_abc_64468_n753_bF_buf3), .B(sqrto_66_), .Y(_auto_iopadmap_cc_313_execute_65414_102_) );
  AND2X2 AND2X2_670 ( .A(u2__abc_44228_n3287), .B(u2__abc_44228_n3292), .Y(u2__abc_44228_n3293) );
  AND2X2 AND2X2_6700 ( .A(u2__abc_44228_n3062_bF_buf22), .B(u2_remHi_442_), .Y(u2__abc_44228_n15111) );
  AND2X2 AND2X2_6701 ( .A(u2__abc_44228_n15081), .B(u2__abc_44228_n7490), .Y(u2__abc_44228_n15112) );
  AND2X2 AND2X2_6702 ( .A(u2__abc_44228_n15114_1), .B(u2__abc_44228_n6907), .Y(u2__abc_44228_n15115) );
  AND2X2 AND2X2_6703 ( .A(u2__abc_44228_n15116), .B(u2__abc_44228_n15117), .Y(u2__abc_44228_n15118) );
  AND2X2 AND2X2_6704 ( .A(u2__abc_44228_n15118), .B(u2__abc_44228_n7547_bF_buf20), .Y(u2__abc_44228_n15119) );
  AND2X2 AND2X2_6705 ( .A(u2__abc_44228_n7548_1_bF_buf21), .B(u2_remHi_440_), .Y(u2__abc_44228_n15120) );
  AND2X2 AND2X2_6706 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n6889), .Y(u2__abc_44228_n15123) );
  AND2X2 AND2X2_6707 ( .A(u2__abc_44228_n15124), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n15125) );
  AND2X2 AND2X2_6708 ( .A(u2__abc_44228_n15122_1), .B(u2__abc_44228_n15125), .Y(u2__abc_44228_n15126) );
  AND2X2 AND2X2_6709 ( .A(u2__abc_44228_n15127), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_remHi_442__FF_INPUT) );
  AND2X2 AND2X2_671 ( .A(u2__abc_44228_n3294), .B(u2_remHi_15_), .Y(u2__abc_44228_n3295) );
  AND2X2 AND2X2_6710 ( .A(u2__abc_44228_n3062_bF_buf21), .B(u2_remHi_443_), .Y(u2__abc_44228_n15129) );
  AND2X2 AND2X2_6711 ( .A(u2__abc_44228_n15134), .B(u2__abc_44228_n7547_bF_buf19), .Y(u2__abc_44228_n15135) );
  AND2X2 AND2X2_6712 ( .A(u2__abc_44228_n15135), .B(u2__abc_44228_n15133), .Y(u2__abc_44228_n15136) );
  AND2X2 AND2X2_6713 ( .A(u2__abc_44228_n7548_1_bF_buf20), .B(u2_remHi_441_), .Y(u2__abc_44228_n15137) );
  AND2X2 AND2X2_6714 ( .A(u2__abc_44228_n2983_bF_buf62), .B(u2__abc_44228_n6883), .Y(u2__abc_44228_n15140_1) );
  AND2X2 AND2X2_6715 ( .A(u2__abc_44228_n15141), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n15142) );
  AND2X2 AND2X2_6716 ( .A(u2__abc_44228_n15139), .B(u2__abc_44228_n15142), .Y(u2__abc_44228_n15143) );
  AND2X2 AND2X2_6717 ( .A(u2__abc_44228_n15144), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_remHi_443__FF_INPUT) );
  AND2X2 AND2X2_6718 ( .A(u2__abc_44228_n3062_bF_buf20), .B(u2_remHi_444_), .Y(u2__abc_44228_n15146) );
  AND2X2 AND2X2_6719 ( .A(u2__abc_44228_n15079), .B(u2__abc_44228_n6923), .Y(u2__abc_44228_n15147) );
  AND2X2 AND2X2_672 ( .A(u2__abc_44228_n3297), .B(sqrto_15_), .Y(u2__abc_44228_n3298) );
  AND2X2 AND2X2_6720 ( .A(u2__abc_44228_n15148), .B(u2__abc_44228_n6892), .Y(u2__abc_44228_n15150) );
  AND2X2 AND2X2_6721 ( .A(u2__abc_44228_n15151), .B(u2__abc_44228_n15149_1), .Y(u2__abc_44228_n15152) );
  AND2X2 AND2X2_6722 ( .A(u2__abc_44228_n15152), .B(u2__abc_44228_n7547_bF_buf18), .Y(u2__abc_44228_n15153) );
  AND2X2 AND2X2_6723 ( .A(u2__abc_44228_n7548_1_bF_buf19), .B(u2_remHi_442_), .Y(u2__abc_44228_n15154) );
  AND2X2 AND2X2_6724 ( .A(u2__abc_44228_n2983_bF_buf61), .B(u2__abc_44228_n6875), .Y(u2__abc_44228_n15157_1) );
  AND2X2 AND2X2_6725 ( .A(u2__abc_44228_n15158), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n15159) );
  AND2X2 AND2X2_6726 ( .A(u2__abc_44228_n15156), .B(u2__abc_44228_n15159), .Y(u2__abc_44228_n15160) );
  AND2X2 AND2X2_6727 ( .A(u2__abc_44228_n15161), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_remHi_444__FF_INPUT) );
  AND2X2 AND2X2_6728 ( .A(u2__abc_44228_n3062_bF_buf19), .B(u2_remHi_445_), .Y(u2__abc_44228_n15163) );
  AND2X2 AND2X2_6729 ( .A(u2__abc_44228_n15151), .B(u2__abc_44228_n7496), .Y(u2__abc_44228_n15165) );
  AND2X2 AND2X2_673 ( .A(u2__abc_44228_n3296), .B(u2__abc_44228_n3299), .Y(u2__abc_44228_n3300) );
  AND2X2 AND2X2_6730 ( .A(u2__abc_44228_n15168), .B(u2__abc_44228_n15166), .Y(u2__abc_44228_n15169) );
  AND2X2 AND2X2_6731 ( .A(u2__abc_44228_n15169), .B(u2__abc_44228_n7547_bF_buf17), .Y(u2__abc_44228_n15170_1) );
  AND2X2 AND2X2_6732 ( .A(u2__abc_44228_n7548_1_bF_buf18), .B(u2_remHi_443_), .Y(u2__abc_44228_n15171) );
  AND2X2 AND2X2_6733 ( .A(u2__abc_44228_n2983_bF_buf59), .B(u2__abc_44228_n6869_1), .Y(u2__abc_44228_n15174) );
  AND2X2 AND2X2_6734 ( .A(u2__abc_44228_n15175), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n15176) );
  AND2X2 AND2X2_6735 ( .A(u2__abc_44228_n15173), .B(u2__abc_44228_n15176), .Y(u2__abc_44228_n15177) );
  AND2X2 AND2X2_6736 ( .A(u2__abc_44228_n15178_1), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_remHi_445__FF_INPUT) );
  AND2X2 AND2X2_6737 ( .A(u2__abc_44228_n3062_bF_buf18), .B(u2_remHi_446_), .Y(u2__abc_44228_n15180) );
  AND2X2 AND2X2_6738 ( .A(u2__abc_44228_n15148), .B(u2__abc_44228_n6893), .Y(u2__abc_44228_n15181) );
  AND2X2 AND2X2_6739 ( .A(u2__abc_44228_n15182), .B(u2__abc_44228_n6878_1), .Y(u2__abc_44228_n15183) );
  AND2X2 AND2X2_674 ( .A(u2__abc_44228_n3301), .B(u2_remHi_14_), .Y(u2__abc_44228_n3302) );
  AND2X2 AND2X2_6740 ( .A(u2__abc_44228_n15185), .B(u2__abc_44228_n7547_bF_buf16), .Y(u2__abc_44228_n15186) );
  AND2X2 AND2X2_6741 ( .A(u2__abc_44228_n15186), .B(u2__abc_44228_n15184), .Y(u2__abc_44228_n15187_1) );
  AND2X2 AND2X2_6742 ( .A(u2__abc_44228_n7548_1_bF_buf17), .B(u2_remHi_444_), .Y(u2__abc_44228_n15188) );
  AND2X2 AND2X2_6743 ( .A(u2__abc_44228_n2983_bF_buf57), .B(u2__abc_44228_n7525), .Y(u2__abc_44228_n15191) );
  AND2X2 AND2X2_6744 ( .A(u2__abc_44228_n15192), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n15193) );
  AND2X2 AND2X2_6745 ( .A(u2__abc_44228_n15190), .B(u2__abc_44228_n15193), .Y(u2__abc_44228_n15194) );
  AND2X2 AND2X2_6746 ( .A(u2__abc_44228_n15195_1), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_remHi_446__FF_INPUT) );
  AND2X2 AND2X2_6747 ( .A(u2__abc_44228_n3062_bF_buf17), .B(u2_remHi_447_), .Y(u2__abc_44228_n15197) );
  AND2X2 AND2X2_6748 ( .A(u2__abc_44228_n15202), .B(u2__abc_44228_n7547_bF_buf15), .Y(u2__abc_44228_n15203) );
  AND2X2 AND2X2_6749 ( .A(u2__abc_44228_n15203), .B(u2__abc_44228_n15201), .Y(u2__abc_44228_n15204) );
  AND2X2 AND2X2_675 ( .A(u2__abc_44228_n3303), .B(sqrto_14_), .Y(u2__abc_44228_n3304) );
  AND2X2 AND2X2_6750 ( .A(u2__abc_44228_n7548_1_bF_buf16), .B(u2_remHi_445_), .Y(u2__abc_44228_n15205_1) );
  AND2X2 AND2X2_6751 ( .A(u2__abc_44228_n2983_bF_buf55), .B(u2__abc_44228_n7532), .Y(u2__abc_44228_n15208) );
  AND2X2 AND2X2_6752 ( .A(u2__abc_44228_n15209), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n15210) );
  AND2X2 AND2X2_6753 ( .A(u2__abc_44228_n15207), .B(u2__abc_44228_n15210), .Y(u2__abc_44228_n15211) );
  AND2X2 AND2X2_6754 ( .A(u2__abc_44228_n15212), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_remHi_447__FF_INPUT) );
  AND2X2 AND2X2_6755 ( .A(u2__abc_44228_n3062_bF_buf16), .B(u2_remHi_448_), .Y(u2__abc_44228_n15214) );
  AND2X2 AND2X2_6756 ( .A(u2__abc_44228_n7508), .B(u2__abc_44228_n7528), .Y(u2__abc_44228_n15216) );
  AND2X2 AND2X2_6757 ( .A(u2__abc_44228_n15217), .B(u2__abc_44228_n15215), .Y(u2__abc_44228_n15218) );
  AND2X2 AND2X2_6758 ( .A(u2__abc_44228_n15219), .B(u2__abc_44228_n15220), .Y(u2__abc_44228_n15221) );
  AND2X2 AND2X2_6759 ( .A(u2__abc_44228_n2983_bF_buf53), .B(u2__abc_44228_n7518), .Y(u2__abc_44228_n15223) );
  AND2X2 AND2X2_676 ( .A(u2__abc_44228_n3306), .B(u2__abc_44228_n3300), .Y(u2__abc_44228_n3307) );
  AND2X2 AND2X2_6760 ( .A(u2__abc_44228_n15224), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n15225) );
  AND2X2 AND2X2_6761 ( .A(u2__abc_44228_n15222_1), .B(u2__abc_44228_n15225), .Y(u2__abc_44228_n15226) );
  AND2X2 AND2X2_6762 ( .A(u2__abc_44228_n15227), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_remHi_448__FF_INPUT) );
  AND2X2 AND2X2_6763 ( .A(u2__abc_44228_n3062_bF_buf15), .B(u2_remHi_449_), .Y(u2__abc_44228_n15229) );
  AND2X2 AND2X2_6764 ( .A(u2__abc_44228_n15217), .B(u2__abc_44228_n7539), .Y(u2__abc_44228_n15231) );
  AND2X2 AND2X2_6765 ( .A(u2__abc_44228_n15234), .B(u2__abc_44228_n15232), .Y(u2__abc_44228_n15235) );
  AND2X2 AND2X2_6766 ( .A(u2__abc_44228_n15235), .B(u2__abc_44228_n7547_bF_buf13), .Y(u2__abc_44228_n15236) );
  AND2X2 AND2X2_6767 ( .A(u2__abc_44228_n7548_1_bF_buf14), .B(u2_remHi_447_), .Y(u2__abc_44228_n15237) );
  AND2X2 AND2X2_6768 ( .A(u2__abc_44228_n2983_bF_buf51), .B(u2__abc_44228_n7512), .Y(u2__abc_44228_n15240) );
  AND2X2 AND2X2_6769 ( .A(u2__abc_44228_n15241_1), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n15242) );
  AND2X2 AND2X2_677 ( .A(u2__abc_44228_n3307), .B(u2__abc_44228_n3293), .Y(u2__abc_44228_n3308) );
  AND2X2 AND2X2_6770 ( .A(u2__abc_44228_n15239), .B(u2__abc_44228_n15242), .Y(u2__abc_44228_n15243) );
  AND2X2 AND2X2_6771 ( .A(u2__abc_44228_n15244), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_remHi_449__FF_INPUT) );
  AND2X2 AND2X2_6772 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2_state_2_), .Y(u2__abc_44228_n15246) );
  AND2X2 AND2X2_6773 ( .A(u2__abc_44228_n2966_bF_buf86), .B(u2_remLo_0_), .Y(u2__abc_44228_n15248) );
  AND2X2 AND2X2_6774 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2__abc_44228_n15248), .Y(u2_remLo_0__FF_INPUT) );
  AND2X2 AND2X2_6775 ( .A(u2__abc_44228_n2966_bF_buf85), .B(u2_remLo_1_), .Y(u2__abc_44228_n15250) );
  AND2X2 AND2X2_6776 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2__abc_44228_n15250), .Y(u2_remLo_1__FF_INPUT) );
  AND2X2 AND2X2_6777 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_2_), .Y(u2__abc_44228_n15252) );
  AND2X2 AND2X2_6778 ( .A(u2__abc_44228_n2972_bF_buf87), .B(u2_remLo_0_), .Y(u2__abc_44228_n15253) );
  AND2X2 AND2X2_6779 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n15253), .Y(u2__abc_44228_n15254) );
  AND2X2 AND2X2_678 ( .A(u2__abc_44228_n3282), .B(u2__abc_44228_n3308), .Y(u2__abc_44228_n3309) );
  AND2X2 AND2X2_6780 ( .A(u2__abc_44228_n15255), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_remLo_2__FF_INPUT) );
  AND2X2 AND2X2_6781 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_3_), .Y(u2__abc_44228_n15257) );
  AND2X2 AND2X2_6782 ( .A(u2__abc_44228_n2972_bF_buf86), .B(u2_remLo_1_), .Y(u2__abc_44228_n15258_1) );
  AND2X2 AND2X2_6783 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n15258_1), .Y(u2__abc_44228_n15259) );
  AND2X2 AND2X2_6784 ( .A(u2__abc_44228_n15260), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_remLo_3__FF_INPUT) );
  AND2X2 AND2X2_6785 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_4_), .Y(u2__abc_44228_n15262) );
  AND2X2 AND2X2_6786 ( .A(u2__abc_44228_n2972_bF_buf85), .B(u2_remLo_2_), .Y(u2__abc_44228_n15263) );
  AND2X2 AND2X2_6787 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n15263), .Y(u2__abc_44228_n15264) );
  AND2X2 AND2X2_6788 ( .A(u2__abc_44228_n15265), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_remLo_4__FF_INPUT) );
  AND2X2 AND2X2_6789 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_5_), .Y(u2__abc_44228_n15267) );
  AND2X2 AND2X2_679 ( .A(u2__abc_44228_n3253), .B(u2__abc_44228_n3309), .Y(u2__abc_44228_n3310) );
  AND2X2 AND2X2_6790 ( .A(u2__abc_44228_n2972_bF_buf84), .B(u2_remLo_3_), .Y(u2__abc_44228_n15268) );
  AND2X2 AND2X2_6791 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n15268), .Y(u2__abc_44228_n15269) );
  AND2X2 AND2X2_6792 ( .A(u2__abc_44228_n15270), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_remLo_5__FF_INPUT) );
  AND2X2 AND2X2_6793 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_6_), .Y(u2__abc_44228_n15272) );
  AND2X2 AND2X2_6794 ( .A(u2__abc_44228_n2972_bF_buf83), .B(u2_remLo_4_), .Y(u2__abc_44228_n15273) );
  AND2X2 AND2X2_6795 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n15273), .Y(u2__abc_44228_n15274) );
  AND2X2 AND2X2_6796 ( .A(u2__abc_44228_n15275), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_remLo_6__FF_INPUT) );
  AND2X2 AND2X2_6797 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_7_), .Y(u2__abc_44228_n15277) );
  AND2X2 AND2X2_6798 ( .A(u2__abc_44228_n2972_bF_buf82), .B(u2_remLo_5_), .Y(u2__abc_44228_n15278) );
  AND2X2 AND2X2_6799 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n15278), .Y(u2__abc_44228_n15279) );
  AND2X2 AND2X2_68 ( .A(_abc_64468_n753_bF_buf2), .B(sqrto_67_), .Y(_auto_iopadmap_cc_313_execute_65414_103_) );
  AND2X2 AND2X2_680 ( .A(u2__abc_44228_n3194), .B(u2__abc_44228_n3310), .Y(u2__abc_44228_n3311) );
  AND2X2 AND2X2_6800 ( .A(u2__abc_44228_n15280), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_remLo_7__FF_INPUT) );
  AND2X2 AND2X2_6801 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_8_), .Y(u2__abc_44228_n15282) );
  AND2X2 AND2X2_6802 ( .A(u2__abc_44228_n2972_bF_buf81), .B(u2_remLo_6_), .Y(u2__abc_44228_n15283) );
  AND2X2 AND2X2_6803 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n15283), .Y(u2__abc_44228_n15284_1) );
  AND2X2 AND2X2_6804 ( .A(u2__abc_44228_n15285), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_remLo_8__FF_INPUT) );
  AND2X2 AND2X2_6805 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_9_), .Y(u2__abc_44228_n15287) );
  AND2X2 AND2X2_6806 ( .A(u2__abc_44228_n2972_bF_buf80), .B(u2_remLo_7_), .Y(u2__abc_44228_n15288) );
  AND2X2 AND2X2_6807 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n15288), .Y(u2__abc_44228_n15289) );
  AND2X2 AND2X2_6808 ( .A(u2__abc_44228_n15290), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_remLo_9__FF_INPUT) );
  AND2X2 AND2X2_6809 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_10_), .Y(u2__abc_44228_n15292) );
  AND2X2 AND2X2_681 ( .A(u2__abc_44228_n3312), .B(u2__abc_44228_n3299), .Y(u2__abc_44228_n3313) );
  AND2X2 AND2X2_6810 ( .A(u2__abc_44228_n2972_bF_buf79), .B(u2_remLo_8_), .Y(u2__abc_44228_n15293_1) );
  AND2X2 AND2X2_6811 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n15293_1), .Y(u2__abc_44228_n15294) );
  AND2X2 AND2X2_6812 ( .A(u2__abc_44228_n15295), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_remLo_10__FF_INPUT) );
  AND2X2 AND2X2_6813 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_11_), .Y(u2__abc_44228_n15297) );
  AND2X2 AND2X2_6814 ( .A(u2__abc_44228_n2972_bF_buf78), .B(u2_remLo_9_), .Y(u2__abc_44228_n15298) );
  AND2X2 AND2X2_6815 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n15298), .Y(u2__abc_44228_n15299) );
  AND2X2 AND2X2_6816 ( .A(u2__abc_44228_n15300), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_remLo_11__FF_INPUT) );
  AND2X2 AND2X2_6817 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_12_), .Y(u2__abc_44228_n15302) );
  AND2X2 AND2X2_6818 ( .A(u2__abc_44228_n2972_bF_buf77), .B(u2_remLo_10_), .Y(u2__abc_44228_n15303) );
  AND2X2 AND2X2_6819 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n15303), .Y(u2__abc_44228_n15304) );
  AND2X2 AND2X2_682 ( .A(u2__abc_44228_n3313), .B(u2__abc_44228_n3293), .Y(u2__abc_44228_n3314) );
  AND2X2 AND2X2_6820 ( .A(u2__abc_44228_n15305), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_remLo_12__FF_INPUT) );
  AND2X2 AND2X2_6821 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_13_), .Y(u2__abc_44228_n15307) );
  AND2X2 AND2X2_6822 ( .A(u2__abc_44228_n2972_bF_buf76), .B(u2_remLo_11_), .Y(u2__abc_44228_n15308) );
  AND2X2 AND2X2_6823 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n15308), .Y(u2__abc_44228_n15309) );
  AND2X2 AND2X2_6824 ( .A(u2__abc_44228_n15310), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_remLo_13__FF_INPUT) );
  AND2X2 AND2X2_6825 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_14_), .Y(u2__abc_44228_n15312) );
  AND2X2 AND2X2_6826 ( .A(u2__abc_44228_n2972_bF_buf75), .B(u2_remLo_12_), .Y(u2__abc_44228_n15313_1) );
  AND2X2 AND2X2_6827 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n15313_1), .Y(u2__abc_44228_n15314) );
  AND2X2 AND2X2_6828 ( .A(u2__abc_44228_n15315), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_remLo_14__FF_INPUT) );
  AND2X2 AND2X2_6829 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_15_), .Y(u2__abc_44228_n15317) );
  AND2X2 AND2X2_683 ( .A(u2__abc_44228_n3316), .B(u2__abc_44228_n3286), .Y(u2__abc_44228_n3317) );
  AND2X2 AND2X2_6830 ( .A(u2__abc_44228_n2972_bF_buf74), .B(u2_remLo_13_), .Y(u2__abc_44228_n15318) );
  AND2X2 AND2X2_6831 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n15318), .Y(u2__abc_44228_n15319) );
  AND2X2 AND2X2_6832 ( .A(u2__abc_44228_n15320), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_remLo_15__FF_INPUT) );
  AND2X2 AND2X2_6833 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_16_), .Y(u2__abc_44228_n15322) );
  AND2X2 AND2X2_6834 ( .A(u2__abc_44228_n2972_bF_buf73), .B(u2_remLo_14_), .Y(u2__abc_44228_n15323) );
  AND2X2 AND2X2_6835 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n15323), .Y(u2__abc_44228_n15324) );
  AND2X2 AND2X2_6836 ( .A(u2__abc_44228_n15325), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_remLo_16__FF_INPUT) );
  AND2X2 AND2X2_6837 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_17_), .Y(u2__abc_44228_n15327) );
  AND2X2 AND2X2_6838 ( .A(u2__abc_44228_n2972_bF_buf72), .B(u2_remLo_15_), .Y(u2__abc_44228_n15328) );
  AND2X2 AND2X2_6839 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n15328), .Y(u2__abc_44228_n15329) );
  AND2X2 AND2X2_684 ( .A(u2__abc_44228_n3319), .B(u2__abc_44228_n3282), .Y(u2__abc_44228_n3320) );
  AND2X2 AND2X2_6840 ( .A(u2__abc_44228_n15330_1), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_remLo_17__FF_INPUT) );
  AND2X2 AND2X2_6841 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_18_), .Y(u2__abc_44228_n15332) );
  AND2X2 AND2X2_6842 ( .A(u2__abc_44228_n2972_bF_buf71), .B(u2_remLo_16_), .Y(u2__abc_44228_n15333) );
  AND2X2 AND2X2_6843 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n15333), .Y(u2__abc_44228_n15334) );
  AND2X2 AND2X2_6844 ( .A(u2__abc_44228_n15335), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_remLo_18__FF_INPUT) );
  AND2X2 AND2X2_6845 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_19_), .Y(u2__abc_44228_n15337) );
  AND2X2 AND2X2_6846 ( .A(u2__abc_44228_n2972_bF_buf70), .B(u2_remLo_17_), .Y(u2__abc_44228_n15338_1) );
  AND2X2 AND2X2_6847 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n15338_1), .Y(u2__abc_44228_n15339) );
  AND2X2 AND2X2_6848 ( .A(u2__abc_44228_n15340), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_remLo_19__FF_INPUT) );
  AND2X2 AND2X2_6849 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_20_), .Y(u2__abc_44228_n15342) );
  AND2X2 AND2X2_685 ( .A(u2__abc_44228_n3321), .B(u2__abc_44228_n3279), .Y(u2__abc_44228_n3322) );
  AND2X2 AND2X2_6850 ( .A(u2__abc_44228_n2972_bF_buf69), .B(u2_remLo_18_), .Y(u2__abc_44228_n15343) );
  AND2X2 AND2X2_6851 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n15343), .Y(u2__abc_44228_n15344) );
  AND2X2 AND2X2_6852 ( .A(u2__abc_44228_n15345), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_remLo_20__FF_INPUT) );
  AND2X2 AND2X2_6853 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_21_), .Y(u2__abc_44228_n15347) );
  AND2X2 AND2X2_6854 ( .A(u2__abc_44228_n2972_bF_buf68), .B(u2_remLo_19_), .Y(u2__abc_44228_n15348_1) );
  AND2X2 AND2X2_6855 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n15348_1), .Y(u2__abc_44228_n15349) );
  AND2X2 AND2X2_6856 ( .A(u2__abc_44228_n15350), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_remLo_21__FF_INPUT) );
  AND2X2 AND2X2_6857 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_22_), .Y(u2__abc_44228_n15352) );
  AND2X2 AND2X2_6858 ( .A(u2__abc_44228_n2972_bF_buf67), .B(u2_remLo_20_), .Y(u2__abc_44228_n15353) );
  AND2X2 AND2X2_6859 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n15353), .Y(u2__abc_44228_n15354) );
  AND2X2 AND2X2_686 ( .A(u2__abc_44228_n3267), .B(u2__abc_44228_n3322), .Y(u2__abc_44228_n3323) );
  AND2X2 AND2X2_6860 ( .A(u2__abc_44228_n15355), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_remLo_22__FF_INPUT) );
  AND2X2 AND2X2_6861 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_23_), .Y(u2__abc_44228_n15357) );
  AND2X2 AND2X2_6862 ( .A(u2__abc_44228_n2972_bF_buf66), .B(u2_remLo_21_), .Y(u2__abc_44228_n15358) );
  AND2X2 AND2X2_6863 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n15358), .Y(u2__abc_44228_n15359) );
  AND2X2 AND2X2_6864 ( .A(u2__abc_44228_n15360), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_remLo_23__FF_INPUT) );
  AND2X2 AND2X2_6865 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_24_), .Y(u2__abc_44228_n15362) );
  AND2X2 AND2X2_6866 ( .A(u2__abc_44228_n2972_bF_buf65), .B(u2_remLo_22_), .Y(u2__abc_44228_n15363) );
  AND2X2 AND2X2_6867 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n15363), .Y(u2__abc_44228_n15364) );
  AND2X2 AND2X2_6868 ( .A(u2__abc_44228_n15365_1), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_remLo_24__FF_INPUT) );
  AND2X2 AND2X2_6869 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_25_), .Y(u2__abc_44228_n15367) );
  AND2X2 AND2X2_687 ( .A(u2__abc_44228_n3259), .B(u2__abc_44228_n3262), .Y(u2__abc_44228_n3324) );
  AND2X2 AND2X2_6870 ( .A(u2__abc_44228_n2972_bF_buf64), .B(u2_remLo_23_), .Y(u2__abc_44228_n15368) );
  AND2X2 AND2X2_6871 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n15368), .Y(u2__abc_44228_n15369) );
  AND2X2 AND2X2_6872 ( .A(u2__abc_44228_n15370), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_remLo_25__FF_INPUT) );
  AND2X2 AND2X2_6873 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_26_), .Y(u2__abc_44228_n15372) );
  AND2X2 AND2X2_6874 ( .A(u2__abc_44228_n2972_bF_buf63), .B(u2_remLo_24_), .Y(u2__abc_44228_n15373_1) );
  AND2X2 AND2X2_6875 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n15373_1), .Y(u2__abc_44228_n15374) );
  AND2X2 AND2X2_6876 ( .A(u2__abc_44228_n15375), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_remLo_26__FF_INPUT) );
  AND2X2 AND2X2_6877 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_27_), .Y(u2__abc_44228_n15377) );
  AND2X2 AND2X2_6878 ( .A(u2__abc_44228_n2972_bF_buf62), .B(u2_remLo_25_), .Y(u2__abc_44228_n15378) );
  AND2X2 AND2X2_6879 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n15378), .Y(u2__abc_44228_n15379) );
  AND2X2 AND2X2_688 ( .A(u2__abc_44228_n3327), .B(u2__abc_44228_n3253), .Y(u2__abc_44228_n3328) );
  AND2X2 AND2X2_6880 ( .A(u2__abc_44228_n15380), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_remLo_27__FF_INPUT) );
  AND2X2 AND2X2_6881 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_28_), .Y(u2__abc_44228_n15382) );
  AND2X2 AND2X2_6882 ( .A(u2__abc_44228_n2972_bF_buf61), .B(u2_remLo_26_), .Y(u2__abc_44228_n15383) );
  AND2X2 AND2X2_6883 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n15383), .Y(u2__abc_44228_n15384_1) );
  AND2X2 AND2X2_6884 ( .A(u2__abc_44228_n15385), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_remLo_28__FF_INPUT) );
  AND2X2 AND2X2_6885 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_29_), .Y(u2__abc_44228_n15387) );
  AND2X2 AND2X2_6886 ( .A(u2__abc_44228_n2972_bF_buf60), .B(u2_remLo_27_), .Y(u2__abc_44228_n15388) );
  AND2X2 AND2X2_6887 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n15388), .Y(u2__abc_44228_n15389) );
  AND2X2 AND2X2_6888 ( .A(u2__abc_44228_n15390), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_remLo_29__FF_INPUT) );
  AND2X2 AND2X2_6889 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_30_), .Y(u2__abc_44228_n15392_1) );
  AND2X2 AND2X2_689 ( .A(u2__abc_44228_n3329), .B(u2__abc_44228_n3229), .Y(u2__abc_44228_n3330) );
  AND2X2 AND2X2_6890 ( .A(u2__abc_44228_n2972_bF_buf59), .B(u2_remLo_28_), .Y(u2__abc_44228_n15393) );
  AND2X2 AND2X2_6891 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n15393), .Y(u2__abc_44228_n15394) );
  AND2X2 AND2X2_6892 ( .A(u2__abc_44228_n15395), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_remLo_30__FF_INPUT) );
  AND2X2 AND2X2_6893 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_31_), .Y(u2__abc_44228_n15397) );
  AND2X2 AND2X2_6894 ( .A(u2__abc_44228_n2972_bF_buf58), .B(u2_remLo_29_), .Y(u2__abc_44228_n15398) );
  AND2X2 AND2X2_6895 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n15398), .Y(u2__abc_44228_n15399) );
  AND2X2 AND2X2_6896 ( .A(u2__abc_44228_n15400), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_remLo_31__FF_INPUT) );
  AND2X2 AND2X2_6897 ( .A(u2__abc_44228_n3061), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2__abc_44228_n15402) );
  AND2X2 AND2X2_6898 ( .A(u2__abc_44228_n15403_bF_buf3), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n15404) );
  AND2X2 AND2X2_6899 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_32_), .Y(u2__abc_44228_n15406) );
  AND2X2 AND2X2_69 ( .A(_abc_64468_n753_bF_buf1), .B(sqrto_68_), .Y(_auto_iopadmap_cc_313_execute_65414_104_) );
  AND2X2 AND2X2_690 ( .A(u2__abc_44228_n3251), .B(u2__abc_44228_n3330), .Y(u2__abc_44228_n3331) );
  AND2X2 AND2X2_6900 ( .A(u2__abc_44228_n2988_bF_buf11), .B(1'b0), .Y(u2__abc_44228_n15407) );
  AND2X2 AND2X2_6901 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2_state_2_), .Y(u2__abc_44228_n15408) );
  AND2X2 AND2X2_6902 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_30_), .Y(u2__abc_44228_n15409_1) );
  AND2X2 AND2X2_6903 ( .A(u2__abc_44228_n15410), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n15411) );
  AND2X2 AND2X2_6904 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_33_), .Y(u2__abc_44228_n15413) );
  AND2X2 AND2X2_6905 ( .A(u2__abc_44228_n2988_bF_buf10), .B(1'b0), .Y(u2__abc_44228_n15414) );
  AND2X2 AND2X2_6906 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_31_), .Y(u2__abc_44228_n15415) );
  AND2X2 AND2X2_6907 ( .A(u2__abc_44228_n15416), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n15417) );
  AND2X2 AND2X2_6908 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_34_), .Y(u2__abc_44228_n15419_1) );
  AND2X2 AND2X2_6909 ( .A(u2__abc_44228_n2988_bF_buf9), .B(1'b0), .Y(u2__abc_44228_n15420) );
  AND2X2 AND2X2_691 ( .A(u2__abc_44228_n3240), .B(u2__abc_44228_n3332), .Y(u2__abc_44228_n3333) );
  AND2X2 AND2X2_6910 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_32_), .Y(u2__abc_44228_n15421) );
  AND2X2 AND2X2_6911 ( .A(u2__abc_44228_n15422), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n15423) );
  AND2X2 AND2X2_6912 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_35_), .Y(u2__abc_44228_n15425) );
  AND2X2 AND2X2_6913 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_33_), .Y(u2__abc_44228_n15426) );
  AND2X2 AND2X2_6914 ( .A(u2__abc_44228_n2988_bF_buf8), .B(1'b0), .Y(u2__abc_44228_n15427_1) );
  AND2X2 AND2X2_6915 ( .A(u2__abc_44228_n15428), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n15429) );
  AND2X2 AND2X2_6916 ( .A(u2__abc_44228_n15403_bF_buf2), .B(u2_remLo_36_), .Y(u2__abc_44228_n15431) );
  AND2X2 AND2X2_6917 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_34_), .Y(u2__abc_44228_n15432) );
  AND2X2 AND2X2_6918 ( .A(u2__abc_44228_n15433), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n15434) );
  AND2X2 AND2X2_6919 ( .A(u2__abc_44228_n15402_bF_buf2), .B(u2_remLo_36_), .Y(u2__abc_44228_n15435_1) );
  AND2X2 AND2X2_692 ( .A(u2__abc_44228_n3334), .B(u2__abc_44228_n3243), .Y(u2__abc_44228_n3335) );
  AND2X2 AND2X2_6920 ( .A(u2__abc_44228_n2989_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n15436) );
  AND2X2 AND2X2_6921 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_37_), .Y(u2__abc_44228_n15439) );
  AND2X2 AND2X2_6922 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_35_), .Y(u2__abc_44228_n15440) );
  AND2X2 AND2X2_6923 ( .A(u2__abc_44228_n2988_bF_buf7), .B(1'b0), .Y(u2__abc_44228_n15441) );
  AND2X2 AND2X2_6924 ( .A(u2__abc_44228_n15442_1), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n15443) );
  AND2X2 AND2X2_6925 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_38_), .Y(u2__abc_44228_n15445) );
  AND2X2 AND2X2_6926 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_36_), .Y(u2__abc_44228_n15446) );
  AND2X2 AND2X2_6927 ( .A(u2__abc_44228_n2988_bF_buf6), .B(1'b0), .Y(u2__abc_44228_n15447) );
  AND2X2 AND2X2_6928 ( .A(u2__abc_44228_n15448), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n15449) );
  AND2X2 AND2X2_6929 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_39_), .Y(u2__abc_44228_n15451) );
  AND2X2 AND2X2_693 ( .A(u2__abc_44228_n3336), .B(u2__abc_44228_n3223), .Y(u2__abc_44228_n3337) );
  AND2X2 AND2X2_6930 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_37_), .Y(u2__abc_44228_n15452) );
  AND2X2 AND2X2_6931 ( .A(u2__abc_44228_n2988_bF_buf5), .B(1'b0), .Y(u2__abc_44228_n15453) );
  AND2X2 AND2X2_6932 ( .A(u2__abc_44228_n15454), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n15455_1) );
  AND2X2 AND2X2_6933 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_40_), .Y(u2__abc_44228_n15457) );
  AND2X2 AND2X2_6934 ( .A(u2__abc_44228_n2988_bF_buf4), .B(1'b0), .Y(u2__abc_44228_n15458) );
  AND2X2 AND2X2_6935 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_38_), .Y(u2__abc_44228_n15459) );
  AND2X2 AND2X2_6936 ( .A(u2__abc_44228_n15460), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n15461) );
  AND2X2 AND2X2_6937 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_41_), .Y(u2__abc_44228_n15463_1) );
  AND2X2 AND2X2_6938 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_39_), .Y(u2__abc_44228_n15464) );
  AND2X2 AND2X2_6939 ( .A(u2__abc_44228_n2988_bF_buf3), .B(1'b0), .Y(u2__abc_44228_n15465) );
  AND2X2 AND2X2_694 ( .A(u2__abc_44228_n3338), .B(u2__abc_44228_n3217), .Y(u2__abc_44228_n3339) );
  AND2X2 AND2X2_6940 ( .A(u2__abc_44228_n15466), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n15467) );
  AND2X2 AND2X2_6941 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_42_), .Y(u2__abc_44228_n15469) );
  AND2X2 AND2X2_6942 ( .A(u2__abc_44228_n2988_bF_buf2), .B(1'b0), .Y(u2__abc_44228_n15470) );
  AND2X2 AND2X2_6943 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_40_), .Y(u2__abc_44228_n15471) );
  AND2X2 AND2X2_6944 ( .A(u2__abc_44228_n15472_1), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n15473_1) );
  AND2X2 AND2X2_6945 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_43_), .Y(u2__abc_44228_n15475) );
  AND2X2 AND2X2_6946 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_41_), .Y(u2__abc_44228_n15476) );
  AND2X2 AND2X2_6947 ( .A(u2__abc_44228_n2988_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n15477) );
  AND2X2 AND2X2_6948 ( .A(u2__abc_44228_n15478), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n15479) );
  AND2X2 AND2X2_6949 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_44_), .Y(u2__abc_44228_n15481_1) );
  AND2X2 AND2X2_695 ( .A(u2__abc_44228_n3340), .B(u2__abc_44228_n3220), .Y(u2__abc_44228_n3341) );
  AND2X2 AND2X2_6950 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_42_), .Y(u2__abc_44228_n15482) );
  AND2X2 AND2X2_6951 ( .A(u2__abc_44228_n2988_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n15483) );
  AND2X2 AND2X2_6952 ( .A(u2__abc_44228_n15484), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n15485) );
  AND2X2 AND2X2_6953 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_45_), .Y(u2__abc_44228_n15487) );
  AND2X2 AND2X2_6954 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_43_), .Y(u2__abc_44228_n15488) );
  AND2X2 AND2X2_6955 ( .A(u2__abc_44228_n2988_bF_buf13), .B(1'b0), .Y(u2__abc_44228_n15489) );
  AND2X2 AND2X2_6956 ( .A(u2__abc_44228_n15490), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n15491) );
  AND2X2 AND2X2_6957 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_46_), .Y(u2__abc_44228_n15493) );
  AND2X2 AND2X2_6958 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_44_), .Y(u2__abc_44228_n15494) );
  AND2X2 AND2X2_6959 ( .A(u2__abc_44228_n2988_bF_buf12), .B(1'b0), .Y(u2__abc_44228_n15495) );
  AND2X2 AND2X2_696 ( .A(u2__abc_44228_n3341), .B(u2__abc_44228_n3208), .Y(u2__abc_44228_n3342) );
  AND2X2 AND2X2_6960 ( .A(u2__abc_44228_n15496), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n15497) );
  AND2X2 AND2X2_6961 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_47_), .Y(u2__abc_44228_n15499) );
  AND2X2 AND2X2_6962 ( .A(u2__abc_44228_n2988_bF_buf11), .B(1'b0), .Y(u2__abc_44228_n15500) );
  AND2X2 AND2X2_6963 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_45_), .Y(u2__abc_44228_n15501) );
  AND2X2 AND2X2_6964 ( .A(u2__abc_44228_n15502), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n15503) );
  AND2X2 AND2X2_6965 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_48_), .Y(u2__abc_44228_n15505) );
  AND2X2 AND2X2_6966 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_46_), .Y(u2__abc_44228_n15506) );
  AND2X2 AND2X2_6967 ( .A(u2__abc_44228_n2988_bF_buf10), .B(1'b0), .Y(u2__abc_44228_n15507) );
  AND2X2 AND2X2_6968 ( .A(u2__abc_44228_n15508), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n15509) );
  AND2X2 AND2X2_6969 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_49_), .Y(u2__abc_44228_n15511) );
  AND2X2 AND2X2_697 ( .A(u2__abc_44228_n3200), .B(u2__abc_44228_n3203), .Y(u2__abc_44228_n3343) );
  AND2X2 AND2X2_6970 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_47_), .Y(u2__abc_44228_n15512) );
  AND2X2 AND2X2_6971 ( .A(u2__abc_44228_n2988_bF_buf9), .B(1'b0), .Y(u2__abc_44228_n15513) );
  AND2X2 AND2X2_6972 ( .A(u2__abc_44228_n15514), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n15515) );
  AND2X2 AND2X2_6973 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_50_), .Y(u2__abc_44228_n15517) );
  AND2X2 AND2X2_6974 ( .A(u2__abc_44228_n2988_bF_buf8), .B(1'b0), .Y(u2__abc_44228_n15518) );
  AND2X2 AND2X2_6975 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_48_), .Y(u2__abc_44228_n15519) );
  AND2X2 AND2X2_6976 ( .A(u2__abc_44228_n15520), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n15521) );
  AND2X2 AND2X2_6977 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_51_), .Y(u2__abc_44228_n15523) );
  AND2X2 AND2X2_6978 ( .A(u2__abc_44228_n2988_bF_buf7), .B(1'b0), .Y(u2__abc_44228_n15524) );
  AND2X2 AND2X2_6979 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_49_), .Y(u2__abc_44228_n15525) );
  AND2X2 AND2X2_698 ( .A(u2__abc_44228_n3349), .B(u2_remHi_61_), .Y(u2__abc_44228_n3350) );
  AND2X2 AND2X2_6980 ( .A(u2__abc_44228_n15526), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n15527) );
  AND2X2 AND2X2_6981 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_52_), .Y(u2__abc_44228_n15529) );
  AND2X2 AND2X2_6982 ( .A(u2__abc_44228_n2988_bF_buf6), .B(1'b0), .Y(u2__abc_44228_n15530) );
  AND2X2 AND2X2_6983 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_50_), .Y(u2__abc_44228_n15531) );
  AND2X2 AND2X2_6984 ( .A(u2__abc_44228_n15532), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n15533) );
  AND2X2 AND2X2_6985 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_53_), .Y(u2__abc_44228_n15535) );
  AND2X2 AND2X2_6986 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_51_), .Y(u2__abc_44228_n15536) );
  AND2X2 AND2X2_6987 ( .A(u2__abc_44228_n2988_bF_buf5), .B(1'b0), .Y(u2__abc_44228_n15537) );
  AND2X2 AND2X2_6988 ( .A(u2__abc_44228_n15538), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n15539) );
  AND2X2 AND2X2_6989 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_52_), .Y(u2__abc_44228_n15541) );
  AND2X2 AND2X2_699 ( .A(u2__abc_44228_n3352), .B(sqrto_61_), .Y(u2__abc_44228_n3353) );
  AND2X2 AND2X2_6990 ( .A(u2__abc_44228_n15403_bF_buf1), .B(u2_remLo_54_), .Y(u2__abc_44228_n15542) );
  AND2X2 AND2X2_6991 ( .A(u2__abc_44228_n15543), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n15544) );
  AND2X2 AND2X2_6992 ( .A(u2__abc_44228_n15402_bF_buf1), .B(u2_remLo_54_), .Y(u2__abc_44228_n15545) );
  AND2X2 AND2X2_6993 ( .A(u2__abc_44228_n2989_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n15546) );
  AND2X2 AND2X2_6994 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_55_), .Y(u2__abc_44228_n15549) );
  AND2X2 AND2X2_6995 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_53_), .Y(u2__abc_44228_n15550) );
  AND2X2 AND2X2_6996 ( .A(u2__abc_44228_n2988_bF_buf4), .B(1'b0), .Y(u2__abc_44228_n15551) );
  AND2X2 AND2X2_6997 ( .A(u2__abc_44228_n15552), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n15553) );
  AND2X2 AND2X2_6998 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_56_), .Y(u2__abc_44228_n15555) );
  AND2X2 AND2X2_6999 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_54_), .Y(u2__abc_44228_n15556) );
  AND2X2 AND2X2_7 ( .A(_abc_64468_n753_bF_buf7), .B(sqrto_6_), .Y(_auto_iopadmap_cc_313_execute_65414_42_) );
  AND2X2 AND2X2_70 ( .A(_abc_64468_n753_bF_buf0), .B(sqrto_69_), .Y(_auto_iopadmap_cc_313_execute_65414_105_) );
  AND2X2 AND2X2_700 ( .A(u2__abc_44228_n3351), .B(u2__abc_44228_n3354), .Y(u2__abc_44228_n3355) );
  AND2X2 AND2X2_7000 ( .A(u2__abc_44228_n2988_bF_buf3), .B(1'b0), .Y(u2__abc_44228_n15557) );
  AND2X2 AND2X2_7001 ( .A(u2__abc_44228_n15558), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n15559) );
  AND2X2 AND2X2_7002 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_57_), .Y(u2__abc_44228_n15561) );
  AND2X2 AND2X2_7003 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_55_), .Y(u2__abc_44228_n15562) );
  AND2X2 AND2X2_7004 ( .A(u2__abc_44228_n2988_bF_buf2), .B(1'b0), .Y(u2__abc_44228_n15563) );
  AND2X2 AND2X2_7005 ( .A(u2__abc_44228_n15564), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n15565) );
  AND2X2 AND2X2_7006 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_58_), .Y(u2__abc_44228_n15567) );
  AND2X2 AND2X2_7007 ( .A(u2__abc_44228_n2988_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n15568) );
  AND2X2 AND2X2_7008 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_56_), .Y(u2__abc_44228_n15569) );
  AND2X2 AND2X2_7009 ( .A(u2__abc_44228_n15570), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n15571) );
  AND2X2 AND2X2_701 ( .A(u2__abc_44228_n3356), .B(u2_remHi_60_), .Y(u2__abc_44228_n3357) );
  AND2X2 AND2X2_7010 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_59_), .Y(u2__abc_44228_n15573) );
  AND2X2 AND2X2_7011 ( .A(u2__abc_44228_n2988_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n15574) );
  AND2X2 AND2X2_7012 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_57_), .Y(u2__abc_44228_n15575) );
  AND2X2 AND2X2_7013 ( .A(u2__abc_44228_n15576), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n15577) );
  AND2X2 AND2X2_7014 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_60_), .Y(u2__abc_44228_n15579) );
  AND2X2 AND2X2_7015 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_58_), .Y(u2__abc_44228_n15580) );
  AND2X2 AND2X2_7016 ( .A(u2__abc_44228_n2988_bF_buf13), .B(1'b0), .Y(u2__abc_44228_n15581) );
  AND2X2 AND2X2_7017 ( .A(u2__abc_44228_n15582), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n15583) );
  AND2X2 AND2X2_7018 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_61_), .Y(u2__abc_44228_n15585) );
  AND2X2 AND2X2_7019 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_59_), .Y(u2__abc_44228_n15586) );
  AND2X2 AND2X2_702 ( .A(u2__abc_44228_n3358), .B(sqrto_60_), .Y(u2__abc_44228_n3359) );
  AND2X2 AND2X2_7020 ( .A(u2__abc_44228_n2988_bF_buf12), .B(1'b0), .Y(u2__abc_44228_n15587) );
  AND2X2 AND2X2_7021 ( .A(u2__abc_44228_n15588), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n15589) );
  AND2X2 AND2X2_7022 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_62_), .Y(u2__abc_44228_n15591) );
  AND2X2 AND2X2_7023 ( .A(u2__abc_44228_n2988_bF_buf11), .B(1'b0), .Y(u2__abc_44228_n15592) );
  AND2X2 AND2X2_7024 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_60_), .Y(u2__abc_44228_n15593) );
  AND2X2 AND2X2_7025 ( .A(u2__abc_44228_n15594), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n15595) );
  AND2X2 AND2X2_7026 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_63_), .Y(u2__abc_44228_n15597) );
  AND2X2 AND2X2_7027 ( .A(u2__abc_44228_n2988_bF_buf10), .B(1'b0), .Y(u2__abc_44228_n15598) );
  AND2X2 AND2X2_7028 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_61_), .Y(u2__abc_44228_n15599) );
  AND2X2 AND2X2_7029 ( .A(u2__abc_44228_n15600), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n15601) );
  AND2X2 AND2X2_703 ( .A(u2__abc_44228_n3361), .B(u2__abc_44228_n3355), .Y(u2__abc_44228_n3362) );
  AND2X2 AND2X2_7030 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_64_), .Y(u2__abc_44228_n15603) );
  AND2X2 AND2X2_7031 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_62_), .Y(u2__abc_44228_n15604) );
  AND2X2 AND2X2_7032 ( .A(u2__abc_44228_n2988_bF_buf9), .B(1'b0), .Y(u2__abc_44228_n15605) );
  AND2X2 AND2X2_7033 ( .A(u2__abc_44228_n15606), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n15607) );
  AND2X2 AND2X2_7034 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_65_), .Y(u2__abc_44228_n15609) );
  AND2X2 AND2X2_7035 ( .A(u2__abc_44228_n2988_bF_buf8), .B(1'b0), .Y(u2__abc_44228_n15610) );
  AND2X2 AND2X2_7036 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_63_), .Y(u2__abc_44228_n15611) );
  AND2X2 AND2X2_7037 ( .A(u2__abc_44228_n15612), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n15613) );
  AND2X2 AND2X2_7038 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_66_), .Y(u2__abc_44228_n15615) );
  AND2X2 AND2X2_7039 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_64_), .Y(u2__abc_44228_n15616) );
  AND2X2 AND2X2_704 ( .A(u2__abc_44228_n3363), .B(u2_remHi_58_), .Y(u2__abc_44228_n3364) );
  AND2X2 AND2X2_7040 ( .A(u2__abc_44228_n2988_bF_buf7), .B(1'b0), .Y(u2__abc_44228_n15617) );
  AND2X2 AND2X2_7041 ( .A(u2__abc_44228_n15618), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n15619) );
  AND2X2 AND2X2_7042 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_67_), .Y(u2__abc_44228_n15621) );
  AND2X2 AND2X2_7043 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_65_), .Y(u2__abc_44228_n15622) );
  AND2X2 AND2X2_7044 ( .A(u2__abc_44228_n2988_bF_buf6), .B(1'b0), .Y(u2__abc_44228_n15623) );
  AND2X2 AND2X2_7045 ( .A(u2__abc_44228_n15624), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n15625) );
  AND2X2 AND2X2_7046 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_68_), .Y(u2__abc_44228_n15627) );
  AND2X2 AND2X2_7047 ( .A(u2__abc_44228_n2988_bF_buf5), .B(1'b0), .Y(u2__abc_44228_n15628) );
  AND2X2 AND2X2_7048 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_66_), .Y(u2__abc_44228_n15629) );
  AND2X2 AND2X2_7049 ( .A(u2__abc_44228_n15630), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n15631) );
  AND2X2 AND2X2_705 ( .A(u2__abc_44228_n3365), .B(sqrto_58_), .Y(u2__abc_44228_n3366) );
  AND2X2 AND2X2_7050 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_69_), .Y(u2__abc_44228_n15633) );
  AND2X2 AND2X2_7051 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_67_), .Y(u2__abc_44228_n15634) );
  AND2X2 AND2X2_7052 ( .A(u2__abc_44228_n2988_bF_buf4), .B(1'b0), .Y(u2__abc_44228_n15635) );
  AND2X2 AND2X2_7053 ( .A(u2__abc_44228_n15636), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n15637) );
  AND2X2 AND2X2_7054 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_70_), .Y(u2__abc_44228_n15639) );
  AND2X2 AND2X2_7055 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_68_), .Y(u2__abc_44228_n15640) );
  AND2X2 AND2X2_7056 ( .A(u2__abc_44228_n2988_bF_buf3), .B(1'b0), .Y(u2__abc_44228_n15641) );
  AND2X2 AND2X2_7057 ( .A(u2__abc_44228_n15642), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n15643) );
  AND2X2 AND2X2_7058 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_71_), .Y(u2__abc_44228_n15645) );
  AND2X2 AND2X2_7059 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_69_), .Y(u2__abc_44228_n15646) );
  AND2X2 AND2X2_706 ( .A(u2__abc_44228_n3369), .B(u2_remHi_59_), .Y(u2__abc_44228_n3370) );
  AND2X2 AND2X2_7060 ( .A(u2__abc_44228_n2988_bF_buf2), .B(1'b0), .Y(u2__abc_44228_n15647) );
  AND2X2 AND2X2_7061 ( .A(u2__abc_44228_n15648), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n15649) );
  AND2X2 AND2X2_7062 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_72_), .Y(u2__abc_44228_n15651) );
  AND2X2 AND2X2_7063 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_70_), .Y(u2__abc_44228_n15652) );
  AND2X2 AND2X2_7064 ( .A(u2__abc_44228_n2988_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n15653) );
  AND2X2 AND2X2_7065 ( .A(u2__abc_44228_n15654), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n15655) );
  AND2X2 AND2X2_7066 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_73_), .Y(u2__abc_44228_n15657) );
  AND2X2 AND2X2_7067 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_71_), .Y(u2__abc_44228_n15658) );
  AND2X2 AND2X2_7068 ( .A(u2__abc_44228_n2988_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n15659) );
  AND2X2 AND2X2_7069 ( .A(u2__abc_44228_n15660), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n15661) );
  AND2X2 AND2X2_707 ( .A(u2__abc_44228_n3372), .B(sqrto_59_), .Y(u2__abc_44228_n3373) );
  AND2X2 AND2X2_7070 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_74_), .Y(u2__abc_44228_n15663) );
  AND2X2 AND2X2_7071 ( .A(u2__abc_44228_n2988_bF_buf13), .B(1'b0), .Y(u2__abc_44228_n15664) );
  AND2X2 AND2X2_7072 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_72_), .Y(u2__abc_44228_n15665) );
  AND2X2 AND2X2_7073 ( .A(u2__abc_44228_n15666), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n15667) );
  AND2X2 AND2X2_7074 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_75_), .Y(u2__abc_44228_n15669) );
  AND2X2 AND2X2_7075 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_73_), .Y(u2__abc_44228_n15670) );
  AND2X2 AND2X2_7076 ( .A(u2__abc_44228_n2988_bF_buf12), .B(1'b0), .Y(u2__abc_44228_n15671) );
  AND2X2 AND2X2_7077 ( .A(u2__abc_44228_n15672), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n15673) );
  AND2X2 AND2X2_7078 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_76_), .Y(u2__abc_44228_n15675) );
  AND2X2 AND2X2_7079 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_74_), .Y(u2__abc_44228_n15676) );
  AND2X2 AND2X2_708 ( .A(u2__abc_44228_n3371), .B(u2__abc_44228_n3374), .Y(u2__abc_44228_n3375) );
  AND2X2 AND2X2_7080 ( .A(u2__abc_44228_n2988_bF_buf11), .B(1'b0), .Y(u2__abc_44228_n15677) );
  AND2X2 AND2X2_7081 ( .A(u2__abc_44228_n15678), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n15679) );
  AND2X2 AND2X2_7082 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_77_), .Y(u2__abc_44228_n15681) );
  AND2X2 AND2X2_7083 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_75_), .Y(u2__abc_44228_n15682) );
  AND2X2 AND2X2_7084 ( .A(u2__abc_44228_n2988_bF_buf10), .B(1'b0), .Y(u2__abc_44228_n15683) );
  AND2X2 AND2X2_7085 ( .A(u2__abc_44228_n15684), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n15685) );
  AND2X2 AND2X2_7086 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_78_), .Y(u2__abc_44228_n15687) );
  AND2X2 AND2X2_7087 ( .A(u2__abc_44228_n2988_bF_buf9), .B(1'b0), .Y(u2__abc_44228_n15688) );
  AND2X2 AND2X2_7088 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_76_), .Y(u2__abc_44228_n15689) );
  AND2X2 AND2X2_7089 ( .A(u2__abc_44228_n15690), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n15691) );
  AND2X2 AND2X2_709 ( .A(u2__abc_44228_n3368), .B(u2__abc_44228_n3375), .Y(u2__abc_44228_n3376) );
  AND2X2 AND2X2_7090 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_79_), .Y(u2__abc_44228_n15693) );
  AND2X2 AND2X2_7091 ( .A(u2__abc_44228_n2988_bF_buf8), .B(1'b0), .Y(u2__abc_44228_n15694) );
  AND2X2 AND2X2_7092 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_77_), .Y(u2__abc_44228_n15695) );
  AND2X2 AND2X2_7093 ( .A(u2__abc_44228_n15696), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n15697) );
  AND2X2 AND2X2_7094 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_80_), .Y(u2__abc_44228_n15699) );
  AND2X2 AND2X2_7095 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_78_), .Y(u2__abc_44228_n15700) );
  AND2X2 AND2X2_7096 ( .A(u2__abc_44228_n2988_bF_buf7), .B(1'b0), .Y(u2__abc_44228_n15701) );
  AND2X2 AND2X2_7097 ( .A(u2__abc_44228_n15702), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n15703) );
  AND2X2 AND2X2_7098 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_81_), .Y(u2__abc_44228_n15705) );
  AND2X2 AND2X2_7099 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_79_), .Y(u2__abc_44228_n15706) );
  AND2X2 AND2X2_71 ( .A(_abc_64468_n753_bF_buf13), .B(sqrto_70_), .Y(_auto_iopadmap_cc_313_execute_65414_106_) );
  AND2X2 AND2X2_710 ( .A(u2__abc_44228_n3362), .B(u2__abc_44228_n3376), .Y(u2__abc_44228_n3377) );
  AND2X2 AND2X2_7100 ( .A(u2__abc_44228_n2988_bF_buf6), .B(1'b0), .Y(u2__abc_44228_n15707) );
  AND2X2 AND2X2_7101 ( .A(u2__abc_44228_n15708), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n15709) );
  AND2X2 AND2X2_7102 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_82_), .Y(u2__abc_44228_n15711) );
  AND2X2 AND2X2_7103 ( .A(u2__abc_44228_n2988_bF_buf5), .B(1'b0), .Y(u2__abc_44228_n15712) );
  AND2X2 AND2X2_7104 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_80_), .Y(u2__abc_44228_n15713) );
  AND2X2 AND2X2_7105 ( .A(u2__abc_44228_n15714), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n15715) );
  AND2X2 AND2X2_7106 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_83_), .Y(u2__abc_44228_n15717) );
  AND2X2 AND2X2_7107 ( .A(u2__abc_44228_n2988_bF_buf4), .B(1'b0), .Y(u2__abc_44228_n15718) );
  AND2X2 AND2X2_7108 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_81_), .Y(u2__abc_44228_n15719) );
  AND2X2 AND2X2_7109 ( .A(u2__abc_44228_n15720), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n15721) );
  AND2X2 AND2X2_711 ( .A(u2__abc_44228_n3378), .B(u2_remHi_57_), .Y(u2__abc_44228_n3379) );
  AND2X2 AND2X2_7110 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_84_), .Y(u2__abc_44228_n15723) );
  AND2X2 AND2X2_7111 ( .A(u2__abc_44228_n2988_bF_buf3), .B(1'b0), .Y(u2__abc_44228_n15724) );
  AND2X2 AND2X2_7112 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_82_), .Y(u2__abc_44228_n15725) );
  AND2X2 AND2X2_7113 ( .A(u2__abc_44228_n15726), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n15727) );
  AND2X2 AND2X2_7114 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_85_), .Y(u2__abc_44228_n15729) );
  AND2X2 AND2X2_7115 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_83_), .Y(u2__abc_44228_n15730) );
  AND2X2 AND2X2_7116 ( .A(u2__abc_44228_n2988_bF_buf2), .B(1'b0), .Y(u2__abc_44228_n15731) );
  AND2X2 AND2X2_7117 ( .A(u2__abc_44228_n15732), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n15733) );
  AND2X2 AND2X2_7118 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_84_), .Y(u2__abc_44228_n15735) );
  AND2X2 AND2X2_7119 ( .A(u2__abc_44228_n15403_bF_buf0), .B(u2_remLo_86_), .Y(u2__abc_44228_n15736) );
  AND2X2 AND2X2_712 ( .A(u2__abc_44228_n3381), .B(sqrto_57_), .Y(u2__abc_44228_n3382) );
  AND2X2 AND2X2_7120 ( .A(u2__abc_44228_n15737), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n15738) );
  AND2X2 AND2X2_7121 ( .A(u2__abc_44228_n15402_bF_buf0), .B(u2_remLo_86_), .Y(u2__abc_44228_n15739) );
  AND2X2 AND2X2_7122 ( .A(u2__abc_44228_n2989_bF_buf3), .B(1'b0), .Y(u2__abc_44228_n15740) );
  AND2X2 AND2X2_7123 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_87_), .Y(u2__abc_44228_n15743) );
  AND2X2 AND2X2_7124 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_85_), .Y(u2__abc_44228_n15744) );
  AND2X2 AND2X2_7125 ( .A(u2__abc_44228_n2988_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n15745) );
  AND2X2 AND2X2_7126 ( .A(u2__abc_44228_n15746), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n15747) );
  AND2X2 AND2X2_7127 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_88_), .Y(u2__abc_44228_n15749) );
  AND2X2 AND2X2_7128 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_86_), .Y(u2__abc_44228_n15750) );
  AND2X2 AND2X2_7129 ( .A(u2__abc_44228_n2988_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n15751) );
  AND2X2 AND2X2_713 ( .A(u2__abc_44228_n3380), .B(u2__abc_44228_n3383), .Y(u2__abc_44228_n3384) );
  AND2X2 AND2X2_7130 ( .A(u2__abc_44228_n15752), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n15753) );
  AND2X2 AND2X2_7131 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_89_), .Y(u2__abc_44228_n15755) );
  AND2X2 AND2X2_7132 ( .A(u2__abc_44228_n2988_bF_buf13), .B(1'b0), .Y(u2__abc_44228_n15756) );
  AND2X2 AND2X2_7133 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_87_), .Y(u2__abc_44228_n15757) );
  AND2X2 AND2X2_7134 ( .A(u2__abc_44228_n15758), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n15759) );
  AND2X2 AND2X2_7135 ( .A(u2__abc_44228_n15403_bF_buf3), .B(u2_remLo_90_), .Y(u2__abc_44228_n15761) );
  AND2X2 AND2X2_7136 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_88_), .Y(u2__abc_44228_n15762) );
  AND2X2 AND2X2_7137 ( .A(u2__abc_44228_n15763), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n15764) );
  AND2X2 AND2X2_7138 ( .A(u2__abc_44228_n15402_bF_buf3), .B(u2_remLo_90_), .Y(u2__abc_44228_n15765) );
  AND2X2 AND2X2_7139 ( .A(u2__abc_44228_n2989_bF_buf2), .B(1'b0), .Y(u2__abc_44228_n15766) );
  AND2X2 AND2X2_714 ( .A(u2__abc_44228_n3385), .B(u2_remHi_56_), .Y(u2__abc_44228_n3386) );
  AND2X2 AND2X2_7140 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_91_), .Y(u2__abc_44228_n15769) );
  AND2X2 AND2X2_7141 ( .A(u2__abc_44228_n2988_bF_buf12), .B(1'b0), .Y(u2__abc_44228_n15770) );
  AND2X2 AND2X2_7142 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_89_), .Y(u2__abc_44228_n15771) );
  AND2X2 AND2X2_7143 ( .A(u2__abc_44228_n15772), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n15773) );
  AND2X2 AND2X2_7144 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_92_), .Y(u2__abc_44228_n15775) );
  AND2X2 AND2X2_7145 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_90_), .Y(u2__abc_44228_n15776) );
  AND2X2 AND2X2_7146 ( .A(u2__abc_44228_n2988_bF_buf11), .B(1'b0), .Y(u2__abc_44228_n15777) );
  AND2X2 AND2X2_7147 ( .A(u2__abc_44228_n15778), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n15779) );
  AND2X2 AND2X2_7148 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_93_), .Y(u2__abc_44228_n15781) );
  AND2X2 AND2X2_7149 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_91_), .Y(u2__abc_44228_n15782) );
  AND2X2 AND2X2_715 ( .A(u2__abc_44228_n3387), .B(sqrto_56_), .Y(u2__abc_44228_n3388) );
  AND2X2 AND2X2_7150 ( .A(u2__abc_44228_n2988_bF_buf10), .B(1'b0), .Y(u2__abc_44228_n15783) );
  AND2X2 AND2X2_7151 ( .A(u2__abc_44228_n15784), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n15785) );
  AND2X2 AND2X2_7152 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_94_), .Y(u2__abc_44228_n15787) );
  AND2X2 AND2X2_7153 ( .A(u2__abc_44228_n2988_bF_buf9), .B(1'b0), .Y(u2__abc_44228_n15788) );
  AND2X2 AND2X2_7154 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_92_), .Y(u2__abc_44228_n15789) );
  AND2X2 AND2X2_7155 ( .A(u2__abc_44228_n15790), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n15791) );
  AND2X2 AND2X2_7156 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_95_), .Y(u2__abc_44228_n15793) );
  AND2X2 AND2X2_7157 ( .A(u2__abc_44228_n2988_bF_buf8), .B(1'b0), .Y(u2__abc_44228_n15794) );
  AND2X2 AND2X2_7158 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_93_), .Y(u2__abc_44228_n15795) );
  AND2X2 AND2X2_7159 ( .A(u2__abc_44228_n15796), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n15797) );
  AND2X2 AND2X2_716 ( .A(u2__abc_44228_n3390), .B(u2__abc_44228_n3384), .Y(u2__abc_44228_n3391) );
  AND2X2 AND2X2_7160 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_96_), .Y(u2__abc_44228_n15799) );
  AND2X2 AND2X2_7161 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_94_), .Y(u2__abc_44228_n15800) );
  AND2X2 AND2X2_7162 ( .A(u2__abc_44228_n2988_bF_buf7), .B(1'b0), .Y(u2__abc_44228_n15801) );
  AND2X2 AND2X2_7163 ( .A(u2__abc_44228_n15802), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n15803) );
  AND2X2 AND2X2_7164 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_97_), .Y(u2__abc_44228_n15805) );
  AND2X2 AND2X2_7165 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_95_), .Y(u2__abc_44228_n15806) );
  AND2X2 AND2X2_7166 ( .A(u2__abc_44228_n2988_bF_buf6), .B(1'b0), .Y(u2__abc_44228_n15807) );
  AND2X2 AND2X2_7167 ( .A(u2__abc_44228_n15808), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n15809) );
  AND2X2 AND2X2_7168 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_98_), .Y(u2__abc_44228_n15811) );
  AND2X2 AND2X2_7169 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_96_), .Y(u2__abc_44228_n15812) );
  AND2X2 AND2X2_717 ( .A(u2__abc_44228_n3392), .B(u2_remHi_55_), .Y(u2__abc_44228_n3393) );
  AND2X2 AND2X2_7170 ( .A(u2__abc_44228_n2988_bF_buf5), .B(1'b0), .Y(u2__abc_44228_n15813) );
  AND2X2 AND2X2_7171 ( .A(u2__abc_44228_n15814), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n15815) );
  AND2X2 AND2X2_7172 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_99_), .Y(u2__abc_44228_n15817) );
  AND2X2 AND2X2_7173 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_97_), .Y(u2__abc_44228_n15818) );
  AND2X2 AND2X2_7174 ( .A(u2__abc_44228_n2988_bF_buf4), .B(1'b0), .Y(u2__abc_44228_n15819) );
  AND2X2 AND2X2_7175 ( .A(u2__abc_44228_n15820), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n15821) );
  AND2X2 AND2X2_7176 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_100_), .Y(u2__abc_44228_n15823) );
  AND2X2 AND2X2_7177 ( .A(u2__abc_44228_n2988_bF_buf3), .B(1'b0), .Y(u2__abc_44228_n15824) );
  AND2X2 AND2X2_7178 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_98_), .Y(u2__abc_44228_n15825) );
  AND2X2 AND2X2_7179 ( .A(u2__abc_44228_n15826), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n15827) );
  AND2X2 AND2X2_718 ( .A(u2__abc_44228_n3395), .B(sqrto_55_), .Y(u2__abc_44228_n3396) );
  AND2X2 AND2X2_7180 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_101_), .Y(u2__abc_44228_n15829) );
  AND2X2 AND2X2_7181 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_99_), .Y(u2__abc_44228_n15830) );
  AND2X2 AND2X2_7182 ( .A(u2__abc_44228_n2988_bF_buf2), .B(1'b0), .Y(u2__abc_44228_n15831) );
  AND2X2 AND2X2_7183 ( .A(u2__abc_44228_n15832), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n15833) );
  AND2X2 AND2X2_7184 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_102_), .Y(u2__abc_44228_n15835) );
  AND2X2 AND2X2_7185 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_100_), .Y(u2__abc_44228_n15836) );
  AND2X2 AND2X2_7186 ( .A(u2__abc_44228_n2988_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n15837) );
  AND2X2 AND2X2_7187 ( .A(u2__abc_44228_n15838), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n15839) );
  AND2X2 AND2X2_7188 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_103_), .Y(u2__abc_44228_n15841) );
  AND2X2 AND2X2_7189 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_101_), .Y(u2__abc_44228_n15842) );
  AND2X2 AND2X2_719 ( .A(u2__abc_44228_n3394), .B(u2__abc_44228_n3397), .Y(u2__abc_44228_n3398) );
  AND2X2 AND2X2_7190 ( .A(u2__abc_44228_n2988_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n15843) );
  AND2X2 AND2X2_7191 ( .A(u2__abc_44228_n15844), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n15845) );
  AND2X2 AND2X2_7192 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_104_), .Y(u2__abc_44228_n15847) );
  AND2X2 AND2X2_7193 ( .A(u2__abc_44228_n2988_bF_buf13), .B(1'b0), .Y(u2__abc_44228_n15848) );
  AND2X2 AND2X2_7194 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_102_), .Y(u2__abc_44228_n15849) );
  AND2X2 AND2X2_7195 ( .A(u2__abc_44228_n15850), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n15851) );
  AND2X2 AND2X2_7196 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_105_), .Y(u2__abc_44228_n15853) );
  AND2X2 AND2X2_7197 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_103_), .Y(u2__abc_44228_n15854) );
  AND2X2 AND2X2_7198 ( .A(u2__abc_44228_n2988_bF_buf12), .B(1'b0), .Y(u2__abc_44228_n15855) );
  AND2X2 AND2X2_7199 ( .A(u2__abc_44228_n15856), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n15857) );
  AND2X2 AND2X2_72 ( .A(_abc_64468_n753_bF_buf12), .B(sqrto_71_), .Y(_auto_iopadmap_cc_313_execute_65414_107_) );
  AND2X2 AND2X2_720 ( .A(u2__abc_44228_n3399), .B(u2_remHi_54_), .Y(u2__abc_44228_n3400) );
  AND2X2 AND2X2_7200 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_106_), .Y(u2__abc_44228_n15859) );
  AND2X2 AND2X2_7201 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_104_), .Y(u2__abc_44228_n15860) );
  AND2X2 AND2X2_7202 ( .A(u2__abc_44228_n2988_bF_buf11), .B(1'b0), .Y(u2__abc_44228_n15861) );
  AND2X2 AND2X2_7203 ( .A(u2__abc_44228_n15862), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n15863) );
  AND2X2 AND2X2_7204 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_107_), .Y(u2__abc_44228_n15865) );
  AND2X2 AND2X2_7205 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_105_), .Y(u2__abc_44228_n15866) );
  AND2X2 AND2X2_7206 ( .A(u2__abc_44228_n2988_bF_buf10), .B(1'b0), .Y(u2__abc_44228_n15867) );
  AND2X2 AND2X2_7207 ( .A(u2__abc_44228_n15868), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n15869) );
  AND2X2 AND2X2_7208 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_108_), .Y(u2__abc_44228_n15871) );
  AND2X2 AND2X2_7209 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_106_), .Y(u2__abc_44228_n15872) );
  AND2X2 AND2X2_721 ( .A(u2__abc_44228_n3401), .B(sqrto_54_), .Y(u2__abc_44228_n3402) );
  AND2X2 AND2X2_7210 ( .A(u2__abc_44228_n2988_bF_buf9), .B(1'b0), .Y(u2__abc_44228_n15873) );
  AND2X2 AND2X2_7211 ( .A(u2__abc_44228_n15874), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n15875) );
  AND2X2 AND2X2_7212 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_109_), .Y(u2__abc_44228_n15877) );
  AND2X2 AND2X2_7213 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_107_), .Y(u2__abc_44228_n15878) );
  AND2X2 AND2X2_7214 ( .A(u2__abc_44228_n2988_bF_buf8), .B(1'b0), .Y(u2__abc_44228_n15879) );
  AND2X2 AND2X2_7215 ( .A(u2__abc_44228_n15880), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n15881) );
  AND2X2 AND2X2_7216 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_110_), .Y(u2__abc_44228_n15883) );
  AND2X2 AND2X2_7217 ( .A(u2__abc_44228_n2988_bF_buf7), .B(1'b0), .Y(u2__abc_44228_n15884) );
  AND2X2 AND2X2_7218 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_108_), .Y(u2__abc_44228_n15885) );
  AND2X2 AND2X2_7219 ( .A(u2__abc_44228_n15886), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n15887) );
  AND2X2 AND2X2_722 ( .A(u2__abc_44228_n3404), .B(u2__abc_44228_n3398), .Y(u2__abc_44228_n3405) );
  AND2X2 AND2X2_7220 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_111_), .Y(u2__abc_44228_n15889) );
  AND2X2 AND2X2_7221 ( .A(u2__abc_44228_n2988_bF_buf6), .B(1'b0), .Y(u2__abc_44228_n15890) );
  AND2X2 AND2X2_7222 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_109_), .Y(u2__abc_44228_n15891) );
  AND2X2 AND2X2_7223 ( .A(u2__abc_44228_n15892), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n15893) );
  AND2X2 AND2X2_7224 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_112_), .Y(u2__abc_44228_n15895) );
  AND2X2 AND2X2_7225 ( .A(u2__abc_44228_n2988_bF_buf5), .B(1'b0), .Y(u2__abc_44228_n15896) );
  AND2X2 AND2X2_7226 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_110_), .Y(u2__abc_44228_n15897) );
  AND2X2 AND2X2_7227 ( .A(u2__abc_44228_n15898), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n15899) );
  AND2X2 AND2X2_7228 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_113_), .Y(u2__abc_44228_n15901) );
  AND2X2 AND2X2_7229 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_111_), .Y(u2__abc_44228_n15902) );
  AND2X2 AND2X2_723 ( .A(u2__abc_44228_n3391), .B(u2__abc_44228_n3405), .Y(u2__abc_44228_n3406) );
  AND2X2 AND2X2_7230 ( .A(u2__abc_44228_n2988_bF_buf4), .B(1'b0), .Y(u2__abc_44228_n15903) );
  AND2X2 AND2X2_7231 ( .A(u2__abc_44228_n15904), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n15905) );
  AND2X2 AND2X2_7232 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_114_), .Y(u2__abc_44228_n15907) );
  AND2X2 AND2X2_7233 ( .A(u2__abc_44228_n2988_bF_buf3), .B(1'b0), .Y(u2__abc_44228_n15908) );
  AND2X2 AND2X2_7234 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_112_), .Y(u2__abc_44228_n15909) );
  AND2X2 AND2X2_7235 ( .A(u2__abc_44228_n15910), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n15911) );
  AND2X2 AND2X2_7236 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_115_), .Y(u2__abc_44228_n15913) );
  AND2X2 AND2X2_7237 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_113_), .Y(u2__abc_44228_n15914) );
  AND2X2 AND2X2_7238 ( .A(u2__abc_44228_n2988_bF_buf2), .B(1'b0), .Y(u2__abc_44228_n15915) );
  AND2X2 AND2X2_7239 ( .A(u2__abc_44228_n15916), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n15917) );
  AND2X2 AND2X2_724 ( .A(u2__abc_44228_n3377), .B(u2__abc_44228_n3406), .Y(u2__abc_44228_n3407) );
  AND2X2 AND2X2_7240 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_116_), .Y(u2__abc_44228_n15919) );
  AND2X2 AND2X2_7241 ( .A(u2__abc_44228_n2988_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n15920) );
  AND2X2 AND2X2_7242 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_114_), .Y(u2__abc_44228_n15921) );
  AND2X2 AND2X2_7243 ( .A(u2__abc_44228_n15922), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n15923) );
  AND2X2 AND2X2_7244 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_117_), .Y(u2__abc_44228_n15925) );
  AND2X2 AND2X2_7245 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_115_), .Y(u2__abc_44228_n15926) );
  AND2X2 AND2X2_7246 ( .A(u2__abc_44228_n2988_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n15927) );
  AND2X2 AND2X2_7247 ( .A(u2__abc_44228_n15928), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n15929) );
  AND2X2 AND2X2_7248 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_116_), .Y(u2__abc_44228_n15931) );
  AND2X2 AND2X2_7249 ( .A(u2__abc_44228_n15403_bF_buf2), .B(u2_remLo_118_), .Y(u2__abc_44228_n15932) );
  AND2X2 AND2X2_725 ( .A(u2__abc_44228_n3408), .B(u2_remHi_53_), .Y(u2__abc_44228_n3409) );
  AND2X2 AND2X2_7250 ( .A(u2__abc_44228_n15933), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n15934) );
  AND2X2 AND2X2_7251 ( .A(u2__abc_44228_n15402_bF_buf2), .B(u2_remLo_118_), .Y(u2__abc_44228_n15935) );
  AND2X2 AND2X2_7252 ( .A(u2__abc_44228_n2989_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n15936) );
  AND2X2 AND2X2_7253 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_119_), .Y(u2__abc_44228_n15939) );
  AND2X2 AND2X2_7254 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_117_), .Y(u2__abc_44228_n15940) );
  AND2X2 AND2X2_7255 ( .A(u2__abc_44228_n2988_bF_buf13), .B(1'b0), .Y(u2__abc_44228_n15941) );
  AND2X2 AND2X2_7256 ( .A(u2__abc_44228_n15942), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n15943) );
  AND2X2 AND2X2_7257 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_120_), .Y(u2__abc_44228_n15945) );
  AND2X2 AND2X2_7258 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_118_), .Y(u2__abc_44228_n15946) );
  AND2X2 AND2X2_7259 ( .A(u2__abc_44228_n2988_bF_buf12), .B(1'b0), .Y(u2__abc_44228_n15947) );
  AND2X2 AND2X2_726 ( .A(u2__abc_44228_n3411), .B(sqrto_53_), .Y(u2__abc_44228_n3412) );
  AND2X2 AND2X2_7260 ( .A(u2__abc_44228_n15948), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n15949) );
  AND2X2 AND2X2_7261 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_121_), .Y(u2__abc_44228_n15951) );
  AND2X2 AND2X2_7262 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_119_), .Y(u2__abc_44228_n15952) );
  AND2X2 AND2X2_7263 ( .A(u2__abc_44228_n2988_bF_buf11), .B(1'b0), .Y(u2__abc_44228_n15953) );
  AND2X2 AND2X2_7264 ( .A(u2__abc_44228_n15954), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n15955) );
  AND2X2 AND2X2_7265 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_122_), .Y(u2__abc_44228_n15957) );
  AND2X2 AND2X2_7266 ( .A(u2__abc_44228_n2988_bF_buf10), .B(1'b0), .Y(u2__abc_44228_n15958) );
  AND2X2 AND2X2_7267 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_120_), .Y(u2__abc_44228_n15959) );
  AND2X2 AND2X2_7268 ( .A(u2__abc_44228_n15960), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n15961) );
  AND2X2 AND2X2_7269 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_123_), .Y(u2__abc_44228_n15963) );
  AND2X2 AND2X2_727 ( .A(u2__abc_44228_n3410), .B(u2__abc_44228_n3413), .Y(u2__abc_44228_n3414) );
  AND2X2 AND2X2_7270 ( .A(u2__abc_44228_n2988_bF_buf9), .B(1'b0), .Y(u2__abc_44228_n15964) );
  AND2X2 AND2X2_7271 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_121_), .Y(u2__abc_44228_n15965) );
  AND2X2 AND2X2_7272 ( .A(u2__abc_44228_n15966), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n15967) );
  AND2X2 AND2X2_7273 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_124_), .Y(u2__abc_44228_n15969) );
  AND2X2 AND2X2_7274 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_122_), .Y(u2__abc_44228_n15970) );
  AND2X2 AND2X2_7275 ( .A(u2__abc_44228_n2988_bF_buf8), .B(1'b0), .Y(u2__abc_44228_n15971) );
  AND2X2 AND2X2_7276 ( .A(u2__abc_44228_n15972), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n15973) );
  AND2X2 AND2X2_7277 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_125_), .Y(u2__abc_44228_n15975) );
  AND2X2 AND2X2_7278 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_123_), .Y(u2__abc_44228_n15976) );
  AND2X2 AND2X2_7279 ( .A(u2__abc_44228_n2988_bF_buf7), .B(1'b0), .Y(u2__abc_44228_n15977) );
  AND2X2 AND2X2_728 ( .A(u2__abc_44228_n3415), .B(u2_remHi_52_), .Y(u2__abc_44228_n3416) );
  AND2X2 AND2X2_7280 ( .A(u2__abc_44228_n15978), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n15979) );
  AND2X2 AND2X2_7281 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_126_), .Y(u2__abc_44228_n15981) );
  AND2X2 AND2X2_7282 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_124_), .Y(u2__abc_44228_n15982) );
  AND2X2 AND2X2_7283 ( .A(u2__abc_44228_n2988_bF_buf6), .B(1'b0), .Y(u2__abc_44228_n15983) );
  AND2X2 AND2X2_7284 ( .A(u2__abc_44228_n15984), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n15985) );
  AND2X2 AND2X2_7285 ( .A(u2__abc_44228_n15403_bF_buf1), .B(u2_remLo_127_), .Y(u2__abc_44228_n15987) );
  AND2X2 AND2X2_7286 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_125_), .Y(u2__abc_44228_n15988) );
  AND2X2 AND2X2_7287 ( .A(u2__abc_44228_n15989), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n15990) );
  AND2X2 AND2X2_7288 ( .A(u2__abc_44228_n15402_bF_buf1), .B(u2_remLo_127_), .Y(u2__abc_44228_n15991) );
  AND2X2 AND2X2_7289 ( .A(u2__abc_44228_n2989_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n15992) );
  AND2X2 AND2X2_729 ( .A(u2__abc_44228_n3417), .B(sqrto_52_), .Y(u2__abc_44228_n3418) );
  AND2X2 AND2X2_7290 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_128_), .Y(u2__abc_44228_n15995) );
  AND2X2 AND2X2_7291 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_126_), .Y(u2__abc_44228_n15996) );
  AND2X2 AND2X2_7292 ( .A(u2__abc_44228_n2988_bF_buf5), .B(1'b0), .Y(u2__abc_44228_n15997) );
  AND2X2 AND2X2_7293 ( .A(u2__abc_44228_n15998), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n15999) );
  AND2X2 AND2X2_7294 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_129_), .Y(u2__abc_44228_n16001) );
  AND2X2 AND2X2_7295 ( .A(u2__abc_44228_n2988_bF_buf4), .B(1'b0), .Y(u2__abc_44228_n16002) );
  AND2X2 AND2X2_7296 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_127_), .Y(u2__abc_44228_n16003) );
  AND2X2 AND2X2_7297 ( .A(u2__abc_44228_n16004), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16005) );
  AND2X2 AND2X2_7298 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_130_), .Y(u2__abc_44228_n16007) );
  AND2X2 AND2X2_7299 ( .A(u2__abc_44228_n2988_bF_buf3), .B(1'b0), .Y(u2__abc_44228_n16008) );
  AND2X2 AND2X2_73 ( .A(_abc_64468_n753_bF_buf11), .B(sqrto_72_), .Y(_auto_iopadmap_cc_313_execute_65414_108_) );
  AND2X2 AND2X2_730 ( .A(u2__abc_44228_n3420), .B(u2__abc_44228_n3414), .Y(u2__abc_44228_n3421) );
  AND2X2 AND2X2_7300 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_128_), .Y(u2__abc_44228_n16009) );
  AND2X2 AND2X2_7301 ( .A(u2__abc_44228_n16010), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16011) );
  AND2X2 AND2X2_7302 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_131_), .Y(u2__abc_44228_n16013) );
  AND2X2 AND2X2_7303 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_129_), .Y(u2__abc_44228_n16014) );
  AND2X2 AND2X2_7304 ( .A(u2__abc_44228_n2988_bF_buf2), .B(1'b0), .Y(u2__abc_44228_n16015) );
  AND2X2 AND2X2_7305 ( .A(u2__abc_44228_n16016), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16017) );
  AND2X2 AND2X2_7306 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_132_), .Y(u2__abc_44228_n16019) );
  AND2X2 AND2X2_7307 ( .A(u2__abc_44228_n2988_bF_buf1), .B(1'b0), .Y(u2__abc_44228_n16020) );
  AND2X2 AND2X2_7308 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_130_), .Y(u2__abc_44228_n16021) );
  AND2X2 AND2X2_7309 ( .A(u2__abc_44228_n16022), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16023) );
  AND2X2 AND2X2_731 ( .A(u2__abc_44228_n3422), .B(u2_remHi_50_), .Y(u2__abc_44228_n3423) );
  AND2X2 AND2X2_7310 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_133_), .Y(u2__abc_44228_n16025) );
  AND2X2 AND2X2_7311 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_131_), .Y(u2__abc_44228_n16026) );
  AND2X2 AND2X2_7312 ( .A(u2__abc_44228_n2988_bF_buf0), .B(1'b0), .Y(u2__abc_44228_n16027) );
  AND2X2 AND2X2_7313 ( .A(u2__abc_44228_n16028), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16029) );
  AND2X2 AND2X2_7314 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_134_), .Y(u2__abc_44228_n16031) );
  AND2X2 AND2X2_7315 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_132_), .Y(u2__abc_44228_n16032) );
  AND2X2 AND2X2_7316 ( .A(u2__abc_44228_n2988_bF_buf13), .B(1'b0), .Y(u2__abc_44228_n16033) );
  AND2X2 AND2X2_7317 ( .A(u2__abc_44228_n16034), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16035) );
  AND2X2 AND2X2_7318 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_135_), .Y(u2__abc_44228_n16037) );
  AND2X2 AND2X2_7319 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_133_), .Y(u2__abc_44228_n16038) );
  AND2X2 AND2X2_732 ( .A(u2__abc_44228_n3424), .B(sqrto_50_), .Y(u2__abc_44228_n3425) );
  AND2X2 AND2X2_7320 ( .A(u2__abc_44228_n2988_bF_buf12), .B(1'b0), .Y(u2__abc_44228_n16039) );
  AND2X2 AND2X2_7321 ( .A(u2__abc_44228_n16040), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16041) );
  AND2X2 AND2X2_7322 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_136_), .Y(u2__abc_44228_n16043) );
  AND2X2 AND2X2_7323 ( .A(u2__abc_44228_n2988_bF_buf11), .B(1'b0), .Y(u2__abc_44228_n16044) );
  AND2X2 AND2X2_7324 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_134_), .Y(u2__abc_44228_n16045) );
  AND2X2 AND2X2_7325 ( .A(u2__abc_44228_n16046), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16047) );
  AND2X2 AND2X2_7326 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_137_), .Y(u2__abc_44228_n16049) );
  AND2X2 AND2X2_7327 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_135_), .Y(u2__abc_44228_n16050) );
  AND2X2 AND2X2_7328 ( .A(u2__abc_44228_n2988_bF_buf10), .B(1'b0), .Y(u2__abc_44228_n16051) );
  AND2X2 AND2X2_7329 ( .A(u2__abc_44228_n16052), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16053) );
  AND2X2 AND2X2_733 ( .A(u2__abc_44228_n3428), .B(u2_remHi_51_), .Y(u2__abc_44228_n3429) );
  AND2X2 AND2X2_7330 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_138_), .Y(u2__abc_44228_n16055) );
  AND2X2 AND2X2_7331 ( .A(u2__abc_44228_n2988_bF_buf9), .B(1'b0), .Y(u2__abc_44228_n16056) );
  AND2X2 AND2X2_7332 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_136_), .Y(u2__abc_44228_n16057) );
  AND2X2 AND2X2_7333 ( .A(u2__abc_44228_n16058), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n16059) );
  AND2X2 AND2X2_7334 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_139_), .Y(u2__abc_44228_n16061) );
  AND2X2 AND2X2_7335 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_137_), .Y(u2__abc_44228_n16062) );
  AND2X2 AND2X2_7336 ( .A(u2__abc_44228_n2988_bF_buf8), .B(1'b0), .Y(u2__abc_44228_n16063) );
  AND2X2 AND2X2_7337 ( .A(u2__abc_44228_n16064), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n16065) );
  AND2X2 AND2X2_7338 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_140_), .Y(u2__abc_44228_n16067) );
  AND2X2 AND2X2_7339 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_138_), .Y(u2__abc_44228_n16068) );
  AND2X2 AND2X2_734 ( .A(u2__abc_44228_n3431), .B(sqrto_51_), .Y(u2__abc_44228_n3432) );
  AND2X2 AND2X2_7340 ( .A(u2__abc_44228_n2988_bF_buf7), .B(1'b0), .Y(u2__abc_44228_n16069) );
  AND2X2 AND2X2_7341 ( .A(u2__abc_44228_n16070), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n16071) );
  AND2X2 AND2X2_7342 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_141_), .Y(u2__abc_44228_n16073) );
  AND2X2 AND2X2_7343 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_139_), .Y(u2__abc_44228_n16074) );
  AND2X2 AND2X2_7344 ( .A(u2__abc_44228_n2988_bF_buf6), .B(1'b0), .Y(u2__abc_44228_n16075) );
  AND2X2 AND2X2_7345 ( .A(u2__abc_44228_n16076), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n16077) );
  AND2X2 AND2X2_7346 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_142_), .Y(u2__abc_44228_n16079) );
  AND2X2 AND2X2_7347 ( .A(u2__abc_44228_n2988_bF_buf5), .B(1'b0), .Y(u2__abc_44228_n16080) );
  AND2X2 AND2X2_7348 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_140_), .Y(u2__abc_44228_n16081) );
  AND2X2 AND2X2_7349 ( .A(u2__abc_44228_n16082), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n16083) );
  AND2X2 AND2X2_735 ( .A(u2__abc_44228_n3430), .B(u2__abc_44228_n3433), .Y(u2__abc_44228_n3434) );
  AND2X2 AND2X2_7350 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_143_), .Y(u2__abc_44228_n16085) );
  AND2X2 AND2X2_7351 ( .A(u2__abc_44228_n2988_bF_buf4), .B(1'b0), .Y(u2__abc_44228_n16086) );
  AND2X2 AND2X2_7352 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_141_), .Y(u2__abc_44228_n16087) );
  AND2X2 AND2X2_7353 ( .A(u2__abc_44228_n16088), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n16089) );
  AND2X2 AND2X2_7354 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_144_), .Y(u2__abc_44228_n16091) );
  AND2X2 AND2X2_7355 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_142_), .Y(u2__abc_44228_n16092) );
  AND2X2 AND2X2_7356 ( .A(u2__abc_44228_n2988_bF_buf3), .B(fracta1_0_), .Y(u2__abc_44228_n16093) );
  AND2X2 AND2X2_7357 ( .A(u2__abc_44228_n16094), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16095) );
  AND2X2 AND2X2_7358 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_143_), .Y(u2__abc_44228_n16097) );
  AND2X2 AND2X2_7359 ( .A(u2__abc_44228_n15403_bF_buf0), .B(u2_remLo_145_), .Y(u2__abc_44228_n16098) );
  AND2X2 AND2X2_736 ( .A(u2__abc_44228_n3427), .B(u2__abc_44228_n3434), .Y(u2__abc_44228_n3435) );
  AND2X2 AND2X2_7360 ( .A(u2__abc_44228_n16099), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16100) );
  AND2X2 AND2X2_7361 ( .A(u2__abc_44228_n15402_bF_buf0), .B(u2_remLo_145_), .Y(u2__abc_44228_n16101) );
  AND2X2 AND2X2_7362 ( .A(u2__abc_44228_n2989_bF_buf3), .B(fracta1_1_), .Y(u2__abc_44228_n16102) );
  AND2X2 AND2X2_7363 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_144_), .Y(u2__abc_44228_n16105) );
  AND2X2 AND2X2_7364 ( .A(u2__abc_44228_n15403_bF_buf3), .B(u2_remLo_146_), .Y(u2__abc_44228_n16106) );
  AND2X2 AND2X2_7365 ( .A(u2__abc_44228_n16107), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16108) );
  AND2X2 AND2X2_7366 ( .A(u2__abc_44228_n15402_bF_buf3), .B(u2_remLo_146_), .Y(u2__abc_44228_n16109) );
  AND2X2 AND2X2_7367 ( .A(u2__abc_44228_n2989_bF_buf2), .B(fracta1_2_), .Y(u2__abc_44228_n16110) );
  AND2X2 AND2X2_7368 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_147_), .Y(u2__abc_44228_n16113) );
  AND2X2 AND2X2_7369 ( .A(u2__abc_44228_n2988_bF_buf2), .B(fracta1_3_), .Y(u2__abc_44228_n16114) );
  AND2X2 AND2X2_737 ( .A(u2__abc_44228_n3421), .B(u2__abc_44228_n3435), .Y(u2__abc_44228_n3436) );
  AND2X2 AND2X2_7370 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_145_), .Y(u2__abc_44228_n16115) );
  AND2X2 AND2X2_7371 ( .A(u2__abc_44228_n16116), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16117) );
  AND2X2 AND2X2_7372 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_148_), .Y(u2__abc_44228_n16119) );
  AND2X2 AND2X2_7373 ( .A(u2__abc_44228_n2988_bF_buf1), .B(fracta1_4_), .Y(u2__abc_44228_n16120) );
  AND2X2 AND2X2_7374 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_146_), .Y(u2__abc_44228_n16121) );
  AND2X2 AND2X2_7375 ( .A(u2__abc_44228_n16122), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16123) );
  AND2X2 AND2X2_7376 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_149_), .Y(u2__abc_44228_n16125) );
  AND2X2 AND2X2_7377 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_147_), .Y(u2__abc_44228_n16126) );
  AND2X2 AND2X2_7378 ( .A(u2__abc_44228_n2988_bF_buf0), .B(fracta1_5_), .Y(u2__abc_44228_n16127) );
  AND2X2 AND2X2_7379 ( .A(u2__abc_44228_n16128), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16129) );
  AND2X2 AND2X2_738 ( .A(u2__abc_44228_n3437), .B(u2_remHi_49_), .Y(u2__abc_44228_n3438) );
  AND2X2 AND2X2_7380 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_148_), .Y(u2__abc_44228_n16131) );
  AND2X2 AND2X2_7381 ( .A(u2__abc_44228_n15403_bF_buf2), .B(u2_remLo_150_), .Y(u2__abc_44228_n16132) );
  AND2X2 AND2X2_7382 ( .A(u2__abc_44228_n16133), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16134) );
  AND2X2 AND2X2_7383 ( .A(u2__abc_44228_n15402_bF_buf2), .B(u2_remLo_150_), .Y(u2__abc_44228_n16135) );
  AND2X2 AND2X2_7384 ( .A(u2__abc_44228_n2989_bF_buf1), .B(fracta1_6_), .Y(u2__abc_44228_n16136) );
  AND2X2 AND2X2_7385 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_151_), .Y(u2__abc_44228_n16139) );
  AND2X2 AND2X2_7386 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_149_), .Y(u2__abc_44228_n16140) );
  AND2X2 AND2X2_7387 ( .A(u2__abc_44228_n2988_bF_buf13), .B(fracta1_7_), .Y(u2__abc_44228_n16141) );
  AND2X2 AND2X2_7388 ( .A(u2__abc_44228_n16142), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16143) );
  AND2X2 AND2X2_7389 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_152_), .Y(u2__abc_44228_n16145) );
  AND2X2 AND2X2_739 ( .A(u2__abc_44228_n3440), .B(sqrto_49_), .Y(u2__abc_44228_n3441) );
  AND2X2 AND2X2_7390 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_150_), .Y(u2__abc_44228_n16146) );
  AND2X2 AND2X2_7391 ( .A(u2__abc_44228_n2988_bF_buf12), .B(fracta1_8_), .Y(u2__abc_44228_n16147) );
  AND2X2 AND2X2_7392 ( .A(u2__abc_44228_n16148), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16149) );
  AND2X2 AND2X2_7393 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_153_), .Y(u2__abc_44228_n16151) );
  AND2X2 AND2X2_7394 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_151_), .Y(u2__abc_44228_n16152) );
  AND2X2 AND2X2_7395 ( .A(u2__abc_44228_n2988_bF_buf11), .B(fracta1_9_), .Y(u2__abc_44228_n16153) );
  AND2X2 AND2X2_7396 ( .A(u2__abc_44228_n16154), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n16155) );
  AND2X2 AND2X2_7397 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_154_), .Y(u2__abc_44228_n16157) );
  AND2X2 AND2X2_7398 ( .A(u2__abc_44228_n2988_bF_buf10), .B(fracta1_10_), .Y(u2__abc_44228_n16158) );
  AND2X2 AND2X2_7399 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_152_), .Y(u2__abc_44228_n16159) );
  AND2X2 AND2X2_74 ( .A(_abc_64468_n753_bF_buf10), .B(sqrto_73_), .Y(_auto_iopadmap_cc_313_execute_65414_109_) );
  AND2X2 AND2X2_740 ( .A(u2__abc_44228_n3439_1), .B(u2__abc_44228_n3442), .Y(u2__abc_44228_n3443) );
  AND2X2 AND2X2_7400 ( .A(u2__abc_44228_n16160), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n16161) );
  AND2X2 AND2X2_7401 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_155_), .Y(u2__abc_44228_n16163) );
  AND2X2 AND2X2_7402 ( .A(u2__abc_44228_n2988_bF_buf9), .B(fracta1_11_), .Y(u2__abc_44228_n16164) );
  AND2X2 AND2X2_7403 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_153_), .Y(u2__abc_44228_n16165) );
  AND2X2 AND2X2_7404 ( .A(u2__abc_44228_n16166), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n16167) );
  AND2X2 AND2X2_7405 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_156_), .Y(u2__abc_44228_n16169) );
  AND2X2 AND2X2_7406 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_154_), .Y(u2__abc_44228_n16170) );
  AND2X2 AND2X2_7407 ( .A(u2__abc_44228_n2988_bF_buf8), .B(fracta1_12_), .Y(u2__abc_44228_n16171) );
  AND2X2 AND2X2_7408 ( .A(u2__abc_44228_n16172), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n16173) );
  AND2X2 AND2X2_7409 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_157_), .Y(u2__abc_44228_n16175) );
  AND2X2 AND2X2_741 ( .A(u2__abc_44228_n3444), .B(u2_remHi_48_), .Y(u2__abc_44228_n3445) );
  AND2X2 AND2X2_7410 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_155_), .Y(u2__abc_44228_n16176) );
  AND2X2 AND2X2_7411 ( .A(u2__abc_44228_n2988_bF_buf7), .B(fracta1_13_), .Y(u2__abc_44228_n16177) );
  AND2X2 AND2X2_7412 ( .A(u2__abc_44228_n16178), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n16179) );
  AND2X2 AND2X2_7413 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_158_), .Y(u2__abc_44228_n16181) );
  AND2X2 AND2X2_7414 ( .A(u2__abc_44228_n2988_bF_buf6), .B(fracta1_14_), .Y(u2__abc_44228_n16182) );
  AND2X2 AND2X2_7415 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_156_), .Y(u2__abc_44228_n16183) );
  AND2X2 AND2X2_7416 ( .A(u2__abc_44228_n16184), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n16185) );
  AND2X2 AND2X2_7417 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_159_), .Y(u2__abc_44228_n16187) );
  AND2X2 AND2X2_7418 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_157_), .Y(u2__abc_44228_n16188) );
  AND2X2 AND2X2_7419 ( .A(u2__abc_44228_n2988_bF_buf5), .B(fracta1_15_), .Y(u2__abc_44228_n16189) );
  AND2X2 AND2X2_742 ( .A(u2__abc_44228_n3446), .B(sqrto_48_), .Y(u2__abc_44228_n3447) );
  AND2X2 AND2X2_7420 ( .A(u2__abc_44228_n16190), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16191) );
  AND2X2 AND2X2_7421 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_160_), .Y(u2__abc_44228_n16193) );
  AND2X2 AND2X2_7422 ( .A(u2__abc_44228_n2988_bF_buf4), .B(fracta1_16_), .Y(u2__abc_44228_n16194) );
  AND2X2 AND2X2_7423 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_158_), .Y(u2__abc_44228_n16195) );
  AND2X2 AND2X2_7424 ( .A(u2__abc_44228_n16196), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16197) );
  AND2X2 AND2X2_7425 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_161_), .Y(u2__abc_44228_n16199) );
  AND2X2 AND2X2_7426 ( .A(u2__abc_44228_n2988_bF_buf3), .B(fracta1_17_), .Y(u2__abc_44228_n16200) );
  AND2X2 AND2X2_7427 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_159_), .Y(u2__abc_44228_n16201) );
  AND2X2 AND2X2_7428 ( .A(u2__abc_44228_n16202), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16203) );
  AND2X2 AND2X2_7429 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_162_), .Y(u2__abc_44228_n16205) );
  AND2X2 AND2X2_743 ( .A(u2__abc_44228_n3449_1), .B(u2__abc_44228_n3443), .Y(u2__abc_44228_n3450) );
  AND2X2 AND2X2_7430 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_160_), .Y(u2__abc_44228_n16206) );
  AND2X2 AND2X2_7431 ( .A(u2__abc_44228_n2988_bF_buf2), .B(fracta1_18_), .Y(u2__abc_44228_n16207) );
  AND2X2 AND2X2_7432 ( .A(u2__abc_44228_n16208), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16209) );
  AND2X2 AND2X2_7433 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_163_), .Y(u2__abc_44228_n16211) );
  AND2X2 AND2X2_7434 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_161_), .Y(u2__abc_44228_n16212) );
  AND2X2 AND2X2_7435 ( .A(u2__abc_44228_n2988_bF_buf1), .B(fracta1_19_), .Y(u2__abc_44228_n16213) );
  AND2X2 AND2X2_7436 ( .A(u2__abc_44228_n16214), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16215) );
  AND2X2 AND2X2_7437 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_164_), .Y(u2__abc_44228_n16217) );
  AND2X2 AND2X2_7438 ( .A(u2__abc_44228_n2988_bF_buf0), .B(fracta1_20_), .Y(u2__abc_44228_n16218) );
  AND2X2 AND2X2_7439 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_162_), .Y(u2__abc_44228_n16219) );
  AND2X2 AND2X2_744 ( .A(u2__abc_44228_n3451), .B(u2_remHi_47_), .Y(u2__abc_44228_n3452) );
  AND2X2 AND2X2_7440 ( .A(u2__abc_44228_n16220), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16221) );
  AND2X2 AND2X2_7441 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_165_), .Y(u2__abc_44228_n16223) );
  AND2X2 AND2X2_7442 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_163_), .Y(u2__abc_44228_n16224) );
  AND2X2 AND2X2_7443 ( .A(u2__abc_44228_n2988_bF_buf13), .B(fracta1_21_), .Y(u2__abc_44228_n16225) );
  AND2X2 AND2X2_7444 ( .A(u2__abc_44228_n16226), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16227) );
  AND2X2 AND2X2_7445 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_166_), .Y(u2__abc_44228_n16229) );
  AND2X2 AND2X2_7446 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_164_), .Y(u2__abc_44228_n16230) );
  AND2X2 AND2X2_7447 ( .A(u2__abc_44228_n2988_bF_buf12), .B(fracta1_22_), .Y(u2__abc_44228_n16231) );
  AND2X2 AND2X2_7448 ( .A(u2__abc_44228_n16232), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16233) );
  AND2X2 AND2X2_7449 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_167_), .Y(u2__abc_44228_n16235) );
  AND2X2 AND2X2_745 ( .A(u2__abc_44228_n3454), .B(sqrto_47_), .Y(u2__abc_44228_n3455) );
  AND2X2 AND2X2_7450 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_165_), .Y(u2__abc_44228_n16236) );
  AND2X2 AND2X2_7451 ( .A(u2__abc_44228_n2988_bF_buf11), .B(fracta1_23_), .Y(u2__abc_44228_n16237) );
  AND2X2 AND2X2_7452 ( .A(u2__abc_44228_n16238), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16239) );
  AND2X2 AND2X2_7453 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_168_), .Y(u2__abc_44228_n16241) );
  AND2X2 AND2X2_7454 ( .A(u2__abc_44228_n2988_bF_buf10), .B(fracta1_24_), .Y(u2__abc_44228_n16242) );
  AND2X2 AND2X2_7455 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_166_), .Y(u2__abc_44228_n16243) );
  AND2X2 AND2X2_7456 ( .A(u2__abc_44228_n16244), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n16245) );
  AND2X2 AND2X2_7457 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_169_), .Y(u2__abc_44228_n16247) );
  AND2X2 AND2X2_7458 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_167_), .Y(u2__abc_44228_n16248) );
  AND2X2 AND2X2_7459 ( .A(u2__abc_44228_n2988_bF_buf9), .B(fracta1_25_), .Y(u2__abc_44228_n16249) );
  AND2X2 AND2X2_746 ( .A(u2__abc_44228_n3453), .B(u2__abc_44228_n3456), .Y(u2__abc_44228_n3457_1) );
  AND2X2 AND2X2_7460 ( .A(u2__abc_44228_n16250), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n16251) );
  AND2X2 AND2X2_7461 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_170_), .Y(u2__abc_44228_n16253) );
  AND2X2 AND2X2_7462 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_168_), .Y(u2__abc_44228_n16254) );
  AND2X2 AND2X2_7463 ( .A(u2__abc_44228_n2988_bF_buf8), .B(fracta1_26_), .Y(u2__abc_44228_n16255) );
  AND2X2 AND2X2_7464 ( .A(u2__abc_44228_n16256), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n16257) );
  AND2X2 AND2X2_7465 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_171_), .Y(u2__abc_44228_n16259) );
  AND2X2 AND2X2_7466 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_169_), .Y(u2__abc_44228_n16260) );
  AND2X2 AND2X2_7467 ( .A(u2__abc_44228_n2988_bF_buf7), .B(fracta1_27_), .Y(u2__abc_44228_n16261) );
  AND2X2 AND2X2_7468 ( .A(u2__abc_44228_n16262), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n16263) );
  AND2X2 AND2X2_7469 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_172_), .Y(u2__abc_44228_n16265) );
  AND2X2 AND2X2_747 ( .A(u2__abc_44228_n3458), .B(u2_remHi_46_), .Y(u2__abc_44228_n3459) );
  AND2X2 AND2X2_7470 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_170_), .Y(u2__abc_44228_n16266) );
  AND2X2 AND2X2_7471 ( .A(u2__abc_44228_n2988_bF_buf6), .B(fracta1_28_), .Y(u2__abc_44228_n16267) );
  AND2X2 AND2X2_7472 ( .A(u2__abc_44228_n16268), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n16269) );
  AND2X2 AND2X2_7473 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_173_), .Y(u2__abc_44228_n16271) );
  AND2X2 AND2X2_7474 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_171_), .Y(u2__abc_44228_n16272) );
  AND2X2 AND2X2_7475 ( .A(u2__abc_44228_n2988_bF_buf5), .B(fracta1_29_), .Y(u2__abc_44228_n16273) );
  AND2X2 AND2X2_7476 ( .A(u2__abc_44228_n16274), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n16275) );
  AND2X2 AND2X2_7477 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_174_), .Y(u2__abc_44228_n16277) );
  AND2X2 AND2X2_7478 ( .A(u2__abc_44228_n2988_bF_buf4), .B(fracta1_30_), .Y(u2__abc_44228_n16278) );
  AND2X2 AND2X2_7479 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_172_), .Y(u2__abc_44228_n16279) );
  AND2X2 AND2X2_748 ( .A(u2__abc_44228_n3460), .B(sqrto_46_), .Y(u2__abc_44228_n3461) );
  AND2X2 AND2X2_7480 ( .A(u2__abc_44228_n16280), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16281) );
  AND2X2 AND2X2_7481 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_173_), .Y(u2__abc_44228_n16283) );
  AND2X2 AND2X2_7482 ( .A(u2__abc_44228_n15403_bF_buf1), .B(u2_remLo_175_), .Y(u2__abc_44228_n16284) );
  AND2X2 AND2X2_7483 ( .A(u2__abc_44228_n16285), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16286) );
  AND2X2 AND2X2_7484 ( .A(u2__abc_44228_n15402_bF_buf1), .B(u2_remLo_175_), .Y(u2__abc_44228_n16287) );
  AND2X2 AND2X2_7485 ( .A(u2__abc_44228_n2989_bF_buf0), .B(fracta1_31_), .Y(u2__abc_44228_n16288) );
  AND2X2 AND2X2_7486 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_176_), .Y(u2__abc_44228_n16291) );
  AND2X2 AND2X2_7487 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_174_), .Y(u2__abc_44228_n16292) );
  AND2X2 AND2X2_7488 ( .A(u2__abc_44228_n2988_bF_buf3), .B(fracta1_32_), .Y(u2__abc_44228_n16293) );
  AND2X2 AND2X2_7489 ( .A(u2__abc_44228_n16294), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16295) );
  AND2X2 AND2X2_749 ( .A(u2__abc_44228_n3463), .B(u2__abc_44228_n3457_1), .Y(u2__abc_44228_n3464) );
  AND2X2 AND2X2_7490 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_175_), .Y(u2__abc_44228_n16297) );
  AND2X2 AND2X2_7491 ( .A(u2__abc_44228_n15403_bF_buf0), .B(u2_remLo_177_), .Y(u2__abc_44228_n16298) );
  AND2X2 AND2X2_7492 ( .A(u2__abc_44228_n16299), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16300) );
  AND2X2 AND2X2_7493 ( .A(u2__abc_44228_n15402_bF_buf0), .B(u2_remLo_177_), .Y(u2__abc_44228_n16301) );
  AND2X2 AND2X2_7494 ( .A(u2__abc_44228_n2989_bF_buf3), .B(fracta1_33_), .Y(u2__abc_44228_n16302) );
  AND2X2 AND2X2_7495 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_176_), .Y(u2__abc_44228_n16305) );
  AND2X2 AND2X2_7496 ( .A(u2__abc_44228_n15403_bF_buf3), .B(u2_remLo_178_), .Y(u2__abc_44228_n16306) );
  AND2X2 AND2X2_7497 ( .A(u2__abc_44228_n16307), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16308) );
  AND2X2 AND2X2_7498 ( .A(u2__abc_44228_n15402_bF_buf3), .B(u2_remLo_178_), .Y(u2__abc_44228_n16309) );
  AND2X2 AND2X2_7499 ( .A(u2__abc_44228_n2989_bF_buf2), .B(fracta1_34_), .Y(u2__abc_44228_n16310) );
  AND2X2 AND2X2_75 ( .A(_abc_64468_n753_bF_buf9), .B(sqrto_74_), .Y(_auto_iopadmap_cc_313_execute_65414_110_) );
  AND2X2 AND2X2_750 ( .A(u2__abc_44228_n3450), .B(u2__abc_44228_n3464), .Y(u2__abc_44228_n3465) );
  AND2X2 AND2X2_7500 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_179_), .Y(u2__abc_44228_n16313) );
  AND2X2 AND2X2_7501 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_177_), .Y(u2__abc_44228_n16314) );
  AND2X2 AND2X2_7502 ( .A(u2__abc_44228_n2988_bF_buf2), .B(fracta1_35_), .Y(u2__abc_44228_n16315) );
  AND2X2 AND2X2_7503 ( .A(u2__abc_44228_n16316), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16317) );
  AND2X2 AND2X2_7504 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_180_), .Y(u2__abc_44228_n16319) );
  AND2X2 AND2X2_7505 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_178_), .Y(u2__abc_44228_n16320) );
  AND2X2 AND2X2_7506 ( .A(u2__abc_44228_n2988_bF_buf1), .B(fracta1_36_), .Y(u2__abc_44228_n16321) );
  AND2X2 AND2X2_7507 ( .A(u2__abc_44228_n16322), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16323) );
  AND2X2 AND2X2_7508 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_181_), .Y(u2__abc_44228_n16325) );
  AND2X2 AND2X2_7509 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_179_), .Y(u2__abc_44228_n16326) );
  AND2X2 AND2X2_751 ( .A(u2__abc_44228_n3436), .B(u2__abc_44228_n3465), .Y(u2__abc_44228_n3466) );
  AND2X2 AND2X2_7510 ( .A(u2__abc_44228_n2988_bF_buf0), .B(fracta1_37_), .Y(u2__abc_44228_n16327) );
  AND2X2 AND2X2_7511 ( .A(u2__abc_44228_n16328), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16329) );
  AND2X2 AND2X2_7512 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_180_), .Y(u2__abc_44228_n16331) );
  AND2X2 AND2X2_7513 ( .A(u2__abc_44228_n15403_bF_buf2), .B(u2_remLo_182_), .Y(u2__abc_44228_n16332) );
  AND2X2 AND2X2_7514 ( .A(u2__abc_44228_n16333), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16334) );
  AND2X2 AND2X2_7515 ( .A(u2__abc_44228_n15402_bF_buf2), .B(u2_remLo_182_), .Y(u2__abc_44228_n16335) );
  AND2X2 AND2X2_7516 ( .A(u2__abc_44228_n2989_bF_buf1), .B(fracta1_38_), .Y(u2__abc_44228_n16336) );
  AND2X2 AND2X2_7517 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_183_), .Y(u2__abc_44228_n16339) );
  AND2X2 AND2X2_7518 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_181_), .Y(u2__abc_44228_n16340) );
  AND2X2 AND2X2_7519 ( .A(u2__abc_44228_n2988_bF_buf13), .B(fracta1_39_), .Y(u2__abc_44228_n16341) );
  AND2X2 AND2X2_752 ( .A(u2__abc_44228_n3407), .B(u2__abc_44228_n3466), .Y(u2__abc_44228_n3467_1) );
  AND2X2 AND2X2_7520 ( .A(u2__abc_44228_n16342), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n16343) );
  AND2X2 AND2X2_7521 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_184_), .Y(u2__abc_44228_n16345) );
  AND2X2 AND2X2_7522 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_182_), .Y(u2__abc_44228_n16346) );
  AND2X2 AND2X2_7523 ( .A(u2__abc_44228_n2988_bF_buf12), .B(fracta1_40_), .Y(u2__abc_44228_n16347) );
  AND2X2 AND2X2_7524 ( .A(u2__abc_44228_n16348), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n16349) );
  AND2X2 AND2X2_7525 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_185_), .Y(u2__abc_44228_n16351) );
  AND2X2 AND2X2_7526 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_183_), .Y(u2__abc_44228_n16352) );
  AND2X2 AND2X2_7527 ( .A(u2__abc_44228_n2988_bF_buf11), .B(fracta1_41_), .Y(u2__abc_44228_n16353) );
  AND2X2 AND2X2_7528 ( .A(u2__abc_44228_n16354), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n16355) );
  AND2X2 AND2X2_7529 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_186_), .Y(u2__abc_44228_n16357) );
  AND2X2 AND2X2_753 ( .A(u2__abc_44228_n3468), .B(u2_remHi_45_), .Y(u2__abc_44228_n3469) );
  AND2X2 AND2X2_7530 ( .A(u2__abc_44228_n2988_bF_buf10), .B(fracta1_42_), .Y(u2__abc_44228_n16358) );
  AND2X2 AND2X2_7531 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_184_), .Y(u2__abc_44228_n16359) );
  AND2X2 AND2X2_7532 ( .A(u2__abc_44228_n16360), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n16361) );
  AND2X2 AND2X2_7533 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_187_), .Y(u2__abc_44228_n16363) );
  AND2X2 AND2X2_7534 ( .A(u2__abc_44228_n2988_bF_buf9), .B(fracta1_43_), .Y(u2__abc_44228_n16364) );
  AND2X2 AND2X2_7535 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_185_), .Y(u2__abc_44228_n16365) );
  AND2X2 AND2X2_7536 ( .A(u2__abc_44228_n16366), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n16367) );
  AND2X2 AND2X2_7537 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_188_), .Y(u2__abc_44228_n16369) );
  AND2X2 AND2X2_7538 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_186_), .Y(u2__abc_44228_n16370) );
  AND2X2 AND2X2_7539 ( .A(u2__abc_44228_n2988_bF_buf8), .B(fracta1_44_), .Y(u2__abc_44228_n16371) );
  AND2X2 AND2X2_754 ( .A(u2__abc_44228_n3471), .B(sqrto_45_), .Y(u2__abc_44228_n3472) );
  AND2X2 AND2X2_7540 ( .A(u2__abc_44228_n16372), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n16373) );
  AND2X2 AND2X2_7541 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_189_), .Y(u2__abc_44228_n16375) );
  AND2X2 AND2X2_7542 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_187_), .Y(u2__abc_44228_n16376) );
  AND2X2 AND2X2_7543 ( .A(u2__abc_44228_n2988_bF_buf7), .B(fracta1_45_), .Y(u2__abc_44228_n16377) );
  AND2X2 AND2X2_7544 ( .A(u2__abc_44228_n16378), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16379) );
  AND2X2 AND2X2_7545 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_190_), .Y(u2__abc_44228_n16381) );
  AND2X2 AND2X2_7546 ( .A(u2__abc_44228_n2988_bF_buf6), .B(fracta1_46_), .Y(u2__abc_44228_n16382) );
  AND2X2 AND2X2_7547 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_188_), .Y(u2__abc_44228_n16383) );
  AND2X2 AND2X2_7548 ( .A(u2__abc_44228_n16384), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16385) );
  AND2X2 AND2X2_7549 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_191_), .Y(u2__abc_44228_n16387) );
  AND2X2 AND2X2_755 ( .A(u2__abc_44228_n3470), .B(u2__abc_44228_n3473), .Y(u2__abc_44228_n3474) );
  AND2X2 AND2X2_7550 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_189_), .Y(u2__abc_44228_n16388) );
  AND2X2 AND2X2_7551 ( .A(u2__abc_44228_n2988_bF_buf5), .B(fracta1_47_), .Y(u2__abc_44228_n16389) );
  AND2X2 AND2X2_7552 ( .A(u2__abc_44228_n16390), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16391) );
  AND2X2 AND2X2_7553 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_192_), .Y(u2__abc_44228_n16393) );
  AND2X2 AND2X2_7554 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_190_), .Y(u2__abc_44228_n16394) );
  AND2X2 AND2X2_7555 ( .A(u2__abc_44228_n2988_bF_buf4), .B(fracta1_48_), .Y(u2__abc_44228_n16395) );
  AND2X2 AND2X2_7556 ( .A(u2__abc_44228_n16396), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16397) );
  AND2X2 AND2X2_7557 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_193_), .Y(u2__abc_44228_n16399) );
  AND2X2 AND2X2_7558 ( .A(u2__abc_44228_n2988_bF_buf3), .B(fracta1_49_), .Y(u2__abc_44228_n16400) );
  AND2X2 AND2X2_7559 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_191_), .Y(u2__abc_44228_n16401) );
  AND2X2 AND2X2_756 ( .A(u2__abc_44228_n3475_1), .B(u2_remHi_44_), .Y(u2__abc_44228_n3476) );
  AND2X2 AND2X2_7560 ( .A(u2__abc_44228_n16402), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16403) );
  AND2X2 AND2X2_7561 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_194_), .Y(u2__abc_44228_n16405) );
  AND2X2 AND2X2_7562 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_192_), .Y(u2__abc_44228_n16406) );
  AND2X2 AND2X2_7563 ( .A(u2__abc_44228_n2988_bF_buf2), .B(fracta1_50_), .Y(u2__abc_44228_n16407) );
  AND2X2 AND2X2_7564 ( .A(u2__abc_44228_n16408), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16409) );
  AND2X2 AND2X2_7565 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_195_), .Y(u2__abc_44228_n16411) );
  AND2X2 AND2X2_7566 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_193_), .Y(u2__abc_44228_n16412) );
  AND2X2 AND2X2_7567 ( .A(u2__abc_44228_n2988_bF_buf1), .B(fracta1_51_), .Y(u2__abc_44228_n16413) );
  AND2X2 AND2X2_7568 ( .A(u2__abc_44228_n16414), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16415) );
  AND2X2 AND2X2_7569 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_196_), .Y(u2__abc_44228_n16417) );
  AND2X2 AND2X2_757 ( .A(u2__abc_44228_n3477), .B(sqrto_44_), .Y(u2__abc_44228_n3478) );
  AND2X2 AND2X2_7570 ( .A(u2__abc_44228_n2988_bF_buf0), .B(fracta1_52_), .Y(u2__abc_44228_n16418) );
  AND2X2 AND2X2_7571 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_194_), .Y(u2__abc_44228_n16419) );
  AND2X2 AND2X2_7572 ( .A(u2__abc_44228_n16420), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16421) );
  AND2X2 AND2X2_7573 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_197_), .Y(u2__abc_44228_n16423) );
  AND2X2 AND2X2_7574 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_195_), .Y(u2__abc_44228_n16424) );
  AND2X2 AND2X2_7575 ( .A(u2__abc_44228_n2988_bF_buf13), .B(fracta1_53_), .Y(u2__abc_44228_n16425) );
  AND2X2 AND2X2_7576 ( .A(u2__abc_44228_n16426), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16427) );
  AND2X2 AND2X2_7577 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_198_), .Y(u2__abc_44228_n16429) );
  AND2X2 AND2X2_7578 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_196_), .Y(u2__abc_44228_n16430) );
  AND2X2 AND2X2_7579 ( .A(u2__abc_44228_n2988_bF_buf12), .B(fracta1_54_), .Y(u2__abc_44228_n16431) );
  AND2X2 AND2X2_758 ( .A(u2__abc_44228_n3480), .B(u2__abc_44228_n3474), .Y(u2__abc_44228_n3481) );
  AND2X2 AND2X2_7580 ( .A(u2__abc_44228_n16432), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n16433) );
  AND2X2 AND2X2_7581 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_199_), .Y(u2__abc_44228_n16435) );
  AND2X2 AND2X2_7582 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_197_), .Y(u2__abc_44228_n16436) );
  AND2X2 AND2X2_7583 ( .A(u2__abc_44228_n2988_bF_buf11), .B(fracta1_55_), .Y(u2__abc_44228_n16437) );
  AND2X2 AND2X2_7584 ( .A(u2__abc_44228_n16438), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n16439) );
  AND2X2 AND2X2_7585 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_200_), .Y(u2__abc_44228_n16441) );
  AND2X2 AND2X2_7586 ( .A(u2__abc_44228_n2988_bF_buf10), .B(fracta1_56_), .Y(u2__abc_44228_n16442) );
  AND2X2 AND2X2_7587 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_198_), .Y(u2__abc_44228_n16443) );
  AND2X2 AND2X2_7588 ( .A(u2__abc_44228_n16444), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n16445) );
  AND2X2 AND2X2_7589 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_201_), .Y(u2__abc_44228_n16447) );
  AND2X2 AND2X2_759 ( .A(u2__abc_44228_n3482), .B(u2_remHi_42_), .Y(u2__abc_44228_n3483) );
  AND2X2 AND2X2_7590 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_199_), .Y(u2__abc_44228_n16448) );
  AND2X2 AND2X2_7591 ( .A(u2__abc_44228_n2988_bF_buf9), .B(fracta1_57_), .Y(u2__abc_44228_n16449) );
  AND2X2 AND2X2_7592 ( .A(u2__abc_44228_n16450), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n16451) );
  AND2X2 AND2X2_7593 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_202_), .Y(u2__abc_44228_n16453) );
  AND2X2 AND2X2_7594 ( .A(u2__abc_44228_n2988_bF_buf8), .B(fracta1_58_), .Y(u2__abc_44228_n16454) );
  AND2X2 AND2X2_7595 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_200_), .Y(u2__abc_44228_n16455) );
  AND2X2 AND2X2_7596 ( .A(u2__abc_44228_n16456), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n16457) );
  AND2X2 AND2X2_7597 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_203_), .Y(u2__abc_44228_n16459) );
  AND2X2 AND2X2_7598 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_201_), .Y(u2__abc_44228_n16460) );
  AND2X2 AND2X2_7599 ( .A(u2__abc_44228_n2988_bF_buf7), .B(fracta1_59_), .Y(u2__abc_44228_n16461) );
  AND2X2 AND2X2_76 ( .A(_abc_64468_n753_bF_buf8), .B(sqrto_75_), .Y(_auto_iopadmap_cc_313_execute_65414_111_) );
  AND2X2 AND2X2_760 ( .A(u2__abc_44228_n3484_1), .B(sqrto_42_), .Y(u2__abc_44228_n3485) );
  AND2X2 AND2X2_7600 ( .A(u2__abc_44228_n16462), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n16463) );
  AND2X2 AND2X2_7601 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_204_), .Y(u2__abc_44228_n16465) );
  AND2X2 AND2X2_7602 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_202_), .Y(u2__abc_44228_n16466) );
  AND2X2 AND2X2_7603 ( .A(u2__abc_44228_n2988_bF_buf6), .B(fracta1_60_), .Y(u2__abc_44228_n16467) );
  AND2X2 AND2X2_7604 ( .A(u2__abc_44228_n16468), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16469) );
  AND2X2 AND2X2_7605 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_205_), .Y(u2__abc_44228_n16471) );
  AND2X2 AND2X2_7606 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_203_), .Y(u2__abc_44228_n16472) );
  AND2X2 AND2X2_7607 ( .A(u2__abc_44228_n2988_bF_buf5), .B(fracta1_61_), .Y(u2__abc_44228_n16473) );
  AND2X2 AND2X2_7608 ( .A(u2__abc_44228_n16474), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16475) );
  AND2X2 AND2X2_7609 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_206_), .Y(u2__abc_44228_n16477) );
  AND2X2 AND2X2_761 ( .A(u2__abc_44228_n3488), .B(u2_remHi_43_), .Y(u2__abc_44228_n3489) );
  AND2X2 AND2X2_7610 ( .A(u2__abc_44228_n2988_bF_buf4), .B(fracta1_62_), .Y(u2__abc_44228_n16478) );
  AND2X2 AND2X2_7611 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_204_), .Y(u2__abc_44228_n16479) );
  AND2X2 AND2X2_7612 ( .A(u2__abc_44228_n16480), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16481) );
  AND2X2 AND2X2_7613 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_207_), .Y(u2__abc_44228_n16483) );
  AND2X2 AND2X2_7614 ( .A(u2__abc_44228_n2988_bF_buf3), .B(fracta1_63_), .Y(u2__abc_44228_n16484) );
  AND2X2 AND2X2_7615 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_205_), .Y(u2__abc_44228_n16485) );
  AND2X2 AND2X2_7616 ( .A(u2__abc_44228_n16486), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16487) );
  AND2X2 AND2X2_7617 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_208_), .Y(u2__abc_44228_n16489) );
  AND2X2 AND2X2_7618 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_206_), .Y(u2__abc_44228_n16490) );
  AND2X2 AND2X2_7619 ( .A(u2__abc_44228_n2988_bF_buf2), .B(fracta1_64_), .Y(u2__abc_44228_n16491) );
  AND2X2 AND2X2_762 ( .A(u2__abc_44228_n3491), .B(sqrto_43_), .Y(u2__abc_44228_n3492) );
  AND2X2 AND2X2_7620 ( .A(u2__abc_44228_n16492), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16493) );
  AND2X2 AND2X2_7621 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_209_), .Y(u2__abc_44228_n16495) );
  AND2X2 AND2X2_7622 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_207_), .Y(u2__abc_44228_n16496) );
  AND2X2 AND2X2_7623 ( .A(u2__abc_44228_n2988_bF_buf1), .B(fracta1_65_), .Y(u2__abc_44228_n16497) );
  AND2X2 AND2X2_7624 ( .A(u2__abc_44228_n16498), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16499) );
  AND2X2 AND2X2_7625 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_208_), .Y(u2__abc_44228_n16501) );
  AND2X2 AND2X2_7626 ( .A(u2__abc_44228_n15403_bF_buf1), .B(u2_remLo_210_), .Y(u2__abc_44228_n16502) );
  AND2X2 AND2X2_7627 ( .A(u2__abc_44228_n16503), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16504) );
  AND2X2 AND2X2_7628 ( .A(u2__abc_44228_n15402_bF_buf1), .B(u2_remLo_210_), .Y(u2__abc_44228_n16505) );
  AND2X2 AND2X2_7629 ( .A(u2__abc_44228_n2989_bF_buf0), .B(fracta1_66_), .Y(u2__abc_44228_n16506) );
  AND2X2 AND2X2_763 ( .A(u2__abc_44228_n3490), .B(u2__abc_44228_n3493), .Y(u2__abc_44228_n3494) );
  AND2X2 AND2X2_7630 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_211_), .Y(u2__abc_44228_n16509) );
  AND2X2 AND2X2_7631 ( .A(u2__abc_44228_n2988_bF_buf0), .B(fracta1_67_), .Y(u2__abc_44228_n16510) );
  AND2X2 AND2X2_7632 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_209_), .Y(u2__abc_44228_n16511) );
  AND2X2 AND2X2_7633 ( .A(u2__abc_44228_n16512), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16513) );
  AND2X2 AND2X2_7634 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_212_), .Y(u2__abc_44228_n16515) );
  AND2X2 AND2X2_7635 ( .A(u2__abc_44228_n2988_bF_buf13), .B(fracta1_68_), .Y(u2__abc_44228_n16516) );
  AND2X2 AND2X2_7636 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_210_), .Y(u2__abc_44228_n16517) );
  AND2X2 AND2X2_7637 ( .A(u2__abc_44228_n16518), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16519) );
  AND2X2 AND2X2_7638 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_213_), .Y(u2__abc_44228_n16521) );
  AND2X2 AND2X2_7639 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_211_), .Y(u2__abc_44228_n16522) );
  AND2X2 AND2X2_764 ( .A(u2__abc_44228_n3487), .B(u2__abc_44228_n3494), .Y(u2__abc_44228_n3495_1) );
  AND2X2 AND2X2_7640 ( .A(u2__abc_44228_n2988_bF_buf12), .B(fracta1_69_), .Y(u2__abc_44228_n16523) );
  AND2X2 AND2X2_7641 ( .A(u2__abc_44228_n16524), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n16525) );
  AND2X2 AND2X2_7642 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_212_), .Y(u2__abc_44228_n16527) );
  AND2X2 AND2X2_7643 ( .A(u2__abc_44228_n15403_bF_buf0), .B(u2_remLo_214_), .Y(u2__abc_44228_n16528) );
  AND2X2 AND2X2_7644 ( .A(u2__abc_44228_n16529), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n16530) );
  AND2X2 AND2X2_7645 ( .A(u2__abc_44228_n15402_bF_buf0), .B(u2_remLo_214_), .Y(u2__abc_44228_n16531) );
  AND2X2 AND2X2_7646 ( .A(u2__abc_44228_n2989_bF_buf3), .B(fracta1_70_), .Y(u2__abc_44228_n16532) );
  AND2X2 AND2X2_7647 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_215_), .Y(u2__abc_44228_n16535) );
  AND2X2 AND2X2_7648 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_213_), .Y(u2__abc_44228_n16536) );
  AND2X2 AND2X2_7649 ( .A(u2__abc_44228_n2988_bF_buf11), .B(fracta1_71_), .Y(u2__abc_44228_n16537) );
  AND2X2 AND2X2_765 ( .A(u2__abc_44228_n3481), .B(u2__abc_44228_n3495_1), .Y(u2__abc_44228_n3496) );
  AND2X2 AND2X2_7650 ( .A(u2__abc_44228_n16538), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n16539) );
  AND2X2 AND2X2_7651 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_216_), .Y(u2__abc_44228_n16541) );
  AND2X2 AND2X2_7652 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_214_), .Y(u2__abc_44228_n16542) );
  AND2X2 AND2X2_7653 ( .A(u2__abc_44228_n2988_bF_buf10), .B(fracta1_72_), .Y(u2__abc_44228_n16543) );
  AND2X2 AND2X2_7654 ( .A(u2__abc_44228_n16544), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n16545) );
  AND2X2 AND2X2_7655 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_217_), .Y(u2__abc_44228_n16547) );
  AND2X2 AND2X2_7656 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_215_), .Y(u2__abc_44228_n16548) );
  AND2X2 AND2X2_7657 ( .A(u2__abc_44228_n2988_bF_buf9), .B(fracta1_73_), .Y(u2__abc_44228_n16549) );
  AND2X2 AND2X2_7658 ( .A(u2__abc_44228_n16550), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n16551) );
  AND2X2 AND2X2_7659 ( .A(u2__abc_44228_n15403_bF_buf3), .B(u2_remLo_218_), .Y(u2__abc_44228_n16553) );
  AND2X2 AND2X2_766 ( .A(u2__abc_44228_n3497), .B(u2_remHi_39_), .Y(u2__abc_44228_n3498) );
  AND2X2 AND2X2_7660 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_216_), .Y(u2__abc_44228_n16554) );
  AND2X2 AND2X2_7661 ( .A(u2__abc_44228_n16555), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n16556) );
  AND2X2 AND2X2_7662 ( .A(u2__abc_44228_n15402_bF_buf3), .B(u2_remLo_218_), .Y(u2__abc_44228_n16557) );
  AND2X2 AND2X2_7663 ( .A(u2__abc_44228_n2989_bF_buf2), .B(fracta1_74_), .Y(u2__abc_44228_n16558) );
  AND2X2 AND2X2_7664 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_219_), .Y(u2__abc_44228_n16561) );
  AND2X2 AND2X2_7665 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_217_), .Y(u2__abc_44228_n16562) );
  AND2X2 AND2X2_7666 ( .A(u2__abc_44228_n2988_bF_buf8), .B(fracta1_75_), .Y(u2__abc_44228_n16563) );
  AND2X2 AND2X2_7667 ( .A(u2__abc_44228_n16564), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16565) );
  AND2X2 AND2X2_7668 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_220_), .Y(u2__abc_44228_n16567) );
  AND2X2 AND2X2_7669 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_218_), .Y(u2__abc_44228_n16568) );
  AND2X2 AND2X2_767 ( .A(u2__abc_44228_n3500), .B(sqrto_39_), .Y(u2__abc_44228_n3501) );
  AND2X2 AND2X2_7670 ( .A(u2__abc_44228_n2988_bF_buf7), .B(fracta1_76_), .Y(u2__abc_44228_n16569) );
  AND2X2 AND2X2_7671 ( .A(u2__abc_44228_n16570), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16571) );
  AND2X2 AND2X2_7672 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_221_), .Y(u2__abc_44228_n16573) );
  AND2X2 AND2X2_7673 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_219_), .Y(u2__abc_44228_n16574) );
  AND2X2 AND2X2_7674 ( .A(u2__abc_44228_n2988_bF_buf6), .B(fracta1_77_), .Y(u2__abc_44228_n16575) );
  AND2X2 AND2X2_7675 ( .A(u2__abc_44228_n16576), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16577) );
  AND2X2 AND2X2_7676 ( .A(u2__abc_44228_n15403_bF_buf2), .B(u2_remLo_222_), .Y(u2__abc_44228_n16579) );
  AND2X2 AND2X2_7677 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_220_), .Y(u2__abc_44228_n16580) );
  AND2X2 AND2X2_7678 ( .A(u2__abc_44228_n16581), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16582) );
  AND2X2 AND2X2_7679 ( .A(u2__abc_44228_n15402_bF_buf2), .B(u2_remLo_222_), .Y(u2__abc_44228_n16583) );
  AND2X2 AND2X2_768 ( .A(u2__abc_44228_n3499), .B(u2__abc_44228_n3502), .Y(u2__abc_44228_n3503) );
  AND2X2 AND2X2_7680 ( .A(u2__abc_44228_n2989_bF_buf1), .B(fracta1_78_), .Y(u2__abc_44228_n16584) );
  AND2X2 AND2X2_7681 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_223_), .Y(u2__abc_44228_n16587) );
  AND2X2 AND2X2_7682 ( .A(u2__abc_44228_n2988_bF_buf5), .B(fracta1_79_), .Y(u2__abc_44228_n16588) );
  AND2X2 AND2X2_7683 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_221_), .Y(u2__abc_44228_n16589) );
  AND2X2 AND2X2_7684 ( .A(u2__abc_44228_n16590), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16591) );
  AND2X2 AND2X2_7685 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_224_), .Y(u2__abc_44228_n16593) );
  AND2X2 AND2X2_7686 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_222_), .Y(u2__abc_44228_n16594) );
  AND2X2 AND2X2_7687 ( .A(u2__abc_44228_n2988_bF_buf4), .B(fracta1_80_), .Y(u2__abc_44228_n16595) );
  AND2X2 AND2X2_7688 ( .A(u2__abc_44228_n16596), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16597) );
  AND2X2 AND2X2_7689 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_225_), .Y(u2__abc_44228_n16599) );
  AND2X2 AND2X2_769 ( .A(u2__abc_44228_n3504), .B(u2_remHi_38_), .Y(u2__abc_44228_n3505_1) );
  AND2X2 AND2X2_7690 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_223_), .Y(u2__abc_44228_n16600) );
  AND2X2 AND2X2_7691 ( .A(u2__abc_44228_n2988_bF_buf3), .B(fracta1_81_), .Y(u2__abc_44228_n16601) );
  AND2X2 AND2X2_7692 ( .A(u2__abc_44228_n16602), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16603) );
  AND2X2 AND2X2_7693 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_226_), .Y(u2__abc_44228_n16605) );
  AND2X2 AND2X2_7694 ( .A(u2__abc_44228_n2988_bF_buf2), .B(fracta1_82_), .Y(u2__abc_44228_n16606) );
  AND2X2 AND2X2_7695 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_224_), .Y(u2__abc_44228_n16607) );
  AND2X2 AND2X2_7696 ( .A(u2__abc_44228_n16608), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16609) );
  AND2X2 AND2X2_7697 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_227_), .Y(u2__abc_44228_n16611) );
  AND2X2 AND2X2_7698 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_225_), .Y(u2__abc_44228_n16612) );
  AND2X2 AND2X2_7699 ( .A(u2__abc_44228_n2988_bF_buf1), .B(fracta1_83_), .Y(u2__abc_44228_n16613) );
  AND2X2 AND2X2_77 ( .A(_abc_64468_n831_1), .B(_abc_64468_n830), .Y(_auto_iopadmap_cc_313_execute_65414_112_) );
  AND2X2 AND2X2_770 ( .A(u2__abc_44228_n3506), .B(sqrto_38_), .Y(u2__abc_44228_n3507) );
  AND2X2 AND2X2_7700 ( .A(u2__abc_44228_n16614), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16615) );
  AND2X2 AND2X2_7701 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_228_), .Y(u2__abc_44228_n16617) );
  AND2X2 AND2X2_7702 ( .A(u2__abc_44228_n2988_bF_buf0), .B(fracta1_84_), .Y(u2__abc_44228_n16618) );
  AND2X2 AND2X2_7703 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_226_), .Y(u2__abc_44228_n16619) );
  AND2X2 AND2X2_7704 ( .A(u2__abc_44228_n16620), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n16621) );
  AND2X2 AND2X2_7705 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_229_), .Y(u2__abc_44228_n16623) );
  AND2X2 AND2X2_7706 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_227_), .Y(u2__abc_44228_n16624) );
  AND2X2 AND2X2_7707 ( .A(u2__abc_44228_n2988_bF_buf13), .B(fracta1_85_), .Y(u2__abc_44228_n16625) );
  AND2X2 AND2X2_7708 ( .A(u2__abc_44228_n16626), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n16627) );
  AND2X2 AND2X2_7709 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_230_), .Y(u2__abc_44228_n16629) );
  AND2X2 AND2X2_771 ( .A(u2__abc_44228_n3509), .B(u2__abc_44228_n3503), .Y(u2__abc_44228_n3510) );
  AND2X2 AND2X2_7710 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_228_), .Y(u2__abc_44228_n16630) );
  AND2X2 AND2X2_7711 ( .A(u2__abc_44228_n2988_bF_buf12), .B(fracta1_86_), .Y(u2__abc_44228_n16631) );
  AND2X2 AND2X2_7712 ( .A(u2__abc_44228_n16632), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n16633) );
  AND2X2 AND2X2_7713 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_231_), .Y(u2__abc_44228_n16635) );
  AND2X2 AND2X2_7714 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_229_), .Y(u2__abc_44228_n16636) );
  AND2X2 AND2X2_7715 ( .A(u2__abc_44228_n2988_bF_buf11), .B(fracta1_87_), .Y(u2__abc_44228_n16637) );
  AND2X2 AND2X2_7716 ( .A(u2__abc_44228_n16638), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n16639) );
  AND2X2 AND2X2_7717 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_232_), .Y(u2__abc_44228_n16641) );
  AND2X2 AND2X2_7718 ( .A(u2__abc_44228_n2988_bF_buf10), .B(fracta1_88_), .Y(u2__abc_44228_n16642) );
  AND2X2 AND2X2_7719 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_230_), .Y(u2__abc_44228_n16643) );
  AND2X2 AND2X2_772 ( .A(u2__abc_44228_n3511), .B(u2_remHi_41_), .Y(u2__abc_44228_n3512) );
  AND2X2 AND2X2_7720 ( .A(u2__abc_44228_n16644), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n16645) );
  AND2X2 AND2X2_7721 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_233_), .Y(u2__abc_44228_n16647) );
  AND2X2 AND2X2_7722 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_231_), .Y(u2__abc_44228_n16648) );
  AND2X2 AND2X2_7723 ( .A(u2__abc_44228_n2988_bF_buf9), .B(fracta1_89_), .Y(u2__abc_44228_n16649) );
  AND2X2 AND2X2_7724 ( .A(u2__abc_44228_n16650), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n16651) );
  AND2X2 AND2X2_7725 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_234_), .Y(u2__abc_44228_n16653) );
  AND2X2 AND2X2_7726 ( .A(u2__abc_44228_n2988_bF_buf8), .B(fracta1_90_), .Y(u2__abc_44228_n16654) );
  AND2X2 AND2X2_7727 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_232_), .Y(u2__abc_44228_n16655) );
  AND2X2 AND2X2_7728 ( .A(u2__abc_44228_n16656), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16657) );
  AND2X2 AND2X2_7729 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_235_), .Y(u2__abc_44228_n16659) );
  AND2X2 AND2X2_773 ( .A(u2__abc_44228_n3514), .B(sqrto_41_), .Y(u2__abc_44228_n3515) );
  AND2X2 AND2X2_7730 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_233_), .Y(u2__abc_44228_n16660) );
  AND2X2 AND2X2_7731 ( .A(u2__abc_44228_n2988_bF_buf7), .B(fracta1_91_), .Y(u2__abc_44228_n16661) );
  AND2X2 AND2X2_7732 ( .A(u2__abc_44228_n16662), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16663) );
  AND2X2 AND2X2_7733 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_236_), .Y(u2__abc_44228_n16665) );
  AND2X2 AND2X2_7734 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_234_), .Y(u2__abc_44228_n16666) );
  AND2X2 AND2X2_7735 ( .A(u2__abc_44228_n2988_bF_buf6), .B(fracta1_92_), .Y(u2__abc_44228_n16667) );
  AND2X2 AND2X2_7736 ( .A(u2__abc_44228_n16668), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16669) );
  AND2X2 AND2X2_7737 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_237_), .Y(u2__abc_44228_n16671) );
  AND2X2 AND2X2_7738 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_235_), .Y(u2__abc_44228_n16672) );
  AND2X2 AND2X2_7739 ( .A(u2__abc_44228_n2988_bF_buf5), .B(fracta1_93_), .Y(u2__abc_44228_n16673) );
  AND2X2 AND2X2_774 ( .A(u2__abc_44228_n3513_1), .B(u2__abc_44228_n3516), .Y(u2__abc_44228_n3517) );
  AND2X2 AND2X2_7740 ( .A(u2__abc_44228_n16674), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16675) );
  AND2X2 AND2X2_7741 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_238_), .Y(u2__abc_44228_n16677) );
  AND2X2 AND2X2_7742 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_236_), .Y(u2__abc_44228_n16678) );
  AND2X2 AND2X2_7743 ( .A(u2__abc_44228_n2988_bF_buf4), .B(fracta1_94_), .Y(u2__abc_44228_n16679) );
  AND2X2 AND2X2_7744 ( .A(u2__abc_44228_n16680), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16681) );
  AND2X2 AND2X2_7745 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_239_), .Y(u2__abc_44228_n16683) );
  AND2X2 AND2X2_7746 ( .A(u2__abc_44228_n2988_bF_buf3), .B(fracta1_95_), .Y(u2__abc_44228_n16684) );
  AND2X2 AND2X2_7747 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_237_), .Y(u2__abc_44228_n16685) );
  AND2X2 AND2X2_7748 ( .A(u2__abc_44228_n16686), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16687) );
  AND2X2 AND2X2_7749 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_240_), .Y(u2__abc_44228_n16689) );
  AND2X2 AND2X2_775 ( .A(u2__abc_44228_n3518), .B(u2_remHi_40_), .Y(u2__abc_44228_n3519) );
  AND2X2 AND2X2_7750 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_238_), .Y(u2__abc_44228_n16690) );
  AND2X2 AND2X2_7751 ( .A(u2__abc_44228_n2988_bF_buf2), .B(fracta1_96_), .Y(u2__abc_44228_n16691) );
  AND2X2 AND2X2_7752 ( .A(u2__abc_44228_n16692), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16693) );
  AND2X2 AND2X2_7753 ( .A(u2__abc_44228_n15405_bF_buf3), .B(u2_remLo_241_), .Y(u2__abc_44228_n16695) );
  AND2X2 AND2X2_7754 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_239_), .Y(u2__abc_44228_n16696) );
  AND2X2 AND2X2_7755 ( .A(u2__abc_44228_n2988_bF_buf1), .B(fracta1_97_), .Y(u2__abc_44228_n16697) );
  AND2X2 AND2X2_7756 ( .A(u2__abc_44228_n16698), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16699) );
  AND2X2 AND2X2_7757 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_240_), .Y(u2__abc_44228_n16701) );
  AND2X2 AND2X2_7758 ( .A(u2__abc_44228_n15403_bF_buf1), .B(u2_remLo_242_), .Y(u2__abc_44228_n16702) );
  AND2X2 AND2X2_7759 ( .A(u2__abc_44228_n16703), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16704) );
  AND2X2 AND2X2_776 ( .A(u2__abc_44228_n3520), .B(sqrto_40_), .Y(u2__abc_44228_n3521) );
  AND2X2 AND2X2_7760 ( .A(u2__abc_44228_n15402_bF_buf1), .B(u2_remLo_242_), .Y(u2__abc_44228_n16705) );
  AND2X2 AND2X2_7761 ( .A(u2__abc_44228_n2989_bF_buf0), .B(fracta1_98_), .Y(u2__abc_44228_n16706) );
  AND2X2 AND2X2_7762 ( .A(u2__abc_44228_n15405_bF_buf2), .B(u2_remLo_243_), .Y(u2__abc_44228_n16709) );
  AND2X2 AND2X2_7763 ( .A(u2__abc_44228_n2988_bF_buf0), .B(fracta1_99_), .Y(u2__abc_44228_n16710) );
  AND2X2 AND2X2_7764 ( .A(u2__abc_44228_n15408_bF_buf13), .B(u2_remLo_241_), .Y(u2__abc_44228_n16711) );
  AND2X2 AND2X2_7765 ( .A(u2__abc_44228_n16712), .B(u2__abc_44228_n2987_bF_buf9), .Y(u2__abc_44228_n16713) );
  AND2X2 AND2X2_7766 ( .A(u2__abc_44228_n15405_bF_buf1), .B(u2_remLo_244_), .Y(u2__abc_44228_n16715) );
  AND2X2 AND2X2_7767 ( .A(u2__abc_44228_n2988_bF_buf13), .B(fracta1_100_), .Y(u2__abc_44228_n16716) );
  AND2X2 AND2X2_7768 ( .A(u2__abc_44228_n15408_bF_buf12), .B(u2_remLo_242_), .Y(u2__abc_44228_n16717) );
  AND2X2 AND2X2_7769 ( .A(u2__abc_44228_n16718), .B(u2__abc_44228_n2987_bF_buf8), .Y(u2__abc_44228_n16719) );
  AND2X2 AND2X2_777 ( .A(u2__abc_44228_n3523_1), .B(u2__abc_44228_n3517), .Y(u2__abc_44228_n3524) );
  AND2X2 AND2X2_7770 ( .A(u2__abc_44228_n15405_bF_buf0), .B(u2_remLo_245_), .Y(u2__abc_44228_n16721) );
  AND2X2 AND2X2_7771 ( .A(u2__abc_44228_n15408_bF_buf11), .B(u2_remLo_243_), .Y(u2__abc_44228_n16722) );
  AND2X2 AND2X2_7772 ( .A(u2__abc_44228_n2988_bF_buf12), .B(fracta1_101_), .Y(u2__abc_44228_n16723) );
  AND2X2 AND2X2_7773 ( .A(u2__abc_44228_n16724), .B(u2__abc_44228_n2987_bF_buf7), .Y(u2__abc_44228_n16725) );
  AND2X2 AND2X2_7774 ( .A(u2__abc_44228_n15408_bF_buf10), .B(u2_remLo_244_), .Y(u2__abc_44228_n16727) );
  AND2X2 AND2X2_7775 ( .A(u2__abc_44228_n15403_bF_buf0), .B(u2_remLo_246_), .Y(u2__abc_44228_n16728) );
  AND2X2 AND2X2_7776 ( .A(u2__abc_44228_n16729), .B(u2__abc_44228_n2987_bF_buf6), .Y(u2__abc_44228_n16730) );
  AND2X2 AND2X2_7777 ( .A(u2__abc_44228_n15402_bF_buf0), .B(u2_remLo_246_), .Y(u2__abc_44228_n16731) );
  AND2X2 AND2X2_7778 ( .A(u2__abc_44228_n2989_bF_buf3), .B(fracta1_102_), .Y(u2__abc_44228_n16732) );
  AND2X2 AND2X2_7779 ( .A(u2__abc_44228_n15405_bF_buf13), .B(u2_remLo_247_), .Y(u2__abc_44228_n16735) );
  AND2X2 AND2X2_778 ( .A(u2__abc_44228_n3510), .B(u2__abc_44228_n3524), .Y(u2__abc_44228_n3525) );
  AND2X2 AND2X2_7780 ( .A(u2__abc_44228_n15408_bF_buf9), .B(u2_remLo_245_), .Y(u2__abc_44228_n16736) );
  AND2X2 AND2X2_7781 ( .A(u2__abc_44228_n2988_bF_buf11), .B(fracta1_103_), .Y(u2__abc_44228_n16737) );
  AND2X2 AND2X2_7782 ( .A(u2__abc_44228_n16738), .B(u2__abc_44228_n2987_bF_buf5), .Y(u2__abc_44228_n16739) );
  AND2X2 AND2X2_7783 ( .A(u2__abc_44228_n15405_bF_buf12), .B(u2_remLo_248_), .Y(u2__abc_44228_n16741) );
  AND2X2 AND2X2_7784 ( .A(u2__abc_44228_n15408_bF_buf8), .B(u2_remLo_246_), .Y(u2__abc_44228_n16742) );
  AND2X2 AND2X2_7785 ( .A(u2__abc_44228_n2988_bF_buf10), .B(fracta1_104_), .Y(u2__abc_44228_n16743) );
  AND2X2 AND2X2_7786 ( .A(u2__abc_44228_n16744), .B(u2__abc_44228_n2987_bF_buf4), .Y(u2__abc_44228_n16745) );
  AND2X2 AND2X2_7787 ( .A(u2__abc_44228_n15405_bF_buf11), .B(u2_remLo_249_), .Y(u2__abc_44228_n16747) );
  AND2X2 AND2X2_7788 ( .A(u2__abc_44228_n15408_bF_buf7), .B(u2_remLo_247_), .Y(u2__abc_44228_n16748) );
  AND2X2 AND2X2_7789 ( .A(u2__abc_44228_n2988_bF_buf9), .B(fracta1_105_), .Y(u2__abc_44228_n16749) );
  AND2X2 AND2X2_779 ( .A(u2__abc_44228_n3496), .B(u2__abc_44228_n3525), .Y(u2__abc_44228_n3526) );
  AND2X2 AND2X2_7790 ( .A(u2__abc_44228_n16750), .B(u2__abc_44228_n2987_bF_buf3), .Y(u2__abc_44228_n16751) );
  AND2X2 AND2X2_7791 ( .A(u2__abc_44228_n15405_bF_buf10), .B(u2_remLo_250_), .Y(u2__abc_44228_n16753) );
  AND2X2 AND2X2_7792 ( .A(u2__abc_44228_n2988_bF_buf8), .B(fracta1_106_), .Y(u2__abc_44228_n16754) );
  AND2X2 AND2X2_7793 ( .A(u2__abc_44228_n15408_bF_buf6), .B(u2_remLo_248_), .Y(u2__abc_44228_n16755) );
  AND2X2 AND2X2_7794 ( .A(u2__abc_44228_n16756), .B(u2__abc_44228_n2987_bF_buf2), .Y(u2__abc_44228_n16757) );
  AND2X2 AND2X2_7795 ( .A(u2__abc_44228_n15403_bF_buf3), .B(u2_remLo_251_), .Y(u2__abc_44228_n16759) );
  AND2X2 AND2X2_7796 ( .A(u2__abc_44228_n15408_bF_buf5), .B(u2_remLo_249_), .Y(u2__abc_44228_n16760) );
  AND2X2 AND2X2_7797 ( .A(u2__abc_44228_n16761), .B(u2__abc_44228_n2987_bF_buf1), .Y(u2__abc_44228_n16762) );
  AND2X2 AND2X2_7798 ( .A(u2__abc_44228_n15402_bF_buf3), .B(u2_remLo_251_), .Y(u2__abc_44228_n16763) );
  AND2X2 AND2X2_7799 ( .A(u2__abc_44228_n2989_bF_buf2), .B(fracta1_107_), .Y(u2__abc_44228_n16764) );
  AND2X2 AND2X2_78 ( .A(_abc_64468_n834), .B(_abc_64468_n833), .Y(_auto_iopadmap_cc_313_execute_65414_113_) );
  AND2X2 AND2X2_780 ( .A(u2__abc_44228_n3527), .B(u2_remHi_37_), .Y(u2__abc_44228_n3528) );
  AND2X2 AND2X2_7800 ( .A(u2__abc_44228_n15405_bF_buf9), .B(u2_remLo_252_), .Y(u2__abc_44228_n16767) );
  AND2X2 AND2X2_7801 ( .A(u2__abc_44228_n15408_bF_buf4), .B(u2_remLo_250_), .Y(u2__abc_44228_n16768) );
  AND2X2 AND2X2_7802 ( .A(u2__abc_44228_n2988_bF_buf7), .B(fracta1_108_), .Y(u2__abc_44228_n16769) );
  AND2X2 AND2X2_7803 ( .A(u2__abc_44228_n16770), .B(u2__abc_44228_n2987_bF_buf0), .Y(u2__abc_44228_n16771) );
  AND2X2 AND2X2_7804 ( .A(u2__abc_44228_n15405_bF_buf8), .B(u2_remLo_253_), .Y(u2__abc_44228_n16773) );
  AND2X2 AND2X2_7805 ( .A(u2__abc_44228_n15408_bF_buf3), .B(u2_remLo_251_), .Y(u2__abc_44228_n16774) );
  AND2X2 AND2X2_7806 ( .A(u2__abc_44228_n2988_bF_buf6), .B(fracta1_109_), .Y(u2__abc_44228_n16775) );
  AND2X2 AND2X2_7807 ( .A(u2__abc_44228_n16776), .B(u2__abc_44228_n2987_bF_buf14), .Y(u2__abc_44228_n16777) );
  AND2X2 AND2X2_7808 ( .A(u2__abc_44228_n15405_bF_buf7), .B(u2_remLo_254_), .Y(u2__abc_44228_n16779) );
  AND2X2 AND2X2_7809 ( .A(u2__abc_44228_n2988_bF_buf5), .B(fracta1_110_), .Y(u2__abc_44228_n16780) );
  AND2X2 AND2X2_781 ( .A(u2__abc_44228_n3530), .B(sqrto_37_), .Y(u2__abc_44228_n3531) );
  AND2X2 AND2X2_7810 ( .A(u2__abc_44228_n15408_bF_buf2), .B(u2_remLo_252_), .Y(u2__abc_44228_n16781) );
  AND2X2 AND2X2_7811 ( .A(u2__abc_44228_n16782), .B(u2__abc_44228_n2987_bF_buf13), .Y(u2__abc_44228_n16783) );
  AND2X2 AND2X2_7812 ( .A(u2__abc_44228_n15405_bF_buf6), .B(u2_remLo_255_), .Y(u2__abc_44228_n16785) );
  AND2X2 AND2X2_7813 ( .A(u2__abc_44228_n15408_bF_buf1), .B(u2_remLo_253_), .Y(u2__abc_44228_n16786) );
  AND2X2 AND2X2_7814 ( .A(u2__abc_44228_n2988_bF_buf4), .B(fracta1_111_), .Y(u2__abc_44228_n16787) );
  AND2X2 AND2X2_7815 ( .A(u2__abc_44228_n16788), .B(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n16789) );
  AND2X2 AND2X2_7816 ( .A(u2__abc_44228_n15405_bF_buf5), .B(u2_remLo_256_), .Y(u2__abc_44228_n16791) );
  AND2X2 AND2X2_7817 ( .A(u2__abc_44228_n2988_bF_buf3), .B(fracta1_112_), .Y(u2__abc_44228_n16792) );
  AND2X2 AND2X2_7818 ( .A(u2__abc_44228_n15408_bF_buf0), .B(u2_remLo_254_), .Y(u2__abc_44228_n16793) );
  AND2X2 AND2X2_7819 ( .A(u2__abc_44228_n16794), .B(u2__abc_44228_n2987_bF_buf11), .Y(u2__abc_44228_n16795) );
  AND2X2 AND2X2_782 ( .A(u2__abc_44228_n3529), .B(u2__abc_44228_n3532_1), .Y(u2__abc_44228_n3533) );
  AND2X2 AND2X2_7820 ( .A(u2__abc_44228_n15405_bF_buf4), .B(u2_remLo_257_), .Y(u2__abc_44228_n16797) );
  AND2X2 AND2X2_7821 ( .A(u2__abc_44228_n2988_bF_buf2), .B(fracta1_113_), .Y(u2__abc_44228_n16798) );
  AND2X2 AND2X2_7822 ( .A(u2__abc_44228_n15408_bF_buf14), .B(u2_remLo_255_), .Y(u2__abc_44228_n16799) );
  AND2X2 AND2X2_7823 ( .A(u2__abc_44228_n16800), .B(u2__abc_44228_n2987_bF_buf10), .Y(u2__abc_44228_n16801) );
  AND2X2 AND2X2_7824 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_258_), .Y(u2__abc_44228_n16803) );
  AND2X2 AND2X2_7825 ( .A(u2__abc_44228_n2972_bF_buf57), .B(u2_remLo_256_), .Y(u2__abc_44228_n16804) );
  AND2X2 AND2X2_7826 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n16804), .Y(u2__abc_44228_n16805) );
  AND2X2 AND2X2_7827 ( .A(u2__abc_44228_n16806), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_remLo_258__FF_INPUT) );
  AND2X2 AND2X2_7828 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_259_), .Y(u2__abc_44228_n16808) );
  AND2X2 AND2X2_7829 ( .A(u2__abc_44228_n2972_bF_buf56), .B(u2_remLo_257_), .Y(u2__abc_44228_n16809) );
  AND2X2 AND2X2_783 ( .A(u2__abc_44228_n3534), .B(u2_remHi_36_), .Y(u2__abc_44228_n3535) );
  AND2X2 AND2X2_7830 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n16809), .Y(u2__abc_44228_n16810) );
  AND2X2 AND2X2_7831 ( .A(u2__abc_44228_n16811), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_remLo_259__FF_INPUT) );
  AND2X2 AND2X2_7832 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_260_), .Y(u2__abc_44228_n16813) );
  AND2X2 AND2X2_7833 ( .A(u2__abc_44228_n2972_bF_buf55), .B(u2_remLo_258_), .Y(u2__abc_44228_n16814) );
  AND2X2 AND2X2_7834 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n16814), .Y(u2__abc_44228_n16815) );
  AND2X2 AND2X2_7835 ( .A(u2__abc_44228_n16816), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_remLo_260__FF_INPUT) );
  AND2X2 AND2X2_7836 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_261_), .Y(u2__abc_44228_n16818) );
  AND2X2 AND2X2_7837 ( .A(u2__abc_44228_n2972_bF_buf54), .B(u2_remLo_259_), .Y(u2__abc_44228_n16819) );
  AND2X2 AND2X2_7838 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n16819), .Y(u2__abc_44228_n16820) );
  AND2X2 AND2X2_7839 ( .A(u2__abc_44228_n16821), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_remLo_261__FF_INPUT) );
  AND2X2 AND2X2_784 ( .A(u2__abc_44228_n3536), .B(sqrto_36_), .Y(u2__abc_44228_n3537) );
  AND2X2 AND2X2_7840 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_262_), .Y(u2__abc_44228_n16823) );
  AND2X2 AND2X2_7841 ( .A(u2__abc_44228_n2972_bF_buf53), .B(u2_remLo_260_), .Y(u2__abc_44228_n16824) );
  AND2X2 AND2X2_7842 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n16824), .Y(u2__abc_44228_n16825) );
  AND2X2 AND2X2_7843 ( .A(u2__abc_44228_n16826), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_remLo_262__FF_INPUT) );
  AND2X2 AND2X2_7844 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_263_), .Y(u2__abc_44228_n16828) );
  AND2X2 AND2X2_7845 ( .A(u2__abc_44228_n2972_bF_buf52), .B(u2_remLo_261_), .Y(u2__abc_44228_n16829) );
  AND2X2 AND2X2_7846 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n16829), .Y(u2__abc_44228_n16830) );
  AND2X2 AND2X2_7847 ( .A(u2__abc_44228_n16831), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_remLo_263__FF_INPUT) );
  AND2X2 AND2X2_7848 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_264_), .Y(u2__abc_44228_n16833) );
  AND2X2 AND2X2_7849 ( .A(u2__abc_44228_n2972_bF_buf51), .B(u2_remLo_262_), .Y(u2__abc_44228_n16834) );
  AND2X2 AND2X2_785 ( .A(u2__abc_44228_n3539), .B(u2__abc_44228_n3533), .Y(u2__abc_44228_n3540) );
  AND2X2 AND2X2_7850 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n16834), .Y(u2__abc_44228_n16835) );
  AND2X2 AND2X2_7851 ( .A(u2__abc_44228_n16836), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_remLo_264__FF_INPUT) );
  AND2X2 AND2X2_7852 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_265_), .Y(u2__abc_44228_n16838) );
  AND2X2 AND2X2_7853 ( .A(u2__abc_44228_n2972_bF_buf50), .B(u2_remLo_263_), .Y(u2__abc_44228_n16839) );
  AND2X2 AND2X2_7854 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n16839), .Y(u2__abc_44228_n16840) );
  AND2X2 AND2X2_7855 ( .A(u2__abc_44228_n16841), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_remLo_265__FF_INPUT) );
  AND2X2 AND2X2_7856 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_266_), .Y(u2__abc_44228_n16843) );
  AND2X2 AND2X2_7857 ( .A(u2__abc_44228_n2972_bF_buf49), .B(u2_remLo_264_), .Y(u2__abc_44228_n16844) );
  AND2X2 AND2X2_7858 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n16844), .Y(u2__abc_44228_n16845) );
  AND2X2 AND2X2_7859 ( .A(u2__abc_44228_n16846), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_remLo_266__FF_INPUT) );
  AND2X2 AND2X2_786 ( .A(u2__abc_44228_n3541_1), .B(u2_remHi_34_), .Y(u2__abc_44228_n3542) );
  AND2X2 AND2X2_7860 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_267_), .Y(u2__abc_44228_n16848) );
  AND2X2 AND2X2_7861 ( .A(u2__abc_44228_n2972_bF_buf48), .B(u2_remLo_265_), .Y(u2__abc_44228_n16849) );
  AND2X2 AND2X2_7862 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n16849), .Y(u2__abc_44228_n16850) );
  AND2X2 AND2X2_7863 ( .A(u2__abc_44228_n16851), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_remLo_267__FF_INPUT) );
  AND2X2 AND2X2_7864 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_268_), .Y(u2__abc_44228_n16853) );
  AND2X2 AND2X2_7865 ( .A(u2__abc_44228_n2972_bF_buf47), .B(u2_remLo_266_), .Y(u2__abc_44228_n16854) );
  AND2X2 AND2X2_7866 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n16854), .Y(u2__abc_44228_n16855) );
  AND2X2 AND2X2_7867 ( .A(u2__abc_44228_n16856), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_remLo_268__FF_INPUT) );
  AND2X2 AND2X2_7868 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_269_), .Y(u2__abc_44228_n16858) );
  AND2X2 AND2X2_7869 ( .A(u2__abc_44228_n2972_bF_buf46), .B(u2_remLo_267_), .Y(u2__abc_44228_n16859) );
  AND2X2 AND2X2_787 ( .A(u2__abc_44228_n3543), .B(sqrto_34_), .Y(u2__abc_44228_n3544) );
  AND2X2 AND2X2_7870 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n16859), .Y(u2__abc_44228_n16860) );
  AND2X2 AND2X2_7871 ( .A(u2__abc_44228_n16861), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_remLo_269__FF_INPUT) );
  AND2X2 AND2X2_7872 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_270_), .Y(u2__abc_44228_n16863) );
  AND2X2 AND2X2_7873 ( .A(u2__abc_44228_n2972_bF_buf45), .B(u2_remLo_268_), .Y(u2__abc_44228_n16864) );
  AND2X2 AND2X2_7874 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n16864), .Y(u2__abc_44228_n16865) );
  AND2X2 AND2X2_7875 ( .A(u2__abc_44228_n16866), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_remLo_270__FF_INPUT) );
  AND2X2 AND2X2_7876 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_271_), .Y(u2__abc_44228_n16868) );
  AND2X2 AND2X2_7877 ( .A(u2__abc_44228_n2972_bF_buf44), .B(u2_remLo_269_), .Y(u2__abc_44228_n16869) );
  AND2X2 AND2X2_7878 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n16869), .Y(u2__abc_44228_n16870) );
  AND2X2 AND2X2_7879 ( .A(u2__abc_44228_n16871), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_remLo_271__FF_INPUT) );
  AND2X2 AND2X2_788 ( .A(u2__abc_44228_n3547), .B(u2_remHi_35_), .Y(u2__abc_44228_n3548) );
  AND2X2 AND2X2_7880 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_272_), .Y(u2__abc_44228_n16873) );
  AND2X2 AND2X2_7881 ( .A(u2__abc_44228_n2972_bF_buf43), .B(u2_remLo_270_), .Y(u2__abc_44228_n16874) );
  AND2X2 AND2X2_7882 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n16874), .Y(u2__abc_44228_n16875) );
  AND2X2 AND2X2_7883 ( .A(u2__abc_44228_n16876), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_remLo_272__FF_INPUT) );
  AND2X2 AND2X2_7884 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_273_), .Y(u2__abc_44228_n16878) );
  AND2X2 AND2X2_7885 ( .A(u2__abc_44228_n2972_bF_buf42), .B(u2_remLo_271_), .Y(u2__abc_44228_n16879) );
  AND2X2 AND2X2_7886 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n16879), .Y(u2__abc_44228_n16880) );
  AND2X2 AND2X2_7887 ( .A(u2__abc_44228_n16881), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_remLo_273__FF_INPUT) );
  AND2X2 AND2X2_7888 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_274_), .Y(u2__abc_44228_n16883) );
  AND2X2 AND2X2_7889 ( .A(u2__abc_44228_n2972_bF_buf41), .B(u2_remLo_272_), .Y(u2__abc_44228_n16884) );
  AND2X2 AND2X2_789 ( .A(u2__abc_44228_n3550), .B(sqrto_35_), .Y(u2__abc_44228_n3551) );
  AND2X2 AND2X2_7890 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n16884), .Y(u2__abc_44228_n16885) );
  AND2X2 AND2X2_7891 ( .A(u2__abc_44228_n16886), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_remLo_274__FF_INPUT) );
  AND2X2 AND2X2_7892 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_275_), .Y(u2__abc_44228_n16888) );
  AND2X2 AND2X2_7893 ( .A(u2__abc_44228_n2972_bF_buf40), .B(u2_remLo_273_), .Y(u2__abc_44228_n16889) );
  AND2X2 AND2X2_7894 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n16889), .Y(u2__abc_44228_n16890) );
  AND2X2 AND2X2_7895 ( .A(u2__abc_44228_n16891), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_remLo_275__FF_INPUT) );
  AND2X2 AND2X2_7896 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_276_), .Y(u2__abc_44228_n16893) );
  AND2X2 AND2X2_7897 ( .A(u2__abc_44228_n2972_bF_buf39), .B(u2_remLo_274_), .Y(u2__abc_44228_n16894) );
  AND2X2 AND2X2_7898 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n16894), .Y(u2__abc_44228_n16895) );
  AND2X2 AND2X2_7899 ( .A(u2__abc_44228_n16896), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_remLo_276__FF_INPUT) );
  AND2X2 AND2X2_79 ( .A(_abc_64468_n837), .B(_abc_64468_n836), .Y(_auto_iopadmap_cc_313_execute_65414_114_) );
  AND2X2 AND2X2_790 ( .A(u2__abc_44228_n3549), .B(u2__abc_44228_n3552_1), .Y(u2__abc_44228_n3553) );
  AND2X2 AND2X2_7900 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_277_), .Y(u2__abc_44228_n16898) );
  AND2X2 AND2X2_7901 ( .A(u2__abc_44228_n2972_bF_buf38), .B(u2_remLo_275_), .Y(u2__abc_44228_n16899) );
  AND2X2 AND2X2_7902 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n16899), .Y(u2__abc_44228_n16900) );
  AND2X2 AND2X2_7903 ( .A(u2__abc_44228_n16901), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_remLo_277__FF_INPUT) );
  AND2X2 AND2X2_7904 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_278_), .Y(u2__abc_44228_n16903) );
  AND2X2 AND2X2_7905 ( .A(u2__abc_44228_n2972_bF_buf37), .B(u2_remLo_276_), .Y(u2__abc_44228_n16904) );
  AND2X2 AND2X2_7906 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n16904), .Y(u2__abc_44228_n16905) );
  AND2X2 AND2X2_7907 ( .A(u2__abc_44228_n16906), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_remLo_278__FF_INPUT) );
  AND2X2 AND2X2_7908 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_279_), .Y(u2__abc_44228_n16908) );
  AND2X2 AND2X2_7909 ( .A(u2__abc_44228_n2972_bF_buf36), .B(u2_remLo_277_), .Y(u2__abc_44228_n16909) );
  AND2X2 AND2X2_791 ( .A(u2__abc_44228_n3546), .B(u2__abc_44228_n3553), .Y(u2__abc_44228_n3554) );
  AND2X2 AND2X2_7910 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n16909), .Y(u2__abc_44228_n16910) );
  AND2X2 AND2X2_7911 ( .A(u2__abc_44228_n16911), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_remLo_279__FF_INPUT) );
  AND2X2 AND2X2_7912 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_280_), .Y(u2__abc_44228_n16913) );
  AND2X2 AND2X2_7913 ( .A(u2__abc_44228_n2972_bF_buf35), .B(u2_remLo_278_), .Y(u2__abc_44228_n16914) );
  AND2X2 AND2X2_7914 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n16914), .Y(u2__abc_44228_n16915) );
  AND2X2 AND2X2_7915 ( .A(u2__abc_44228_n16916), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_remLo_280__FF_INPUT) );
  AND2X2 AND2X2_7916 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_281_), .Y(u2__abc_44228_n16918) );
  AND2X2 AND2X2_7917 ( .A(u2__abc_44228_n2972_bF_buf34), .B(u2_remLo_279_), .Y(u2__abc_44228_n16919) );
  AND2X2 AND2X2_7918 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n16919), .Y(u2__abc_44228_n16920) );
  AND2X2 AND2X2_7919 ( .A(u2__abc_44228_n16921), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_remLo_281__FF_INPUT) );
  AND2X2 AND2X2_792 ( .A(u2__abc_44228_n3540), .B(u2__abc_44228_n3554), .Y(u2__abc_44228_n3555) );
  AND2X2 AND2X2_7920 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_282_), .Y(u2__abc_44228_n16923) );
  AND2X2 AND2X2_7921 ( .A(u2__abc_44228_n2972_bF_buf33), .B(u2_remLo_280_), .Y(u2__abc_44228_n16924) );
  AND2X2 AND2X2_7922 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n16924), .Y(u2__abc_44228_n16925) );
  AND2X2 AND2X2_7923 ( .A(u2__abc_44228_n16926), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_remLo_282__FF_INPUT) );
  AND2X2 AND2X2_7924 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_283_), .Y(u2__abc_44228_n16928) );
  AND2X2 AND2X2_7925 ( .A(u2__abc_44228_n2972_bF_buf32), .B(u2_remLo_281_), .Y(u2__abc_44228_n16929) );
  AND2X2 AND2X2_7926 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n16929), .Y(u2__abc_44228_n16930) );
  AND2X2 AND2X2_7927 ( .A(u2__abc_44228_n16931), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_remLo_283__FF_INPUT) );
  AND2X2 AND2X2_7928 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_284_), .Y(u2__abc_44228_n16933) );
  AND2X2 AND2X2_7929 ( .A(u2__abc_44228_n2972_bF_buf31), .B(u2_remLo_282_), .Y(u2__abc_44228_n16934) );
  AND2X2 AND2X2_793 ( .A(u2__abc_44228_n3557), .B(u2__abc_44228_n3559), .Y(u2__abc_44228_n3560) );
  AND2X2 AND2X2_7930 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n16934), .Y(u2__abc_44228_n16935) );
  AND2X2 AND2X2_7931 ( .A(u2__abc_44228_n16936), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_remLo_284__FF_INPUT) );
  AND2X2 AND2X2_7932 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_285_), .Y(u2__abc_44228_n16938) );
  AND2X2 AND2X2_7933 ( .A(u2__abc_44228_n2972_bF_buf30), .B(u2_remLo_283_), .Y(u2__abc_44228_n16939) );
  AND2X2 AND2X2_7934 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n16939), .Y(u2__abc_44228_n16940) );
  AND2X2 AND2X2_7935 ( .A(u2__abc_44228_n16941), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_remLo_285__FF_INPUT) );
  AND2X2 AND2X2_7936 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_286_), .Y(u2__abc_44228_n16943) );
  AND2X2 AND2X2_7937 ( .A(u2__abc_44228_n2972_bF_buf29), .B(u2_remLo_284_), .Y(u2__abc_44228_n16944) );
  AND2X2 AND2X2_7938 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n16944), .Y(u2__abc_44228_n16945) );
  AND2X2 AND2X2_7939 ( .A(u2__abc_44228_n16946), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_remLo_286__FF_INPUT) );
  AND2X2 AND2X2_794 ( .A(u2__abc_44228_n3562_1), .B(u2__abc_44228_n3564), .Y(u2__abc_44228_n3565) );
  AND2X2 AND2X2_7940 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_287_), .Y(u2__abc_44228_n16948) );
  AND2X2 AND2X2_7941 ( .A(u2__abc_44228_n2972_bF_buf28), .B(u2_remLo_285_), .Y(u2__abc_44228_n16949) );
  AND2X2 AND2X2_7942 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n16949), .Y(u2__abc_44228_n16950) );
  AND2X2 AND2X2_7943 ( .A(u2__abc_44228_n16951), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_remLo_287__FF_INPUT) );
  AND2X2 AND2X2_7944 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_288_), .Y(u2__abc_44228_n16953) );
  AND2X2 AND2X2_7945 ( .A(u2__abc_44228_n2972_bF_buf27), .B(u2_remLo_286_), .Y(u2__abc_44228_n16954) );
  AND2X2 AND2X2_7946 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n16954), .Y(u2__abc_44228_n16955) );
  AND2X2 AND2X2_7947 ( .A(u2__abc_44228_n16956), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_remLo_288__FF_INPUT) );
  AND2X2 AND2X2_7948 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_289_), .Y(u2__abc_44228_n16958) );
  AND2X2 AND2X2_7949 ( .A(u2__abc_44228_n2972_bF_buf26), .B(u2_remLo_287_), .Y(u2__abc_44228_n16959) );
  AND2X2 AND2X2_795 ( .A(u2__abc_44228_n3560), .B(u2__abc_44228_n3565), .Y(u2__abc_44228_n3566) );
  AND2X2 AND2X2_7950 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n16959), .Y(u2__abc_44228_n16960) );
  AND2X2 AND2X2_7951 ( .A(u2__abc_44228_n16961), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_remLo_289__FF_INPUT) );
  AND2X2 AND2X2_7952 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_290_), .Y(u2__abc_44228_n16963) );
  AND2X2 AND2X2_7953 ( .A(u2__abc_44228_n2972_bF_buf25), .B(u2_remLo_288_), .Y(u2__abc_44228_n16964) );
  AND2X2 AND2X2_7954 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n16964), .Y(u2__abc_44228_n16965) );
  AND2X2 AND2X2_7955 ( .A(u2__abc_44228_n16966), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_remLo_290__FF_INPUT) );
  AND2X2 AND2X2_7956 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_291_), .Y(u2__abc_44228_n16968) );
  AND2X2 AND2X2_7957 ( .A(u2__abc_44228_n2972_bF_buf24), .B(u2_remLo_289_), .Y(u2__abc_44228_n16969) );
  AND2X2 AND2X2_7958 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n16969), .Y(u2__abc_44228_n16970) );
  AND2X2 AND2X2_7959 ( .A(u2__abc_44228_n16971), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_remLo_291__FF_INPUT) );
  AND2X2 AND2X2_796 ( .A(u2__abc_44228_n3567), .B(u2_remHi_30_), .Y(u2__abc_44228_n3568) );
  AND2X2 AND2X2_7960 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_292_), .Y(u2__abc_44228_n16973) );
  AND2X2 AND2X2_7961 ( .A(u2__abc_44228_n2972_bF_buf23), .B(u2_remLo_290_), .Y(u2__abc_44228_n16974) );
  AND2X2 AND2X2_7962 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n16974), .Y(u2__abc_44228_n16975) );
  AND2X2 AND2X2_7963 ( .A(u2__abc_44228_n16976), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_remLo_292__FF_INPUT) );
  AND2X2 AND2X2_7964 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_293_), .Y(u2__abc_44228_n16978) );
  AND2X2 AND2X2_7965 ( .A(u2__abc_44228_n2972_bF_buf22), .B(u2_remLo_291_), .Y(u2__abc_44228_n16979) );
  AND2X2 AND2X2_7966 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n16979), .Y(u2__abc_44228_n16980) );
  AND2X2 AND2X2_7967 ( .A(u2__abc_44228_n16981), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_remLo_293__FF_INPUT) );
  AND2X2 AND2X2_7968 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_294_), .Y(u2__abc_44228_n16983) );
  AND2X2 AND2X2_7969 ( .A(u2__abc_44228_n2972_bF_buf21), .B(u2_remLo_292_), .Y(u2__abc_44228_n16984) );
  AND2X2 AND2X2_797 ( .A(u2__abc_44228_n3569), .B(sqrto_30_), .Y(u2__abc_44228_n3570) );
  AND2X2 AND2X2_7970 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n16984), .Y(u2__abc_44228_n16985) );
  AND2X2 AND2X2_7971 ( .A(u2__abc_44228_n16986), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_remLo_294__FF_INPUT) );
  AND2X2 AND2X2_7972 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_295_), .Y(u2__abc_44228_n16988) );
  AND2X2 AND2X2_7973 ( .A(u2__abc_44228_n2972_bF_buf20), .B(u2_remLo_293_), .Y(u2__abc_44228_n16989) );
  AND2X2 AND2X2_7974 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n16989), .Y(u2__abc_44228_n16990) );
  AND2X2 AND2X2_7975 ( .A(u2__abc_44228_n16991), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_remLo_295__FF_INPUT) );
  AND2X2 AND2X2_7976 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_296_), .Y(u2__abc_44228_n16993) );
  AND2X2 AND2X2_7977 ( .A(u2__abc_44228_n2972_bF_buf19), .B(u2_remLo_294_), .Y(u2__abc_44228_n16994) );
  AND2X2 AND2X2_7978 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n16994), .Y(u2__abc_44228_n16995) );
  AND2X2 AND2X2_7979 ( .A(u2__abc_44228_n16996), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_remLo_296__FF_INPUT) );
  AND2X2 AND2X2_798 ( .A(u2__abc_44228_n3573), .B(u2_remHi_31_), .Y(u2__abc_44228_n3574) );
  AND2X2 AND2X2_7980 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_297_), .Y(u2__abc_44228_n16998) );
  AND2X2 AND2X2_7981 ( .A(u2__abc_44228_n2972_bF_buf18), .B(u2_remLo_295_), .Y(u2__abc_44228_n16999) );
  AND2X2 AND2X2_7982 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n16999), .Y(u2__abc_44228_n17000) );
  AND2X2 AND2X2_7983 ( .A(u2__abc_44228_n17001), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_remLo_297__FF_INPUT) );
  AND2X2 AND2X2_7984 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_298_), .Y(u2__abc_44228_n17003) );
  AND2X2 AND2X2_7985 ( .A(u2__abc_44228_n2972_bF_buf17), .B(u2_remLo_296_), .Y(u2__abc_44228_n17004) );
  AND2X2 AND2X2_7986 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17004), .Y(u2__abc_44228_n17005) );
  AND2X2 AND2X2_7987 ( .A(u2__abc_44228_n17006), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_remLo_298__FF_INPUT) );
  AND2X2 AND2X2_7988 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_299_), .Y(u2__abc_44228_n17008) );
  AND2X2 AND2X2_7989 ( .A(u2__abc_44228_n2972_bF_buf16), .B(u2_remLo_297_), .Y(u2__abc_44228_n17009) );
  AND2X2 AND2X2_799 ( .A(u2__abc_44228_n3576), .B(sqrto_31_), .Y(u2__abc_44228_n3577) );
  AND2X2 AND2X2_7990 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17009), .Y(u2__abc_44228_n17010) );
  AND2X2 AND2X2_7991 ( .A(u2__abc_44228_n17011), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_remLo_299__FF_INPUT) );
  AND2X2 AND2X2_7992 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_300_), .Y(u2__abc_44228_n17013) );
  AND2X2 AND2X2_7993 ( .A(u2__abc_44228_n2972_bF_buf15), .B(u2_remLo_298_), .Y(u2__abc_44228_n17014) );
  AND2X2 AND2X2_7994 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17014), .Y(u2__abc_44228_n17015) );
  AND2X2 AND2X2_7995 ( .A(u2__abc_44228_n17016), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_remLo_300__FF_INPUT) );
  AND2X2 AND2X2_7996 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_301_), .Y(u2__abc_44228_n17018) );
  AND2X2 AND2X2_7997 ( .A(u2__abc_44228_n2972_bF_buf14), .B(u2_remLo_299_), .Y(u2__abc_44228_n17019) );
  AND2X2 AND2X2_7998 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17019), .Y(u2__abc_44228_n17020) );
  AND2X2 AND2X2_7999 ( .A(u2__abc_44228_n17021), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_remLo_301__FF_INPUT) );
  AND2X2 AND2X2_8 ( .A(_abc_64468_n753_bF_buf6), .B(sqrto_7_), .Y(_auto_iopadmap_cc_313_execute_65414_43_) );
  AND2X2 AND2X2_80 ( .A(_abc_64468_n840_1), .B(_abc_64468_n839_1), .Y(_auto_iopadmap_cc_313_execute_65414_115_) );
  AND2X2 AND2X2_800 ( .A(u2__abc_44228_n3575), .B(u2__abc_44228_n3578), .Y(u2__abc_44228_n3579) );
  AND2X2 AND2X2_8000 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_302_), .Y(u2__abc_44228_n17023) );
  AND2X2 AND2X2_8001 ( .A(u2__abc_44228_n2972_bF_buf13), .B(u2_remLo_300_), .Y(u2__abc_44228_n17024) );
  AND2X2 AND2X2_8002 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17024), .Y(u2__abc_44228_n17025) );
  AND2X2 AND2X2_8003 ( .A(u2__abc_44228_n17026), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_remLo_302__FF_INPUT) );
  AND2X2 AND2X2_8004 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_303_), .Y(u2__abc_44228_n17028) );
  AND2X2 AND2X2_8005 ( .A(u2__abc_44228_n2972_bF_buf12), .B(u2_remLo_301_), .Y(u2__abc_44228_n17029) );
  AND2X2 AND2X2_8006 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17029), .Y(u2__abc_44228_n17030) );
  AND2X2 AND2X2_8007 ( .A(u2__abc_44228_n17031), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_remLo_303__FF_INPUT) );
  AND2X2 AND2X2_8008 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_304_), .Y(u2__abc_44228_n17033) );
  AND2X2 AND2X2_8009 ( .A(u2__abc_44228_n2972_bF_buf11), .B(u2_remLo_302_), .Y(u2__abc_44228_n17034) );
  AND2X2 AND2X2_801 ( .A(u2__abc_44228_n3572), .B(u2__abc_44228_n3579), .Y(u2__abc_44228_n3580_1) );
  AND2X2 AND2X2_8010 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17034), .Y(u2__abc_44228_n17035) );
  AND2X2 AND2X2_8011 ( .A(u2__abc_44228_n17036), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_remLo_304__FF_INPUT) );
  AND2X2 AND2X2_8012 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_305_), .Y(u2__abc_44228_n17038) );
  AND2X2 AND2X2_8013 ( .A(u2__abc_44228_n2972_bF_buf10), .B(u2_remLo_303_), .Y(u2__abc_44228_n17039) );
  AND2X2 AND2X2_8014 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17039), .Y(u2__abc_44228_n17040) );
  AND2X2 AND2X2_8015 ( .A(u2__abc_44228_n17041), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_remLo_305__FF_INPUT) );
  AND2X2 AND2X2_8016 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_306_), .Y(u2__abc_44228_n17043) );
  AND2X2 AND2X2_8017 ( .A(u2__abc_44228_n2972_bF_buf9), .B(u2_remLo_304_), .Y(u2__abc_44228_n17044) );
  AND2X2 AND2X2_8018 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17044), .Y(u2__abc_44228_n17045) );
  AND2X2 AND2X2_8019 ( .A(u2__abc_44228_n17046), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_remLo_306__FF_INPUT) );
  AND2X2 AND2X2_802 ( .A(u2__abc_44228_n3580_1), .B(u2__abc_44228_n3566), .Y(u2__abc_44228_n3581) );
  AND2X2 AND2X2_8020 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_307_), .Y(u2__abc_44228_n17048) );
  AND2X2 AND2X2_8021 ( .A(u2__abc_44228_n2972_bF_buf8), .B(u2_remLo_305_), .Y(u2__abc_44228_n17049) );
  AND2X2 AND2X2_8022 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17049), .Y(u2__abc_44228_n17050) );
  AND2X2 AND2X2_8023 ( .A(u2__abc_44228_n17051), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_remLo_307__FF_INPUT) );
  AND2X2 AND2X2_8024 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_308_), .Y(u2__abc_44228_n17053) );
  AND2X2 AND2X2_8025 ( .A(u2__abc_44228_n2972_bF_buf7), .B(u2_remLo_306_), .Y(u2__abc_44228_n17054) );
  AND2X2 AND2X2_8026 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17054), .Y(u2__abc_44228_n17055) );
  AND2X2 AND2X2_8027 ( .A(u2__abc_44228_n17056), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_remLo_308__FF_INPUT) );
  AND2X2 AND2X2_8028 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_309_), .Y(u2__abc_44228_n17058) );
  AND2X2 AND2X2_8029 ( .A(u2__abc_44228_n2972_bF_buf6), .B(u2_remLo_307_), .Y(u2__abc_44228_n17059) );
  AND2X2 AND2X2_803 ( .A(u2__abc_44228_n3555), .B(u2__abc_44228_n3581), .Y(u2__abc_44228_n3582) );
  AND2X2 AND2X2_8030 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17059), .Y(u2__abc_44228_n17060) );
  AND2X2 AND2X2_8031 ( .A(u2__abc_44228_n17061), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_remLo_309__FF_INPUT) );
  AND2X2 AND2X2_8032 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_310_), .Y(u2__abc_44228_n17063) );
  AND2X2 AND2X2_8033 ( .A(u2__abc_44228_n2972_bF_buf5), .B(u2_remLo_308_), .Y(u2__abc_44228_n17064) );
  AND2X2 AND2X2_8034 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17064), .Y(u2__abc_44228_n17065) );
  AND2X2 AND2X2_8035 ( .A(u2__abc_44228_n17066), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_remLo_310__FF_INPUT) );
  AND2X2 AND2X2_8036 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_311_), .Y(u2__abc_44228_n17068) );
  AND2X2 AND2X2_8037 ( .A(u2__abc_44228_n2972_bF_buf4), .B(u2_remLo_309_), .Y(u2__abc_44228_n17069) );
  AND2X2 AND2X2_8038 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17069), .Y(u2__abc_44228_n17070) );
  AND2X2 AND2X2_8039 ( .A(u2__abc_44228_n17071), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_remLo_311__FF_INPUT) );
  AND2X2 AND2X2_804 ( .A(u2__abc_44228_n3526), .B(u2__abc_44228_n3582), .Y(u2__abc_44228_n3583) );
  AND2X2 AND2X2_8040 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_312_), .Y(u2__abc_44228_n17073) );
  AND2X2 AND2X2_8041 ( .A(u2__abc_44228_n2972_bF_buf3), .B(u2_remLo_310_), .Y(u2__abc_44228_n17074) );
  AND2X2 AND2X2_8042 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17074), .Y(u2__abc_44228_n17075) );
  AND2X2 AND2X2_8043 ( .A(u2__abc_44228_n17076), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_remLo_312__FF_INPUT) );
  AND2X2 AND2X2_8044 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_313_), .Y(u2__abc_44228_n17078) );
  AND2X2 AND2X2_8045 ( .A(u2__abc_44228_n2972_bF_buf2), .B(u2_remLo_311_), .Y(u2__abc_44228_n17079) );
  AND2X2 AND2X2_8046 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17079), .Y(u2__abc_44228_n17080) );
  AND2X2 AND2X2_8047 ( .A(u2__abc_44228_n17081), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_remLo_313__FF_INPUT) );
  AND2X2 AND2X2_8048 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_314_), .Y(u2__abc_44228_n17083) );
  AND2X2 AND2X2_8049 ( .A(u2__abc_44228_n2972_bF_buf1), .B(u2_remLo_312_), .Y(u2__abc_44228_n17084) );
  AND2X2 AND2X2_805 ( .A(u2__abc_44228_n3467_1), .B(u2__abc_44228_n3583), .Y(u2__abc_44228_n3584) );
  AND2X2 AND2X2_8050 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17084), .Y(u2__abc_44228_n17085) );
  AND2X2 AND2X2_8051 ( .A(u2__abc_44228_n17086), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_remLo_314__FF_INPUT) );
  AND2X2 AND2X2_8052 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_315_), .Y(u2__abc_44228_n17088) );
  AND2X2 AND2X2_8053 ( .A(u2__abc_44228_n2972_bF_buf0), .B(u2_remLo_313_), .Y(u2__abc_44228_n17089) );
  AND2X2 AND2X2_8054 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17089), .Y(u2__abc_44228_n17090) );
  AND2X2 AND2X2_8055 ( .A(u2__abc_44228_n17091), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_remLo_315__FF_INPUT) );
  AND2X2 AND2X2_8056 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_316_), .Y(u2__abc_44228_n17093) );
  AND2X2 AND2X2_8057 ( .A(u2__abc_44228_n2972_bF_buf107), .B(u2_remLo_314_), .Y(u2__abc_44228_n17094) );
  AND2X2 AND2X2_8058 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17094), .Y(u2__abc_44228_n17095) );
  AND2X2 AND2X2_8059 ( .A(u2__abc_44228_n17096), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_remLo_316__FF_INPUT) );
  AND2X2 AND2X2_806 ( .A(u2__abc_44228_n3348), .B(u2__abc_44228_n3584), .Y(u2__abc_44228_n3585) );
  AND2X2 AND2X2_8060 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_317_), .Y(u2__abc_44228_n17098) );
  AND2X2 AND2X2_8061 ( .A(u2__abc_44228_n2972_bF_buf106), .B(u2_remLo_315_), .Y(u2__abc_44228_n17099) );
  AND2X2 AND2X2_8062 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17099), .Y(u2__abc_44228_n17100) );
  AND2X2 AND2X2_8063 ( .A(u2__abc_44228_n17101), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_remLo_317__FF_INPUT) );
  AND2X2 AND2X2_8064 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_318_), .Y(u2__abc_44228_n17103) );
  AND2X2 AND2X2_8065 ( .A(u2__abc_44228_n2972_bF_buf105), .B(u2_remLo_316_), .Y(u2__abc_44228_n17104) );
  AND2X2 AND2X2_8066 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17104), .Y(u2__abc_44228_n17105) );
  AND2X2 AND2X2_8067 ( .A(u2__abc_44228_n17106), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_remLo_318__FF_INPUT) );
  AND2X2 AND2X2_8068 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_319_), .Y(u2__abc_44228_n17108) );
  AND2X2 AND2X2_8069 ( .A(u2__abc_44228_n2972_bF_buf104), .B(u2_remLo_317_), .Y(u2__abc_44228_n17109) );
  AND2X2 AND2X2_807 ( .A(u2__abc_44228_n3586), .B(u2__abc_44228_n3578), .Y(u2__abc_44228_n3587) );
  AND2X2 AND2X2_8070 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17109), .Y(u2__abc_44228_n17110) );
  AND2X2 AND2X2_8071 ( .A(u2__abc_44228_n17111), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_remLo_319__FF_INPUT) );
  AND2X2 AND2X2_8072 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_320_), .Y(u2__abc_44228_n17113) );
  AND2X2 AND2X2_8073 ( .A(u2__abc_44228_n2972_bF_buf103), .B(u2_remLo_318_), .Y(u2__abc_44228_n17114) );
  AND2X2 AND2X2_8074 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17114), .Y(u2__abc_44228_n17115) );
  AND2X2 AND2X2_8075 ( .A(u2__abc_44228_n17116), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_remLo_320__FF_INPUT) );
  AND2X2 AND2X2_8076 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_321_), .Y(u2__abc_44228_n17118) );
  AND2X2 AND2X2_8077 ( .A(u2__abc_44228_n2972_bF_buf102), .B(u2_remLo_319_), .Y(u2__abc_44228_n17119) );
  AND2X2 AND2X2_8078 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17119), .Y(u2__abc_44228_n17120) );
  AND2X2 AND2X2_8079 ( .A(u2__abc_44228_n17121), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_remLo_321__FF_INPUT) );
  AND2X2 AND2X2_808 ( .A(u2__abc_44228_n3587), .B(u2__abc_44228_n3566), .Y(u2__abc_44228_n3588_1) );
  AND2X2 AND2X2_8080 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_322_), .Y(u2__abc_44228_n17123) );
  AND2X2 AND2X2_8081 ( .A(u2__abc_44228_n2972_bF_buf101), .B(u2_remLo_320_), .Y(u2__abc_44228_n17124) );
  AND2X2 AND2X2_8082 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17124), .Y(u2__abc_44228_n17125) );
  AND2X2 AND2X2_8083 ( .A(u2__abc_44228_n17126), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_remLo_322__FF_INPUT) );
  AND2X2 AND2X2_8084 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_323_), .Y(u2__abc_44228_n17128) );
  AND2X2 AND2X2_8085 ( .A(u2__abc_44228_n2972_bF_buf100), .B(u2_remLo_321_), .Y(u2__abc_44228_n17129) );
  AND2X2 AND2X2_8086 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17129), .Y(u2__abc_44228_n17130) );
  AND2X2 AND2X2_8087 ( .A(u2__abc_44228_n17131), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_remLo_323__FF_INPUT) );
  AND2X2 AND2X2_8088 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_324_), .Y(u2__abc_44228_n17133) );
  AND2X2 AND2X2_8089 ( .A(u2__abc_44228_n2972_bF_buf99), .B(u2_remLo_322_), .Y(u2__abc_44228_n17134) );
  AND2X2 AND2X2_809 ( .A(u2__abc_44228_n3590), .B(u2__abc_44228_n3559), .Y(u2__abc_44228_n3591) );
  AND2X2 AND2X2_8090 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17134), .Y(u2__abc_44228_n17135) );
  AND2X2 AND2X2_8091 ( .A(u2__abc_44228_n17136), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_remLo_324__FF_INPUT) );
  AND2X2 AND2X2_8092 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_325_), .Y(u2__abc_44228_n17138) );
  AND2X2 AND2X2_8093 ( .A(u2__abc_44228_n2972_bF_buf98), .B(u2_remLo_323_), .Y(u2__abc_44228_n17139) );
  AND2X2 AND2X2_8094 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17139), .Y(u2__abc_44228_n17140) );
  AND2X2 AND2X2_8095 ( .A(u2__abc_44228_n17141), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_remLo_325__FF_INPUT) );
  AND2X2 AND2X2_8096 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_326_), .Y(u2__abc_44228_n17143) );
  AND2X2 AND2X2_8097 ( .A(u2__abc_44228_n2972_bF_buf97), .B(u2_remLo_324_), .Y(u2__abc_44228_n17144) );
  AND2X2 AND2X2_8098 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17144), .Y(u2__abc_44228_n17145) );
  AND2X2 AND2X2_8099 ( .A(u2__abc_44228_n17146), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_remLo_326__FF_INPUT) );
  AND2X2 AND2X2_81 ( .A(_abc_64468_n843), .B(_abc_64468_n842), .Y(_auto_iopadmap_cc_313_execute_65414_116_) );
  AND2X2 AND2X2_810 ( .A(u2__abc_44228_n3593), .B(u2__abc_44228_n3555), .Y(u2__abc_44228_n3594) );
  AND2X2 AND2X2_8100 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_327_), .Y(u2__abc_44228_n17148) );
  AND2X2 AND2X2_8101 ( .A(u2__abc_44228_n2972_bF_buf96), .B(u2_remLo_325_), .Y(u2__abc_44228_n17149) );
  AND2X2 AND2X2_8102 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17149), .Y(u2__abc_44228_n17150) );
  AND2X2 AND2X2_8103 ( .A(u2__abc_44228_n17151), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_remLo_327__FF_INPUT) );
  AND2X2 AND2X2_8104 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_328_), .Y(u2__abc_44228_n17153) );
  AND2X2 AND2X2_8105 ( .A(u2__abc_44228_n2972_bF_buf95), .B(u2_remLo_326_), .Y(u2__abc_44228_n17154) );
  AND2X2 AND2X2_8106 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17154), .Y(u2__abc_44228_n17155) );
  AND2X2 AND2X2_8107 ( .A(u2__abc_44228_n17156), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_remLo_328__FF_INPUT) );
  AND2X2 AND2X2_8108 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_329_), .Y(u2__abc_44228_n17158) );
  AND2X2 AND2X2_8109 ( .A(u2__abc_44228_n2972_bF_buf94), .B(u2_remLo_327_), .Y(u2__abc_44228_n17159) );
  AND2X2 AND2X2_811 ( .A(u2__abc_44228_n3595), .B(u2__abc_44228_n3549), .Y(u2__abc_44228_n3596) );
  AND2X2 AND2X2_8110 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17159), .Y(u2__abc_44228_n17160) );
  AND2X2 AND2X2_8111 ( .A(u2__abc_44228_n17161), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_remLo_329__FF_INPUT) );
  AND2X2 AND2X2_8112 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_330_), .Y(u2__abc_44228_n17163) );
  AND2X2 AND2X2_8113 ( .A(u2__abc_44228_n2972_bF_buf93), .B(u2_remLo_328_), .Y(u2__abc_44228_n17164) );
  AND2X2 AND2X2_8114 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17164), .Y(u2__abc_44228_n17165) );
  AND2X2 AND2X2_8115 ( .A(u2__abc_44228_n17166), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_remLo_330__FF_INPUT) );
  AND2X2 AND2X2_8116 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_331_), .Y(u2__abc_44228_n17168) );
  AND2X2 AND2X2_8117 ( .A(u2__abc_44228_n2972_bF_buf92), .B(u2_remLo_329_), .Y(u2__abc_44228_n17169) );
  AND2X2 AND2X2_8118 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17169), .Y(u2__abc_44228_n17170) );
  AND2X2 AND2X2_8119 ( .A(u2__abc_44228_n17171), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_remLo_331__FF_INPUT) );
  AND2X2 AND2X2_812 ( .A(u2__abc_44228_n3597_1), .B(u2__abc_44228_n3552_1), .Y(u2__abc_44228_n3598) );
  AND2X2 AND2X2_8120 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_332_), .Y(u2__abc_44228_n17173) );
  AND2X2 AND2X2_8121 ( .A(u2__abc_44228_n2972_bF_buf91), .B(u2_remLo_330_), .Y(u2__abc_44228_n17174) );
  AND2X2 AND2X2_8122 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17174), .Y(u2__abc_44228_n17175) );
  AND2X2 AND2X2_8123 ( .A(u2__abc_44228_n17176), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_remLo_332__FF_INPUT) );
  AND2X2 AND2X2_8124 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_333_), .Y(u2__abc_44228_n17178) );
  AND2X2 AND2X2_8125 ( .A(u2__abc_44228_n2972_bF_buf90), .B(u2_remLo_331_), .Y(u2__abc_44228_n17179) );
  AND2X2 AND2X2_8126 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17179), .Y(u2__abc_44228_n17180) );
  AND2X2 AND2X2_8127 ( .A(u2__abc_44228_n17181), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_remLo_333__FF_INPUT) );
  AND2X2 AND2X2_8128 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_334_), .Y(u2__abc_44228_n17183) );
  AND2X2 AND2X2_8129 ( .A(u2__abc_44228_n2972_bF_buf89), .B(u2_remLo_332_), .Y(u2__abc_44228_n17184) );
  AND2X2 AND2X2_813 ( .A(u2__abc_44228_n3598), .B(u2__abc_44228_n3540), .Y(u2__abc_44228_n3599) );
  AND2X2 AND2X2_8130 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17184), .Y(u2__abc_44228_n17185) );
  AND2X2 AND2X2_8131 ( .A(u2__abc_44228_n17186), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_remLo_334__FF_INPUT) );
  AND2X2 AND2X2_8132 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_335_), .Y(u2__abc_44228_n17188) );
  AND2X2 AND2X2_8133 ( .A(u2__abc_44228_n2972_bF_buf88), .B(u2_remLo_333_), .Y(u2__abc_44228_n17189) );
  AND2X2 AND2X2_8134 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17189), .Y(u2__abc_44228_n17190) );
  AND2X2 AND2X2_8135 ( .A(u2__abc_44228_n17191), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_remLo_335__FF_INPUT) );
  AND2X2 AND2X2_8136 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_336_), .Y(u2__abc_44228_n17193) );
  AND2X2 AND2X2_8137 ( .A(u2__abc_44228_n2972_bF_buf87), .B(u2_remLo_334_), .Y(u2__abc_44228_n17194) );
  AND2X2 AND2X2_8138 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17194), .Y(u2__abc_44228_n17195) );
  AND2X2 AND2X2_8139 ( .A(u2__abc_44228_n17196), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_remLo_336__FF_INPUT) );
  AND2X2 AND2X2_814 ( .A(u2__abc_44228_n3600), .B(u2__abc_44228_n3532_1), .Y(u2__abc_44228_n3601) );
  AND2X2 AND2X2_8140 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_337_), .Y(u2__abc_44228_n17198) );
  AND2X2 AND2X2_8141 ( .A(u2__abc_44228_n2972_bF_buf86), .B(u2_remLo_335_), .Y(u2__abc_44228_n17199) );
  AND2X2 AND2X2_8142 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17199), .Y(u2__abc_44228_n17200) );
  AND2X2 AND2X2_8143 ( .A(u2__abc_44228_n17201), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_remLo_337__FF_INPUT) );
  AND2X2 AND2X2_8144 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_338_), .Y(u2__abc_44228_n17203) );
  AND2X2 AND2X2_8145 ( .A(u2__abc_44228_n2972_bF_buf85), .B(u2_remLo_336_), .Y(u2__abc_44228_n17204) );
  AND2X2 AND2X2_8146 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17204), .Y(u2__abc_44228_n17205) );
  AND2X2 AND2X2_8147 ( .A(u2__abc_44228_n17206), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_remLo_338__FF_INPUT) );
  AND2X2 AND2X2_8148 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_339_), .Y(u2__abc_44228_n17208) );
  AND2X2 AND2X2_8149 ( .A(u2__abc_44228_n2972_bF_buf84), .B(u2_remLo_337_), .Y(u2__abc_44228_n17209) );
  AND2X2 AND2X2_815 ( .A(u2__abc_44228_n3603), .B(u2__abc_44228_n3526), .Y(u2__abc_44228_n3604) );
  AND2X2 AND2X2_8150 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17209), .Y(u2__abc_44228_n17210) );
  AND2X2 AND2X2_8151 ( .A(u2__abc_44228_n17211), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_remLo_339__FF_INPUT) );
  AND2X2 AND2X2_8152 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_340_), .Y(u2__abc_44228_n17213) );
  AND2X2 AND2X2_8153 ( .A(u2__abc_44228_n2972_bF_buf83), .B(u2_remLo_338_), .Y(u2__abc_44228_n17214) );
  AND2X2 AND2X2_8154 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17214), .Y(u2__abc_44228_n17215) );
  AND2X2 AND2X2_8155 ( .A(u2__abc_44228_n17216), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_remLo_340__FF_INPUT) );
  AND2X2 AND2X2_8156 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_341_), .Y(u2__abc_44228_n17218) );
  AND2X2 AND2X2_8157 ( .A(u2__abc_44228_n2972_bF_buf82), .B(u2_remLo_339_), .Y(u2__abc_44228_n17219) );
  AND2X2 AND2X2_8158 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17219), .Y(u2__abc_44228_n17220) );
  AND2X2 AND2X2_8159 ( .A(u2__abc_44228_n17221), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_remLo_341__FF_INPUT) );
  AND2X2 AND2X2_816 ( .A(u2__abc_44228_n3605), .B(u2__abc_44228_n3502), .Y(u2__abc_44228_n3606) );
  AND2X2 AND2X2_8160 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_342_), .Y(u2__abc_44228_n17223) );
  AND2X2 AND2X2_8161 ( .A(u2__abc_44228_n2972_bF_buf81), .B(u2_remLo_340_), .Y(u2__abc_44228_n17224) );
  AND2X2 AND2X2_8162 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17224), .Y(u2__abc_44228_n17225) );
  AND2X2 AND2X2_8163 ( .A(u2__abc_44228_n17226), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_remLo_342__FF_INPUT) );
  AND2X2 AND2X2_8164 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_343_), .Y(u2__abc_44228_n17228) );
  AND2X2 AND2X2_8165 ( .A(u2__abc_44228_n2972_bF_buf80), .B(u2_remLo_341_), .Y(u2__abc_44228_n17229) );
  AND2X2 AND2X2_8166 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17229), .Y(u2__abc_44228_n17230) );
  AND2X2 AND2X2_8167 ( .A(u2__abc_44228_n17231), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_remLo_343__FF_INPUT) );
  AND2X2 AND2X2_8168 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_344_), .Y(u2__abc_44228_n17233) );
  AND2X2 AND2X2_8169 ( .A(u2__abc_44228_n2972_bF_buf79), .B(u2_remLo_342_), .Y(u2__abc_44228_n17234) );
  AND2X2 AND2X2_817 ( .A(u2__abc_44228_n3524), .B(u2__abc_44228_n3606), .Y(u2__abc_44228_n3607) );
  AND2X2 AND2X2_8170 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17234), .Y(u2__abc_44228_n17235) );
  AND2X2 AND2X2_8171 ( .A(u2__abc_44228_n17236), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_remLo_344__FF_INPUT) );
  AND2X2 AND2X2_8172 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_345_), .Y(u2__abc_44228_n17238) );
  AND2X2 AND2X2_8173 ( .A(u2__abc_44228_n2972_bF_buf78), .B(u2_remLo_343_), .Y(u2__abc_44228_n17239) );
  AND2X2 AND2X2_8174 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17239), .Y(u2__abc_44228_n17240) );
  AND2X2 AND2X2_8175 ( .A(u2__abc_44228_n17241), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_remLo_345__FF_INPUT) );
  AND2X2 AND2X2_8176 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_346_), .Y(u2__abc_44228_n17243) );
  AND2X2 AND2X2_8177 ( .A(u2__abc_44228_n2972_bF_buf77), .B(u2_remLo_344_), .Y(u2__abc_44228_n17244) );
  AND2X2 AND2X2_8178 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17244), .Y(u2__abc_44228_n17245) );
  AND2X2 AND2X2_8179 ( .A(u2__abc_44228_n17246), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_remLo_346__FF_INPUT) );
  AND2X2 AND2X2_818 ( .A(u2__abc_44228_n3513_1), .B(u2__abc_44228_n3608_1), .Y(u2__abc_44228_n3609) );
  AND2X2 AND2X2_8180 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_347_), .Y(u2__abc_44228_n17248) );
  AND2X2 AND2X2_8181 ( .A(u2__abc_44228_n2972_bF_buf76), .B(u2_remLo_345_), .Y(u2__abc_44228_n17249) );
  AND2X2 AND2X2_8182 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17249), .Y(u2__abc_44228_n17250) );
  AND2X2 AND2X2_8183 ( .A(u2__abc_44228_n17251), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_remLo_347__FF_INPUT) );
  AND2X2 AND2X2_8184 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_348_), .Y(u2__abc_44228_n17253) );
  AND2X2 AND2X2_8185 ( .A(u2__abc_44228_n2972_bF_buf75), .B(u2_remLo_346_), .Y(u2__abc_44228_n17254) );
  AND2X2 AND2X2_8186 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17254), .Y(u2__abc_44228_n17255) );
  AND2X2 AND2X2_8187 ( .A(u2__abc_44228_n17256), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_remLo_348__FF_INPUT) );
  AND2X2 AND2X2_8188 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_349_), .Y(u2__abc_44228_n17258) );
  AND2X2 AND2X2_8189 ( .A(u2__abc_44228_n2972_bF_buf74), .B(u2_remLo_347_), .Y(u2__abc_44228_n17259) );
  AND2X2 AND2X2_819 ( .A(u2__abc_44228_n3610), .B(u2__abc_44228_n3516), .Y(u2__abc_44228_n3611) );
  AND2X2 AND2X2_8190 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17259), .Y(u2__abc_44228_n17260) );
  AND2X2 AND2X2_8191 ( .A(u2__abc_44228_n17261), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_remLo_349__FF_INPUT) );
  AND2X2 AND2X2_8192 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_350_), .Y(u2__abc_44228_n17263) );
  AND2X2 AND2X2_8193 ( .A(u2__abc_44228_n2972_bF_buf73), .B(u2_remLo_348_), .Y(u2__abc_44228_n17264) );
  AND2X2 AND2X2_8194 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17264), .Y(u2__abc_44228_n17265) );
  AND2X2 AND2X2_8195 ( .A(u2__abc_44228_n17266), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_remLo_350__FF_INPUT) );
  AND2X2 AND2X2_8196 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_351_), .Y(u2__abc_44228_n17268) );
  AND2X2 AND2X2_8197 ( .A(u2__abc_44228_n2972_bF_buf72), .B(u2_remLo_349_), .Y(u2__abc_44228_n17269) );
  AND2X2 AND2X2_8198 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17269), .Y(u2__abc_44228_n17270) );
  AND2X2 AND2X2_8199 ( .A(u2__abc_44228_n17271), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_remLo_351__FF_INPUT) );
  AND2X2 AND2X2_82 ( .A(_abc_64468_n846), .B(_abc_64468_n845), .Y(_auto_iopadmap_cc_313_execute_65414_117_) );
  AND2X2 AND2X2_820 ( .A(u2__abc_44228_n3612), .B(u2__abc_44228_n3496), .Y(u2__abc_44228_n3613) );
  AND2X2 AND2X2_8200 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_352_), .Y(u2__abc_44228_n17273) );
  AND2X2 AND2X2_8201 ( .A(u2__abc_44228_n2972_bF_buf71), .B(u2_remLo_350_), .Y(u2__abc_44228_n17274) );
  AND2X2 AND2X2_8202 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17274), .Y(u2__abc_44228_n17275) );
  AND2X2 AND2X2_8203 ( .A(u2__abc_44228_n17276), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_remLo_352__FF_INPUT) );
  AND2X2 AND2X2_8204 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_353_), .Y(u2__abc_44228_n17278) );
  AND2X2 AND2X2_8205 ( .A(u2__abc_44228_n2972_bF_buf70), .B(u2_remLo_351_), .Y(u2__abc_44228_n17279) );
  AND2X2 AND2X2_8206 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17279), .Y(u2__abc_44228_n17280) );
  AND2X2 AND2X2_8207 ( .A(u2__abc_44228_n17281), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_remLo_353__FF_INPUT) );
  AND2X2 AND2X2_8208 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_354_), .Y(u2__abc_44228_n17283) );
  AND2X2 AND2X2_8209 ( .A(u2__abc_44228_n2972_bF_buf69), .B(u2_remLo_352_), .Y(u2__abc_44228_n17284) );
  AND2X2 AND2X2_821 ( .A(u2__abc_44228_n3473), .B(u2__abc_44228_n3476), .Y(u2__abc_44228_n3614) );
  AND2X2 AND2X2_8210 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17284), .Y(u2__abc_44228_n17285) );
  AND2X2 AND2X2_8211 ( .A(u2__abc_44228_n17286), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_remLo_354__FF_INPUT) );
  AND2X2 AND2X2_8212 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_355_), .Y(u2__abc_44228_n17288) );
  AND2X2 AND2X2_8213 ( .A(u2__abc_44228_n2972_bF_buf68), .B(u2_remLo_353_), .Y(u2__abc_44228_n17289) );
  AND2X2 AND2X2_8214 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17289), .Y(u2__abc_44228_n17290) );
  AND2X2 AND2X2_8215 ( .A(u2__abc_44228_n17291), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_remLo_355__FF_INPUT) );
  AND2X2 AND2X2_8216 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_356_), .Y(u2__abc_44228_n17293) );
  AND2X2 AND2X2_8217 ( .A(u2__abc_44228_n2972_bF_buf67), .B(u2_remLo_354_), .Y(u2__abc_44228_n17294) );
  AND2X2 AND2X2_8218 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17294), .Y(u2__abc_44228_n17295) );
  AND2X2 AND2X2_8219 ( .A(u2__abc_44228_n17296), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_remLo_356__FF_INPUT) );
  AND2X2 AND2X2_822 ( .A(u2__abc_44228_n3616), .B(u2__abc_44228_n3490), .Y(u2__abc_44228_n3617_1) );
  AND2X2 AND2X2_8220 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_357_), .Y(u2__abc_44228_n17298) );
  AND2X2 AND2X2_8221 ( .A(u2__abc_44228_n2972_bF_buf66), .B(u2_remLo_355_), .Y(u2__abc_44228_n17299) );
  AND2X2 AND2X2_8222 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17299), .Y(u2__abc_44228_n17300) );
  AND2X2 AND2X2_8223 ( .A(u2__abc_44228_n17301), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_remLo_357__FF_INPUT) );
  AND2X2 AND2X2_8224 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_358_), .Y(u2__abc_44228_n17303) );
  AND2X2 AND2X2_8225 ( .A(u2__abc_44228_n2972_bF_buf65), .B(u2_remLo_356_), .Y(u2__abc_44228_n17304) );
  AND2X2 AND2X2_8226 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17304), .Y(u2__abc_44228_n17305) );
  AND2X2 AND2X2_8227 ( .A(u2__abc_44228_n17306), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_remLo_358__FF_INPUT) );
  AND2X2 AND2X2_8228 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_359_), .Y(u2__abc_44228_n17308) );
  AND2X2 AND2X2_8229 ( .A(u2__abc_44228_n2972_bF_buf64), .B(u2_remLo_357_), .Y(u2__abc_44228_n17309) );
  AND2X2 AND2X2_823 ( .A(u2__abc_44228_n3618), .B(u2__abc_44228_n3493), .Y(u2__abc_44228_n3619) );
  AND2X2 AND2X2_8230 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17309), .Y(u2__abc_44228_n17310) );
  AND2X2 AND2X2_8231 ( .A(u2__abc_44228_n17311), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_remLo_359__FF_INPUT) );
  AND2X2 AND2X2_8232 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_360_), .Y(u2__abc_44228_n17313) );
  AND2X2 AND2X2_8233 ( .A(u2__abc_44228_n2972_bF_buf63), .B(u2_remLo_358_), .Y(u2__abc_44228_n17314) );
  AND2X2 AND2X2_8234 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17314), .Y(u2__abc_44228_n17315) );
  AND2X2 AND2X2_8235 ( .A(u2__abc_44228_n17316), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_remLo_360__FF_INPUT) );
  AND2X2 AND2X2_8236 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_361_), .Y(u2__abc_44228_n17318) );
  AND2X2 AND2X2_8237 ( .A(u2__abc_44228_n2972_bF_buf62), .B(u2_remLo_359_), .Y(u2__abc_44228_n17319) );
  AND2X2 AND2X2_8238 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17319), .Y(u2__abc_44228_n17320) );
  AND2X2 AND2X2_8239 ( .A(u2__abc_44228_n17321), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_remLo_361__FF_INPUT) );
  AND2X2 AND2X2_824 ( .A(u2__abc_44228_n3619), .B(u2__abc_44228_n3481), .Y(u2__abc_44228_n3620) );
  AND2X2 AND2X2_8240 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_362_), .Y(u2__abc_44228_n17323) );
  AND2X2 AND2X2_8241 ( .A(u2__abc_44228_n2972_bF_buf61), .B(u2_remLo_360_), .Y(u2__abc_44228_n17324) );
  AND2X2 AND2X2_8242 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17324), .Y(u2__abc_44228_n17325) );
  AND2X2 AND2X2_8243 ( .A(u2__abc_44228_n17326), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_remLo_362__FF_INPUT) );
  AND2X2 AND2X2_8244 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_363_), .Y(u2__abc_44228_n17328) );
  AND2X2 AND2X2_8245 ( .A(u2__abc_44228_n2972_bF_buf60), .B(u2_remLo_361_), .Y(u2__abc_44228_n17329) );
  AND2X2 AND2X2_8246 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17329), .Y(u2__abc_44228_n17330) );
  AND2X2 AND2X2_8247 ( .A(u2__abc_44228_n17331), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_remLo_363__FF_INPUT) );
  AND2X2 AND2X2_8248 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_364_), .Y(u2__abc_44228_n17333) );
  AND2X2 AND2X2_8249 ( .A(u2__abc_44228_n2972_bF_buf59), .B(u2_remLo_362_), .Y(u2__abc_44228_n17334) );
  AND2X2 AND2X2_825 ( .A(u2__abc_44228_n3623), .B(u2__abc_44228_n3467_1), .Y(u2__abc_44228_n3624) );
  AND2X2 AND2X2_8250 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17334), .Y(u2__abc_44228_n17335) );
  AND2X2 AND2X2_8251 ( .A(u2__abc_44228_n17336), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_remLo_364__FF_INPUT) );
  AND2X2 AND2X2_8252 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_365_), .Y(u2__abc_44228_n17338) );
  AND2X2 AND2X2_8253 ( .A(u2__abc_44228_n2972_bF_buf58), .B(u2_remLo_363_), .Y(u2__abc_44228_n17339) );
  AND2X2 AND2X2_8254 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17339), .Y(u2__abc_44228_n17340) );
  AND2X2 AND2X2_8255 ( .A(u2__abc_44228_n17341), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_remLo_365__FF_INPUT) );
  AND2X2 AND2X2_8256 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_366_), .Y(u2__abc_44228_n17343) );
  AND2X2 AND2X2_8257 ( .A(u2__abc_44228_n2972_bF_buf57), .B(u2_remLo_364_), .Y(u2__abc_44228_n17344) );
  AND2X2 AND2X2_8258 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17344), .Y(u2__abc_44228_n17345) );
  AND2X2 AND2X2_8259 ( .A(u2__abc_44228_n17346), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_remLo_366__FF_INPUT) );
  AND2X2 AND2X2_826 ( .A(u2__abc_44228_n3625), .B(u2__abc_44228_n3456), .Y(u2__abc_44228_n3626) );
  AND2X2 AND2X2_8260 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_367_), .Y(u2__abc_44228_n17348) );
  AND2X2 AND2X2_8261 ( .A(u2__abc_44228_n2972_bF_buf56), .B(u2_remLo_365_), .Y(u2__abc_44228_n17349) );
  AND2X2 AND2X2_8262 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17349), .Y(u2__abc_44228_n17350) );
  AND2X2 AND2X2_8263 ( .A(u2__abc_44228_n17351), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_remLo_367__FF_INPUT) );
  AND2X2 AND2X2_8264 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_368_), .Y(u2__abc_44228_n17353) );
  AND2X2 AND2X2_8265 ( .A(u2__abc_44228_n2972_bF_buf55), .B(u2_remLo_366_), .Y(u2__abc_44228_n17354) );
  AND2X2 AND2X2_8266 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17354), .Y(u2__abc_44228_n17355) );
  AND2X2 AND2X2_8267 ( .A(u2__abc_44228_n17356), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_remLo_368__FF_INPUT) );
  AND2X2 AND2X2_8268 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_369_), .Y(u2__abc_44228_n17358) );
  AND2X2 AND2X2_8269 ( .A(u2__abc_44228_n2972_bF_buf54), .B(u2_remLo_367_), .Y(u2__abc_44228_n17359) );
  AND2X2 AND2X2_827 ( .A(u2__abc_44228_n3450), .B(u2__abc_44228_n3626), .Y(u2__abc_44228_n3627_1) );
  AND2X2 AND2X2_8270 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17359), .Y(u2__abc_44228_n17360) );
  AND2X2 AND2X2_8271 ( .A(u2__abc_44228_n17361), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_remLo_369__FF_INPUT) );
  AND2X2 AND2X2_8272 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_370_), .Y(u2__abc_44228_n17363) );
  AND2X2 AND2X2_8273 ( .A(u2__abc_44228_n2972_bF_buf53), .B(u2_remLo_368_), .Y(u2__abc_44228_n17364) );
  AND2X2 AND2X2_8274 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17364), .Y(u2__abc_44228_n17365) );
  AND2X2 AND2X2_8275 ( .A(u2__abc_44228_n17366), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_remLo_370__FF_INPUT) );
  AND2X2 AND2X2_8276 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_371_), .Y(u2__abc_44228_n17368) );
  AND2X2 AND2X2_8277 ( .A(u2__abc_44228_n2972_bF_buf52), .B(u2_remLo_369_), .Y(u2__abc_44228_n17369) );
  AND2X2 AND2X2_8278 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17369), .Y(u2__abc_44228_n17370) );
  AND2X2 AND2X2_8279 ( .A(u2__abc_44228_n17371), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_remLo_371__FF_INPUT) );
  AND2X2 AND2X2_828 ( .A(u2__abc_44228_n3442), .B(u2__abc_44228_n3445), .Y(u2__abc_44228_n3628) );
  AND2X2 AND2X2_8280 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_372_), .Y(u2__abc_44228_n17373) );
  AND2X2 AND2X2_8281 ( .A(u2__abc_44228_n2972_bF_buf51), .B(u2_remLo_370_), .Y(u2__abc_44228_n17374) );
  AND2X2 AND2X2_8282 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17374), .Y(u2__abc_44228_n17375) );
  AND2X2 AND2X2_8283 ( .A(u2__abc_44228_n17376), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_remLo_372__FF_INPUT) );
  AND2X2 AND2X2_8284 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_373_), .Y(u2__abc_44228_n17378) );
  AND2X2 AND2X2_8285 ( .A(u2__abc_44228_n2972_bF_buf50), .B(u2_remLo_371_), .Y(u2__abc_44228_n17379) );
  AND2X2 AND2X2_8286 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17379), .Y(u2__abc_44228_n17380) );
  AND2X2 AND2X2_8287 ( .A(u2__abc_44228_n17381), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_remLo_373__FF_INPUT) );
  AND2X2 AND2X2_8288 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_374_), .Y(u2__abc_44228_n17383) );
  AND2X2 AND2X2_8289 ( .A(u2__abc_44228_n2972_bF_buf49), .B(u2_remLo_372_), .Y(u2__abc_44228_n17384) );
  AND2X2 AND2X2_829 ( .A(u2__abc_44228_n3630), .B(u2__abc_44228_n3436), .Y(u2__abc_44228_n3631) );
  AND2X2 AND2X2_8290 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17384), .Y(u2__abc_44228_n17385) );
  AND2X2 AND2X2_8291 ( .A(u2__abc_44228_n17386), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_remLo_374__FF_INPUT) );
  AND2X2 AND2X2_8292 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_375_), .Y(u2__abc_44228_n17388) );
  AND2X2 AND2X2_8293 ( .A(u2__abc_44228_n2972_bF_buf48), .B(u2_remLo_373_), .Y(u2__abc_44228_n17389) );
  AND2X2 AND2X2_8294 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17389), .Y(u2__abc_44228_n17390) );
  AND2X2 AND2X2_8295 ( .A(u2__abc_44228_n17391), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_remLo_375__FF_INPUT) );
  AND2X2 AND2X2_8296 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_376_), .Y(u2__abc_44228_n17393) );
  AND2X2 AND2X2_8297 ( .A(u2__abc_44228_n2972_bF_buf47), .B(u2_remLo_374_), .Y(u2__abc_44228_n17394) );
  AND2X2 AND2X2_8298 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17394), .Y(u2__abc_44228_n17395) );
  AND2X2 AND2X2_8299 ( .A(u2__abc_44228_n17396), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_remLo_376__FF_INPUT) );
  AND2X2 AND2X2_83 ( .A(_abc_64468_n849), .B(_abc_64468_n848), .Y(_auto_iopadmap_cc_313_execute_65414_118_) );
  AND2X2 AND2X2_830 ( .A(u2__abc_44228_n3632), .B(u2__abc_44228_n3430), .Y(u2__abc_44228_n3633) );
  AND2X2 AND2X2_8300 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_377_), .Y(u2__abc_44228_n17398) );
  AND2X2 AND2X2_8301 ( .A(u2__abc_44228_n2972_bF_buf46), .B(u2_remLo_375_), .Y(u2__abc_44228_n17399) );
  AND2X2 AND2X2_8302 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17399), .Y(u2__abc_44228_n17400) );
  AND2X2 AND2X2_8303 ( .A(u2__abc_44228_n17401), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_remLo_377__FF_INPUT) );
  AND2X2 AND2X2_8304 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_378_), .Y(u2__abc_44228_n17403) );
  AND2X2 AND2X2_8305 ( .A(u2__abc_44228_n2972_bF_buf45), .B(u2_remLo_376_), .Y(u2__abc_44228_n17404) );
  AND2X2 AND2X2_8306 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17404), .Y(u2__abc_44228_n17405) );
  AND2X2 AND2X2_8307 ( .A(u2__abc_44228_n17406), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_remLo_378__FF_INPUT) );
  AND2X2 AND2X2_8308 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_379_), .Y(u2__abc_44228_n17408) );
  AND2X2 AND2X2_8309 ( .A(u2__abc_44228_n2972_bF_buf44), .B(u2_remLo_377_), .Y(u2__abc_44228_n17409) );
  AND2X2 AND2X2_831 ( .A(u2__abc_44228_n3634), .B(u2__abc_44228_n3433), .Y(u2__abc_44228_n3635) );
  AND2X2 AND2X2_8310 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17409), .Y(u2__abc_44228_n17410) );
  AND2X2 AND2X2_8311 ( .A(u2__abc_44228_n17411), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_remLo_379__FF_INPUT) );
  AND2X2 AND2X2_8312 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_380_), .Y(u2__abc_44228_n17413) );
  AND2X2 AND2X2_8313 ( .A(u2__abc_44228_n2972_bF_buf43), .B(u2_remLo_378_), .Y(u2__abc_44228_n17414) );
  AND2X2 AND2X2_8314 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17414), .Y(u2__abc_44228_n17415) );
  AND2X2 AND2X2_8315 ( .A(u2__abc_44228_n17416), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_remLo_380__FF_INPUT) );
  AND2X2 AND2X2_8316 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_381_), .Y(u2__abc_44228_n17418) );
  AND2X2 AND2X2_8317 ( .A(u2__abc_44228_n2972_bF_buf42), .B(u2_remLo_379_), .Y(u2__abc_44228_n17419) );
  AND2X2 AND2X2_8318 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17419), .Y(u2__abc_44228_n17420) );
  AND2X2 AND2X2_8319 ( .A(u2__abc_44228_n17421), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_remLo_381__FF_INPUT) );
  AND2X2 AND2X2_832 ( .A(u2__abc_44228_n3635), .B(u2__abc_44228_n3421), .Y(u2__abc_44228_n3636) );
  AND2X2 AND2X2_8320 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_382_), .Y(u2__abc_44228_n17423) );
  AND2X2 AND2X2_8321 ( .A(u2__abc_44228_n2972_bF_buf41), .B(u2_remLo_380_), .Y(u2__abc_44228_n17424) );
  AND2X2 AND2X2_8322 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17424), .Y(u2__abc_44228_n17425) );
  AND2X2 AND2X2_8323 ( .A(u2__abc_44228_n17426), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_remLo_382__FF_INPUT) );
  AND2X2 AND2X2_8324 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_383_), .Y(u2__abc_44228_n17428) );
  AND2X2 AND2X2_8325 ( .A(u2__abc_44228_n2972_bF_buf40), .B(u2_remLo_381_), .Y(u2__abc_44228_n17429) );
  AND2X2 AND2X2_8326 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17429), .Y(u2__abc_44228_n17430) );
  AND2X2 AND2X2_8327 ( .A(u2__abc_44228_n17431), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_remLo_383__FF_INPUT) );
  AND2X2 AND2X2_8328 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_384_), .Y(u2__abc_44228_n17433) );
  AND2X2 AND2X2_8329 ( .A(u2__abc_44228_n2972_bF_buf39), .B(u2_remLo_382_), .Y(u2__abc_44228_n17434) );
  AND2X2 AND2X2_833 ( .A(u2__abc_44228_n3413), .B(u2__abc_44228_n3416), .Y(u2__abc_44228_n3637_1) );
  AND2X2 AND2X2_8330 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17434), .Y(u2__abc_44228_n17435) );
  AND2X2 AND2X2_8331 ( .A(u2__abc_44228_n17436), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_remLo_384__FF_INPUT) );
  AND2X2 AND2X2_8332 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_385_), .Y(u2__abc_44228_n17438) );
  AND2X2 AND2X2_8333 ( .A(u2__abc_44228_n2972_bF_buf38), .B(u2_remLo_383_), .Y(u2__abc_44228_n17439) );
  AND2X2 AND2X2_8334 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17439), .Y(u2__abc_44228_n17440) );
  AND2X2 AND2X2_8335 ( .A(u2__abc_44228_n17441), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_remLo_385__FF_INPUT) );
  AND2X2 AND2X2_8336 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_386_), .Y(u2__abc_44228_n17443) );
  AND2X2 AND2X2_8337 ( .A(u2__abc_44228_n2972_bF_buf37), .B(u2_remLo_384_), .Y(u2__abc_44228_n17444) );
  AND2X2 AND2X2_8338 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17444), .Y(u2__abc_44228_n17445) );
  AND2X2 AND2X2_8339 ( .A(u2__abc_44228_n17446), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_remLo_386__FF_INPUT) );
  AND2X2 AND2X2_834 ( .A(u2__abc_44228_n3640), .B(u2__abc_44228_n3407), .Y(u2__abc_44228_n3641) );
  AND2X2 AND2X2_8340 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_387_), .Y(u2__abc_44228_n17448) );
  AND2X2 AND2X2_8341 ( .A(u2__abc_44228_n2972_bF_buf36), .B(u2_remLo_385_), .Y(u2__abc_44228_n17449) );
  AND2X2 AND2X2_8342 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17449), .Y(u2__abc_44228_n17450) );
  AND2X2 AND2X2_8343 ( .A(u2__abc_44228_n17451), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_remLo_387__FF_INPUT) );
  AND2X2 AND2X2_8344 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_388_), .Y(u2__abc_44228_n17453) );
  AND2X2 AND2X2_8345 ( .A(u2__abc_44228_n2972_bF_buf35), .B(u2_remLo_386_), .Y(u2__abc_44228_n17454) );
  AND2X2 AND2X2_8346 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17454), .Y(u2__abc_44228_n17455) );
  AND2X2 AND2X2_8347 ( .A(u2__abc_44228_n17456), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_remLo_388__FF_INPUT) );
  AND2X2 AND2X2_8348 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_389_), .Y(u2__abc_44228_n17458) );
  AND2X2 AND2X2_8349 ( .A(u2__abc_44228_n2972_bF_buf34), .B(u2_remLo_387_), .Y(u2__abc_44228_n17459) );
  AND2X2 AND2X2_835 ( .A(u2__abc_44228_n3643), .B(u2__abc_44228_n3394), .Y(u2__abc_44228_n3644) );
  AND2X2 AND2X2_8350 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17459), .Y(u2__abc_44228_n17460) );
  AND2X2 AND2X2_8351 ( .A(u2__abc_44228_n17461), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_remLo_389__FF_INPUT) );
  AND2X2 AND2X2_8352 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_390_), .Y(u2__abc_44228_n17463) );
  AND2X2 AND2X2_8353 ( .A(u2__abc_44228_n2972_bF_buf33), .B(u2_remLo_388_), .Y(u2__abc_44228_n17464) );
  AND2X2 AND2X2_8354 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17464), .Y(u2__abc_44228_n17465) );
  AND2X2 AND2X2_8355 ( .A(u2__abc_44228_n17466), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_remLo_390__FF_INPUT) );
  AND2X2 AND2X2_8356 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_391_), .Y(u2__abc_44228_n17468) );
  AND2X2 AND2X2_8357 ( .A(u2__abc_44228_n2972_bF_buf32), .B(u2_remLo_389_), .Y(u2__abc_44228_n17469) );
  AND2X2 AND2X2_8358 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17469), .Y(u2__abc_44228_n17470) );
  AND2X2 AND2X2_8359 ( .A(u2__abc_44228_n17471), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_remLo_391__FF_INPUT) );
  AND2X2 AND2X2_836 ( .A(u2__abc_44228_n3645), .B(u2__abc_44228_n3391), .Y(u2__abc_44228_n3646) );
  AND2X2 AND2X2_8360 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_392_), .Y(u2__abc_44228_n17473) );
  AND2X2 AND2X2_8361 ( .A(u2__abc_44228_n2972_bF_buf31), .B(u2_remLo_390_), .Y(u2__abc_44228_n17474) );
  AND2X2 AND2X2_8362 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17474), .Y(u2__abc_44228_n17475) );
  AND2X2 AND2X2_8363 ( .A(u2__abc_44228_n17476), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_remLo_392__FF_INPUT) );
  AND2X2 AND2X2_8364 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_393_), .Y(u2__abc_44228_n17478) );
  AND2X2 AND2X2_8365 ( .A(u2__abc_44228_n2972_bF_buf30), .B(u2_remLo_391_), .Y(u2__abc_44228_n17479) );
  AND2X2 AND2X2_8366 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17479), .Y(u2__abc_44228_n17480) );
  AND2X2 AND2X2_8367 ( .A(u2__abc_44228_n17481), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_remLo_393__FF_INPUT) );
  AND2X2 AND2X2_8368 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_394_), .Y(u2__abc_44228_n17483) );
  AND2X2 AND2X2_8369 ( .A(u2__abc_44228_n2972_bF_buf29), .B(u2_remLo_392_), .Y(u2__abc_44228_n17484) );
  AND2X2 AND2X2_837 ( .A(u2__abc_44228_n3380), .B(u2__abc_44228_n3647_1), .Y(u2__abc_44228_n3648) );
  AND2X2 AND2X2_8370 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17484), .Y(u2__abc_44228_n17485) );
  AND2X2 AND2X2_8371 ( .A(u2__abc_44228_n17486), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_remLo_394__FF_INPUT) );
  AND2X2 AND2X2_8372 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_395_), .Y(u2__abc_44228_n17488) );
  AND2X2 AND2X2_8373 ( .A(u2__abc_44228_n2972_bF_buf28), .B(u2_remLo_393_), .Y(u2__abc_44228_n17489) );
  AND2X2 AND2X2_8374 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17489), .Y(u2__abc_44228_n17490) );
  AND2X2 AND2X2_8375 ( .A(u2__abc_44228_n17491), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_remLo_395__FF_INPUT) );
  AND2X2 AND2X2_8376 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_396_), .Y(u2__abc_44228_n17493) );
  AND2X2 AND2X2_8377 ( .A(u2__abc_44228_n2972_bF_buf27), .B(u2_remLo_394_), .Y(u2__abc_44228_n17494) );
  AND2X2 AND2X2_8378 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17494), .Y(u2__abc_44228_n17495) );
  AND2X2 AND2X2_8379 ( .A(u2__abc_44228_n17496), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_remLo_396__FF_INPUT) );
  AND2X2 AND2X2_838 ( .A(u2__abc_44228_n3649), .B(u2__abc_44228_n3383), .Y(u2__abc_44228_n3650) );
  AND2X2 AND2X2_8380 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_397_), .Y(u2__abc_44228_n17498) );
  AND2X2 AND2X2_8381 ( .A(u2__abc_44228_n2972_bF_buf26), .B(u2_remLo_395_), .Y(u2__abc_44228_n17499) );
  AND2X2 AND2X2_8382 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17499), .Y(u2__abc_44228_n17500) );
  AND2X2 AND2X2_8383 ( .A(u2__abc_44228_n17501), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_remLo_397__FF_INPUT) );
  AND2X2 AND2X2_8384 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_398_), .Y(u2__abc_44228_n17503) );
  AND2X2 AND2X2_8385 ( .A(u2__abc_44228_n2972_bF_buf25), .B(u2_remLo_396_), .Y(u2__abc_44228_n17504) );
  AND2X2 AND2X2_8386 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17504), .Y(u2__abc_44228_n17505) );
  AND2X2 AND2X2_8387 ( .A(u2__abc_44228_n17506), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_remLo_398__FF_INPUT) );
  AND2X2 AND2X2_8388 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_399_), .Y(u2__abc_44228_n17508) );
  AND2X2 AND2X2_8389 ( .A(u2__abc_44228_n2972_bF_buf24), .B(u2_remLo_397_), .Y(u2__abc_44228_n17509) );
  AND2X2 AND2X2_839 ( .A(u2__abc_44228_n3651), .B(u2__abc_44228_n3377), .Y(u2__abc_44228_n3652) );
  AND2X2 AND2X2_8390 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17509), .Y(u2__abc_44228_n17510) );
  AND2X2 AND2X2_8391 ( .A(u2__abc_44228_n17511), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_remLo_399__FF_INPUT) );
  AND2X2 AND2X2_8392 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_400_), .Y(u2__abc_44228_n17513) );
  AND2X2 AND2X2_8393 ( .A(u2__abc_44228_n2972_bF_buf23), .B(u2_remLo_398_), .Y(u2__abc_44228_n17514) );
  AND2X2 AND2X2_8394 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17514), .Y(u2__abc_44228_n17515) );
  AND2X2 AND2X2_8395 ( .A(u2__abc_44228_n17516), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_remLo_400__FF_INPUT) );
  AND2X2 AND2X2_8396 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_401_), .Y(u2__abc_44228_n17518) );
  AND2X2 AND2X2_8397 ( .A(u2__abc_44228_n2972_bF_buf22), .B(u2_remLo_399_), .Y(u2__abc_44228_n17519) );
  AND2X2 AND2X2_8398 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17519), .Y(u2__abc_44228_n17520) );
  AND2X2 AND2X2_8399 ( .A(u2__abc_44228_n17521), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_remLo_401__FF_INPUT) );
  AND2X2 AND2X2_84 ( .A(_abc_64468_n852), .B(_abc_64468_n851), .Y(_auto_iopadmap_cc_313_execute_65414_119_) );
  AND2X2 AND2X2_840 ( .A(u2__abc_44228_n3354), .B(u2__abc_44228_n3357), .Y(u2__abc_44228_n3653) );
  AND2X2 AND2X2_8400 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_402_), .Y(u2__abc_44228_n17523) );
  AND2X2 AND2X2_8401 ( .A(u2__abc_44228_n2972_bF_buf21), .B(u2_remLo_400_), .Y(u2__abc_44228_n17524) );
  AND2X2 AND2X2_8402 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17524), .Y(u2__abc_44228_n17525) );
  AND2X2 AND2X2_8403 ( .A(u2__abc_44228_n17526), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_remLo_402__FF_INPUT) );
  AND2X2 AND2X2_8404 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_403_), .Y(u2__abc_44228_n17528) );
  AND2X2 AND2X2_8405 ( .A(u2__abc_44228_n2972_bF_buf20), .B(u2_remLo_401_), .Y(u2__abc_44228_n17529) );
  AND2X2 AND2X2_8406 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17529), .Y(u2__abc_44228_n17530) );
  AND2X2 AND2X2_8407 ( .A(u2__abc_44228_n17531), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_remLo_403__FF_INPUT) );
  AND2X2 AND2X2_8408 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_404_), .Y(u2__abc_44228_n17533) );
  AND2X2 AND2X2_8409 ( .A(u2__abc_44228_n2972_bF_buf19), .B(u2_remLo_402_), .Y(u2__abc_44228_n17534) );
  AND2X2 AND2X2_841 ( .A(u2__abc_44228_n3655), .B(u2__abc_44228_n3371), .Y(u2__abc_44228_n3656_1) );
  AND2X2 AND2X2_8410 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17534), .Y(u2__abc_44228_n17535) );
  AND2X2 AND2X2_8411 ( .A(u2__abc_44228_n17536), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_remLo_404__FF_INPUT) );
  AND2X2 AND2X2_8412 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_405_), .Y(u2__abc_44228_n17538) );
  AND2X2 AND2X2_8413 ( .A(u2__abc_44228_n2972_bF_buf18), .B(u2_remLo_403_), .Y(u2__abc_44228_n17539) );
  AND2X2 AND2X2_8414 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17539), .Y(u2__abc_44228_n17540) );
  AND2X2 AND2X2_8415 ( .A(u2__abc_44228_n17541), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_remLo_405__FF_INPUT) );
  AND2X2 AND2X2_8416 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_406_), .Y(u2__abc_44228_n17543) );
  AND2X2 AND2X2_8417 ( .A(u2__abc_44228_n2972_bF_buf17), .B(u2_remLo_404_), .Y(u2__abc_44228_n17544) );
  AND2X2 AND2X2_8418 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17544), .Y(u2__abc_44228_n17545) );
  AND2X2 AND2X2_8419 ( .A(u2__abc_44228_n17546), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_remLo_406__FF_INPUT) );
  AND2X2 AND2X2_842 ( .A(u2__abc_44228_n3657), .B(u2__abc_44228_n3374), .Y(u2__abc_44228_n3658) );
  AND2X2 AND2X2_8420 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_407_), .Y(u2__abc_44228_n17548) );
  AND2X2 AND2X2_8421 ( .A(u2__abc_44228_n2972_bF_buf16), .B(u2_remLo_405_), .Y(u2__abc_44228_n17549) );
  AND2X2 AND2X2_8422 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17549), .Y(u2__abc_44228_n17550) );
  AND2X2 AND2X2_8423 ( .A(u2__abc_44228_n17551), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_remLo_407__FF_INPUT) );
  AND2X2 AND2X2_8424 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_408_), .Y(u2__abc_44228_n17553) );
  AND2X2 AND2X2_8425 ( .A(u2__abc_44228_n2972_bF_buf15), .B(u2_remLo_406_), .Y(u2__abc_44228_n17554) );
  AND2X2 AND2X2_8426 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17554), .Y(u2__abc_44228_n17555) );
  AND2X2 AND2X2_8427 ( .A(u2__abc_44228_n17556), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_remLo_408__FF_INPUT) );
  AND2X2 AND2X2_8428 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_409_), .Y(u2__abc_44228_n17558) );
  AND2X2 AND2X2_8429 ( .A(u2__abc_44228_n2972_bF_buf14), .B(u2_remLo_407_), .Y(u2__abc_44228_n17559) );
  AND2X2 AND2X2_843 ( .A(u2__abc_44228_n3658), .B(u2__abc_44228_n3362), .Y(u2__abc_44228_n3659) );
  AND2X2 AND2X2_8430 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17559), .Y(u2__abc_44228_n17560) );
  AND2X2 AND2X2_8431 ( .A(u2__abc_44228_n17561), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_remLo_409__FF_INPUT) );
  AND2X2 AND2X2_8432 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_410_), .Y(u2__abc_44228_n17563) );
  AND2X2 AND2X2_8433 ( .A(u2__abc_44228_n2972_bF_buf13), .B(u2_remLo_408_), .Y(u2__abc_44228_n17564) );
  AND2X2 AND2X2_8434 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17564), .Y(u2__abc_44228_n17565) );
  AND2X2 AND2X2_8435 ( .A(u2__abc_44228_n17566), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_remLo_410__FF_INPUT) );
  AND2X2 AND2X2_8436 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_411_), .Y(u2__abc_44228_n17568) );
  AND2X2 AND2X2_8437 ( .A(u2__abc_44228_n2972_bF_buf12), .B(u2_remLo_409_), .Y(u2__abc_44228_n17569) );
  AND2X2 AND2X2_8438 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17569), .Y(u2__abc_44228_n17570) );
  AND2X2 AND2X2_8439 ( .A(u2__abc_44228_n17571), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_remLo_411__FF_INPUT) );
  AND2X2 AND2X2_844 ( .A(u2__abc_44228_n3665), .B(u2_remHi_125_), .Y(u2__abc_44228_n3666_1) );
  AND2X2 AND2X2_8440 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_412_), .Y(u2__abc_44228_n17573) );
  AND2X2 AND2X2_8441 ( .A(u2__abc_44228_n2972_bF_buf11), .B(u2_remLo_410_), .Y(u2__abc_44228_n17574) );
  AND2X2 AND2X2_8442 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17574), .Y(u2__abc_44228_n17575) );
  AND2X2 AND2X2_8443 ( .A(u2__abc_44228_n17576), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_remLo_412__FF_INPUT) );
  AND2X2 AND2X2_8444 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_413_), .Y(u2__abc_44228_n17578) );
  AND2X2 AND2X2_8445 ( .A(u2__abc_44228_n2972_bF_buf10), .B(u2_remLo_411_), .Y(u2__abc_44228_n17579) );
  AND2X2 AND2X2_8446 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17579), .Y(u2__abc_44228_n17580) );
  AND2X2 AND2X2_8447 ( .A(u2__abc_44228_n17581), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_remLo_413__FF_INPUT) );
  AND2X2 AND2X2_8448 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_414_), .Y(u2__abc_44228_n17583) );
  AND2X2 AND2X2_8449 ( .A(u2__abc_44228_n2972_bF_buf9), .B(u2_remLo_412_), .Y(u2__abc_44228_n17584) );
  AND2X2 AND2X2_845 ( .A(u2__abc_44228_n3668), .B(sqrto_125_), .Y(u2__abc_44228_n3669) );
  AND2X2 AND2X2_8450 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17584), .Y(u2__abc_44228_n17585) );
  AND2X2 AND2X2_8451 ( .A(u2__abc_44228_n17586), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_remLo_414__FF_INPUT) );
  AND2X2 AND2X2_8452 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_415_), .Y(u2__abc_44228_n17588) );
  AND2X2 AND2X2_8453 ( .A(u2__abc_44228_n2972_bF_buf8), .B(u2_remLo_413_), .Y(u2__abc_44228_n17589) );
  AND2X2 AND2X2_8454 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17589), .Y(u2__abc_44228_n17590) );
  AND2X2 AND2X2_8455 ( .A(u2__abc_44228_n17591), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_remLo_415__FF_INPUT) );
  AND2X2 AND2X2_8456 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_416_), .Y(u2__abc_44228_n17593) );
  AND2X2 AND2X2_8457 ( .A(u2__abc_44228_n2972_bF_buf7), .B(u2_remLo_414_), .Y(u2__abc_44228_n17594) );
  AND2X2 AND2X2_8458 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17594), .Y(u2__abc_44228_n17595) );
  AND2X2 AND2X2_8459 ( .A(u2__abc_44228_n17596), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_remLo_416__FF_INPUT) );
  AND2X2 AND2X2_846 ( .A(u2__abc_44228_n3667), .B(u2__abc_44228_n3670), .Y(u2__abc_44228_n3671) );
  AND2X2 AND2X2_8460 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_417_), .Y(u2__abc_44228_n17598) );
  AND2X2 AND2X2_8461 ( .A(u2__abc_44228_n2972_bF_buf6), .B(u2_remLo_415_), .Y(u2__abc_44228_n17599) );
  AND2X2 AND2X2_8462 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17599), .Y(u2__abc_44228_n17600) );
  AND2X2 AND2X2_8463 ( .A(u2__abc_44228_n17601), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_remLo_417__FF_INPUT) );
  AND2X2 AND2X2_8464 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_418_), .Y(u2__abc_44228_n17603) );
  AND2X2 AND2X2_8465 ( .A(u2__abc_44228_n2972_bF_buf5), .B(u2_remLo_416_), .Y(u2__abc_44228_n17604) );
  AND2X2 AND2X2_8466 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17604), .Y(u2__abc_44228_n17605) );
  AND2X2 AND2X2_8467 ( .A(u2__abc_44228_n17606), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_remLo_418__FF_INPUT) );
  AND2X2 AND2X2_8468 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_419_), .Y(u2__abc_44228_n17608) );
  AND2X2 AND2X2_8469 ( .A(u2__abc_44228_n2972_bF_buf4), .B(u2_remLo_417_), .Y(u2__abc_44228_n17609) );
  AND2X2 AND2X2_847 ( .A(u2__abc_44228_n3672), .B(u2_remHi_124_), .Y(u2__abc_44228_n3673) );
  AND2X2 AND2X2_8470 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17609), .Y(u2__abc_44228_n17610) );
  AND2X2 AND2X2_8471 ( .A(u2__abc_44228_n17611), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_remLo_419__FF_INPUT) );
  AND2X2 AND2X2_8472 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_420_), .Y(u2__abc_44228_n17613) );
  AND2X2 AND2X2_8473 ( .A(u2__abc_44228_n2972_bF_buf3), .B(u2_remLo_418_), .Y(u2__abc_44228_n17614) );
  AND2X2 AND2X2_8474 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17614), .Y(u2__abc_44228_n17615) );
  AND2X2 AND2X2_8475 ( .A(u2__abc_44228_n17616), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_remLo_420__FF_INPUT) );
  AND2X2 AND2X2_8476 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_421_), .Y(u2__abc_44228_n17618) );
  AND2X2 AND2X2_8477 ( .A(u2__abc_44228_n2972_bF_buf2), .B(u2_remLo_419_), .Y(u2__abc_44228_n17619) );
  AND2X2 AND2X2_8478 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17619), .Y(u2__abc_44228_n17620) );
  AND2X2 AND2X2_8479 ( .A(u2__abc_44228_n17621), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_remLo_421__FF_INPUT) );
  AND2X2 AND2X2_848 ( .A(u2__abc_44228_n3674), .B(sqrto_124_), .Y(u2__abc_44228_n3675_1) );
  AND2X2 AND2X2_8480 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_422_), .Y(u2__abc_44228_n17623) );
  AND2X2 AND2X2_8481 ( .A(u2__abc_44228_n2972_bF_buf1), .B(u2_remLo_420_), .Y(u2__abc_44228_n17624) );
  AND2X2 AND2X2_8482 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17624), .Y(u2__abc_44228_n17625) );
  AND2X2 AND2X2_8483 ( .A(u2__abc_44228_n17626), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_remLo_422__FF_INPUT) );
  AND2X2 AND2X2_8484 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_423_), .Y(u2__abc_44228_n17628) );
  AND2X2 AND2X2_8485 ( .A(u2__abc_44228_n2972_bF_buf0), .B(u2_remLo_421_), .Y(u2__abc_44228_n17629) );
  AND2X2 AND2X2_8486 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17629), .Y(u2__abc_44228_n17630) );
  AND2X2 AND2X2_8487 ( .A(u2__abc_44228_n17631), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_remLo_423__FF_INPUT) );
  AND2X2 AND2X2_8488 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_424_), .Y(u2__abc_44228_n17633) );
  AND2X2 AND2X2_8489 ( .A(u2__abc_44228_n2972_bF_buf107), .B(u2_remLo_422_), .Y(u2__abc_44228_n17634) );
  AND2X2 AND2X2_849 ( .A(u2__abc_44228_n3677), .B(u2__abc_44228_n3671), .Y(u2__abc_44228_n3678) );
  AND2X2 AND2X2_8490 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17634), .Y(u2__abc_44228_n17635) );
  AND2X2 AND2X2_8491 ( .A(u2__abc_44228_n17636), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_remLo_424__FF_INPUT) );
  AND2X2 AND2X2_8492 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_425_), .Y(u2__abc_44228_n17638) );
  AND2X2 AND2X2_8493 ( .A(u2__abc_44228_n2972_bF_buf106), .B(u2_remLo_423_), .Y(u2__abc_44228_n17639) );
  AND2X2 AND2X2_8494 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17639), .Y(u2__abc_44228_n17640) );
  AND2X2 AND2X2_8495 ( .A(u2__abc_44228_n17641), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_remLo_425__FF_INPUT) );
  AND2X2 AND2X2_8496 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_426_), .Y(u2__abc_44228_n17643) );
  AND2X2 AND2X2_8497 ( .A(u2__abc_44228_n2972_bF_buf105), .B(u2_remLo_424_), .Y(u2__abc_44228_n17644) );
  AND2X2 AND2X2_8498 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17644), .Y(u2__abc_44228_n17645) );
  AND2X2 AND2X2_8499 ( .A(u2__abc_44228_n17646), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_remLo_426__FF_INPUT) );
  AND2X2 AND2X2_85 ( .A(_abc_64468_n855), .B(_abc_64468_n854), .Y(_auto_iopadmap_cc_313_execute_65414_120_) );
  AND2X2 AND2X2_850 ( .A(u2__abc_44228_n3679), .B(u2_remHi_122_), .Y(u2__abc_44228_n3680) );
  AND2X2 AND2X2_8500 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_427_), .Y(u2__abc_44228_n17648) );
  AND2X2 AND2X2_8501 ( .A(u2__abc_44228_n2972_bF_buf104), .B(u2_remLo_425_), .Y(u2__abc_44228_n17649) );
  AND2X2 AND2X2_8502 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17649), .Y(u2__abc_44228_n17650) );
  AND2X2 AND2X2_8503 ( .A(u2__abc_44228_n17651), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_remLo_427__FF_INPUT) );
  AND2X2 AND2X2_8504 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_428_), .Y(u2__abc_44228_n17653) );
  AND2X2 AND2X2_8505 ( .A(u2__abc_44228_n2972_bF_buf103), .B(u2_remLo_426_), .Y(u2__abc_44228_n17654) );
  AND2X2 AND2X2_8506 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17654), .Y(u2__abc_44228_n17655) );
  AND2X2 AND2X2_8507 ( .A(u2__abc_44228_n17656), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_remLo_428__FF_INPUT) );
  AND2X2 AND2X2_8508 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_429_), .Y(u2__abc_44228_n17658) );
  AND2X2 AND2X2_8509 ( .A(u2__abc_44228_n2972_bF_buf102), .B(u2_remLo_427_), .Y(u2__abc_44228_n17659) );
  AND2X2 AND2X2_851 ( .A(u2__abc_44228_n3681), .B(sqrto_122_), .Y(u2__abc_44228_n3682) );
  AND2X2 AND2X2_8510 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17659), .Y(u2__abc_44228_n17660) );
  AND2X2 AND2X2_8511 ( .A(u2__abc_44228_n17661), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_remLo_429__FF_INPUT) );
  AND2X2 AND2X2_8512 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_430_), .Y(u2__abc_44228_n17663) );
  AND2X2 AND2X2_8513 ( .A(u2__abc_44228_n2972_bF_buf101), .B(u2_remLo_428_), .Y(u2__abc_44228_n17664) );
  AND2X2 AND2X2_8514 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17664), .Y(u2__abc_44228_n17665) );
  AND2X2 AND2X2_8515 ( .A(u2__abc_44228_n17666), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_remLo_430__FF_INPUT) );
  AND2X2 AND2X2_8516 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_431_), .Y(u2__abc_44228_n17668) );
  AND2X2 AND2X2_8517 ( .A(u2__abc_44228_n2972_bF_buf100), .B(u2_remLo_429_), .Y(u2__abc_44228_n17669) );
  AND2X2 AND2X2_8518 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17669), .Y(u2__abc_44228_n17670) );
  AND2X2 AND2X2_8519 ( .A(u2__abc_44228_n17671), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_remLo_431__FF_INPUT) );
  AND2X2 AND2X2_852 ( .A(u2__abc_44228_n3685_1), .B(u2_remHi_123_), .Y(u2__abc_44228_n3686) );
  AND2X2 AND2X2_8520 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_432_), .Y(u2__abc_44228_n17673) );
  AND2X2 AND2X2_8521 ( .A(u2__abc_44228_n2972_bF_buf99), .B(u2_remLo_430_), .Y(u2__abc_44228_n17674) );
  AND2X2 AND2X2_8522 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17674), .Y(u2__abc_44228_n17675) );
  AND2X2 AND2X2_8523 ( .A(u2__abc_44228_n17676), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_remLo_432__FF_INPUT) );
  AND2X2 AND2X2_8524 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_433_), .Y(u2__abc_44228_n17678) );
  AND2X2 AND2X2_8525 ( .A(u2__abc_44228_n2972_bF_buf98), .B(u2_remLo_431_), .Y(u2__abc_44228_n17679) );
  AND2X2 AND2X2_8526 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17679), .Y(u2__abc_44228_n17680) );
  AND2X2 AND2X2_8527 ( .A(u2__abc_44228_n17681), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_remLo_433__FF_INPUT) );
  AND2X2 AND2X2_8528 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_434_), .Y(u2__abc_44228_n17683) );
  AND2X2 AND2X2_8529 ( .A(u2__abc_44228_n2972_bF_buf97), .B(u2_remLo_432_), .Y(u2__abc_44228_n17684) );
  AND2X2 AND2X2_853 ( .A(u2__abc_44228_n3688), .B(sqrto_123_), .Y(u2__abc_44228_n3689) );
  AND2X2 AND2X2_8530 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17684), .Y(u2__abc_44228_n17685) );
  AND2X2 AND2X2_8531 ( .A(u2__abc_44228_n17686), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_remLo_434__FF_INPUT) );
  AND2X2 AND2X2_8532 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remLo_435_), .Y(u2__abc_44228_n17688) );
  AND2X2 AND2X2_8533 ( .A(u2__abc_44228_n2972_bF_buf96), .B(u2_remLo_433_), .Y(u2__abc_44228_n17689) );
  AND2X2 AND2X2_8534 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17689), .Y(u2__abc_44228_n17690) );
  AND2X2 AND2X2_8535 ( .A(u2__abc_44228_n17691), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_remLo_435__FF_INPUT) );
  AND2X2 AND2X2_8536 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remLo_436_), .Y(u2__abc_44228_n17693) );
  AND2X2 AND2X2_8537 ( .A(u2__abc_44228_n2972_bF_buf95), .B(u2_remLo_434_), .Y(u2__abc_44228_n17694) );
  AND2X2 AND2X2_8538 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17694), .Y(u2__abc_44228_n17695) );
  AND2X2 AND2X2_8539 ( .A(u2__abc_44228_n17696), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_remLo_436__FF_INPUT) );
  AND2X2 AND2X2_854 ( .A(u2__abc_44228_n3687), .B(u2__abc_44228_n3690), .Y(u2__abc_44228_n3691) );
  AND2X2 AND2X2_8540 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2_remLo_437_), .Y(u2__abc_44228_n17698) );
  AND2X2 AND2X2_8541 ( .A(u2__abc_44228_n2972_bF_buf94), .B(u2_remLo_435_), .Y(u2__abc_44228_n17699) );
  AND2X2 AND2X2_8542 ( .A(u2__abc_44228_n2984_bF_buf12), .B(u2__abc_44228_n17699), .Y(u2__abc_44228_n17700) );
  AND2X2 AND2X2_8543 ( .A(u2__abc_44228_n17701), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_remLo_437__FF_INPUT) );
  AND2X2 AND2X2_8544 ( .A(u2__abc_44228_n15247_bF_buf12), .B(u2_remLo_438_), .Y(u2__abc_44228_n17703) );
  AND2X2 AND2X2_8545 ( .A(u2__abc_44228_n2972_bF_buf93), .B(u2_remLo_436_), .Y(u2__abc_44228_n17704) );
  AND2X2 AND2X2_8546 ( .A(u2__abc_44228_n2984_bF_buf11), .B(u2__abc_44228_n17704), .Y(u2__abc_44228_n17705) );
  AND2X2 AND2X2_8547 ( .A(u2__abc_44228_n17706), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_remLo_438__FF_INPUT) );
  AND2X2 AND2X2_8548 ( .A(u2__abc_44228_n15247_bF_buf11), .B(u2_remLo_439_), .Y(u2__abc_44228_n17708) );
  AND2X2 AND2X2_8549 ( .A(u2__abc_44228_n2972_bF_buf92), .B(u2_remLo_437_), .Y(u2__abc_44228_n17709) );
  AND2X2 AND2X2_855 ( .A(u2__abc_44228_n3684), .B(u2__abc_44228_n3691), .Y(u2__abc_44228_n3692) );
  AND2X2 AND2X2_8550 ( .A(u2__abc_44228_n2984_bF_buf10), .B(u2__abc_44228_n17709), .Y(u2__abc_44228_n17710) );
  AND2X2 AND2X2_8551 ( .A(u2__abc_44228_n17711), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_remLo_439__FF_INPUT) );
  AND2X2 AND2X2_8552 ( .A(u2__abc_44228_n15247_bF_buf10), .B(u2_remLo_440_), .Y(u2__abc_44228_n17713) );
  AND2X2 AND2X2_8553 ( .A(u2__abc_44228_n2972_bF_buf91), .B(u2_remLo_438_), .Y(u2__abc_44228_n17714) );
  AND2X2 AND2X2_8554 ( .A(u2__abc_44228_n2984_bF_buf9), .B(u2__abc_44228_n17714), .Y(u2__abc_44228_n17715) );
  AND2X2 AND2X2_8555 ( .A(u2__abc_44228_n17716), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_remLo_440__FF_INPUT) );
  AND2X2 AND2X2_8556 ( .A(u2__abc_44228_n15247_bF_buf9), .B(u2_remLo_441_), .Y(u2__abc_44228_n17718) );
  AND2X2 AND2X2_8557 ( .A(u2__abc_44228_n2972_bF_buf90), .B(u2_remLo_439_), .Y(u2__abc_44228_n17719) );
  AND2X2 AND2X2_8558 ( .A(u2__abc_44228_n2984_bF_buf8), .B(u2__abc_44228_n17719), .Y(u2__abc_44228_n17720) );
  AND2X2 AND2X2_8559 ( .A(u2__abc_44228_n17721), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_remLo_441__FF_INPUT) );
  AND2X2 AND2X2_856 ( .A(u2__abc_44228_n3678), .B(u2__abc_44228_n3692), .Y(u2__abc_44228_n3693) );
  AND2X2 AND2X2_8560 ( .A(u2__abc_44228_n15247_bF_buf8), .B(u2_remLo_442_), .Y(u2__abc_44228_n17723) );
  AND2X2 AND2X2_8561 ( .A(u2__abc_44228_n2972_bF_buf89), .B(u2_remLo_440_), .Y(u2__abc_44228_n17724) );
  AND2X2 AND2X2_8562 ( .A(u2__abc_44228_n2984_bF_buf7), .B(u2__abc_44228_n17724), .Y(u2__abc_44228_n17725) );
  AND2X2 AND2X2_8563 ( .A(u2__abc_44228_n17726), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_remLo_442__FF_INPUT) );
  AND2X2 AND2X2_8564 ( .A(u2__abc_44228_n15247_bF_buf7), .B(u2_remLo_443_), .Y(u2__abc_44228_n17728) );
  AND2X2 AND2X2_8565 ( .A(u2__abc_44228_n2972_bF_buf88), .B(u2_remLo_441_), .Y(u2__abc_44228_n17729) );
  AND2X2 AND2X2_8566 ( .A(u2__abc_44228_n2984_bF_buf6), .B(u2__abc_44228_n17729), .Y(u2__abc_44228_n17730) );
  AND2X2 AND2X2_8567 ( .A(u2__abc_44228_n17731), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_remLo_443__FF_INPUT) );
  AND2X2 AND2X2_8568 ( .A(u2__abc_44228_n15247_bF_buf6), .B(u2_remLo_444_), .Y(u2__abc_44228_n17733) );
  AND2X2 AND2X2_8569 ( .A(u2__abc_44228_n2972_bF_buf87), .B(u2_remLo_442_), .Y(u2__abc_44228_n17734) );
  AND2X2 AND2X2_857 ( .A(u2__abc_44228_n3694_1), .B(u2_remHi_119_), .Y(u2__abc_44228_n3695) );
  AND2X2 AND2X2_8570 ( .A(u2__abc_44228_n2984_bF_buf5), .B(u2__abc_44228_n17734), .Y(u2__abc_44228_n17735) );
  AND2X2 AND2X2_8571 ( .A(u2__abc_44228_n17736), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_remLo_444__FF_INPUT) );
  AND2X2 AND2X2_8572 ( .A(u2__abc_44228_n15247_bF_buf5), .B(u2_remLo_445_), .Y(u2__abc_44228_n17738) );
  AND2X2 AND2X2_8573 ( .A(u2__abc_44228_n2972_bF_buf86), .B(u2_remLo_443_), .Y(u2__abc_44228_n17739) );
  AND2X2 AND2X2_8574 ( .A(u2__abc_44228_n2984_bF_buf4), .B(u2__abc_44228_n17739), .Y(u2__abc_44228_n17740) );
  AND2X2 AND2X2_8575 ( .A(u2__abc_44228_n17741), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_remLo_445__FF_INPUT) );
  AND2X2 AND2X2_8576 ( .A(u2__abc_44228_n15247_bF_buf4), .B(u2_remLo_446_), .Y(u2__abc_44228_n17743) );
  AND2X2 AND2X2_8577 ( .A(u2__abc_44228_n2972_bF_buf85), .B(u2_remLo_444_), .Y(u2__abc_44228_n17744) );
  AND2X2 AND2X2_8578 ( .A(u2__abc_44228_n2984_bF_buf3), .B(u2__abc_44228_n17744), .Y(u2__abc_44228_n17745) );
  AND2X2 AND2X2_8579 ( .A(u2__abc_44228_n17746), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_remLo_446__FF_INPUT) );
  AND2X2 AND2X2_858 ( .A(u2__abc_44228_n3697), .B(sqrto_119_), .Y(u2__abc_44228_n3698) );
  AND2X2 AND2X2_8580 ( .A(u2__abc_44228_n15247_bF_buf3), .B(u2_remLo_447_), .Y(u2__abc_44228_n17748) );
  AND2X2 AND2X2_8581 ( .A(u2__abc_44228_n2972_bF_buf84), .B(u2_remLo_445_), .Y(u2__abc_44228_n17749) );
  AND2X2 AND2X2_8582 ( .A(u2__abc_44228_n2984_bF_buf2), .B(u2__abc_44228_n17749), .Y(u2__abc_44228_n17750) );
  AND2X2 AND2X2_8583 ( .A(u2__abc_44228_n17751), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_remLo_447__FF_INPUT) );
  AND2X2 AND2X2_8584 ( .A(u2__abc_44228_n15247_bF_buf2), .B(u2_remLo_448_), .Y(u2__abc_44228_n17753) );
  AND2X2 AND2X2_8585 ( .A(u2__abc_44228_n2972_bF_buf83), .B(u2_remLo_446_), .Y(u2__abc_44228_n17754) );
  AND2X2 AND2X2_8586 ( .A(u2__abc_44228_n2984_bF_buf1), .B(u2__abc_44228_n17754), .Y(u2__abc_44228_n17755) );
  AND2X2 AND2X2_8587 ( .A(u2__abc_44228_n17756), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_remLo_448__FF_INPUT) );
  AND2X2 AND2X2_8588 ( .A(u2__abc_44228_n15247_bF_buf1), .B(u2_remLo_449_), .Y(u2__abc_44228_n17758) );
  AND2X2 AND2X2_8589 ( .A(u2__abc_44228_n2972_bF_buf82), .B(u2_remLo_447_), .Y(u2__abc_44228_n17759) );
  AND2X2 AND2X2_859 ( .A(u2__abc_44228_n3696), .B(u2__abc_44228_n3699), .Y(u2__abc_44228_n3700) );
  AND2X2 AND2X2_8590 ( .A(u2__abc_44228_n2984_bF_buf0), .B(u2__abc_44228_n17759), .Y(u2__abc_44228_n17760) );
  AND2X2 AND2X2_8591 ( .A(u2__abc_44228_n17761), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_remLo_449__FF_INPUT) );
  AND2X2 AND2X2_8592 ( .A(u2__abc_44228_n15247_bF_buf0), .B(u2_remHiShift_0_), .Y(u2__abc_44228_n17763) );
  AND2X2 AND2X2_8593 ( .A(u2__abc_44228_n2972_bF_buf81), .B(u2_remLo_448_), .Y(u2__abc_44228_n17764) );
  AND2X2 AND2X2_8594 ( .A(u2__abc_44228_n2984_bF_buf14), .B(u2__abc_44228_n17764), .Y(u2__abc_44228_n17765) );
  AND2X2 AND2X2_8595 ( .A(u2__abc_44228_n17766), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_remLo_450__FF_INPUT) );
  AND2X2 AND2X2_8596 ( .A(u2__abc_44228_n15247_bF_buf14), .B(u2_remHiShift_1_), .Y(u2__abc_44228_n17768) );
  AND2X2 AND2X2_8597 ( .A(u2__abc_44228_n2972_bF_buf80), .B(u2_remLo_449_), .Y(u2__abc_44228_n17769) );
  AND2X2 AND2X2_8598 ( .A(u2__abc_44228_n2984_bF_buf13), .B(u2__abc_44228_n17769), .Y(u2__abc_44228_n17770) );
  AND2X2 AND2X2_8599 ( .A(u2__abc_44228_n17771), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_remLo_451__FF_INPUT) );
  AND2X2 AND2X2_86 ( .A(_abc_64468_n858), .B(_abc_64468_n857), .Y(_auto_iopadmap_cc_313_execute_65414_121_) );
  AND2X2 AND2X2_860 ( .A(u2__abc_44228_n3701), .B(u2_remHi_118_), .Y(u2__abc_44228_n3702) );
  AND2X2 AND2X2_8600 ( .A(u2__abc_44228_n2966_bF_buf75), .B(u2_root_0_), .Y(u2__abc_44228_n17773) );
  AND2X2 AND2X2_8601 ( .A(u2__abc_44228_n15247_bF_buf13), .B(u2__abc_44228_n17773), .Y(u2_root_0__FF_INPUT) );
  AND2X2 AND2X2_8602 ( .A(u2__abc_44228_n3062_bF_buf13), .B(sqrto_0_), .Y(u2__abc_44228_n17775) );
  AND2X2 AND2X2_8603 ( .A(u2__abc_44228_n7547_bF_buf12), .B(u2_root_0_), .Y(u2__abc_44228_n17776) );
  AND2X2 AND2X2_8604 ( .A(u2__abc_44228_n17777), .B(u2__abc_44228_n17778), .Y(u2__abc_44228_n17779) );
  AND2X2 AND2X2_8605 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n3077), .Y(u2__abc_44228_n17781) );
  AND2X2 AND2X2_8606 ( .A(u2__abc_44228_n17782), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n17783) );
  AND2X2 AND2X2_8607 ( .A(u2__abc_44228_n17780), .B(u2__abc_44228_n17783), .Y(u2__abc_44228_n17784) );
  AND2X2 AND2X2_8608 ( .A(u2__abc_44228_n17785), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_root_1__FF_INPUT) );
  AND2X2 AND2X2_8609 ( .A(u2__abc_44228_n3062_bF_buf12), .B(sqrto_1_), .Y(u2__abc_44228_n17787) );
  AND2X2 AND2X2_861 ( .A(u2__abc_44228_n3703), .B(sqrto_118_), .Y(u2__abc_44228_n3704_1) );
  AND2X2 AND2X2_8610 ( .A(u2__abc_44228_n17776), .B(sqrto_0_), .Y(u2__abc_44228_n17789) );
  AND2X2 AND2X2_8611 ( .A(u2__abc_44228_n17790), .B(u2__abc_44228_n17788), .Y(u2__abc_44228_n17791) );
  AND2X2 AND2X2_8612 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n3074), .Y(u2__abc_44228_n17793) );
  AND2X2 AND2X2_8613 ( .A(u2__abc_44228_n17794), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n17795) );
  AND2X2 AND2X2_8614 ( .A(u2__abc_44228_n17792), .B(u2__abc_44228_n17795), .Y(u2__abc_44228_n17796) );
  AND2X2 AND2X2_8615 ( .A(u2__abc_44228_n17797), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_root_2__FF_INPUT) );
  AND2X2 AND2X2_8616 ( .A(u2__abc_44228_n3062_bF_buf11), .B(sqrto_2_), .Y(u2__abc_44228_n17799) );
  AND2X2 AND2X2_8617 ( .A(u2__abc_44228_n17789), .B(sqrto_1_), .Y(u2__abc_44228_n17801) );
  AND2X2 AND2X2_8618 ( .A(u2__abc_44228_n17802), .B(u2__abc_44228_n17800), .Y(u2__abc_44228_n17803) );
  AND2X2 AND2X2_8619 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n3104), .Y(u2__abc_44228_n17805) );
  AND2X2 AND2X2_862 ( .A(u2__abc_44228_n3706), .B(u2__abc_44228_n3700), .Y(u2__abc_44228_n3707) );
  AND2X2 AND2X2_8620 ( .A(u2__abc_44228_n17806), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n17807) );
  AND2X2 AND2X2_8621 ( .A(u2__abc_44228_n17804), .B(u2__abc_44228_n17807), .Y(u2__abc_44228_n17808) );
  AND2X2 AND2X2_8622 ( .A(u2__abc_44228_n17809), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_root_3__FF_INPUT) );
  AND2X2 AND2X2_8623 ( .A(u2__abc_44228_n3062_bF_buf10), .B(sqrto_3_), .Y(u2__abc_44228_n17811) );
  AND2X2 AND2X2_8624 ( .A(u2__abc_44228_n17801), .B(sqrto_2_), .Y(u2__abc_44228_n17813) );
  AND2X2 AND2X2_8625 ( .A(u2__abc_44228_n17814), .B(u2__abc_44228_n17812), .Y(u2__abc_44228_n17815) );
  AND2X2 AND2X2_8626 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n3099), .Y(u2__abc_44228_n17817) );
  AND2X2 AND2X2_8627 ( .A(u2__abc_44228_n17818), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n17819) );
  AND2X2 AND2X2_8628 ( .A(u2__abc_44228_n17816), .B(u2__abc_44228_n17819), .Y(u2__abc_44228_n17820) );
  AND2X2 AND2X2_8629 ( .A(u2__abc_44228_n17821), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_root_4__FF_INPUT) );
  AND2X2 AND2X2_863 ( .A(u2__abc_44228_n3708), .B(u2_remHi_121_), .Y(u2__abc_44228_n3709) );
  AND2X2 AND2X2_8630 ( .A(u2__abc_44228_n3062_bF_buf9), .B(sqrto_4_), .Y(u2__abc_44228_n17823) );
  AND2X2 AND2X2_8631 ( .A(u2__abc_44228_n17813), .B(sqrto_3_), .Y(u2__abc_44228_n17825) );
  AND2X2 AND2X2_8632 ( .A(u2__abc_44228_n17826), .B(u2__abc_44228_n17824), .Y(u2__abc_44228_n17827) );
  AND2X2 AND2X2_8633 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n3095), .Y(u2__abc_44228_n17829) );
  AND2X2 AND2X2_8634 ( .A(u2__abc_44228_n17830), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n17831) );
  AND2X2 AND2X2_8635 ( .A(u2__abc_44228_n17828), .B(u2__abc_44228_n17831), .Y(u2__abc_44228_n17832) );
  AND2X2 AND2X2_8636 ( .A(u2__abc_44228_n17833), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_root_5__FF_INPUT) );
  AND2X2 AND2X2_8637 ( .A(u2__abc_44228_n3062_bF_buf8), .B(sqrto_5_), .Y(u2__abc_44228_n17835) );
  AND2X2 AND2X2_8638 ( .A(u2__abc_44228_n17825), .B(sqrto_4_), .Y(u2__abc_44228_n17837) );
  AND2X2 AND2X2_8639 ( .A(u2__abc_44228_n17838), .B(u2__abc_44228_n17836), .Y(u2__abc_44228_n17839) );
  AND2X2 AND2X2_864 ( .A(u2__abc_44228_n3711), .B(sqrto_121_), .Y(u2__abc_44228_n3712) );
  AND2X2 AND2X2_8640 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n3090), .Y(u2__abc_44228_n17841) );
  AND2X2 AND2X2_8641 ( .A(u2__abc_44228_n17842), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n17843) );
  AND2X2 AND2X2_8642 ( .A(u2__abc_44228_n17840), .B(u2__abc_44228_n17843), .Y(u2__abc_44228_n17844) );
  AND2X2 AND2X2_8643 ( .A(u2__abc_44228_n17845), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_root_6__FF_INPUT) );
  AND2X2 AND2X2_8644 ( .A(u2__abc_44228_n3062_bF_buf7), .B(sqrto_6_), .Y(u2__abc_44228_n17847) );
  AND2X2 AND2X2_8645 ( .A(u2__abc_44228_n17837), .B(sqrto_5_), .Y(u2__abc_44228_n17849) );
  AND2X2 AND2X2_8646 ( .A(u2__abc_44228_n17850), .B(u2__abc_44228_n17848), .Y(u2__abc_44228_n17851) );
  AND2X2 AND2X2_8647 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n3161), .Y(u2__abc_44228_n17853) );
  AND2X2 AND2X2_8648 ( .A(u2__abc_44228_n17854), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n17855) );
  AND2X2 AND2X2_8649 ( .A(u2__abc_44228_n17852), .B(u2__abc_44228_n17855), .Y(u2__abc_44228_n17856) );
  AND2X2 AND2X2_865 ( .A(u2__abc_44228_n3710), .B(u2__abc_44228_n3713), .Y(u2__abc_44228_n3714_1) );
  AND2X2 AND2X2_8650 ( .A(u2__abc_44228_n17857), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_root_7__FF_INPUT) );
  AND2X2 AND2X2_8651 ( .A(u2__abc_44228_n3062_bF_buf6), .B(sqrto_7_), .Y(u2__abc_44228_n17859) );
  AND2X2 AND2X2_8652 ( .A(u2__abc_44228_n17849), .B(sqrto_6_), .Y(u2__abc_44228_n17861) );
  AND2X2 AND2X2_8653 ( .A(u2__abc_44228_n17862), .B(u2__abc_44228_n17860), .Y(u2__abc_44228_n17863) );
  AND2X2 AND2X2_8654 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n3167), .Y(u2__abc_44228_n17865) );
  AND2X2 AND2X2_8655 ( .A(u2__abc_44228_n17866), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n17867) );
  AND2X2 AND2X2_8656 ( .A(u2__abc_44228_n17864), .B(u2__abc_44228_n17867), .Y(u2__abc_44228_n17868) );
  AND2X2 AND2X2_8657 ( .A(u2__abc_44228_n17869), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_root_8__FF_INPUT) );
  AND2X2 AND2X2_8658 ( .A(u2__abc_44228_n3062_bF_buf5), .B(sqrto_8_), .Y(u2__abc_44228_n17871) );
  AND2X2 AND2X2_8659 ( .A(u2__abc_44228_n17861), .B(sqrto_7_), .Y(u2__abc_44228_n17873) );
  AND2X2 AND2X2_866 ( .A(u2__abc_44228_n3715), .B(u2_remHi_120_), .Y(u2__abc_44228_n3716) );
  AND2X2 AND2X2_8660 ( .A(u2__abc_44228_n17874), .B(u2__abc_44228_n17872), .Y(u2__abc_44228_n17875) );
  AND2X2 AND2X2_8661 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n3157), .Y(u2__abc_44228_n17877) );
  AND2X2 AND2X2_8662 ( .A(u2__abc_44228_n17878), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n17879) );
  AND2X2 AND2X2_8663 ( .A(u2__abc_44228_n17876), .B(u2__abc_44228_n17879), .Y(u2__abc_44228_n17880) );
  AND2X2 AND2X2_8664 ( .A(u2__abc_44228_n17881), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_root_9__FF_INPUT) );
  AND2X2 AND2X2_8665 ( .A(u2__abc_44228_n3062_bF_buf4), .B(sqrto_9_), .Y(u2__abc_44228_n17883) );
  AND2X2 AND2X2_8666 ( .A(u2__abc_44228_n17873), .B(sqrto_8_), .Y(u2__abc_44228_n17885) );
  AND2X2 AND2X2_8667 ( .A(u2__abc_44228_n17886), .B(u2__abc_44228_n17884), .Y(u2__abc_44228_n17887) );
  AND2X2 AND2X2_8668 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n3152), .Y(u2__abc_44228_n17889) );
  AND2X2 AND2X2_8669 ( .A(u2__abc_44228_n17890), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n17891) );
  AND2X2 AND2X2_867 ( .A(u2__abc_44228_n3717), .B(sqrto_120_), .Y(u2__abc_44228_n3718) );
  AND2X2 AND2X2_8670 ( .A(u2__abc_44228_n17888), .B(u2__abc_44228_n17891), .Y(u2__abc_44228_n17892) );
  AND2X2 AND2X2_8671 ( .A(u2__abc_44228_n17893), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_root_10__FF_INPUT) );
  AND2X2 AND2X2_8672 ( .A(u2__abc_44228_n3062_bF_buf3), .B(sqrto_10_), .Y(u2__abc_44228_n17895) );
  AND2X2 AND2X2_8673 ( .A(u2__abc_44228_n17885), .B(sqrto_9_), .Y(u2__abc_44228_n17897) );
  AND2X2 AND2X2_8674 ( .A(u2__abc_44228_n17898), .B(u2__abc_44228_n17896), .Y(u2__abc_44228_n17899) );
  AND2X2 AND2X2_8675 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n3142), .Y(u2__abc_44228_n17901) );
  AND2X2 AND2X2_8676 ( .A(u2__abc_44228_n17902), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n17903) );
  AND2X2 AND2X2_8677 ( .A(u2__abc_44228_n17900), .B(u2__abc_44228_n17903), .Y(u2__abc_44228_n17904) );
  AND2X2 AND2X2_8678 ( .A(u2__abc_44228_n17905), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_root_11__FF_INPUT) );
  AND2X2 AND2X2_8679 ( .A(u2__abc_44228_n3062_bF_buf2), .B(sqrto_11_), .Y(u2__abc_44228_n17907) );
  AND2X2 AND2X2_868 ( .A(u2__abc_44228_n3720), .B(u2__abc_44228_n3714_1), .Y(u2__abc_44228_n3721) );
  AND2X2 AND2X2_8680 ( .A(u2__abc_44228_n17897), .B(sqrto_10_), .Y(u2__abc_44228_n17909) );
  AND2X2 AND2X2_8681 ( .A(u2__abc_44228_n17910), .B(u2__abc_44228_n17908), .Y(u2__abc_44228_n17911) );
  AND2X2 AND2X2_8682 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n3135), .Y(u2__abc_44228_n17913) );
  AND2X2 AND2X2_8683 ( .A(u2__abc_44228_n17914), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n17915) );
  AND2X2 AND2X2_8684 ( .A(u2__abc_44228_n17912), .B(u2__abc_44228_n17915), .Y(u2__abc_44228_n17916) );
  AND2X2 AND2X2_8685 ( .A(u2__abc_44228_n17917), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_root_12__FF_INPUT) );
  AND2X2 AND2X2_8686 ( .A(u2__abc_44228_n3062_bF_buf1), .B(sqrto_12_), .Y(u2__abc_44228_n17919) );
  AND2X2 AND2X2_8687 ( .A(u2__abc_44228_n17909), .B(sqrto_11_), .Y(u2__abc_44228_n17921) );
  AND2X2 AND2X2_8688 ( .A(u2__abc_44228_n17922), .B(u2__abc_44228_n17920), .Y(u2__abc_44228_n17923) );
  AND2X2 AND2X2_8689 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n3128), .Y(u2__abc_44228_n17925) );
  AND2X2 AND2X2_869 ( .A(u2__abc_44228_n3707), .B(u2__abc_44228_n3721), .Y(u2__abc_44228_n3722) );
  AND2X2 AND2X2_8690 ( .A(u2__abc_44228_n17926), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n17927) );
  AND2X2 AND2X2_8691 ( .A(u2__abc_44228_n17924), .B(u2__abc_44228_n17927), .Y(u2__abc_44228_n17928) );
  AND2X2 AND2X2_8692 ( .A(u2__abc_44228_n17929), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_root_13__FF_INPUT) );
  AND2X2 AND2X2_8693 ( .A(u2__abc_44228_n3062_bF_buf0), .B(sqrto_13_), .Y(u2__abc_44228_n17931) );
  AND2X2 AND2X2_8694 ( .A(u2__abc_44228_n17921), .B(sqrto_12_), .Y(u2__abc_44228_n17933) );
  AND2X2 AND2X2_8695 ( .A(u2__abc_44228_n17934), .B(u2__abc_44228_n17932), .Y(u2__abc_44228_n17935) );
  AND2X2 AND2X2_8696 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n3121), .Y(u2__abc_44228_n17937) );
  AND2X2 AND2X2_8697 ( .A(u2__abc_44228_n17938), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n17939) );
  AND2X2 AND2X2_8698 ( .A(u2__abc_44228_n17936), .B(u2__abc_44228_n17939), .Y(u2__abc_44228_n17940) );
  AND2X2 AND2X2_8699 ( .A(u2__abc_44228_n17941), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_root_14__FF_INPUT) );
  AND2X2 AND2X2_87 ( .A(_abc_64468_n861), .B(_abc_64468_n860), .Y(_auto_iopadmap_cc_313_execute_65414_122_) );
  AND2X2 AND2X2_870 ( .A(u2__abc_44228_n3693), .B(u2__abc_44228_n3722), .Y(u2__abc_44228_n3723_1) );
  AND2X2 AND2X2_8700 ( .A(u2__abc_44228_n3062_bF_buf92), .B(sqrto_14_), .Y(u2__abc_44228_n17943) );
  AND2X2 AND2X2_8701 ( .A(u2__abc_44228_n17933), .B(sqrto_13_), .Y(u2__abc_44228_n17945) );
  AND2X2 AND2X2_8702 ( .A(u2__abc_44228_n17946), .B(u2__abc_44228_n17944), .Y(u2__abc_44228_n17947) );
  AND2X2 AND2X2_8703 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n3301), .Y(u2__abc_44228_n17949) );
  AND2X2 AND2X2_8704 ( .A(u2__abc_44228_n17950), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n17951) );
  AND2X2 AND2X2_8705 ( .A(u2__abc_44228_n17948), .B(u2__abc_44228_n17951), .Y(u2__abc_44228_n17952) );
  AND2X2 AND2X2_8706 ( .A(u2__abc_44228_n17953), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_root_15__FF_INPUT) );
  AND2X2 AND2X2_8707 ( .A(u2__abc_44228_n3062_bF_buf91), .B(sqrto_15_), .Y(u2__abc_44228_n17955) );
  AND2X2 AND2X2_8708 ( .A(u2__abc_44228_n17945), .B(sqrto_14_), .Y(u2__abc_44228_n17957) );
  AND2X2 AND2X2_8709 ( .A(u2__abc_44228_n17958), .B(u2__abc_44228_n17956), .Y(u2__abc_44228_n17959) );
  AND2X2 AND2X2_871 ( .A(u2__abc_44228_n3724), .B(u2_remHi_117_), .Y(u2__abc_44228_n3725) );
  AND2X2 AND2X2_8710 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n3294), .Y(u2__abc_44228_n17961) );
  AND2X2 AND2X2_8711 ( .A(u2__abc_44228_n17962), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n17963) );
  AND2X2 AND2X2_8712 ( .A(u2__abc_44228_n17960), .B(u2__abc_44228_n17963), .Y(u2__abc_44228_n17964) );
  AND2X2 AND2X2_8713 ( .A(u2__abc_44228_n17965), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_root_16__FF_INPUT) );
  AND2X2 AND2X2_8714 ( .A(u2__abc_44228_n3062_bF_buf90), .B(sqrto_16_), .Y(u2__abc_44228_n17967) );
  AND2X2 AND2X2_8715 ( .A(u2__abc_44228_n17957), .B(sqrto_15_), .Y(u2__abc_44228_n17969) );
  AND2X2 AND2X2_8716 ( .A(u2__abc_44228_n17970), .B(u2__abc_44228_n17968), .Y(u2__abc_44228_n17971) );
  AND2X2 AND2X2_8717 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n3290), .Y(u2__abc_44228_n17973) );
  AND2X2 AND2X2_8718 ( .A(u2__abc_44228_n17974), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n17975) );
  AND2X2 AND2X2_8719 ( .A(u2__abc_44228_n17972), .B(u2__abc_44228_n17975), .Y(u2__abc_44228_n17976) );
  AND2X2 AND2X2_872 ( .A(u2__abc_44228_n3727), .B(sqrto_117_), .Y(u2__abc_44228_n3728) );
  AND2X2 AND2X2_8720 ( .A(u2__abc_44228_n17977), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_root_17__FF_INPUT) );
  AND2X2 AND2X2_8721 ( .A(u2__abc_44228_n3062_bF_buf89), .B(sqrto_17_), .Y(u2__abc_44228_n17979) );
  AND2X2 AND2X2_8722 ( .A(u2__abc_44228_n17969), .B(sqrto_16_), .Y(u2__abc_44228_n17981) );
  AND2X2 AND2X2_8723 ( .A(u2__abc_44228_n17982), .B(u2__abc_44228_n17980), .Y(u2__abc_44228_n17983) );
  AND2X2 AND2X2_8724 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n3285), .Y(u2__abc_44228_n17985) );
  AND2X2 AND2X2_8725 ( .A(u2__abc_44228_n17986), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n17987) );
  AND2X2 AND2X2_8726 ( .A(u2__abc_44228_n17984), .B(u2__abc_44228_n17987), .Y(u2__abc_44228_n17988) );
  AND2X2 AND2X2_8727 ( .A(u2__abc_44228_n17989), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_root_18__FF_INPUT) );
  AND2X2 AND2X2_8728 ( .A(u2__abc_44228_n3062_bF_buf88), .B(sqrto_18_), .Y(u2__abc_44228_n17991) );
  AND2X2 AND2X2_8729 ( .A(u2__abc_44228_n17981), .B(sqrto_17_), .Y(u2__abc_44228_n17993) );
  AND2X2 AND2X2_873 ( .A(u2__abc_44228_n3726), .B(u2__abc_44228_n3729), .Y(u2__abc_44228_n3730) );
  AND2X2 AND2X2_8730 ( .A(u2__abc_44228_n17994), .B(u2__abc_44228_n17992), .Y(u2__abc_44228_n17995) );
  AND2X2 AND2X2_8731 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n3268), .Y(u2__abc_44228_n17997) );
  AND2X2 AND2X2_8732 ( .A(u2__abc_44228_n17998), .B(u2__abc_44228_n2972_bF_buf61), .Y(u2__abc_44228_n17999) );
  AND2X2 AND2X2_8733 ( .A(u2__abc_44228_n17996), .B(u2__abc_44228_n17999), .Y(u2__abc_44228_n18000) );
  AND2X2 AND2X2_8734 ( .A(u2__abc_44228_n18001), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_root_19__FF_INPUT) );
  AND2X2 AND2X2_8735 ( .A(u2__abc_44228_n3062_bF_buf87), .B(sqrto_19_), .Y(u2__abc_44228_n18003) );
  AND2X2 AND2X2_8736 ( .A(u2__abc_44228_n17993), .B(sqrto_18_), .Y(u2__abc_44228_n18005) );
  AND2X2 AND2X2_8737 ( .A(u2__abc_44228_n18006), .B(u2__abc_44228_n18004), .Y(u2__abc_44228_n18007) );
  AND2X2 AND2X2_8738 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n3274), .Y(u2__abc_44228_n18009) );
  AND2X2 AND2X2_8739 ( .A(u2__abc_44228_n18010), .B(u2__abc_44228_n2972_bF_buf60), .Y(u2__abc_44228_n18011) );
  AND2X2 AND2X2_874 ( .A(u2__abc_44228_n3731), .B(u2_remHi_116_), .Y(u2__abc_44228_n3732_1) );
  AND2X2 AND2X2_8740 ( .A(u2__abc_44228_n18008), .B(u2__abc_44228_n18011), .Y(u2__abc_44228_n18012) );
  AND2X2 AND2X2_8741 ( .A(u2__abc_44228_n18013), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_root_20__FF_INPUT) );
  AND2X2 AND2X2_8742 ( .A(u2__abc_44228_n3062_bF_buf86), .B(sqrto_20_), .Y(u2__abc_44228_n18015) );
  AND2X2 AND2X2_8743 ( .A(u2__abc_44228_n18005), .B(sqrto_19_), .Y(u2__abc_44228_n18017) );
  AND2X2 AND2X2_8744 ( .A(u2__abc_44228_n18018), .B(u2__abc_44228_n18016), .Y(u2__abc_44228_n18019) );
  AND2X2 AND2X2_8745 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n3261), .Y(u2__abc_44228_n18021) );
  AND2X2 AND2X2_8746 ( .A(u2__abc_44228_n18022), .B(u2__abc_44228_n2972_bF_buf59), .Y(u2__abc_44228_n18023) );
  AND2X2 AND2X2_8747 ( .A(u2__abc_44228_n18020), .B(u2__abc_44228_n18023), .Y(u2__abc_44228_n18024) );
  AND2X2 AND2X2_8748 ( .A(u2__abc_44228_n18025), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_root_21__FF_INPUT) );
  AND2X2 AND2X2_8749 ( .A(u2__abc_44228_n3062_bF_buf85), .B(sqrto_21_), .Y(u2__abc_44228_n18027) );
  AND2X2 AND2X2_875 ( .A(u2__abc_44228_n3733), .B(sqrto_116_), .Y(u2__abc_44228_n3734) );
  AND2X2 AND2X2_8750 ( .A(u2__abc_44228_n18017), .B(sqrto_20_), .Y(u2__abc_44228_n18029) );
  AND2X2 AND2X2_8751 ( .A(u2__abc_44228_n18030), .B(u2__abc_44228_n18028), .Y(u2__abc_44228_n18031) );
  AND2X2 AND2X2_8752 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n3254), .Y(u2__abc_44228_n18033) );
  AND2X2 AND2X2_8753 ( .A(u2__abc_44228_n18034), .B(u2__abc_44228_n2972_bF_buf58), .Y(u2__abc_44228_n18035) );
  AND2X2 AND2X2_8754 ( .A(u2__abc_44228_n18032), .B(u2__abc_44228_n18035), .Y(u2__abc_44228_n18036) );
  AND2X2 AND2X2_8755 ( .A(u2__abc_44228_n18037), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_root_22__FF_INPUT) );
  AND2X2 AND2X2_8756 ( .A(u2__abc_44228_n3062_bF_buf84), .B(sqrto_22_), .Y(u2__abc_44228_n18039) );
  AND2X2 AND2X2_8757 ( .A(u2__abc_44228_n18029), .B(sqrto_21_), .Y(u2__abc_44228_n18041) );
  AND2X2 AND2X2_8758 ( .A(u2__abc_44228_n18042), .B(u2__abc_44228_n18040), .Y(u2__abc_44228_n18043) );
  AND2X2 AND2X2_8759 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n3231), .Y(u2__abc_44228_n18045) );
  AND2X2 AND2X2_876 ( .A(u2__abc_44228_n3736), .B(u2__abc_44228_n3730), .Y(u2__abc_44228_n3737) );
  AND2X2 AND2X2_8760 ( .A(u2__abc_44228_n18046), .B(u2__abc_44228_n2972_bF_buf57), .Y(u2__abc_44228_n18047) );
  AND2X2 AND2X2_8761 ( .A(u2__abc_44228_n18044), .B(u2__abc_44228_n18047), .Y(u2__abc_44228_n18048) );
  AND2X2 AND2X2_8762 ( .A(u2__abc_44228_n18049), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_root_23__FF_INPUT) );
  AND2X2 AND2X2_8763 ( .A(u2__abc_44228_n3062_bF_buf83), .B(sqrto_23_), .Y(u2__abc_44228_n18051) );
  AND2X2 AND2X2_8764 ( .A(u2__abc_44228_n18041), .B(sqrto_22_), .Y(u2__abc_44228_n18053) );
  AND2X2 AND2X2_8765 ( .A(u2__abc_44228_n18054), .B(u2__abc_44228_n18052), .Y(u2__abc_44228_n18055) );
  AND2X2 AND2X2_8766 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n3224), .Y(u2__abc_44228_n18057) );
  AND2X2 AND2X2_8767 ( .A(u2__abc_44228_n18058), .B(u2__abc_44228_n2972_bF_buf56), .Y(u2__abc_44228_n18059) );
  AND2X2 AND2X2_8768 ( .A(u2__abc_44228_n18056), .B(u2__abc_44228_n18059), .Y(u2__abc_44228_n18060) );
  AND2X2 AND2X2_8769 ( .A(u2__abc_44228_n18061), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_root_24__FF_INPUT) );
  AND2X2 AND2X2_877 ( .A(u2__abc_44228_n3738), .B(u2_remHi_115_), .Y(u2__abc_44228_n3739) );
  AND2X2 AND2X2_8770 ( .A(u2__abc_44228_n3062_bF_buf82), .B(sqrto_24_), .Y(u2__abc_44228_n18063) );
  AND2X2 AND2X2_8771 ( .A(u2__abc_44228_n18053), .B(sqrto_23_), .Y(u2__abc_44228_n18065) );
  AND2X2 AND2X2_8772 ( .A(u2__abc_44228_n18066), .B(u2__abc_44228_n18064), .Y(u2__abc_44228_n18067) );
  AND2X2 AND2X2_8773 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n3245), .Y(u2__abc_44228_n18069) );
  AND2X2 AND2X2_8774 ( .A(u2__abc_44228_n18070), .B(u2__abc_44228_n2972_bF_buf55), .Y(u2__abc_44228_n18071) );
  AND2X2 AND2X2_8775 ( .A(u2__abc_44228_n18068), .B(u2__abc_44228_n18071), .Y(u2__abc_44228_n18072) );
  AND2X2 AND2X2_8776 ( .A(u2__abc_44228_n18073), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_root_25__FF_INPUT) );
  AND2X2 AND2X2_8777 ( .A(u2__abc_44228_n3062_bF_buf81), .B(sqrto_25_), .Y(u2__abc_44228_n18075) );
  AND2X2 AND2X2_8778 ( .A(u2__abc_44228_n18065), .B(sqrto_24_), .Y(u2__abc_44228_n18077) );
  AND2X2 AND2X2_8779 ( .A(u2__abc_44228_n18078), .B(u2__abc_44228_n18076), .Y(u2__abc_44228_n18079) );
  AND2X2 AND2X2_878 ( .A(u2__abc_44228_n3741), .B(sqrto_115_), .Y(u2__abc_44228_n3742) );
  AND2X2 AND2X2_8780 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n3238), .Y(u2__abc_44228_n18081) );
  AND2X2 AND2X2_8781 ( .A(u2__abc_44228_n18082), .B(u2__abc_44228_n2972_bF_buf54), .Y(u2__abc_44228_n18083) );
  AND2X2 AND2X2_8782 ( .A(u2__abc_44228_n18080), .B(u2__abc_44228_n18083), .Y(u2__abc_44228_n18084) );
  AND2X2 AND2X2_8783 ( .A(u2__abc_44228_n18085), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_root_26__FF_INPUT) );
  AND2X2 AND2X2_8784 ( .A(u2__abc_44228_n3062_bF_buf80), .B(sqrto_26_), .Y(u2__abc_44228_n18087) );
  AND2X2 AND2X2_8785 ( .A(u2__abc_44228_n18077), .B(sqrto_25_), .Y(u2__abc_44228_n18089) );
  AND2X2 AND2X2_8786 ( .A(u2__abc_44228_n18090), .B(u2__abc_44228_n18088), .Y(u2__abc_44228_n18091) );
  AND2X2 AND2X2_8787 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n3209), .Y(u2__abc_44228_n18093) );
  AND2X2 AND2X2_8788 ( .A(u2__abc_44228_n18094), .B(u2__abc_44228_n2972_bF_buf53), .Y(u2__abc_44228_n18095) );
  AND2X2 AND2X2_8789 ( .A(u2__abc_44228_n18092), .B(u2__abc_44228_n18095), .Y(u2__abc_44228_n18096) );
  AND2X2 AND2X2_879 ( .A(u2__abc_44228_n3740_1), .B(u2__abc_44228_n3743), .Y(u2__abc_44228_n3744) );
  AND2X2 AND2X2_8790 ( .A(u2__abc_44228_n18097), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_root_27__FF_INPUT) );
  AND2X2 AND2X2_8791 ( .A(u2__abc_44228_n3062_bF_buf79), .B(sqrto_27_), .Y(u2__abc_44228_n18099) );
  AND2X2 AND2X2_8792 ( .A(u2__abc_44228_n18089), .B(sqrto_26_), .Y(u2__abc_44228_n18101) );
  AND2X2 AND2X2_8793 ( .A(u2__abc_44228_n18102), .B(u2__abc_44228_n18100), .Y(u2__abc_44228_n18103) );
  AND2X2 AND2X2_8794 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n3215), .Y(u2__abc_44228_n18105) );
  AND2X2 AND2X2_8795 ( .A(u2__abc_44228_n18106), .B(u2__abc_44228_n2972_bF_buf52), .Y(u2__abc_44228_n18107) );
  AND2X2 AND2X2_8796 ( .A(u2__abc_44228_n18104), .B(u2__abc_44228_n18107), .Y(u2__abc_44228_n18108) );
  AND2X2 AND2X2_8797 ( .A(u2__abc_44228_n18109), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_root_28__FF_INPUT) );
  AND2X2 AND2X2_8798 ( .A(u2__abc_44228_n3062_bF_buf78), .B(sqrto_28_), .Y(u2__abc_44228_n18111) );
  AND2X2 AND2X2_8799 ( .A(u2__abc_44228_n18101), .B(sqrto_27_), .Y(u2__abc_44228_n18113) );
  AND2X2 AND2X2_88 ( .A(_abc_64468_n864), .B(_abc_64468_n863), .Y(_auto_iopadmap_cc_313_execute_65414_123_) );
  AND2X2 AND2X2_880 ( .A(u2__abc_44228_n3745), .B(u2_remHi_114_), .Y(u2__abc_44228_n3746) );
  AND2X2 AND2X2_8800 ( .A(u2__abc_44228_n18114), .B(u2__abc_44228_n18112), .Y(u2__abc_44228_n18115) );
  AND2X2 AND2X2_8801 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n3202), .Y(u2__abc_44228_n18117) );
  AND2X2 AND2X2_8802 ( .A(u2__abc_44228_n18118), .B(u2__abc_44228_n2972_bF_buf51), .Y(u2__abc_44228_n18119) );
  AND2X2 AND2X2_8803 ( .A(u2__abc_44228_n18116), .B(u2__abc_44228_n18119), .Y(u2__abc_44228_n18120) );
  AND2X2 AND2X2_8804 ( .A(u2__abc_44228_n18121), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_root_29__FF_INPUT) );
  AND2X2 AND2X2_8805 ( .A(u2__abc_44228_n3062_bF_buf77), .B(sqrto_29_), .Y(u2__abc_44228_n18123) );
  AND2X2 AND2X2_8806 ( .A(u2__abc_44228_n18113), .B(sqrto_28_), .Y(u2__abc_44228_n18125) );
  AND2X2 AND2X2_8807 ( .A(u2__abc_44228_n18126), .B(u2__abc_44228_n18124), .Y(u2__abc_44228_n18127) );
  AND2X2 AND2X2_8808 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n3195), .Y(u2__abc_44228_n18129) );
  AND2X2 AND2X2_8809 ( .A(u2__abc_44228_n18130), .B(u2__abc_44228_n2972_bF_buf50), .Y(u2__abc_44228_n18131) );
  AND2X2 AND2X2_881 ( .A(u2__abc_44228_n3747), .B(sqrto_114_), .Y(u2__abc_44228_n3748) );
  AND2X2 AND2X2_8810 ( .A(u2__abc_44228_n18128), .B(u2__abc_44228_n18131), .Y(u2__abc_44228_n18132) );
  AND2X2 AND2X2_8811 ( .A(u2__abc_44228_n18133), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_root_30__FF_INPUT) );
  AND2X2 AND2X2_8812 ( .A(u2__abc_44228_n3062_bF_buf76), .B(sqrto_30_), .Y(u2__abc_44228_n18135) );
  AND2X2 AND2X2_8813 ( .A(u2__abc_44228_n18125), .B(sqrto_29_), .Y(u2__abc_44228_n18137) );
  AND2X2 AND2X2_8814 ( .A(u2__abc_44228_n18138), .B(u2__abc_44228_n18136), .Y(u2__abc_44228_n18139) );
  AND2X2 AND2X2_8815 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n3567), .Y(u2__abc_44228_n18141) );
  AND2X2 AND2X2_8816 ( .A(u2__abc_44228_n18142), .B(u2__abc_44228_n2972_bF_buf49), .Y(u2__abc_44228_n18143) );
  AND2X2 AND2X2_8817 ( .A(u2__abc_44228_n18140), .B(u2__abc_44228_n18143), .Y(u2__abc_44228_n18144) );
  AND2X2 AND2X2_8818 ( .A(u2__abc_44228_n18145), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_root_31__FF_INPUT) );
  AND2X2 AND2X2_8819 ( .A(u2__abc_44228_n3062_bF_buf75), .B(sqrto_31_), .Y(u2__abc_44228_n18147) );
  AND2X2 AND2X2_882 ( .A(u2__abc_44228_n3750_1), .B(u2__abc_44228_n3744), .Y(u2__abc_44228_n3751) );
  AND2X2 AND2X2_8820 ( .A(u2__abc_44228_n18137), .B(sqrto_30_), .Y(u2__abc_44228_n18149) );
  AND2X2 AND2X2_8821 ( .A(u2__abc_44228_n18150), .B(u2__abc_44228_n18148), .Y(u2__abc_44228_n18151) );
  AND2X2 AND2X2_8822 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n3573), .Y(u2__abc_44228_n18153) );
  AND2X2 AND2X2_8823 ( .A(u2__abc_44228_n18154), .B(u2__abc_44228_n2972_bF_buf48), .Y(u2__abc_44228_n18155) );
  AND2X2 AND2X2_8824 ( .A(u2__abc_44228_n18152), .B(u2__abc_44228_n18155), .Y(u2__abc_44228_n18156) );
  AND2X2 AND2X2_8825 ( .A(u2__abc_44228_n18157), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_root_32__FF_INPUT) );
  AND2X2 AND2X2_8826 ( .A(u2__abc_44228_n3062_bF_buf74), .B(sqrto_32_), .Y(u2__abc_44228_n18159) );
  AND2X2 AND2X2_8827 ( .A(u2__abc_44228_n18149), .B(sqrto_31_), .Y(u2__abc_44228_n18161) );
  AND2X2 AND2X2_8828 ( .A(u2__abc_44228_n18162), .B(u2__abc_44228_n18160), .Y(u2__abc_44228_n18163) );
  AND2X2 AND2X2_8829 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n3563), .Y(u2__abc_44228_n18165) );
  AND2X2 AND2X2_883 ( .A(u2__abc_44228_n3737), .B(u2__abc_44228_n3751), .Y(u2__abc_44228_n3752) );
  AND2X2 AND2X2_8830 ( .A(u2__abc_44228_n18166), .B(u2__abc_44228_n2972_bF_buf47), .Y(u2__abc_44228_n18167) );
  AND2X2 AND2X2_8831 ( .A(u2__abc_44228_n18164), .B(u2__abc_44228_n18167), .Y(u2__abc_44228_n18168) );
  AND2X2 AND2X2_8832 ( .A(u2__abc_44228_n18169), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_root_33__FF_INPUT) );
  AND2X2 AND2X2_8833 ( .A(u2__abc_44228_n3062_bF_buf73), .B(sqrto_33_), .Y(u2__abc_44228_n18171) );
  AND2X2 AND2X2_8834 ( .A(u2__abc_44228_n18161), .B(sqrto_32_), .Y(u2__abc_44228_n18173) );
  AND2X2 AND2X2_8835 ( .A(u2__abc_44228_n18174), .B(u2__abc_44228_n18172), .Y(u2__abc_44228_n18175) );
  AND2X2 AND2X2_8836 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n3558), .Y(u2__abc_44228_n18177) );
  AND2X2 AND2X2_8837 ( .A(u2__abc_44228_n18178), .B(u2__abc_44228_n2972_bF_buf46), .Y(u2__abc_44228_n18179) );
  AND2X2 AND2X2_8838 ( .A(u2__abc_44228_n18176), .B(u2__abc_44228_n18179), .Y(u2__abc_44228_n18180) );
  AND2X2 AND2X2_8839 ( .A(u2__abc_44228_n18181), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_root_34__FF_INPUT) );
  AND2X2 AND2X2_884 ( .A(u2__abc_44228_n3753), .B(u2_remHi_113_), .Y(u2__abc_44228_n3754) );
  AND2X2 AND2X2_8840 ( .A(u2__abc_44228_n3062_bF_buf72), .B(sqrto_34_), .Y(u2__abc_44228_n18183) );
  AND2X2 AND2X2_8841 ( .A(u2__abc_44228_n18173), .B(sqrto_33_), .Y(u2__abc_44228_n18185) );
  AND2X2 AND2X2_8842 ( .A(u2__abc_44228_n18186), .B(u2__abc_44228_n18184), .Y(u2__abc_44228_n18187) );
  AND2X2 AND2X2_8843 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n3541_1), .Y(u2__abc_44228_n18189) );
  AND2X2 AND2X2_8844 ( .A(u2__abc_44228_n18190), .B(u2__abc_44228_n2972_bF_buf45), .Y(u2__abc_44228_n18191) );
  AND2X2 AND2X2_8845 ( .A(u2__abc_44228_n18188), .B(u2__abc_44228_n18191), .Y(u2__abc_44228_n18192) );
  AND2X2 AND2X2_8846 ( .A(u2__abc_44228_n18193), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_root_35__FF_INPUT) );
  AND2X2 AND2X2_8847 ( .A(u2__abc_44228_n3062_bF_buf71), .B(sqrto_35_), .Y(u2__abc_44228_n18195) );
  AND2X2 AND2X2_8848 ( .A(u2__abc_44228_n18185), .B(sqrto_34_), .Y(u2__abc_44228_n18197) );
  AND2X2 AND2X2_8849 ( .A(u2__abc_44228_n18198), .B(u2__abc_44228_n18196), .Y(u2__abc_44228_n18199) );
  AND2X2 AND2X2_885 ( .A(u2__abc_44228_n3756), .B(sqrto_113_), .Y(u2__abc_44228_n3757) );
  AND2X2 AND2X2_8850 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n3547), .Y(u2__abc_44228_n18201) );
  AND2X2 AND2X2_8851 ( .A(u2__abc_44228_n18202), .B(u2__abc_44228_n2972_bF_buf44), .Y(u2__abc_44228_n18203) );
  AND2X2 AND2X2_8852 ( .A(u2__abc_44228_n18200), .B(u2__abc_44228_n18203), .Y(u2__abc_44228_n18204) );
  AND2X2 AND2X2_8853 ( .A(u2__abc_44228_n18205), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_root_36__FF_INPUT) );
  AND2X2 AND2X2_8854 ( .A(u2__abc_44228_n3062_bF_buf70), .B(sqrto_36_), .Y(u2__abc_44228_n18207) );
  AND2X2 AND2X2_8855 ( .A(u2__abc_44228_n18197), .B(sqrto_35_), .Y(u2__abc_44228_n18209) );
  AND2X2 AND2X2_8856 ( .A(u2__abc_44228_n18210), .B(u2__abc_44228_n18208), .Y(u2__abc_44228_n18211) );
  AND2X2 AND2X2_8857 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n3534), .Y(u2__abc_44228_n18213) );
  AND2X2 AND2X2_8858 ( .A(u2__abc_44228_n18214), .B(u2__abc_44228_n2972_bF_buf43), .Y(u2__abc_44228_n18215) );
  AND2X2 AND2X2_8859 ( .A(u2__abc_44228_n18212), .B(u2__abc_44228_n18215), .Y(u2__abc_44228_n18216) );
  AND2X2 AND2X2_886 ( .A(u2__abc_44228_n3755), .B(u2__abc_44228_n3758), .Y(u2__abc_44228_n3759_1) );
  AND2X2 AND2X2_8860 ( .A(u2__abc_44228_n18217), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_root_37__FF_INPUT) );
  AND2X2 AND2X2_8861 ( .A(u2__abc_44228_n3062_bF_buf69), .B(sqrto_37_), .Y(u2__abc_44228_n18219) );
  AND2X2 AND2X2_8862 ( .A(u2__abc_44228_n18209), .B(sqrto_36_), .Y(u2__abc_44228_n18221) );
  AND2X2 AND2X2_8863 ( .A(u2__abc_44228_n18222), .B(u2__abc_44228_n18220), .Y(u2__abc_44228_n18223) );
  AND2X2 AND2X2_8864 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n3527), .Y(u2__abc_44228_n18225) );
  AND2X2 AND2X2_8865 ( .A(u2__abc_44228_n18226), .B(u2__abc_44228_n2972_bF_buf42), .Y(u2__abc_44228_n18227) );
  AND2X2 AND2X2_8866 ( .A(u2__abc_44228_n18224), .B(u2__abc_44228_n18227), .Y(u2__abc_44228_n18228) );
  AND2X2 AND2X2_8867 ( .A(u2__abc_44228_n18229), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_root_38__FF_INPUT) );
  AND2X2 AND2X2_8868 ( .A(u2__abc_44228_n3062_bF_buf68), .B(sqrto_38_), .Y(u2__abc_44228_n18231) );
  AND2X2 AND2X2_8869 ( .A(u2__abc_44228_n18221), .B(sqrto_37_), .Y(u2__abc_44228_n18233) );
  AND2X2 AND2X2_887 ( .A(u2__abc_44228_n3760), .B(u2_remHi_112_), .Y(u2__abc_44228_n3761) );
  AND2X2 AND2X2_8870 ( .A(u2__abc_44228_n18234), .B(u2__abc_44228_n18232), .Y(u2__abc_44228_n18235) );
  AND2X2 AND2X2_8871 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n3504), .Y(u2__abc_44228_n18237) );
  AND2X2 AND2X2_8872 ( .A(u2__abc_44228_n18238), .B(u2__abc_44228_n2972_bF_buf41), .Y(u2__abc_44228_n18239) );
  AND2X2 AND2X2_8873 ( .A(u2__abc_44228_n18236), .B(u2__abc_44228_n18239), .Y(u2__abc_44228_n18240) );
  AND2X2 AND2X2_8874 ( .A(u2__abc_44228_n18241), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_root_39__FF_INPUT) );
  AND2X2 AND2X2_8875 ( .A(u2__abc_44228_n3062_bF_buf67), .B(sqrto_39_), .Y(u2__abc_44228_n18243) );
  AND2X2 AND2X2_8876 ( .A(u2__abc_44228_n18233), .B(sqrto_38_), .Y(u2__abc_44228_n18245) );
  AND2X2 AND2X2_8877 ( .A(u2__abc_44228_n18246), .B(u2__abc_44228_n18244), .Y(u2__abc_44228_n18247) );
  AND2X2 AND2X2_8878 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n3497), .Y(u2__abc_44228_n18249) );
  AND2X2 AND2X2_8879 ( .A(u2__abc_44228_n18250), .B(u2__abc_44228_n2972_bF_buf40), .Y(u2__abc_44228_n18251) );
  AND2X2 AND2X2_888 ( .A(u2__abc_44228_n3762), .B(sqrto_112_), .Y(u2__abc_44228_n3763) );
  AND2X2 AND2X2_8880 ( .A(u2__abc_44228_n18248), .B(u2__abc_44228_n18251), .Y(u2__abc_44228_n18252) );
  AND2X2 AND2X2_8881 ( .A(u2__abc_44228_n18253), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_root_40__FF_INPUT) );
  AND2X2 AND2X2_8882 ( .A(u2__abc_44228_n3062_bF_buf66), .B(sqrto_40_), .Y(u2__abc_44228_n18255) );
  AND2X2 AND2X2_8883 ( .A(u2__abc_44228_n18245), .B(sqrto_39_), .Y(u2__abc_44228_n18257) );
  AND2X2 AND2X2_8884 ( .A(u2__abc_44228_n18258), .B(u2__abc_44228_n18256), .Y(u2__abc_44228_n18259) );
  AND2X2 AND2X2_8885 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n3518), .Y(u2__abc_44228_n18261) );
  AND2X2 AND2X2_8886 ( .A(u2__abc_44228_n18262), .B(u2__abc_44228_n2972_bF_buf39), .Y(u2__abc_44228_n18263) );
  AND2X2 AND2X2_8887 ( .A(u2__abc_44228_n18260), .B(u2__abc_44228_n18263), .Y(u2__abc_44228_n18264) );
  AND2X2 AND2X2_8888 ( .A(u2__abc_44228_n18265), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_root_41__FF_INPUT) );
  AND2X2 AND2X2_8889 ( .A(u2__abc_44228_n3062_bF_buf65), .B(sqrto_41_), .Y(u2__abc_44228_n18267) );
  AND2X2 AND2X2_889 ( .A(u2__abc_44228_n3765), .B(u2__abc_44228_n3759_1), .Y(u2__abc_44228_n3766) );
  AND2X2 AND2X2_8890 ( .A(u2__abc_44228_n18257), .B(sqrto_40_), .Y(u2__abc_44228_n18269) );
  AND2X2 AND2X2_8891 ( .A(u2__abc_44228_n18270), .B(u2__abc_44228_n18268), .Y(u2__abc_44228_n18271) );
  AND2X2 AND2X2_8892 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n3511), .Y(u2__abc_44228_n18273) );
  AND2X2 AND2X2_8893 ( .A(u2__abc_44228_n18274), .B(u2__abc_44228_n2972_bF_buf38), .Y(u2__abc_44228_n18275) );
  AND2X2 AND2X2_8894 ( .A(u2__abc_44228_n18272), .B(u2__abc_44228_n18275), .Y(u2__abc_44228_n18276) );
  AND2X2 AND2X2_8895 ( .A(u2__abc_44228_n18277), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_root_42__FF_INPUT) );
  AND2X2 AND2X2_8896 ( .A(u2__abc_44228_n3062_bF_buf64), .B(sqrto_42_), .Y(u2__abc_44228_n18279) );
  AND2X2 AND2X2_8897 ( .A(u2__abc_44228_n18269), .B(sqrto_41_), .Y(u2__abc_44228_n18281) );
  AND2X2 AND2X2_8898 ( .A(u2__abc_44228_n18282), .B(u2__abc_44228_n18280), .Y(u2__abc_44228_n18283) );
  AND2X2 AND2X2_8899 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n3482), .Y(u2__abc_44228_n18285) );
  AND2X2 AND2X2_89 ( .A(_abc_64468_n867), .B(_abc_64468_n866), .Y(_auto_iopadmap_cc_313_execute_65414_124_) );
  AND2X2 AND2X2_890 ( .A(u2__abc_44228_n3767), .B(u2_remHi_110_), .Y(u2__abc_44228_n3768_1) );
  AND2X2 AND2X2_8900 ( .A(u2__abc_44228_n18286), .B(u2__abc_44228_n2972_bF_buf37), .Y(u2__abc_44228_n18287) );
  AND2X2 AND2X2_8901 ( .A(u2__abc_44228_n18284), .B(u2__abc_44228_n18287), .Y(u2__abc_44228_n18288) );
  AND2X2 AND2X2_8902 ( .A(u2__abc_44228_n18289), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_root_43__FF_INPUT) );
  AND2X2 AND2X2_8903 ( .A(u2__abc_44228_n3062_bF_buf63), .B(sqrto_43_), .Y(u2__abc_44228_n18291) );
  AND2X2 AND2X2_8904 ( .A(u2__abc_44228_n18281), .B(sqrto_42_), .Y(u2__abc_44228_n18293) );
  AND2X2 AND2X2_8905 ( .A(u2__abc_44228_n18294), .B(u2__abc_44228_n18292), .Y(u2__abc_44228_n18295) );
  AND2X2 AND2X2_8906 ( .A(u2__abc_44228_n2983_bF_buf104), .B(u2__abc_44228_n3488), .Y(u2__abc_44228_n18297) );
  AND2X2 AND2X2_8907 ( .A(u2__abc_44228_n18298), .B(u2__abc_44228_n2972_bF_buf36), .Y(u2__abc_44228_n18299) );
  AND2X2 AND2X2_8908 ( .A(u2__abc_44228_n18296), .B(u2__abc_44228_n18299), .Y(u2__abc_44228_n18300) );
  AND2X2 AND2X2_8909 ( .A(u2__abc_44228_n18301), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_root_44__FF_INPUT) );
  AND2X2 AND2X2_891 ( .A(u2__abc_44228_n3769), .B(sqrto_110_), .Y(u2__abc_44228_n3770) );
  AND2X2 AND2X2_8910 ( .A(u2__abc_44228_n3062_bF_buf62), .B(sqrto_44_), .Y(u2__abc_44228_n18303) );
  AND2X2 AND2X2_8911 ( .A(u2__abc_44228_n18293), .B(sqrto_43_), .Y(u2__abc_44228_n18305) );
  AND2X2 AND2X2_8912 ( .A(u2__abc_44228_n18306), .B(u2__abc_44228_n18304), .Y(u2__abc_44228_n18307) );
  AND2X2 AND2X2_8913 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n3475_1), .Y(u2__abc_44228_n18309) );
  AND2X2 AND2X2_8914 ( .A(u2__abc_44228_n18310), .B(u2__abc_44228_n2972_bF_buf35), .Y(u2__abc_44228_n18311) );
  AND2X2 AND2X2_8915 ( .A(u2__abc_44228_n18308), .B(u2__abc_44228_n18311), .Y(u2__abc_44228_n18312) );
  AND2X2 AND2X2_8916 ( .A(u2__abc_44228_n18313), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_root_45__FF_INPUT) );
  AND2X2 AND2X2_8917 ( .A(u2__abc_44228_n3062_bF_buf61), .B(sqrto_45_), .Y(u2__abc_44228_n18315) );
  AND2X2 AND2X2_8918 ( .A(u2__abc_44228_n18305), .B(sqrto_44_), .Y(u2__abc_44228_n18317) );
  AND2X2 AND2X2_8919 ( .A(u2__abc_44228_n18318), .B(u2__abc_44228_n18316), .Y(u2__abc_44228_n18319) );
  AND2X2 AND2X2_892 ( .A(u2__abc_44228_n3773), .B(u2_remHi_111_), .Y(u2__abc_44228_n3774) );
  AND2X2 AND2X2_8920 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n3468), .Y(u2__abc_44228_n18321) );
  AND2X2 AND2X2_8921 ( .A(u2__abc_44228_n18322), .B(u2__abc_44228_n2972_bF_buf34), .Y(u2__abc_44228_n18323) );
  AND2X2 AND2X2_8922 ( .A(u2__abc_44228_n18320), .B(u2__abc_44228_n18323), .Y(u2__abc_44228_n18324) );
  AND2X2 AND2X2_8923 ( .A(u2__abc_44228_n18325), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_root_46__FF_INPUT) );
  AND2X2 AND2X2_8924 ( .A(u2__abc_44228_n3062_bF_buf60), .B(sqrto_46_), .Y(u2__abc_44228_n18327) );
  AND2X2 AND2X2_8925 ( .A(u2__abc_44228_n18317), .B(sqrto_45_), .Y(u2__abc_44228_n18329) );
  AND2X2 AND2X2_8926 ( .A(u2__abc_44228_n18330), .B(u2__abc_44228_n18328), .Y(u2__abc_44228_n18331) );
  AND2X2 AND2X2_8927 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n3458), .Y(u2__abc_44228_n18333) );
  AND2X2 AND2X2_8928 ( .A(u2__abc_44228_n18334), .B(u2__abc_44228_n2972_bF_buf33), .Y(u2__abc_44228_n18335) );
  AND2X2 AND2X2_8929 ( .A(u2__abc_44228_n18332), .B(u2__abc_44228_n18335), .Y(u2__abc_44228_n18336) );
  AND2X2 AND2X2_893 ( .A(u2__abc_44228_n3776), .B(sqrto_111_), .Y(u2__abc_44228_n3777) );
  AND2X2 AND2X2_8930 ( .A(u2__abc_44228_n18337), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_root_47__FF_INPUT) );
  AND2X2 AND2X2_8931 ( .A(u2__abc_44228_n3062_bF_buf59), .B(sqrto_47_), .Y(u2__abc_44228_n18339) );
  AND2X2 AND2X2_8932 ( .A(u2__abc_44228_n18329), .B(sqrto_46_), .Y(u2__abc_44228_n18341) );
  AND2X2 AND2X2_8933 ( .A(u2__abc_44228_n18342), .B(u2__abc_44228_n18340), .Y(u2__abc_44228_n18343) );
  AND2X2 AND2X2_8934 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n3451), .Y(u2__abc_44228_n18345) );
  AND2X2 AND2X2_8935 ( .A(u2__abc_44228_n18346), .B(u2__abc_44228_n2972_bF_buf32), .Y(u2__abc_44228_n18347) );
  AND2X2 AND2X2_8936 ( .A(u2__abc_44228_n18344), .B(u2__abc_44228_n18347), .Y(u2__abc_44228_n18348) );
  AND2X2 AND2X2_8937 ( .A(u2__abc_44228_n18349), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_root_48__FF_INPUT) );
  AND2X2 AND2X2_8938 ( .A(u2__abc_44228_n3062_bF_buf58), .B(sqrto_48_), .Y(u2__abc_44228_n18351) );
  AND2X2 AND2X2_8939 ( .A(u2__abc_44228_n18341), .B(sqrto_47_), .Y(u2__abc_44228_n18353) );
  AND2X2 AND2X2_894 ( .A(u2__abc_44228_n3775), .B(u2__abc_44228_n3778), .Y(u2__abc_44228_n3779_1) );
  AND2X2 AND2X2_8940 ( .A(u2__abc_44228_n18354), .B(u2__abc_44228_n18352), .Y(u2__abc_44228_n18355) );
  AND2X2 AND2X2_8941 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n3444), .Y(u2__abc_44228_n18357) );
  AND2X2 AND2X2_8942 ( .A(u2__abc_44228_n18358), .B(u2__abc_44228_n2972_bF_buf31), .Y(u2__abc_44228_n18359) );
  AND2X2 AND2X2_8943 ( .A(u2__abc_44228_n18356), .B(u2__abc_44228_n18359), .Y(u2__abc_44228_n18360) );
  AND2X2 AND2X2_8944 ( .A(u2__abc_44228_n18361), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_root_49__FF_INPUT) );
  AND2X2 AND2X2_8945 ( .A(u2__abc_44228_n3062_bF_buf57), .B(sqrto_49_), .Y(u2__abc_44228_n18363) );
  AND2X2 AND2X2_8946 ( .A(u2__abc_44228_n18353), .B(sqrto_48_), .Y(u2__abc_44228_n18365) );
  AND2X2 AND2X2_8947 ( .A(u2__abc_44228_n18366), .B(u2__abc_44228_n18364), .Y(u2__abc_44228_n18367) );
  AND2X2 AND2X2_8948 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n3437), .Y(u2__abc_44228_n18369) );
  AND2X2 AND2X2_8949 ( .A(u2__abc_44228_n18370), .B(u2__abc_44228_n2972_bF_buf30), .Y(u2__abc_44228_n18371) );
  AND2X2 AND2X2_895 ( .A(u2__abc_44228_n3772), .B(u2__abc_44228_n3779_1), .Y(u2__abc_44228_n3780) );
  AND2X2 AND2X2_8950 ( .A(u2__abc_44228_n18368), .B(u2__abc_44228_n18371), .Y(u2__abc_44228_n18372) );
  AND2X2 AND2X2_8951 ( .A(u2__abc_44228_n18373), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_root_50__FF_INPUT) );
  AND2X2 AND2X2_8952 ( .A(u2__abc_44228_n3062_bF_buf56), .B(sqrto_50_), .Y(u2__abc_44228_n18375) );
  AND2X2 AND2X2_8953 ( .A(u2__abc_44228_n18365), .B(sqrto_49_), .Y(u2__abc_44228_n18377) );
  AND2X2 AND2X2_8954 ( .A(u2__abc_44228_n18378), .B(u2__abc_44228_n18376), .Y(u2__abc_44228_n18379) );
  AND2X2 AND2X2_8955 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n3422), .Y(u2__abc_44228_n18381) );
  AND2X2 AND2X2_8956 ( .A(u2__abc_44228_n18382), .B(u2__abc_44228_n2972_bF_buf29), .Y(u2__abc_44228_n18383) );
  AND2X2 AND2X2_8957 ( .A(u2__abc_44228_n18380), .B(u2__abc_44228_n18383), .Y(u2__abc_44228_n18384) );
  AND2X2 AND2X2_8958 ( .A(u2__abc_44228_n18385), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_root_51__FF_INPUT) );
  AND2X2 AND2X2_8959 ( .A(u2__abc_44228_n3062_bF_buf55), .B(sqrto_51_), .Y(u2__abc_44228_n18387) );
  AND2X2 AND2X2_896 ( .A(u2__abc_44228_n3766), .B(u2__abc_44228_n3780), .Y(u2__abc_44228_n3781) );
  AND2X2 AND2X2_8960 ( .A(u2__abc_44228_n18377), .B(sqrto_50_), .Y(u2__abc_44228_n18389) );
  AND2X2 AND2X2_8961 ( .A(u2__abc_44228_n18390), .B(u2__abc_44228_n18388), .Y(u2__abc_44228_n18391) );
  AND2X2 AND2X2_8962 ( .A(u2__abc_44228_n2983_bF_buf88), .B(u2__abc_44228_n3428), .Y(u2__abc_44228_n18393) );
  AND2X2 AND2X2_8963 ( .A(u2__abc_44228_n18394), .B(u2__abc_44228_n2972_bF_buf28), .Y(u2__abc_44228_n18395) );
  AND2X2 AND2X2_8964 ( .A(u2__abc_44228_n18392), .B(u2__abc_44228_n18395), .Y(u2__abc_44228_n18396) );
  AND2X2 AND2X2_8965 ( .A(u2__abc_44228_n18397), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_root_52__FF_INPUT) );
  AND2X2 AND2X2_8966 ( .A(u2__abc_44228_n3062_bF_buf54), .B(sqrto_52_), .Y(u2__abc_44228_n18399) );
  AND2X2 AND2X2_8967 ( .A(u2__abc_44228_n18389), .B(sqrto_51_), .Y(u2__abc_44228_n18401) );
  AND2X2 AND2X2_8968 ( .A(u2__abc_44228_n18402), .B(u2__abc_44228_n18400), .Y(u2__abc_44228_n18403) );
  AND2X2 AND2X2_8969 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n3415), .Y(u2__abc_44228_n18405) );
  AND2X2 AND2X2_897 ( .A(u2__abc_44228_n3781), .B(u2__abc_44228_n3752), .Y(u2__abc_44228_n3782) );
  AND2X2 AND2X2_8970 ( .A(u2__abc_44228_n18406), .B(u2__abc_44228_n2972_bF_buf27), .Y(u2__abc_44228_n18407) );
  AND2X2 AND2X2_8971 ( .A(u2__abc_44228_n18404), .B(u2__abc_44228_n18407), .Y(u2__abc_44228_n18408) );
  AND2X2 AND2X2_8972 ( .A(u2__abc_44228_n18409), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_root_53__FF_INPUT) );
  AND2X2 AND2X2_8973 ( .A(u2__abc_44228_n3062_bF_buf53), .B(sqrto_53_), .Y(u2__abc_44228_n18411) );
  AND2X2 AND2X2_8974 ( .A(u2__abc_44228_n18401), .B(sqrto_52_), .Y(u2__abc_44228_n18413) );
  AND2X2 AND2X2_8975 ( .A(u2__abc_44228_n18414), .B(u2__abc_44228_n18412), .Y(u2__abc_44228_n18415) );
  AND2X2 AND2X2_8976 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n3408), .Y(u2__abc_44228_n18417) );
  AND2X2 AND2X2_8977 ( .A(u2__abc_44228_n18418), .B(u2__abc_44228_n2972_bF_buf26), .Y(u2__abc_44228_n18419) );
  AND2X2 AND2X2_8978 ( .A(u2__abc_44228_n18416), .B(u2__abc_44228_n18419), .Y(u2__abc_44228_n18420) );
  AND2X2 AND2X2_8979 ( .A(u2__abc_44228_n18421), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_root_54__FF_INPUT) );
  AND2X2 AND2X2_898 ( .A(u2__abc_44228_n3782), .B(u2__abc_44228_n3723_1), .Y(u2__abc_44228_n3783) );
  AND2X2 AND2X2_8980 ( .A(u2__abc_44228_n3062_bF_buf52), .B(sqrto_54_), .Y(u2__abc_44228_n18423) );
  AND2X2 AND2X2_8981 ( .A(u2__abc_44228_n18413), .B(sqrto_53_), .Y(u2__abc_44228_n18425) );
  AND2X2 AND2X2_8982 ( .A(u2__abc_44228_n18426), .B(u2__abc_44228_n18424), .Y(u2__abc_44228_n18427) );
  AND2X2 AND2X2_8983 ( .A(u2__abc_44228_n2983_bF_buf82), .B(u2__abc_44228_n3399), .Y(u2__abc_44228_n18429) );
  AND2X2 AND2X2_8984 ( .A(u2__abc_44228_n18430), .B(u2__abc_44228_n2972_bF_buf25), .Y(u2__abc_44228_n18431) );
  AND2X2 AND2X2_8985 ( .A(u2__abc_44228_n18428), .B(u2__abc_44228_n18431), .Y(u2__abc_44228_n18432) );
  AND2X2 AND2X2_8986 ( .A(u2__abc_44228_n18433), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_root_55__FF_INPUT) );
  AND2X2 AND2X2_8987 ( .A(u2__abc_44228_n3062_bF_buf51), .B(sqrto_55_), .Y(u2__abc_44228_n18435) );
  AND2X2 AND2X2_8988 ( .A(u2__abc_44228_n18425), .B(sqrto_54_), .Y(u2__abc_44228_n18437) );
  AND2X2 AND2X2_8989 ( .A(u2__abc_44228_n18438), .B(u2__abc_44228_n18436), .Y(u2__abc_44228_n18439) );
  AND2X2 AND2X2_899 ( .A(u2__abc_44228_n3784), .B(u2_remHi_109_), .Y(u2__abc_44228_n3785) );
  AND2X2 AND2X2_8990 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n3392), .Y(u2__abc_44228_n18441) );
  AND2X2 AND2X2_8991 ( .A(u2__abc_44228_n18442), .B(u2__abc_44228_n2972_bF_buf24), .Y(u2__abc_44228_n18443) );
  AND2X2 AND2X2_8992 ( .A(u2__abc_44228_n18440), .B(u2__abc_44228_n18443), .Y(u2__abc_44228_n18444) );
  AND2X2 AND2X2_8993 ( .A(u2__abc_44228_n18445), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_root_56__FF_INPUT) );
  AND2X2 AND2X2_8994 ( .A(u2__abc_44228_n3062_bF_buf50), .B(sqrto_56_), .Y(u2__abc_44228_n18447) );
  AND2X2 AND2X2_8995 ( .A(u2__abc_44228_n18437), .B(sqrto_55_), .Y(u2__abc_44228_n18449) );
  AND2X2 AND2X2_8996 ( .A(u2__abc_44228_n18450), .B(u2__abc_44228_n18448), .Y(u2__abc_44228_n18451) );
  AND2X2 AND2X2_8997 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n3385), .Y(u2__abc_44228_n18453) );
  AND2X2 AND2X2_8998 ( .A(u2__abc_44228_n18454), .B(u2__abc_44228_n2972_bF_buf23), .Y(u2__abc_44228_n18455) );
  AND2X2 AND2X2_8999 ( .A(u2__abc_44228_n18452), .B(u2__abc_44228_n18455), .Y(u2__abc_44228_n18456) );
  AND2X2 AND2X2_9 ( .A(_abc_64468_n753_bF_buf5), .B(sqrto_8_), .Y(_auto_iopadmap_cc_313_execute_65414_44_) );
  AND2X2 AND2X2_90 ( .A(_abc_64468_n870), .B(_abc_64468_n869), .Y(_auto_iopadmap_cc_313_execute_65414_125_) );
  AND2X2 AND2X2_900 ( .A(u2__abc_44228_n3787), .B(sqrto_109_), .Y(u2__abc_44228_n3788) );
  AND2X2 AND2X2_9000 ( .A(u2__abc_44228_n18457), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_root_57__FF_INPUT) );
  AND2X2 AND2X2_9001 ( .A(u2__abc_44228_n3062_bF_buf49), .B(sqrto_57_), .Y(u2__abc_44228_n18459) );
  AND2X2 AND2X2_9002 ( .A(u2__abc_44228_n18449), .B(sqrto_56_), .Y(u2__abc_44228_n18461) );
  AND2X2 AND2X2_9003 ( .A(u2__abc_44228_n18462), .B(u2__abc_44228_n18460), .Y(u2__abc_44228_n18463) );
  AND2X2 AND2X2_9004 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n3378), .Y(u2__abc_44228_n18465) );
  AND2X2 AND2X2_9005 ( .A(u2__abc_44228_n18466), .B(u2__abc_44228_n2972_bF_buf22), .Y(u2__abc_44228_n18467) );
  AND2X2 AND2X2_9006 ( .A(u2__abc_44228_n18464), .B(u2__abc_44228_n18467), .Y(u2__abc_44228_n18468) );
  AND2X2 AND2X2_9007 ( .A(u2__abc_44228_n18469), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_root_58__FF_INPUT) );
  AND2X2 AND2X2_9008 ( .A(u2__abc_44228_n3062_bF_buf48), .B(sqrto_58_), .Y(u2__abc_44228_n18471) );
  AND2X2 AND2X2_9009 ( .A(u2__abc_44228_n18461), .B(sqrto_57_), .Y(u2__abc_44228_n18473) );
  AND2X2 AND2X2_901 ( .A(u2__abc_44228_n3786), .B(u2__abc_44228_n3789_1), .Y(u2__abc_44228_n3790) );
  AND2X2 AND2X2_9010 ( .A(u2__abc_44228_n18474), .B(u2__abc_44228_n18472), .Y(u2__abc_44228_n18475) );
  AND2X2 AND2X2_9011 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n3363), .Y(u2__abc_44228_n18477) );
  AND2X2 AND2X2_9012 ( .A(u2__abc_44228_n18478), .B(u2__abc_44228_n2972_bF_buf21), .Y(u2__abc_44228_n18479) );
  AND2X2 AND2X2_9013 ( .A(u2__abc_44228_n18476), .B(u2__abc_44228_n18479), .Y(u2__abc_44228_n18480) );
  AND2X2 AND2X2_9014 ( .A(u2__abc_44228_n18481), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_root_59__FF_INPUT) );
  AND2X2 AND2X2_9015 ( .A(u2__abc_44228_n3062_bF_buf47), .B(sqrto_59_), .Y(u2__abc_44228_n18483) );
  AND2X2 AND2X2_9016 ( .A(u2__abc_44228_n18473), .B(sqrto_58_), .Y(u2__abc_44228_n18485) );
  AND2X2 AND2X2_9017 ( .A(u2__abc_44228_n18486), .B(u2__abc_44228_n18484), .Y(u2__abc_44228_n18487) );
  AND2X2 AND2X2_9018 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n3369), .Y(u2__abc_44228_n18489) );
  AND2X2 AND2X2_9019 ( .A(u2__abc_44228_n18490), .B(u2__abc_44228_n2972_bF_buf20), .Y(u2__abc_44228_n18491) );
  AND2X2 AND2X2_902 ( .A(u2__abc_44228_n3791), .B(u2_remHi_108_), .Y(u2__abc_44228_n3792) );
  AND2X2 AND2X2_9020 ( .A(u2__abc_44228_n18488), .B(u2__abc_44228_n18491), .Y(u2__abc_44228_n18492) );
  AND2X2 AND2X2_9021 ( .A(u2__abc_44228_n18493), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_root_60__FF_INPUT) );
  AND2X2 AND2X2_9022 ( .A(u2__abc_44228_n3062_bF_buf46), .B(sqrto_60_), .Y(u2__abc_44228_n18495) );
  AND2X2 AND2X2_9023 ( .A(u2__abc_44228_n18485), .B(sqrto_59_), .Y(u2__abc_44228_n18497) );
  AND2X2 AND2X2_9024 ( .A(u2__abc_44228_n18498), .B(u2__abc_44228_n18496), .Y(u2__abc_44228_n18499) );
  AND2X2 AND2X2_9025 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n3356), .Y(u2__abc_44228_n18501) );
  AND2X2 AND2X2_9026 ( .A(u2__abc_44228_n18502), .B(u2__abc_44228_n2972_bF_buf19), .Y(u2__abc_44228_n18503) );
  AND2X2 AND2X2_9027 ( .A(u2__abc_44228_n18500), .B(u2__abc_44228_n18503), .Y(u2__abc_44228_n18504) );
  AND2X2 AND2X2_9028 ( .A(u2__abc_44228_n18505), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_root_61__FF_INPUT) );
  AND2X2 AND2X2_9029 ( .A(u2__abc_44228_n3062_bF_buf45), .B(sqrto_61_), .Y(u2__abc_44228_n18507) );
  AND2X2 AND2X2_903 ( .A(u2__abc_44228_n3793), .B(sqrto_108_), .Y(u2__abc_44228_n3794) );
  AND2X2 AND2X2_9030 ( .A(u2__abc_44228_n18497), .B(sqrto_60_), .Y(u2__abc_44228_n18509) );
  AND2X2 AND2X2_9031 ( .A(u2__abc_44228_n18510), .B(u2__abc_44228_n18508), .Y(u2__abc_44228_n18511) );
  AND2X2 AND2X2_9032 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n3349), .Y(u2__abc_44228_n18513) );
  AND2X2 AND2X2_9033 ( .A(u2__abc_44228_n18514), .B(u2__abc_44228_n2972_bF_buf18), .Y(u2__abc_44228_n18515) );
  AND2X2 AND2X2_9034 ( .A(u2__abc_44228_n18512), .B(u2__abc_44228_n18515), .Y(u2__abc_44228_n18516) );
  AND2X2 AND2X2_9035 ( .A(u2__abc_44228_n18517), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_root_62__FF_INPUT) );
  AND2X2 AND2X2_9036 ( .A(u2__abc_44228_n3062_bF_buf44), .B(sqrto_62_), .Y(u2__abc_44228_n18519) );
  AND2X2 AND2X2_9037 ( .A(u2__abc_44228_n18509), .B(sqrto_61_), .Y(u2__abc_44228_n18521) );
  AND2X2 AND2X2_9038 ( .A(u2__abc_44228_n18522), .B(u2__abc_44228_n18520), .Y(u2__abc_44228_n18523) );
  AND2X2 AND2X2_9039 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n4129), .Y(u2__abc_44228_n18525) );
  AND2X2 AND2X2_904 ( .A(u2__abc_44228_n3796), .B(u2__abc_44228_n3790), .Y(u2__abc_44228_n3797) );
  AND2X2 AND2X2_9040 ( .A(u2__abc_44228_n18526), .B(u2__abc_44228_n2972_bF_buf17), .Y(u2__abc_44228_n18527) );
  AND2X2 AND2X2_9041 ( .A(u2__abc_44228_n18524), .B(u2__abc_44228_n18527), .Y(u2__abc_44228_n18528) );
  AND2X2 AND2X2_9042 ( .A(u2__abc_44228_n18529), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_root_63__FF_INPUT) );
  AND2X2 AND2X2_9043 ( .A(u2__abc_44228_n3062_bF_buf43), .B(sqrto_63_), .Y(u2__abc_44228_n18531) );
  AND2X2 AND2X2_9044 ( .A(u2__abc_44228_n18521), .B(sqrto_62_), .Y(u2__abc_44228_n18533) );
  AND2X2 AND2X2_9045 ( .A(u2__abc_44228_n18534), .B(u2__abc_44228_n18532), .Y(u2__abc_44228_n18535) );
  AND2X2 AND2X2_9046 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n4122), .Y(u2__abc_44228_n18537) );
  AND2X2 AND2X2_9047 ( .A(u2__abc_44228_n18538), .B(u2__abc_44228_n2972_bF_buf16), .Y(u2__abc_44228_n18539) );
  AND2X2 AND2X2_9048 ( .A(u2__abc_44228_n18536), .B(u2__abc_44228_n18539), .Y(u2__abc_44228_n18540) );
  AND2X2 AND2X2_9049 ( .A(u2__abc_44228_n18541), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_root_64__FF_INPUT) );
  AND2X2 AND2X2_905 ( .A(u2__abc_44228_n3798_1), .B(u2_remHi_106_), .Y(u2__abc_44228_n3799) );
  AND2X2 AND2X2_9050 ( .A(u2__abc_44228_n3062_bF_buf42), .B(sqrto_64_), .Y(u2__abc_44228_n18543) );
  AND2X2 AND2X2_9051 ( .A(u2__abc_44228_n18533), .B(sqrto_63_), .Y(u2__abc_44228_n18545) );
  AND2X2 AND2X2_9052 ( .A(u2__abc_44228_n18546), .B(u2__abc_44228_n18544), .Y(u2__abc_44228_n18547) );
  AND2X2 AND2X2_9053 ( .A(u2__abc_44228_n2983_bF_buf62), .B(u2__abc_44228_n4118), .Y(u2__abc_44228_n18549) );
  AND2X2 AND2X2_9054 ( .A(u2__abc_44228_n18550), .B(u2__abc_44228_n2972_bF_buf15), .Y(u2__abc_44228_n18551) );
  AND2X2 AND2X2_9055 ( .A(u2__abc_44228_n18548), .B(u2__abc_44228_n18551), .Y(u2__abc_44228_n18552) );
  AND2X2 AND2X2_9056 ( .A(u2__abc_44228_n18553), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_root_65__FF_INPUT) );
  AND2X2 AND2X2_9057 ( .A(u2__abc_44228_n3062_bF_buf41), .B(sqrto_65_), .Y(u2__abc_44228_n18555) );
  AND2X2 AND2X2_9058 ( .A(u2__abc_44228_n18545), .B(sqrto_64_), .Y(u2__abc_44228_n18557) );
  AND2X2 AND2X2_9059 ( .A(u2__abc_44228_n18558), .B(u2__abc_44228_n18556), .Y(u2__abc_44228_n18559) );
  AND2X2 AND2X2_906 ( .A(u2__abc_44228_n3800), .B(sqrto_106_), .Y(u2__abc_44228_n3801) );
  AND2X2 AND2X2_9060 ( .A(u2__abc_44228_n2983_bF_buf60), .B(u2__abc_44228_n4113), .Y(u2__abc_44228_n18561) );
  AND2X2 AND2X2_9061 ( .A(u2__abc_44228_n18562), .B(u2__abc_44228_n2972_bF_buf14), .Y(u2__abc_44228_n18563) );
  AND2X2 AND2X2_9062 ( .A(u2__abc_44228_n18560), .B(u2__abc_44228_n18563), .Y(u2__abc_44228_n18564) );
  AND2X2 AND2X2_9063 ( .A(u2__abc_44228_n18565), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_root_66__FF_INPUT) );
  AND2X2 AND2X2_9064 ( .A(u2__abc_44228_n3062_bF_buf40), .B(sqrto_66_), .Y(u2__abc_44228_n18567) );
  AND2X2 AND2X2_9065 ( .A(u2__abc_44228_n18557), .B(sqrto_65_), .Y(u2__abc_44228_n18569) );
  AND2X2 AND2X2_9066 ( .A(u2__abc_44228_n18570), .B(u2__abc_44228_n18568), .Y(u2__abc_44228_n18571) );
  AND2X2 AND2X2_9067 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n4103), .Y(u2__abc_44228_n18573) );
  AND2X2 AND2X2_9068 ( .A(u2__abc_44228_n18574), .B(u2__abc_44228_n2972_bF_buf13), .Y(u2__abc_44228_n18575) );
  AND2X2 AND2X2_9069 ( .A(u2__abc_44228_n18572), .B(u2__abc_44228_n18575), .Y(u2__abc_44228_n18576) );
  AND2X2 AND2X2_907 ( .A(u2__abc_44228_n3804), .B(u2_remHi_107_), .Y(u2__abc_44228_n3805) );
  AND2X2 AND2X2_9070 ( .A(u2__abc_44228_n18577), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_root_67__FF_INPUT) );
  AND2X2 AND2X2_9071 ( .A(u2__abc_44228_n3062_bF_buf39), .B(sqrto_67_), .Y(u2__abc_44228_n18579) );
  AND2X2 AND2X2_9072 ( .A(u2__abc_44228_n18569), .B(sqrto_66_), .Y(u2__abc_44228_n18581) );
  AND2X2 AND2X2_9073 ( .A(u2__abc_44228_n18582), .B(u2__abc_44228_n18580), .Y(u2__abc_44228_n18583) );
  AND2X2 AND2X2_9074 ( .A(u2__abc_44228_n2983_bF_buf56), .B(u2__abc_44228_n4096), .Y(u2__abc_44228_n18585) );
  AND2X2 AND2X2_9075 ( .A(u2__abc_44228_n18586), .B(u2__abc_44228_n2972_bF_buf12), .Y(u2__abc_44228_n18587) );
  AND2X2 AND2X2_9076 ( .A(u2__abc_44228_n18584), .B(u2__abc_44228_n18587), .Y(u2__abc_44228_n18588) );
  AND2X2 AND2X2_9077 ( .A(u2__abc_44228_n18589), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_root_68__FF_INPUT) );
  AND2X2 AND2X2_9078 ( .A(u2__abc_44228_n3062_bF_buf38), .B(sqrto_68_), .Y(u2__abc_44228_n18591) );
  AND2X2 AND2X2_9079 ( .A(u2__abc_44228_n18581), .B(sqrto_67_), .Y(u2__abc_44228_n18593) );
  AND2X2 AND2X2_908 ( .A(u2__abc_44228_n3807_1), .B(sqrto_107_), .Y(u2__abc_44228_n3808) );
  AND2X2 AND2X2_9080 ( .A(u2__abc_44228_n18594), .B(u2__abc_44228_n18592), .Y(u2__abc_44228_n18595) );
  AND2X2 AND2X2_9081 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n4089), .Y(u2__abc_44228_n18597) );
  AND2X2 AND2X2_9082 ( .A(u2__abc_44228_n18598), .B(u2__abc_44228_n2972_bF_buf11), .Y(u2__abc_44228_n18599) );
  AND2X2 AND2X2_9083 ( .A(u2__abc_44228_n18596), .B(u2__abc_44228_n18599), .Y(u2__abc_44228_n18600) );
  AND2X2 AND2X2_9084 ( .A(u2__abc_44228_n18601), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_root_69__FF_INPUT) );
  AND2X2 AND2X2_9085 ( .A(u2__abc_44228_n3062_bF_buf37), .B(sqrto_69_), .Y(u2__abc_44228_n18603) );
  AND2X2 AND2X2_9086 ( .A(u2__abc_44228_n18593), .B(sqrto_68_), .Y(u2__abc_44228_n18605) );
  AND2X2 AND2X2_9087 ( .A(u2__abc_44228_n18606), .B(u2__abc_44228_n18604), .Y(u2__abc_44228_n18607) );
  AND2X2 AND2X2_9088 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n4082), .Y(u2__abc_44228_n18609) );
  AND2X2 AND2X2_9089 ( .A(u2__abc_44228_n18610), .B(u2__abc_44228_n2972_bF_buf10), .Y(u2__abc_44228_n18611) );
  AND2X2 AND2X2_909 ( .A(u2__abc_44228_n3806), .B(u2__abc_44228_n3809), .Y(u2__abc_44228_n3810) );
  AND2X2 AND2X2_9090 ( .A(u2__abc_44228_n18608), .B(u2__abc_44228_n18611), .Y(u2__abc_44228_n18612) );
  AND2X2 AND2X2_9091 ( .A(u2__abc_44228_n18613), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_root_70__FF_INPUT) );
  AND2X2 AND2X2_9092 ( .A(u2__abc_44228_n3062_bF_buf36), .B(sqrto_70_), .Y(u2__abc_44228_n18615) );
  AND2X2 AND2X2_9093 ( .A(u2__abc_44228_n18605), .B(sqrto_69_), .Y(u2__abc_44228_n18617) );
  AND2X2 AND2X2_9094 ( .A(u2__abc_44228_n18618), .B(u2__abc_44228_n18616), .Y(u2__abc_44228_n18619) );
  AND2X2 AND2X2_9095 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2__abc_44228_n4059), .Y(u2__abc_44228_n18621) );
  AND2X2 AND2X2_9096 ( .A(u2__abc_44228_n18622), .B(u2__abc_44228_n2972_bF_buf9), .Y(u2__abc_44228_n18623) );
  AND2X2 AND2X2_9097 ( .A(u2__abc_44228_n18620), .B(u2__abc_44228_n18623), .Y(u2__abc_44228_n18624) );
  AND2X2 AND2X2_9098 ( .A(u2__abc_44228_n18625), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_root_71__FF_INPUT) );
  AND2X2 AND2X2_9099 ( .A(u2__abc_44228_n3062_bF_buf35), .B(sqrto_71_), .Y(u2__abc_44228_n18627) );
  AND2X2 AND2X2_91 ( .A(_abc_64468_n873), .B(_abc_64468_n872), .Y(_auto_iopadmap_cc_313_execute_65414_126_) );
  AND2X2 AND2X2_910 ( .A(u2__abc_44228_n3803), .B(u2__abc_44228_n3810), .Y(u2__abc_44228_n3811) );
  AND2X2 AND2X2_9100 ( .A(u2__abc_44228_n18617), .B(sqrto_70_), .Y(u2__abc_44228_n18629) );
  AND2X2 AND2X2_9101 ( .A(u2__abc_44228_n18630), .B(u2__abc_44228_n18628), .Y(u2__abc_44228_n18631) );
  AND2X2 AND2X2_9102 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n4052), .Y(u2__abc_44228_n18633) );
  AND2X2 AND2X2_9103 ( .A(u2__abc_44228_n18634), .B(u2__abc_44228_n2972_bF_buf8), .Y(u2__abc_44228_n18635) );
  AND2X2 AND2X2_9104 ( .A(u2__abc_44228_n18632), .B(u2__abc_44228_n18635), .Y(u2__abc_44228_n18636) );
  AND2X2 AND2X2_9105 ( .A(u2__abc_44228_n18637), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_root_72__FF_INPUT) );
  AND2X2 AND2X2_9106 ( .A(u2__abc_44228_n3062_bF_buf34), .B(sqrto_72_), .Y(u2__abc_44228_n18639) );
  AND2X2 AND2X2_9107 ( .A(u2__abc_44228_n18629), .B(sqrto_71_), .Y(u2__abc_44228_n18641) );
  AND2X2 AND2X2_9108 ( .A(u2__abc_44228_n18642), .B(u2__abc_44228_n18640), .Y(u2__abc_44228_n18643) );
  AND2X2 AND2X2_9109 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n4073), .Y(u2__abc_44228_n18645) );
  AND2X2 AND2X2_911 ( .A(u2__abc_44228_n3797), .B(u2__abc_44228_n3811), .Y(u2__abc_44228_n3812) );
  AND2X2 AND2X2_9110 ( .A(u2__abc_44228_n18646), .B(u2__abc_44228_n2972_bF_buf7), .Y(u2__abc_44228_n18647) );
  AND2X2 AND2X2_9111 ( .A(u2__abc_44228_n18644), .B(u2__abc_44228_n18647), .Y(u2__abc_44228_n18648) );
  AND2X2 AND2X2_9112 ( .A(u2__abc_44228_n18649), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_root_73__FF_INPUT) );
  AND2X2 AND2X2_9113 ( .A(u2__abc_44228_n3062_bF_buf33), .B(sqrto_73_), .Y(u2__abc_44228_n18651) );
  AND2X2 AND2X2_9114 ( .A(u2__abc_44228_n18641), .B(sqrto_72_), .Y(u2__abc_44228_n18653) );
  AND2X2 AND2X2_9115 ( .A(u2__abc_44228_n18654), .B(u2__abc_44228_n18652), .Y(u2__abc_44228_n18655) );
  AND2X2 AND2X2_9116 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n4066), .Y(u2__abc_44228_n18657) );
  AND2X2 AND2X2_9117 ( .A(u2__abc_44228_n18658), .B(u2__abc_44228_n2972_bF_buf6), .Y(u2__abc_44228_n18659) );
  AND2X2 AND2X2_9118 ( .A(u2__abc_44228_n18656), .B(u2__abc_44228_n18659), .Y(u2__abc_44228_n18660) );
  AND2X2 AND2X2_9119 ( .A(u2__abc_44228_n18661), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_root_74__FF_INPUT) );
  AND2X2 AND2X2_912 ( .A(u2__abc_44228_n3813), .B(u2_remHi_103_), .Y(u2__abc_44228_n3814) );
  AND2X2 AND2X2_9120 ( .A(u2__abc_44228_n3062_bF_buf32), .B(sqrto_74_), .Y(u2__abc_44228_n18663) );
  AND2X2 AND2X2_9121 ( .A(u2__abc_44228_n18653), .B(sqrto_73_), .Y(u2__abc_44228_n18665) );
  AND2X2 AND2X2_9122 ( .A(u2__abc_44228_n18666), .B(u2__abc_44228_n18664), .Y(u2__abc_44228_n18667) );
  AND2X2 AND2X2_9123 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n4037), .Y(u2__abc_44228_n18669) );
  AND2X2 AND2X2_9124 ( .A(u2__abc_44228_n18670), .B(u2__abc_44228_n2972_bF_buf5), .Y(u2__abc_44228_n18671) );
  AND2X2 AND2X2_9125 ( .A(u2__abc_44228_n18668), .B(u2__abc_44228_n18671), .Y(u2__abc_44228_n18672) );
  AND2X2 AND2X2_9126 ( .A(u2__abc_44228_n18673), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_root_75__FF_INPUT) );
  AND2X2 AND2X2_9127 ( .A(u2__abc_44228_n3062_bF_buf31), .B(sqrto_75_), .Y(u2__abc_44228_n18675) );
  AND2X2 AND2X2_9128 ( .A(u2__abc_44228_n18665), .B(sqrto_74_), .Y(u2__abc_44228_n18677) );
  AND2X2 AND2X2_9129 ( .A(u2__abc_44228_n18678), .B(u2__abc_44228_n18676), .Y(u2__abc_44228_n18679) );
  AND2X2 AND2X2_913 ( .A(u2__abc_44228_n3816_1), .B(sqrto_103_), .Y(u2__abc_44228_n3817) );
  AND2X2 AND2X2_9130 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n4043), .Y(u2__abc_44228_n18681) );
  AND2X2 AND2X2_9131 ( .A(u2__abc_44228_n18682), .B(u2__abc_44228_n2972_bF_buf4), .Y(u2__abc_44228_n18683) );
  AND2X2 AND2X2_9132 ( .A(u2__abc_44228_n18680), .B(u2__abc_44228_n18683), .Y(u2__abc_44228_n18684) );
  AND2X2 AND2X2_9133 ( .A(u2__abc_44228_n18685), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_root_76__FF_INPUT) );
  AND2X2 AND2X2_9134 ( .A(u2__abc_44228_n3062_bF_buf30), .B(sqrto_76_), .Y(u2__abc_44228_n18687) );
  AND2X2 AND2X2_9135 ( .A(u2__abc_44228_n18677), .B(sqrto_75_), .Y(u2__abc_44228_n18689) );
  AND2X2 AND2X2_9136 ( .A(u2__abc_44228_n18690), .B(u2__abc_44228_n18688), .Y(u2__abc_44228_n18691) );
  AND2X2 AND2X2_9137 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n4030), .Y(u2__abc_44228_n18693) );
  AND2X2 AND2X2_9138 ( .A(u2__abc_44228_n18694), .B(u2__abc_44228_n2972_bF_buf3), .Y(u2__abc_44228_n18695) );
  AND2X2 AND2X2_9139 ( .A(u2__abc_44228_n18692), .B(u2__abc_44228_n18695), .Y(u2__abc_44228_n18696) );
  AND2X2 AND2X2_914 ( .A(u2__abc_44228_n3815), .B(u2__abc_44228_n3818), .Y(u2__abc_44228_n3819) );
  AND2X2 AND2X2_9140 ( .A(u2__abc_44228_n18697), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_root_77__FF_INPUT) );
  AND2X2 AND2X2_9141 ( .A(u2__abc_44228_n3062_bF_buf29), .B(sqrto_77_), .Y(u2__abc_44228_n18699) );
  AND2X2 AND2X2_9142 ( .A(u2__abc_44228_n18689), .B(sqrto_76_), .Y(u2__abc_44228_n18701) );
  AND2X2 AND2X2_9143 ( .A(u2__abc_44228_n18702), .B(u2__abc_44228_n18700), .Y(u2__abc_44228_n18703) );
  AND2X2 AND2X2_9144 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n4023), .Y(u2__abc_44228_n18705) );
  AND2X2 AND2X2_9145 ( .A(u2__abc_44228_n18706), .B(u2__abc_44228_n2972_bF_buf2), .Y(u2__abc_44228_n18707) );
  AND2X2 AND2X2_9146 ( .A(u2__abc_44228_n18704), .B(u2__abc_44228_n18707), .Y(u2__abc_44228_n18708) );
  AND2X2 AND2X2_9147 ( .A(u2__abc_44228_n18709), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_root_78__FF_INPUT) );
  AND2X2 AND2X2_9148 ( .A(u2__abc_44228_n3062_bF_buf28), .B(sqrto_78_), .Y(u2__abc_44228_n18711) );
  AND2X2 AND2X2_9149 ( .A(u2__abc_44228_n18701), .B(sqrto_77_), .Y(u2__abc_44228_n18713) );
  AND2X2 AND2X2_915 ( .A(u2__abc_44228_n3820), .B(u2_remHi_102_), .Y(u2__abc_44228_n3821) );
  AND2X2 AND2X2_9150 ( .A(u2__abc_44228_n18714), .B(u2__abc_44228_n18712), .Y(u2__abc_44228_n18715) );
  AND2X2 AND2X2_9151 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n4006), .Y(u2__abc_44228_n18717) );
  AND2X2 AND2X2_9152 ( .A(u2__abc_44228_n18718), .B(u2__abc_44228_n2972_bF_buf1), .Y(u2__abc_44228_n18719) );
  AND2X2 AND2X2_9153 ( .A(u2__abc_44228_n18716), .B(u2__abc_44228_n18719), .Y(u2__abc_44228_n18720) );
  AND2X2 AND2X2_9154 ( .A(u2__abc_44228_n18721), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_root_79__FF_INPUT) );
  AND2X2 AND2X2_9155 ( .A(u2__abc_44228_n3062_bF_buf27), .B(sqrto_79_), .Y(u2__abc_44228_n18723) );
  AND2X2 AND2X2_9156 ( .A(u2__abc_44228_n18713), .B(sqrto_78_), .Y(u2__abc_44228_n18725) );
  AND2X2 AND2X2_9157 ( .A(u2__abc_44228_n18726), .B(u2__abc_44228_n18724), .Y(u2__abc_44228_n18727) );
  AND2X2 AND2X2_9158 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n4012), .Y(u2__abc_44228_n18729) );
  AND2X2 AND2X2_9159 ( .A(u2__abc_44228_n18730), .B(u2__abc_44228_n2972_bF_buf0), .Y(u2__abc_44228_n18731) );
  AND2X2 AND2X2_916 ( .A(u2__abc_44228_n3822), .B(sqrto_102_), .Y(u2__abc_44228_n3823) );
  AND2X2 AND2X2_9160 ( .A(u2__abc_44228_n18728), .B(u2__abc_44228_n18731), .Y(u2__abc_44228_n18732) );
  AND2X2 AND2X2_9161 ( .A(u2__abc_44228_n18733), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_root_80__FF_INPUT) );
  AND2X2 AND2X2_9162 ( .A(u2__abc_44228_n3062_bF_buf26), .B(sqrto_80_), .Y(u2__abc_44228_n18735) );
  AND2X2 AND2X2_9163 ( .A(u2__abc_44228_n18725), .B(sqrto_79_), .Y(u2__abc_44228_n18737) );
  AND2X2 AND2X2_9164 ( .A(u2__abc_44228_n18738), .B(u2__abc_44228_n18736), .Y(u2__abc_44228_n18739) );
  AND2X2 AND2X2_9165 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n3999), .Y(u2__abc_44228_n18741) );
  AND2X2 AND2X2_9166 ( .A(u2__abc_44228_n18742), .B(u2__abc_44228_n2972_bF_buf107), .Y(u2__abc_44228_n18743) );
  AND2X2 AND2X2_9167 ( .A(u2__abc_44228_n18740), .B(u2__abc_44228_n18743), .Y(u2__abc_44228_n18744) );
  AND2X2 AND2X2_9168 ( .A(u2__abc_44228_n18745), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_root_81__FF_INPUT) );
  AND2X2 AND2X2_9169 ( .A(u2__abc_44228_n3062_bF_buf25), .B(sqrto_81_), .Y(u2__abc_44228_n18747) );
  AND2X2 AND2X2_917 ( .A(u2__abc_44228_n3825_1), .B(u2__abc_44228_n3819), .Y(u2__abc_44228_n3826) );
  AND2X2 AND2X2_9170 ( .A(u2__abc_44228_n18737), .B(sqrto_80_), .Y(u2__abc_44228_n18749) );
  AND2X2 AND2X2_9171 ( .A(u2__abc_44228_n18750), .B(u2__abc_44228_n18748), .Y(u2__abc_44228_n18751) );
  AND2X2 AND2X2_9172 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n3992), .Y(u2__abc_44228_n18753) );
  AND2X2 AND2X2_9173 ( .A(u2__abc_44228_n18754), .B(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n18755) );
  AND2X2 AND2X2_9174 ( .A(u2__abc_44228_n18752), .B(u2__abc_44228_n18755), .Y(u2__abc_44228_n18756) );
  AND2X2 AND2X2_9175 ( .A(u2__abc_44228_n18757), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_root_82__FF_INPUT) );
  AND2X2 AND2X2_9176 ( .A(u2__abc_44228_n3062_bF_buf24), .B(sqrto_82_), .Y(u2__abc_44228_n18759) );
  AND2X2 AND2X2_9177 ( .A(u2__abc_44228_n18749), .B(sqrto_81_), .Y(u2__abc_44228_n18761) );
  AND2X2 AND2X2_9178 ( .A(u2__abc_44228_n18762), .B(u2__abc_44228_n18760), .Y(u2__abc_44228_n18763) );
  AND2X2 AND2X2_9179 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n3977), .Y(u2__abc_44228_n18765) );
  AND2X2 AND2X2_918 ( .A(u2__abc_44228_n3827), .B(u2_remHi_105_), .Y(u2__abc_44228_n3828) );
  AND2X2 AND2X2_9180 ( .A(u2__abc_44228_n18766), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n18767) );
  AND2X2 AND2X2_9181 ( .A(u2__abc_44228_n18764), .B(u2__abc_44228_n18767), .Y(u2__abc_44228_n18768) );
  AND2X2 AND2X2_9182 ( .A(u2__abc_44228_n18769), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_root_83__FF_INPUT) );
  AND2X2 AND2X2_9183 ( .A(u2__abc_44228_n3062_bF_buf23), .B(sqrto_83_), .Y(u2__abc_44228_n18771) );
  AND2X2 AND2X2_9184 ( .A(u2__abc_44228_n18761), .B(sqrto_82_), .Y(u2__abc_44228_n18773) );
  AND2X2 AND2X2_9185 ( .A(u2__abc_44228_n18774), .B(u2__abc_44228_n18772), .Y(u2__abc_44228_n18775) );
  AND2X2 AND2X2_9186 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n3983), .Y(u2__abc_44228_n18777) );
  AND2X2 AND2X2_9187 ( .A(u2__abc_44228_n18778), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n18779) );
  AND2X2 AND2X2_9188 ( .A(u2__abc_44228_n18776), .B(u2__abc_44228_n18779), .Y(u2__abc_44228_n18780) );
  AND2X2 AND2X2_9189 ( .A(u2__abc_44228_n18781), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_root_84__FF_INPUT) );
  AND2X2 AND2X2_919 ( .A(u2__abc_44228_n3830), .B(sqrto_105_), .Y(u2__abc_44228_n3831) );
  AND2X2 AND2X2_9190 ( .A(u2__abc_44228_n3062_bF_buf22), .B(sqrto_84_), .Y(u2__abc_44228_n18783) );
  AND2X2 AND2X2_9191 ( .A(u2__abc_44228_n18773), .B(sqrto_83_), .Y(u2__abc_44228_n18785) );
  AND2X2 AND2X2_9192 ( .A(u2__abc_44228_n18786), .B(u2__abc_44228_n18784), .Y(u2__abc_44228_n18787) );
  AND2X2 AND2X2_9193 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n3970), .Y(u2__abc_44228_n18789) );
  AND2X2 AND2X2_9194 ( .A(u2__abc_44228_n18790), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n18791) );
  AND2X2 AND2X2_9195 ( .A(u2__abc_44228_n18788), .B(u2__abc_44228_n18791), .Y(u2__abc_44228_n18792) );
  AND2X2 AND2X2_9196 ( .A(u2__abc_44228_n18793), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_root_85__FF_INPUT) );
  AND2X2 AND2X2_9197 ( .A(u2__abc_44228_n3062_bF_buf21), .B(sqrto_85_), .Y(u2__abc_44228_n18795) );
  AND2X2 AND2X2_9198 ( .A(u2__abc_44228_n18785), .B(sqrto_84_), .Y(u2__abc_44228_n18797) );
  AND2X2 AND2X2_9199 ( .A(u2__abc_44228_n18798), .B(u2__abc_44228_n18796), .Y(u2__abc_44228_n18799) );
  AND2X2 AND2X2_92 ( .A(_abc_64468_n876), .B(_abc_64468_n875), .Y(_auto_iopadmap_cc_313_execute_65414_127_) );
  AND2X2 AND2X2_920 ( .A(u2__abc_44228_n3829), .B(u2__abc_44228_n3832), .Y(u2__abc_44228_n3833) );
  AND2X2 AND2X2_9200 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n3963), .Y(u2__abc_44228_n18801) );
  AND2X2 AND2X2_9201 ( .A(u2__abc_44228_n18802), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n18803) );
  AND2X2 AND2X2_9202 ( .A(u2__abc_44228_n18800), .B(u2__abc_44228_n18803), .Y(u2__abc_44228_n18804) );
  AND2X2 AND2X2_9203 ( .A(u2__abc_44228_n18805), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_root_86__FF_INPUT) );
  AND2X2 AND2X2_9204 ( .A(u2__abc_44228_n3062_bF_buf20), .B(sqrto_86_), .Y(u2__abc_44228_n18807) );
  AND2X2 AND2X2_9205 ( .A(u2__abc_44228_n18797), .B(sqrto_85_), .Y(u2__abc_44228_n18809) );
  AND2X2 AND2X2_9206 ( .A(u2__abc_44228_n18810), .B(u2__abc_44228_n18808), .Y(u2__abc_44228_n18811) );
  AND2X2 AND2X2_9207 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n3947), .Y(u2__abc_44228_n18813) );
  AND2X2 AND2X2_9208 ( .A(u2__abc_44228_n18814), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n18815) );
  AND2X2 AND2X2_9209 ( .A(u2__abc_44228_n18812), .B(u2__abc_44228_n18815), .Y(u2__abc_44228_n18816) );
  AND2X2 AND2X2_921 ( .A(u2__abc_44228_n3834), .B(u2_remHi_104_), .Y(u2__abc_44228_n3835_1) );
  AND2X2 AND2X2_9210 ( .A(u2__abc_44228_n18817), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_root_87__FF_INPUT) );
  AND2X2 AND2X2_9211 ( .A(u2__abc_44228_n3062_bF_buf19), .B(sqrto_87_), .Y(u2__abc_44228_n18819) );
  AND2X2 AND2X2_9212 ( .A(u2__abc_44228_n18809), .B(sqrto_86_), .Y(u2__abc_44228_n18821) );
  AND2X2 AND2X2_9213 ( .A(u2__abc_44228_n18822), .B(u2__abc_44228_n18820), .Y(u2__abc_44228_n18823) );
  AND2X2 AND2X2_9214 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n3953), .Y(u2__abc_44228_n18825) );
  AND2X2 AND2X2_9215 ( .A(u2__abc_44228_n18826), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n18827) );
  AND2X2 AND2X2_9216 ( .A(u2__abc_44228_n18824), .B(u2__abc_44228_n18827), .Y(u2__abc_44228_n18828) );
  AND2X2 AND2X2_9217 ( .A(u2__abc_44228_n18829), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_root_88__FF_INPUT) );
  AND2X2 AND2X2_9218 ( .A(u2__abc_44228_n3062_bF_buf18), .B(sqrto_88_), .Y(u2__abc_44228_n18831) );
  AND2X2 AND2X2_9219 ( .A(u2__abc_44228_n18821), .B(sqrto_87_), .Y(u2__abc_44228_n18833) );
  AND2X2 AND2X2_922 ( .A(u2__abc_44228_n3836), .B(sqrto_104_), .Y(u2__abc_44228_n3837) );
  AND2X2 AND2X2_9220 ( .A(u2__abc_44228_n18834), .B(u2__abc_44228_n18832), .Y(u2__abc_44228_n18835) );
  AND2X2 AND2X2_9221 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n3940_1), .Y(u2__abc_44228_n18837) );
  AND2X2 AND2X2_9222 ( .A(u2__abc_44228_n18838), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n18839) );
  AND2X2 AND2X2_9223 ( .A(u2__abc_44228_n18836), .B(u2__abc_44228_n18839), .Y(u2__abc_44228_n18840) );
  AND2X2 AND2X2_9224 ( .A(u2__abc_44228_n18841), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_root_89__FF_INPUT) );
  AND2X2 AND2X2_9225 ( .A(u2__abc_44228_n3062_bF_buf17), .B(sqrto_89_), .Y(u2__abc_44228_n18843) );
  AND2X2 AND2X2_9226 ( .A(u2__abc_44228_n18833), .B(sqrto_88_), .Y(u2__abc_44228_n18845) );
  AND2X2 AND2X2_9227 ( .A(u2__abc_44228_n18846), .B(u2__abc_44228_n18844), .Y(u2__abc_44228_n18847) );
  AND2X2 AND2X2_9228 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n3933), .Y(u2__abc_44228_n18849) );
  AND2X2 AND2X2_9229 ( .A(u2__abc_44228_n18850), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n18851) );
  AND2X2 AND2X2_923 ( .A(u2__abc_44228_n3839), .B(u2__abc_44228_n3833), .Y(u2__abc_44228_n3840) );
  AND2X2 AND2X2_9230 ( .A(u2__abc_44228_n18848), .B(u2__abc_44228_n18851), .Y(u2__abc_44228_n18852) );
  AND2X2 AND2X2_9231 ( .A(u2__abc_44228_n18853), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_root_90__FF_INPUT) );
  AND2X2 AND2X2_9232 ( .A(u2__abc_44228_n3062_bF_buf16), .B(sqrto_90_), .Y(u2__abc_44228_n18855) );
  AND2X2 AND2X2_9233 ( .A(u2__abc_44228_n18845), .B(sqrto_89_), .Y(u2__abc_44228_n18857) );
  AND2X2 AND2X2_9234 ( .A(u2__abc_44228_n18858), .B(u2__abc_44228_n18856), .Y(u2__abc_44228_n18859) );
  AND2X2 AND2X2_9235 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n3918), .Y(u2__abc_44228_n18861) );
  AND2X2 AND2X2_9236 ( .A(u2__abc_44228_n18862), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n18863) );
  AND2X2 AND2X2_9237 ( .A(u2__abc_44228_n18860), .B(u2__abc_44228_n18863), .Y(u2__abc_44228_n18864) );
  AND2X2 AND2X2_9238 ( .A(u2__abc_44228_n18865), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_root_91__FF_INPUT) );
  AND2X2 AND2X2_9239 ( .A(u2__abc_44228_n3062_bF_buf15), .B(sqrto_91_), .Y(u2__abc_44228_n18867) );
  AND2X2 AND2X2_924 ( .A(u2__abc_44228_n3826), .B(u2__abc_44228_n3840), .Y(u2__abc_44228_n3841) );
  AND2X2 AND2X2_9240 ( .A(u2__abc_44228_n18857), .B(sqrto_90_), .Y(u2__abc_44228_n18869) );
  AND2X2 AND2X2_9241 ( .A(u2__abc_44228_n18870), .B(u2__abc_44228_n18868), .Y(u2__abc_44228_n18871) );
  AND2X2 AND2X2_9242 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n3924), .Y(u2__abc_44228_n18873) );
  AND2X2 AND2X2_9243 ( .A(u2__abc_44228_n18874), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n18875) );
  AND2X2 AND2X2_9244 ( .A(u2__abc_44228_n18872), .B(u2__abc_44228_n18875), .Y(u2__abc_44228_n18876) );
  AND2X2 AND2X2_9245 ( .A(u2__abc_44228_n18877), .B(u2__abc_44228_n2966_bF_buf91), .Y(u2_root_92__FF_INPUT) );
  AND2X2 AND2X2_9246 ( .A(u2__abc_44228_n3062_bF_buf14), .B(sqrto_92_), .Y(u2__abc_44228_n18879) );
  AND2X2 AND2X2_9247 ( .A(u2__abc_44228_n18869), .B(sqrto_91_), .Y(u2__abc_44228_n18881) );
  AND2X2 AND2X2_9248 ( .A(u2__abc_44228_n18882), .B(u2__abc_44228_n18880), .Y(u2__abc_44228_n18883) );
  AND2X2 AND2X2_9249 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n3911), .Y(u2__abc_44228_n18885) );
  AND2X2 AND2X2_925 ( .A(u2__abc_44228_n3812), .B(u2__abc_44228_n3841), .Y(u2__abc_44228_n3842) );
  AND2X2 AND2X2_9250 ( .A(u2__abc_44228_n18886), .B(u2__abc_44228_n2972_bF_buf95), .Y(u2__abc_44228_n18887) );
  AND2X2 AND2X2_9251 ( .A(u2__abc_44228_n18884), .B(u2__abc_44228_n18887), .Y(u2__abc_44228_n18888) );
  AND2X2 AND2X2_9252 ( .A(u2__abc_44228_n18889), .B(u2__abc_44228_n2966_bF_buf90), .Y(u2_root_93__FF_INPUT) );
  AND2X2 AND2X2_9253 ( .A(u2__abc_44228_n3062_bF_buf13), .B(sqrto_93_), .Y(u2__abc_44228_n18891) );
  AND2X2 AND2X2_9254 ( .A(u2__abc_44228_n18881), .B(sqrto_92_), .Y(u2__abc_44228_n18893) );
  AND2X2 AND2X2_9255 ( .A(u2__abc_44228_n18894), .B(u2__abc_44228_n18892), .Y(u2__abc_44228_n18895) );
  AND2X2 AND2X2_9256 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n3904), .Y(u2__abc_44228_n18897) );
  AND2X2 AND2X2_9257 ( .A(u2__abc_44228_n18898), .B(u2__abc_44228_n2972_bF_buf94), .Y(u2__abc_44228_n18899) );
  AND2X2 AND2X2_9258 ( .A(u2__abc_44228_n18896), .B(u2__abc_44228_n18899), .Y(u2__abc_44228_n18900) );
  AND2X2 AND2X2_9259 ( .A(u2__abc_44228_n18901), .B(u2__abc_44228_n2966_bF_buf89), .Y(u2_root_94__FF_INPUT) );
  AND2X2 AND2X2_926 ( .A(u2__abc_44228_n3843), .B(u2_remHi_101_), .Y(u2__abc_44228_n3844_1) );
  AND2X2 AND2X2_9260 ( .A(u2__abc_44228_n3062_bF_buf12), .B(sqrto_94_), .Y(u2__abc_44228_n18903) );
  AND2X2 AND2X2_9261 ( .A(u2__abc_44228_n18893), .B(sqrto_93_), .Y(u2__abc_44228_n18905) );
  AND2X2 AND2X2_9262 ( .A(u2__abc_44228_n18906), .B(u2__abc_44228_n18904), .Y(u2__abc_44228_n18907) );
  AND2X2 AND2X2_9263 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n3886), .Y(u2__abc_44228_n18909) );
  AND2X2 AND2X2_9264 ( .A(u2__abc_44228_n18910), .B(u2__abc_44228_n2972_bF_buf93), .Y(u2__abc_44228_n18911) );
  AND2X2 AND2X2_9265 ( .A(u2__abc_44228_n18908), .B(u2__abc_44228_n18911), .Y(u2__abc_44228_n18912) );
  AND2X2 AND2X2_9266 ( .A(u2__abc_44228_n18913), .B(u2__abc_44228_n2966_bF_buf88), .Y(u2_root_95__FF_INPUT) );
  AND2X2 AND2X2_9267 ( .A(u2__abc_44228_n3062_bF_buf11), .B(sqrto_95_), .Y(u2__abc_44228_n18915) );
  AND2X2 AND2X2_9268 ( .A(u2__abc_44228_n18905), .B(sqrto_94_), .Y(u2__abc_44228_n18917) );
  AND2X2 AND2X2_9269 ( .A(u2__abc_44228_n18918), .B(u2__abc_44228_n18916), .Y(u2__abc_44228_n18919) );
  AND2X2 AND2X2_927 ( .A(u2__abc_44228_n3846), .B(sqrto_101_), .Y(u2__abc_44228_n3847) );
  AND2X2 AND2X2_9270 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n3892), .Y(u2__abc_44228_n18921) );
  AND2X2 AND2X2_9271 ( .A(u2__abc_44228_n18922), .B(u2__abc_44228_n2972_bF_buf92), .Y(u2__abc_44228_n18923) );
  AND2X2 AND2X2_9272 ( .A(u2__abc_44228_n18920), .B(u2__abc_44228_n18923), .Y(u2__abc_44228_n18924) );
  AND2X2 AND2X2_9273 ( .A(u2__abc_44228_n18925), .B(u2__abc_44228_n2966_bF_buf87), .Y(u2_root_96__FF_INPUT) );
  AND2X2 AND2X2_9274 ( .A(u2__abc_44228_n3062_bF_buf10), .B(sqrto_96_), .Y(u2__abc_44228_n18927) );
  AND2X2 AND2X2_9275 ( .A(u2__abc_44228_n18917), .B(sqrto_95_), .Y(u2__abc_44228_n18929) );
  AND2X2 AND2X2_9276 ( .A(u2__abc_44228_n18930), .B(u2__abc_44228_n18928), .Y(u2__abc_44228_n18931) );
  AND2X2 AND2X2_9277 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n3879), .Y(u2__abc_44228_n18933) );
  AND2X2 AND2X2_9278 ( .A(u2__abc_44228_n18934), .B(u2__abc_44228_n2972_bF_buf91), .Y(u2__abc_44228_n18935) );
  AND2X2 AND2X2_9279 ( .A(u2__abc_44228_n18932), .B(u2__abc_44228_n18935), .Y(u2__abc_44228_n18936) );
  AND2X2 AND2X2_928 ( .A(u2__abc_44228_n3845), .B(u2__abc_44228_n3848), .Y(u2__abc_44228_n3849) );
  AND2X2 AND2X2_9280 ( .A(u2__abc_44228_n18937), .B(u2__abc_44228_n2966_bF_buf86), .Y(u2_root_97__FF_INPUT) );
  AND2X2 AND2X2_9281 ( .A(u2__abc_44228_n3062_bF_buf9), .B(sqrto_97_), .Y(u2__abc_44228_n18939) );
  AND2X2 AND2X2_9282 ( .A(u2__abc_44228_n18929), .B(sqrto_96_), .Y(u2__abc_44228_n18941) );
  AND2X2 AND2X2_9283 ( .A(u2__abc_44228_n18942), .B(u2__abc_44228_n18940), .Y(u2__abc_44228_n18943) );
  AND2X2 AND2X2_9284 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n3872), .Y(u2__abc_44228_n18945) );
  AND2X2 AND2X2_9285 ( .A(u2__abc_44228_n18946), .B(u2__abc_44228_n2972_bF_buf90), .Y(u2__abc_44228_n18947) );
  AND2X2 AND2X2_9286 ( .A(u2__abc_44228_n18944), .B(u2__abc_44228_n18947), .Y(u2__abc_44228_n18948) );
  AND2X2 AND2X2_9287 ( .A(u2__abc_44228_n18949), .B(u2__abc_44228_n2966_bF_buf85), .Y(u2_root_98__FF_INPUT) );
  AND2X2 AND2X2_9288 ( .A(u2__abc_44228_n3062_bF_buf8), .B(sqrto_98_), .Y(u2__abc_44228_n18951) );
  AND2X2 AND2X2_9289 ( .A(u2__abc_44228_n18941), .B(sqrto_97_), .Y(u2__abc_44228_n18953) );
  AND2X2 AND2X2_929 ( .A(u2__abc_44228_n3850), .B(u2_remHi_100_), .Y(u2__abc_44228_n3851) );
  AND2X2 AND2X2_9290 ( .A(u2__abc_44228_n18954), .B(u2__abc_44228_n18952), .Y(u2__abc_44228_n18955) );
  AND2X2 AND2X2_9291 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n3857), .Y(u2__abc_44228_n18957) );
  AND2X2 AND2X2_9292 ( .A(u2__abc_44228_n18958), .B(u2__abc_44228_n2972_bF_buf89), .Y(u2__abc_44228_n18959) );
  AND2X2 AND2X2_9293 ( .A(u2__abc_44228_n18956), .B(u2__abc_44228_n18959), .Y(u2__abc_44228_n18960) );
  AND2X2 AND2X2_9294 ( .A(u2__abc_44228_n18961), .B(u2__abc_44228_n2966_bF_buf84), .Y(u2_root_99__FF_INPUT) );
  AND2X2 AND2X2_9295 ( .A(u2__abc_44228_n3062_bF_buf7), .B(sqrto_99_), .Y(u2__abc_44228_n18963) );
  AND2X2 AND2X2_9296 ( .A(u2__abc_44228_n18953), .B(sqrto_98_), .Y(u2__abc_44228_n18965) );
  AND2X2 AND2X2_9297 ( .A(u2__abc_44228_n18966), .B(u2__abc_44228_n18964), .Y(u2__abc_44228_n18967) );
  AND2X2 AND2X2_9298 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n3863), .Y(u2__abc_44228_n18969) );
  AND2X2 AND2X2_9299 ( .A(u2__abc_44228_n18970), .B(u2__abc_44228_n2972_bF_buf88), .Y(u2__abc_44228_n18971) );
  AND2X2 AND2X2_93 ( .A(_abc_64468_n879), .B(_abc_64468_n878), .Y(_auto_iopadmap_cc_313_execute_65414_128_) );
  AND2X2 AND2X2_930 ( .A(u2__abc_44228_n3852), .B(sqrto_100_), .Y(u2__abc_44228_n3853) );
  AND2X2 AND2X2_9300 ( .A(u2__abc_44228_n18968), .B(u2__abc_44228_n18971), .Y(u2__abc_44228_n18972) );
  AND2X2 AND2X2_9301 ( .A(u2__abc_44228_n18973), .B(u2__abc_44228_n2966_bF_buf83), .Y(u2_root_100__FF_INPUT) );
  AND2X2 AND2X2_9302 ( .A(u2__abc_44228_n3062_bF_buf6), .B(sqrto_100_), .Y(u2__abc_44228_n18975) );
  AND2X2 AND2X2_9303 ( .A(u2__abc_44228_n18965), .B(sqrto_99_), .Y(u2__abc_44228_n18977) );
  AND2X2 AND2X2_9304 ( .A(u2__abc_44228_n18978), .B(u2__abc_44228_n18976), .Y(u2__abc_44228_n18979) );
  AND2X2 AND2X2_9305 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n3850), .Y(u2__abc_44228_n18981) );
  AND2X2 AND2X2_9306 ( .A(u2__abc_44228_n18982), .B(u2__abc_44228_n2972_bF_buf87), .Y(u2__abc_44228_n18983) );
  AND2X2 AND2X2_9307 ( .A(u2__abc_44228_n18980), .B(u2__abc_44228_n18983), .Y(u2__abc_44228_n18984) );
  AND2X2 AND2X2_9308 ( .A(u2__abc_44228_n18985), .B(u2__abc_44228_n2966_bF_buf82), .Y(u2_root_101__FF_INPUT) );
  AND2X2 AND2X2_9309 ( .A(u2__abc_44228_n3062_bF_buf5), .B(sqrto_101_), .Y(u2__abc_44228_n18987) );
  AND2X2 AND2X2_931 ( .A(u2__abc_44228_n3855), .B(u2__abc_44228_n3849), .Y(u2__abc_44228_n3856) );
  AND2X2 AND2X2_9310 ( .A(u2__abc_44228_n18977), .B(sqrto_100_), .Y(u2__abc_44228_n18989) );
  AND2X2 AND2X2_9311 ( .A(u2__abc_44228_n18990), .B(u2__abc_44228_n18988), .Y(u2__abc_44228_n18991) );
  AND2X2 AND2X2_9312 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n3843), .Y(u2__abc_44228_n18993) );
  AND2X2 AND2X2_9313 ( .A(u2__abc_44228_n18994), .B(u2__abc_44228_n2972_bF_buf86), .Y(u2__abc_44228_n18995) );
  AND2X2 AND2X2_9314 ( .A(u2__abc_44228_n18992), .B(u2__abc_44228_n18995), .Y(u2__abc_44228_n18996) );
  AND2X2 AND2X2_9315 ( .A(u2__abc_44228_n18997), .B(u2__abc_44228_n2966_bF_buf81), .Y(u2_root_102__FF_INPUT) );
  AND2X2 AND2X2_9316 ( .A(u2__abc_44228_n3062_bF_buf4), .B(sqrto_102_), .Y(u2__abc_44228_n18999) );
  AND2X2 AND2X2_9317 ( .A(u2__abc_44228_n18989), .B(sqrto_101_), .Y(u2__abc_44228_n19001) );
  AND2X2 AND2X2_9318 ( .A(u2__abc_44228_n19002), .B(u2__abc_44228_n19000), .Y(u2__abc_44228_n19003) );
  AND2X2 AND2X2_9319 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n3820), .Y(u2__abc_44228_n19005) );
  AND2X2 AND2X2_932 ( .A(u2__abc_44228_n3857), .B(u2_remHi_98_), .Y(u2__abc_44228_n3858) );
  AND2X2 AND2X2_9320 ( .A(u2__abc_44228_n19006), .B(u2__abc_44228_n2972_bF_buf85), .Y(u2__abc_44228_n19007) );
  AND2X2 AND2X2_9321 ( .A(u2__abc_44228_n19004), .B(u2__abc_44228_n19007), .Y(u2__abc_44228_n19008) );
  AND2X2 AND2X2_9322 ( .A(u2__abc_44228_n19009), .B(u2__abc_44228_n2966_bF_buf80), .Y(u2_root_103__FF_INPUT) );
  AND2X2 AND2X2_9323 ( .A(u2__abc_44228_n3062_bF_buf3), .B(sqrto_103_), .Y(u2__abc_44228_n19011) );
  AND2X2 AND2X2_9324 ( .A(u2__abc_44228_n19001), .B(sqrto_102_), .Y(u2__abc_44228_n19013) );
  AND2X2 AND2X2_9325 ( .A(u2__abc_44228_n19014), .B(u2__abc_44228_n19012), .Y(u2__abc_44228_n19015) );
  AND2X2 AND2X2_9326 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n3813), .Y(u2__abc_44228_n19017) );
  AND2X2 AND2X2_9327 ( .A(u2__abc_44228_n19018), .B(u2__abc_44228_n2972_bF_buf84), .Y(u2__abc_44228_n19019) );
  AND2X2 AND2X2_9328 ( .A(u2__abc_44228_n19016), .B(u2__abc_44228_n19019), .Y(u2__abc_44228_n19020) );
  AND2X2 AND2X2_9329 ( .A(u2__abc_44228_n19021), .B(u2__abc_44228_n2966_bF_buf79), .Y(u2_root_104__FF_INPUT) );
  AND2X2 AND2X2_933 ( .A(u2__abc_44228_n3859), .B(sqrto_98_), .Y(u2__abc_44228_n3860) );
  AND2X2 AND2X2_9330 ( .A(u2__abc_44228_n3062_bF_buf2), .B(sqrto_104_), .Y(u2__abc_44228_n19023) );
  AND2X2 AND2X2_9331 ( .A(u2__abc_44228_n19013), .B(sqrto_103_), .Y(u2__abc_44228_n19025) );
  AND2X2 AND2X2_9332 ( .A(u2__abc_44228_n19026), .B(u2__abc_44228_n19024), .Y(u2__abc_44228_n19027) );
  AND2X2 AND2X2_9333 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n3834), .Y(u2__abc_44228_n19029) );
  AND2X2 AND2X2_9334 ( .A(u2__abc_44228_n19030), .B(u2__abc_44228_n2972_bF_buf83), .Y(u2__abc_44228_n19031) );
  AND2X2 AND2X2_9335 ( .A(u2__abc_44228_n19028), .B(u2__abc_44228_n19031), .Y(u2__abc_44228_n19032) );
  AND2X2 AND2X2_9336 ( .A(u2__abc_44228_n19033), .B(u2__abc_44228_n2966_bF_buf78), .Y(u2_root_105__FF_INPUT) );
  AND2X2 AND2X2_9337 ( .A(u2__abc_44228_n3062_bF_buf1), .B(sqrto_105_), .Y(u2__abc_44228_n19035) );
  AND2X2 AND2X2_9338 ( .A(u2__abc_44228_n19025), .B(sqrto_104_), .Y(u2__abc_44228_n19037) );
  AND2X2 AND2X2_9339 ( .A(u2__abc_44228_n19038), .B(u2__abc_44228_n19036), .Y(u2__abc_44228_n19039) );
  AND2X2 AND2X2_934 ( .A(u2__abc_44228_n3863), .B(u2_remHi_99_), .Y(u2__abc_44228_n3864_1) );
  AND2X2 AND2X2_9340 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n3827), .Y(u2__abc_44228_n19041) );
  AND2X2 AND2X2_9341 ( .A(u2__abc_44228_n19042), .B(u2__abc_44228_n2972_bF_buf82), .Y(u2__abc_44228_n19043) );
  AND2X2 AND2X2_9342 ( .A(u2__abc_44228_n19040), .B(u2__abc_44228_n19043), .Y(u2__abc_44228_n19044) );
  AND2X2 AND2X2_9343 ( .A(u2__abc_44228_n19045), .B(u2__abc_44228_n2966_bF_buf77), .Y(u2_root_106__FF_INPUT) );
  AND2X2 AND2X2_9344 ( .A(u2__abc_44228_n3062_bF_buf0), .B(sqrto_106_), .Y(u2__abc_44228_n19047) );
  AND2X2 AND2X2_9345 ( .A(u2__abc_44228_n19037), .B(sqrto_105_), .Y(u2__abc_44228_n19049) );
  AND2X2 AND2X2_9346 ( .A(u2__abc_44228_n19050), .B(u2__abc_44228_n19048), .Y(u2__abc_44228_n19051) );
  AND2X2 AND2X2_9347 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n3798_1), .Y(u2__abc_44228_n19053) );
  AND2X2 AND2X2_9348 ( .A(u2__abc_44228_n19054), .B(u2__abc_44228_n2972_bF_buf81), .Y(u2__abc_44228_n19055) );
  AND2X2 AND2X2_9349 ( .A(u2__abc_44228_n19052), .B(u2__abc_44228_n19055), .Y(u2__abc_44228_n19056) );
  AND2X2 AND2X2_935 ( .A(u2__abc_44228_n3866), .B(sqrto_99_), .Y(u2__abc_44228_n3867) );
  AND2X2 AND2X2_9350 ( .A(u2__abc_44228_n19057), .B(u2__abc_44228_n2966_bF_buf76), .Y(u2_root_107__FF_INPUT) );
  AND2X2 AND2X2_9351 ( .A(u2__abc_44228_n3062_bF_buf92), .B(sqrto_107_), .Y(u2__abc_44228_n19059) );
  AND2X2 AND2X2_9352 ( .A(u2__abc_44228_n19049), .B(sqrto_106_), .Y(u2__abc_44228_n19061) );
  AND2X2 AND2X2_9353 ( .A(u2__abc_44228_n19062), .B(u2__abc_44228_n19060), .Y(u2__abc_44228_n19063) );
  AND2X2 AND2X2_9354 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n3804), .Y(u2__abc_44228_n19065) );
  AND2X2 AND2X2_9355 ( .A(u2__abc_44228_n19066), .B(u2__abc_44228_n2972_bF_buf80), .Y(u2__abc_44228_n19067) );
  AND2X2 AND2X2_9356 ( .A(u2__abc_44228_n19064), .B(u2__abc_44228_n19067), .Y(u2__abc_44228_n19068) );
  AND2X2 AND2X2_9357 ( .A(u2__abc_44228_n19069), .B(u2__abc_44228_n2966_bF_buf75), .Y(u2_root_108__FF_INPUT) );
  AND2X2 AND2X2_9358 ( .A(u2__abc_44228_n3062_bF_buf91), .B(sqrto_108_), .Y(u2__abc_44228_n19071) );
  AND2X2 AND2X2_9359 ( .A(u2__abc_44228_n19061), .B(sqrto_107_), .Y(u2__abc_44228_n19073) );
  AND2X2 AND2X2_936 ( .A(u2__abc_44228_n3865), .B(u2__abc_44228_n3868), .Y(u2__abc_44228_n3869) );
  AND2X2 AND2X2_9360 ( .A(u2__abc_44228_n19074), .B(u2__abc_44228_n19072), .Y(u2__abc_44228_n19075) );
  AND2X2 AND2X2_9361 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n3791), .Y(u2__abc_44228_n19077) );
  AND2X2 AND2X2_9362 ( .A(u2__abc_44228_n19078), .B(u2__abc_44228_n2972_bF_buf79), .Y(u2__abc_44228_n19079) );
  AND2X2 AND2X2_9363 ( .A(u2__abc_44228_n19076), .B(u2__abc_44228_n19079), .Y(u2__abc_44228_n19080) );
  AND2X2 AND2X2_9364 ( .A(u2__abc_44228_n19081), .B(u2__abc_44228_n2966_bF_buf74), .Y(u2_root_109__FF_INPUT) );
  AND2X2 AND2X2_9365 ( .A(u2__abc_44228_n3062_bF_buf90), .B(sqrto_109_), .Y(u2__abc_44228_n19083) );
  AND2X2 AND2X2_9366 ( .A(u2__abc_44228_n19073), .B(sqrto_108_), .Y(u2__abc_44228_n19085) );
  AND2X2 AND2X2_9367 ( .A(u2__abc_44228_n19086), .B(u2__abc_44228_n19084), .Y(u2__abc_44228_n19087) );
  AND2X2 AND2X2_9368 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n3784), .Y(u2__abc_44228_n19089) );
  AND2X2 AND2X2_9369 ( .A(u2__abc_44228_n19090), .B(u2__abc_44228_n2972_bF_buf78), .Y(u2__abc_44228_n19091) );
  AND2X2 AND2X2_937 ( .A(u2__abc_44228_n3862), .B(u2__abc_44228_n3869), .Y(u2__abc_44228_n3870) );
  AND2X2 AND2X2_9370 ( .A(u2__abc_44228_n19088), .B(u2__abc_44228_n19091), .Y(u2__abc_44228_n19092) );
  AND2X2 AND2X2_9371 ( .A(u2__abc_44228_n19093), .B(u2__abc_44228_n2966_bF_buf73), .Y(u2_root_110__FF_INPUT) );
  AND2X2 AND2X2_9372 ( .A(u2__abc_44228_n3062_bF_buf89), .B(sqrto_110_), .Y(u2__abc_44228_n19095) );
  AND2X2 AND2X2_9373 ( .A(u2__abc_44228_n19085), .B(sqrto_109_), .Y(u2__abc_44228_n19097) );
  AND2X2 AND2X2_9374 ( .A(u2__abc_44228_n19098), .B(u2__abc_44228_n19096), .Y(u2__abc_44228_n19099) );
  AND2X2 AND2X2_9375 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n3767), .Y(u2__abc_44228_n19101) );
  AND2X2 AND2X2_9376 ( .A(u2__abc_44228_n19102), .B(u2__abc_44228_n2972_bF_buf77), .Y(u2__abc_44228_n19103) );
  AND2X2 AND2X2_9377 ( .A(u2__abc_44228_n19100), .B(u2__abc_44228_n19103), .Y(u2__abc_44228_n19104) );
  AND2X2 AND2X2_9378 ( .A(u2__abc_44228_n19105), .B(u2__abc_44228_n2966_bF_buf72), .Y(u2_root_111__FF_INPUT) );
  AND2X2 AND2X2_9379 ( .A(u2__abc_44228_n3062_bF_buf88), .B(sqrto_111_), .Y(u2__abc_44228_n19107) );
  AND2X2 AND2X2_938 ( .A(u2__abc_44228_n3856), .B(u2__abc_44228_n3870), .Y(u2__abc_44228_n3871) );
  AND2X2 AND2X2_9380 ( .A(u2__abc_44228_n19097), .B(sqrto_110_), .Y(u2__abc_44228_n19109) );
  AND2X2 AND2X2_9381 ( .A(u2__abc_44228_n19110), .B(u2__abc_44228_n19108), .Y(u2__abc_44228_n19111) );
  AND2X2 AND2X2_9382 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n3773), .Y(u2__abc_44228_n19113) );
  AND2X2 AND2X2_9383 ( .A(u2__abc_44228_n19114), .B(u2__abc_44228_n2972_bF_buf76), .Y(u2__abc_44228_n19115) );
  AND2X2 AND2X2_9384 ( .A(u2__abc_44228_n19112), .B(u2__abc_44228_n19115), .Y(u2__abc_44228_n19116) );
  AND2X2 AND2X2_9385 ( .A(u2__abc_44228_n19117), .B(u2__abc_44228_n2966_bF_buf71), .Y(u2_root_112__FF_INPUT) );
  AND2X2 AND2X2_9386 ( .A(u2__abc_44228_n3062_bF_buf87), .B(sqrto_112_), .Y(u2__abc_44228_n19119) );
  AND2X2 AND2X2_9387 ( .A(u2__abc_44228_n19109), .B(sqrto_111_), .Y(u2__abc_44228_n19121) );
  AND2X2 AND2X2_9388 ( .A(u2__abc_44228_n19122), .B(u2__abc_44228_n19120), .Y(u2__abc_44228_n19123) );
  AND2X2 AND2X2_9389 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n3760), .Y(u2__abc_44228_n19125) );
  AND2X2 AND2X2_939 ( .A(u2__abc_44228_n3872), .B(u2_remHi_97_), .Y(u2__abc_44228_n3873_1) );
  AND2X2 AND2X2_9390 ( .A(u2__abc_44228_n19126), .B(u2__abc_44228_n2972_bF_buf75), .Y(u2__abc_44228_n19127) );
  AND2X2 AND2X2_9391 ( .A(u2__abc_44228_n19124), .B(u2__abc_44228_n19127), .Y(u2__abc_44228_n19128) );
  AND2X2 AND2X2_9392 ( .A(u2__abc_44228_n19129), .B(u2__abc_44228_n2966_bF_buf70), .Y(u2_root_113__FF_INPUT) );
  AND2X2 AND2X2_9393 ( .A(u2__abc_44228_n3062_bF_buf86), .B(sqrto_113_), .Y(u2__abc_44228_n19131) );
  AND2X2 AND2X2_9394 ( .A(u2__abc_44228_n19121), .B(sqrto_112_), .Y(u2__abc_44228_n19133) );
  AND2X2 AND2X2_9395 ( .A(u2__abc_44228_n19134), .B(u2__abc_44228_n19132), .Y(u2__abc_44228_n19135) );
  AND2X2 AND2X2_9396 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n3753), .Y(u2__abc_44228_n19137) );
  AND2X2 AND2X2_9397 ( .A(u2__abc_44228_n19138), .B(u2__abc_44228_n2972_bF_buf74), .Y(u2__abc_44228_n19139) );
  AND2X2 AND2X2_9398 ( .A(u2__abc_44228_n19136), .B(u2__abc_44228_n19139), .Y(u2__abc_44228_n19140) );
  AND2X2 AND2X2_9399 ( .A(u2__abc_44228_n19141), .B(u2__abc_44228_n2966_bF_buf69), .Y(u2_root_114__FF_INPUT) );
  AND2X2 AND2X2_94 ( .A(_abc_64468_n882), .B(_abc_64468_n881), .Y(_auto_iopadmap_cc_313_execute_65414_129_) );
  AND2X2 AND2X2_940 ( .A(u2__abc_44228_n3875), .B(sqrto_97_), .Y(u2__abc_44228_n3876) );
  AND2X2 AND2X2_9400 ( .A(u2__abc_44228_n3062_bF_buf85), .B(sqrto_114_), .Y(u2__abc_44228_n19143) );
  AND2X2 AND2X2_9401 ( .A(u2__abc_44228_n19133), .B(sqrto_113_), .Y(u2__abc_44228_n19145) );
  AND2X2 AND2X2_9402 ( .A(u2__abc_44228_n19146), .B(u2__abc_44228_n19144), .Y(u2__abc_44228_n19147) );
  AND2X2 AND2X2_9403 ( .A(u2__abc_44228_n2983_bF_buf104), .B(u2__abc_44228_n3745), .Y(u2__abc_44228_n19149) );
  AND2X2 AND2X2_9404 ( .A(u2__abc_44228_n19150), .B(u2__abc_44228_n2972_bF_buf73), .Y(u2__abc_44228_n19151) );
  AND2X2 AND2X2_9405 ( .A(u2__abc_44228_n19148), .B(u2__abc_44228_n19151), .Y(u2__abc_44228_n19152) );
  AND2X2 AND2X2_9406 ( .A(u2__abc_44228_n19153), .B(u2__abc_44228_n2966_bF_buf68), .Y(u2_root_115__FF_INPUT) );
  AND2X2 AND2X2_9407 ( .A(u2__abc_44228_n3062_bF_buf84), .B(sqrto_115_), .Y(u2__abc_44228_n19155) );
  AND2X2 AND2X2_9408 ( .A(u2__abc_44228_n19145), .B(sqrto_114_), .Y(u2__abc_44228_n19157) );
  AND2X2 AND2X2_9409 ( .A(u2__abc_44228_n19158), .B(u2__abc_44228_n19156), .Y(u2__abc_44228_n19159) );
  AND2X2 AND2X2_941 ( .A(u2__abc_44228_n3874), .B(u2__abc_44228_n3877), .Y(u2__abc_44228_n3878) );
  AND2X2 AND2X2_9410 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n3738), .Y(u2__abc_44228_n19161) );
  AND2X2 AND2X2_9411 ( .A(u2__abc_44228_n19162), .B(u2__abc_44228_n2972_bF_buf72), .Y(u2__abc_44228_n19163) );
  AND2X2 AND2X2_9412 ( .A(u2__abc_44228_n19160), .B(u2__abc_44228_n19163), .Y(u2__abc_44228_n19164) );
  AND2X2 AND2X2_9413 ( .A(u2__abc_44228_n19165), .B(u2__abc_44228_n2966_bF_buf67), .Y(u2_root_116__FF_INPUT) );
  AND2X2 AND2X2_9414 ( .A(u2__abc_44228_n3062_bF_buf83), .B(sqrto_116_), .Y(u2__abc_44228_n19167) );
  AND2X2 AND2X2_9415 ( .A(u2__abc_44228_n19157), .B(sqrto_115_), .Y(u2__abc_44228_n19169) );
  AND2X2 AND2X2_9416 ( .A(u2__abc_44228_n19170), .B(u2__abc_44228_n19168), .Y(u2__abc_44228_n19171) );
  AND2X2 AND2X2_9417 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n3731), .Y(u2__abc_44228_n19173) );
  AND2X2 AND2X2_9418 ( .A(u2__abc_44228_n19174), .B(u2__abc_44228_n2972_bF_buf71), .Y(u2__abc_44228_n19175) );
  AND2X2 AND2X2_9419 ( .A(u2__abc_44228_n19172), .B(u2__abc_44228_n19175), .Y(u2__abc_44228_n19176) );
  AND2X2 AND2X2_942 ( .A(u2__abc_44228_n3879), .B(u2_remHi_96_), .Y(u2__abc_44228_n3880) );
  AND2X2 AND2X2_9420 ( .A(u2__abc_44228_n19177), .B(u2__abc_44228_n2966_bF_buf66), .Y(u2_root_117__FF_INPUT) );
  AND2X2 AND2X2_9421 ( .A(u2__abc_44228_n3062_bF_buf82), .B(sqrto_117_), .Y(u2__abc_44228_n19179) );
  AND2X2 AND2X2_9422 ( .A(u2__abc_44228_n19169), .B(sqrto_116_), .Y(u2__abc_44228_n19181) );
  AND2X2 AND2X2_9423 ( .A(u2__abc_44228_n19182), .B(u2__abc_44228_n19180), .Y(u2__abc_44228_n19183) );
  AND2X2 AND2X2_9424 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n3724), .Y(u2__abc_44228_n19185) );
  AND2X2 AND2X2_9425 ( .A(u2__abc_44228_n19186), .B(u2__abc_44228_n2972_bF_buf70), .Y(u2__abc_44228_n19187) );
  AND2X2 AND2X2_9426 ( .A(u2__abc_44228_n19184), .B(u2__abc_44228_n19187), .Y(u2__abc_44228_n19188) );
  AND2X2 AND2X2_9427 ( .A(u2__abc_44228_n19189), .B(u2__abc_44228_n2966_bF_buf65), .Y(u2_root_118__FF_INPUT) );
  AND2X2 AND2X2_9428 ( .A(u2__abc_44228_n3062_bF_buf81), .B(sqrto_118_), .Y(u2__abc_44228_n19191) );
  AND2X2 AND2X2_9429 ( .A(u2__abc_44228_n19181), .B(sqrto_117_), .Y(u2__abc_44228_n19193) );
  AND2X2 AND2X2_943 ( .A(u2__abc_44228_n3881), .B(sqrto_96_), .Y(u2__abc_44228_n3882_1) );
  AND2X2 AND2X2_9430 ( .A(u2__abc_44228_n19194), .B(u2__abc_44228_n19192), .Y(u2__abc_44228_n19195) );
  AND2X2 AND2X2_9431 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n3701), .Y(u2__abc_44228_n19197) );
  AND2X2 AND2X2_9432 ( .A(u2__abc_44228_n19198), .B(u2__abc_44228_n2972_bF_buf69), .Y(u2__abc_44228_n19199) );
  AND2X2 AND2X2_9433 ( .A(u2__abc_44228_n19196), .B(u2__abc_44228_n19199), .Y(u2__abc_44228_n19200) );
  AND2X2 AND2X2_9434 ( .A(u2__abc_44228_n19201), .B(u2__abc_44228_n2966_bF_buf64), .Y(u2_root_119__FF_INPUT) );
  AND2X2 AND2X2_9435 ( .A(u2__abc_44228_n3062_bF_buf80), .B(sqrto_119_), .Y(u2__abc_44228_n19203) );
  AND2X2 AND2X2_9436 ( .A(u2__abc_44228_n19193), .B(sqrto_118_), .Y(u2__abc_44228_n19205) );
  AND2X2 AND2X2_9437 ( .A(u2__abc_44228_n19206), .B(u2__abc_44228_n19204), .Y(u2__abc_44228_n19207) );
  AND2X2 AND2X2_9438 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n3694_1), .Y(u2__abc_44228_n19209) );
  AND2X2 AND2X2_9439 ( .A(u2__abc_44228_n19210), .B(u2__abc_44228_n2972_bF_buf68), .Y(u2__abc_44228_n19211) );
  AND2X2 AND2X2_944 ( .A(u2__abc_44228_n3884), .B(u2__abc_44228_n3878), .Y(u2__abc_44228_n3885) );
  AND2X2 AND2X2_9440 ( .A(u2__abc_44228_n19208), .B(u2__abc_44228_n19211), .Y(u2__abc_44228_n19212) );
  AND2X2 AND2X2_9441 ( .A(u2__abc_44228_n19213), .B(u2__abc_44228_n2966_bF_buf63), .Y(u2_root_120__FF_INPUT) );
  AND2X2 AND2X2_9442 ( .A(u2__abc_44228_n3062_bF_buf79), .B(sqrto_120_), .Y(u2__abc_44228_n19215) );
  AND2X2 AND2X2_9443 ( .A(u2__abc_44228_n19205), .B(sqrto_119_), .Y(u2__abc_44228_n19217) );
  AND2X2 AND2X2_9444 ( .A(u2__abc_44228_n19218), .B(u2__abc_44228_n19216), .Y(u2__abc_44228_n19219) );
  AND2X2 AND2X2_9445 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n3715), .Y(u2__abc_44228_n19221) );
  AND2X2 AND2X2_9446 ( .A(u2__abc_44228_n19222), .B(u2__abc_44228_n2972_bF_buf67), .Y(u2__abc_44228_n19223) );
  AND2X2 AND2X2_9447 ( .A(u2__abc_44228_n19220), .B(u2__abc_44228_n19223), .Y(u2__abc_44228_n19224) );
  AND2X2 AND2X2_9448 ( .A(u2__abc_44228_n19225), .B(u2__abc_44228_n2966_bF_buf62), .Y(u2_root_121__FF_INPUT) );
  AND2X2 AND2X2_9449 ( .A(u2__abc_44228_n3062_bF_buf78), .B(sqrto_121_), .Y(u2__abc_44228_n19227) );
  AND2X2 AND2X2_945 ( .A(u2__abc_44228_n3886), .B(u2_remHi_94_), .Y(u2__abc_44228_n3887) );
  AND2X2 AND2X2_9450 ( .A(u2__abc_44228_n19217), .B(sqrto_120_), .Y(u2__abc_44228_n19229) );
  AND2X2 AND2X2_9451 ( .A(u2__abc_44228_n19230), .B(u2__abc_44228_n19228), .Y(u2__abc_44228_n19231) );
  AND2X2 AND2X2_9452 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n3708), .Y(u2__abc_44228_n19233) );
  AND2X2 AND2X2_9453 ( .A(u2__abc_44228_n19234), .B(u2__abc_44228_n2972_bF_buf66), .Y(u2__abc_44228_n19235) );
  AND2X2 AND2X2_9454 ( .A(u2__abc_44228_n19232), .B(u2__abc_44228_n19235), .Y(u2__abc_44228_n19236) );
  AND2X2 AND2X2_9455 ( .A(u2__abc_44228_n19237), .B(u2__abc_44228_n2966_bF_buf61), .Y(u2_root_122__FF_INPUT) );
  AND2X2 AND2X2_9456 ( .A(u2__abc_44228_n3062_bF_buf77), .B(sqrto_122_), .Y(u2__abc_44228_n19239) );
  AND2X2 AND2X2_9457 ( .A(u2__abc_44228_n19229), .B(sqrto_121_), .Y(u2__abc_44228_n19241) );
  AND2X2 AND2X2_9458 ( .A(u2__abc_44228_n19242), .B(u2__abc_44228_n19240), .Y(u2__abc_44228_n19243) );
  AND2X2 AND2X2_9459 ( .A(u2__abc_44228_n2983_bF_buf88), .B(u2__abc_44228_n3679), .Y(u2__abc_44228_n19245) );
  AND2X2 AND2X2_946 ( .A(u2__abc_44228_n3888), .B(sqrto_94_), .Y(u2__abc_44228_n3889) );
  AND2X2 AND2X2_9460 ( .A(u2__abc_44228_n19246), .B(u2__abc_44228_n2972_bF_buf65), .Y(u2__abc_44228_n19247) );
  AND2X2 AND2X2_9461 ( .A(u2__abc_44228_n19244), .B(u2__abc_44228_n19247), .Y(u2__abc_44228_n19248) );
  AND2X2 AND2X2_9462 ( .A(u2__abc_44228_n19249), .B(u2__abc_44228_n2966_bF_buf60), .Y(u2_root_123__FF_INPUT) );
  AND2X2 AND2X2_9463 ( .A(u2__abc_44228_n3062_bF_buf76), .B(sqrto_123_), .Y(u2__abc_44228_n19251) );
  AND2X2 AND2X2_9464 ( .A(u2__abc_44228_n19241), .B(sqrto_122_), .Y(u2__abc_44228_n19253) );
  AND2X2 AND2X2_9465 ( .A(u2__abc_44228_n19254), .B(u2__abc_44228_n19252), .Y(u2__abc_44228_n19255) );
  AND2X2 AND2X2_9466 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n3685_1), .Y(u2__abc_44228_n19257) );
  AND2X2 AND2X2_9467 ( .A(u2__abc_44228_n19258), .B(u2__abc_44228_n2972_bF_buf64), .Y(u2__abc_44228_n19259) );
  AND2X2 AND2X2_9468 ( .A(u2__abc_44228_n19256), .B(u2__abc_44228_n19259), .Y(u2__abc_44228_n19260) );
  AND2X2 AND2X2_9469 ( .A(u2__abc_44228_n19261), .B(u2__abc_44228_n2966_bF_buf59), .Y(u2_root_124__FF_INPUT) );
  AND2X2 AND2X2_947 ( .A(u2__abc_44228_n3892), .B(u2_remHi_95_), .Y(u2__abc_44228_n3893_1) );
  AND2X2 AND2X2_9470 ( .A(u2__abc_44228_n3062_bF_buf75), .B(sqrto_124_), .Y(u2__abc_44228_n19263) );
  AND2X2 AND2X2_9471 ( .A(u2__abc_44228_n19253), .B(sqrto_123_), .Y(u2__abc_44228_n19265) );
  AND2X2 AND2X2_9472 ( .A(u2__abc_44228_n19266), .B(u2__abc_44228_n19264), .Y(u2__abc_44228_n19267) );
  AND2X2 AND2X2_9473 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n3672), .Y(u2__abc_44228_n19269) );
  AND2X2 AND2X2_9474 ( .A(u2__abc_44228_n19270), .B(u2__abc_44228_n2972_bF_buf63), .Y(u2__abc_44228_n19271) );
  AND2X2 AND2X2_9475 ( .A(u2__abc_44228_n19268), .B(u2__abc_44228_n19271), .Y(u2__abc_44228_n19272) );
  AND2X2 AND2X2_9476 ( .A(u2__abc_44228_n19273), .B(u2__abc_44228_n2966_bF_buf58), .Y(u2_root_125__FF_INPUT) );
  AND2X2 AND2X2_9477 ( .A(u2__abc_44228_n3062_bF_buf74), .B(sqrto_125_), .Y(u2__abc_44228_n19275) );
  AND2X2 AND2X2_9478 ( .A(u2__abc_44228_n19265), .B(sqrto_124_), .Y(u2__abc_44228_n19277) );
  AND2X2 AND2X2_9479 ( .A(u2__abc_44228_n19278), .B(u2__abc_44228_n19276), .Y(u2__abc_44228_n19279) );
  AND2X2 AND2X2_948 ( .A(u2__abc_44228_n3895), .B(sqrto_95_), .Y(u2__abc_44228_n3896) );
  AND2X2 AND2X2_9480 ( .A(u2__abc_44228_n2983_bF_buf82), .B(u2__abc_44228_n3665), .Y(u2__abc_44228_n19281) );
  AND2X2 AND2X2_9481 ( .A(u2__abc_44228_n19282), .B(u2__abc_44228_n2972_bF_buf62), .Y(u2__abc_44228_n19283) );
  AND2X2 AND2X2_9482 ( .A(u2__abc_44228_n19280), .B(u2__abc_44228_n19283), .Y(u2__abc_44228_n19284) );
  AND2X2 AND2X2_9483 ( .A(u2__abc_44228_n19285), .B(u2__abc_44228_n2966_bF_buf57), .Y(u2_root_126__FF_INPUT) );
  AND2X2 AND2X2_9484 ( .A(u2__abc_44228_n3062_bF_buf73), .B(sqrto_126_), .Y(u2__abc_44228_n19287) );
  AND2X2 AND2X2_9485 ( .A(u2__abc_44228_n19277), .B(sqrto_125_), .Y(u2__abc_44228_n19289) );
  AND2X2 AND2X2_9486 ( .A(u2__abc_44228_n19290), .B(u2__abc_44228_n19288), .Y(u2__abc_44228_n19291) );
  AND2X2 AND2X2_9487 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n5244), .Y(u2__abc_44228_n19293) );
  AND2X2 AND2X2_9488 ( .A(u2__abc_44228_n19294), .B(u2__abc_44228_n2972_bF_buf61), .Y(u2__abc_44228_n19295) );
  AND2X2 AND2X2_9489 ( .A(u2__abc_44228_n19292), .B(u2__abc_44228_n19295), .Y(u2__abc_44228_n19296) );
  AND2X2 AND2X2_949 ( .A(u2__abc_44228_n3894), .B(u2__abc_44228_n3897), .Y(u2__abc_44228_n3898) );
  AND2X2 AND2X2_9490 ( .A(u2__abc_44228_n19297), .B(u2__abc_44228_n2966_bF_buf56), .Y(u2_root_127__FF_INPUT) );
  AND2X2 AND2X2_9491 ( .A(u2__abc_44228_n3062_bF_buf72), .B(sqrto_127_), .Y(u2__abc_44228_n19299) );
  AND2X2 AND2X2_9492 ( .A(u2__abc_44228_n19289), .B(sqrto_126_), .Y(u2__abc_44228_n19301) );
  AND2X2 AND2X2_9493 ( .A(u2__abc_44228_n19302), .B(u2__abc_44228_n19300), .Y(u2__abc_44228_n19303) );
  AND2X2 AND2X2_9494 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n5237), .Y(u2__abc_44228_n19305) );
  AND2X2 AND2X2_9495 ( .A(u2__abc_44228_n19306), .B(u2__abc_44228_n2972_bF_buf60), .Y(u2__abc_44228_n19307) );
  AND2X2 AND2X2_9496 ( .A(u2__abc_44228_n19304), .B(u2__abc_44228_n19307), .Y(u2__abc_44228_n19308) );
  AND2X2 AND2X2_9497 ( .A(u2__abc_44228_n19309), .B(u2__abc_44228_n2966_bF_buf55), .Y(u2_root_128__FF_INPUT) );
  AND2X2 AND2X2_9498 ( .A(u2__abc_44228_n3062_bF_buf71), .B(sqrto_128_), .Y(u2__abc_44228_n19311) );
  AND2X2 AND2X2_9499 ( .A(u2__abc_44228_n19301), .B(sqrto_127_), .Y(u2__abc_44228_n19313) );
  AND2X2 AND2X2_95 ( .A(_abc_64468_n885), .B(_abc_64468_n884), .Y(_auto_iopadmap_cc_313_execute_65414_130_) );
  AND2X2 AND2X2_950 ( .A(u2__abc_44228_n3891), .B(u2__abc_44228_n3898), .Y(u2__abc_44228_n3899) );
  AND2X2 AND2X2_9500 ( .A(u2__abc_44228_n19314), .B(u2__abc_44228_n19312), .Y(u2__abc_44228_n19315) );
  AND2X2 AND2X2_9501 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n5233), .Y(u2__abc_44228_n19317) );
  AND2X2 AND2X2_9502 ( .A(u2__abc_44228_n19318), .B(u2__abc_44228_n2972_bF_buf59), .Y(u2__abc_44228_n19319) );
  AND2X2 AND2X2_9503 ( .A(u2__abc_44228_n19316), .B(u2__abc_44228_n19319), .Y(u2__abc_44228_n19320) );
  AND2X2 AND2X2_9504 ( .A(u2__abc_44228_n19321), .B(u2__abc_44228_n2966_bF_buf54), .Y(u2_root_129__FF_INPUT) );
  AND2X2 AND2X2_9505 ( .A(u2__abc_44228_n3062_bF_buf70), .B(sqrto_129_), .Y(u2__abc_44228_n19323) );
  AND2X2 AND2X2_9506 ( .A(u2__abc_44228_n19313), .B(sqrto_128_), .Y(u2__abc_44228_n19325) );
  AND2X2 AND2X2_9507 ( .A(u2__abc_44228_n19326), .B(u2__abc_44228_n19324), .Y(u2__abc_44228_n19327) );
  AND2X2 AND2X2_9508 ( .A(u2__abc_44228_n2983_bF_buf74), .B(u2__abc_44228_n5228), .Y(u2__abc_44228_n19329) );
  AND2X2 AND2X2_9509 ( .A(u2__abc_44228_n19330), .B(u2__abc_44228_n2972_bF_buf58), .Y(u2__abc_44228_n19331) );
  AND2X2 AND2X2_951 ( .A(u2__abc_44228_n3885), .B(u2__abc_44228_n3899), .Y(u2__abc_44228_n3900) );
  AND2X2 AND2X2_9510 ( .A(u2__abc_44228_n19328), .B(u2__abc_44228_n19331), .Y(u2__abc_44228_n19332) );
  AND2X2 AND2X2_9511 ( .A(u2__abc_44228_n19333), .B(u2__abc_44228_n2966_bF_buf53), .Y(u2_root_130__FF_INPUT) );
  AND2X2 AND2X2_9512 ( .A(u2__abc_44228_n3062_bF_buf69), .B(sqrto_130_), .Y(u2__abc_44228_n19335) );
  AND2X2 AND2X2_9513 ( .A(u2__abc_44228_n19325), .B(sqrto_129_), .Y(u2__abc_44228_n19337) );
  AND2X2 AND2X2_9514 ( .A(u2__abc_44228_n19338), .B(u2__abc_44228_n19336), .Y(u2__abc_44228_n19339) );
  AND2X2 AND2X2_9515 ( .A(u2__abc_44228_n2983_bF_buf72), .B(u2__abc_44228_n5218), .Y(u2__abc_44228_n19341) );
  AND2X2 AND2X2_9516 ( .A(u2__abc_44228_n19342), .B(u2__abc_44228_n2972_bF_buf57), .Y(u2__abc_44228_n19343) );
  AND2X2 AND2X2_9517 ( .A(u2__abc_44228_n19340), .B(u2__abc_44228_n19343), .Y(u2__abc_44228_n19344) );
  AND2X2 AND2X2_9518 ( .A(u2__abc_44228_n19345), .B(u2__abc_44228_n2966_bF_buf52), .Y(u2_root_131__FF_INPUT) );
  AND2X2 AND2X2_9519 ( .A(u2__abc_44228_n3062_bF_buf68), .B(sqrto_131_), .Y(u2__abc_44228_n19347) );
  AND2X2 AND2X2_952 ( .A(u2__abc_44228_n3871), .B(u2__abc_44228_n3900), .Y(u2__abc_44228_n3901) );
  AND2X2 AND2X2_9520 ( .A(u2__abc_44228_n19337), .B(sqrto_130_), .Y(u2__abc_44228_n19349) );
  AND2X2 AND2X2_9521 ( .A(u2__abc_44228_n19350), .B(u2__abc_44228_n19348), .Y(u2__abc_44228_n19351) );
  AND2X2 AND2X2_9522 ( .A(u2__abc_44228_n2983_bF_buf70), .B(u2__abc_44228_n5211_1), .Y(u2__abc_44228_n19353) );
  AND2X2 AND2X2_9523 ( .A(u2__abc_44228_n19354), .B(u2__abc_44228_n2972_bF_buf56), .Y(u2__abc_44228_n19355) );
  AND2X2 AND2X2_9524 ( .A(u2__abc_44228_n19352), .B(u2__abc_44228_n19355), .Y(u2__abc_44228_n19356) );
  AND2X2 AND2X2_9525 ( .A(u2__abc_44228_n19357), .B(u2__abc_44228_n2966_bF_buf51), .Y(u2_root_132__FF_INPUT) );
  AND2X2 AND2X2_9526 ( .A(u2__abc_44228_n3062_bF_buf67), .B(sqrto_132_), .Y(u2__abc_44228_n19359) );
  AND2X2 AND2X2_9527 ( .A(u2__abc_44228_n19349), .B(sqrto_131_), .Y(u2__abc_44228_n19361) );
  AND2X2 AND2X2_9528 ( .A(u2__abc_44228_n19362), .B(u2__abc_44228_n19360), .Y(u2__abc_44228_n19363) );
  AND2X2 AND2X2_9529 ( .A(u2__abc_44228_n2983_bF_buf68), .B(u2__abc_44228_n5204), .Y(u2__abc_44228_n19365) );
  AND2X2 AND2X2_953 ( .A(u2__abc_44228_n3842), .B(u2__abc_44228_n3901), .Y(u2__abc_44228_n3902) );
  AND2X2 AND2X2_9530 ( .A(u2__abc_44228_n19366), .B(u2__abc_44228_n2972_bF_buf55), .Y(u2__abc_44228_n19367) );
  AND2X2 AND2X2_9531 ( .A(u2__abc_44228_n19364), .B(u2__abc_44228_n19367), .Y(u2__abc_44228_n19368) );
  AND2X2 AND2X2_9532 ( .A(u2__abc_44228_n19369), .B(u2__abc_44228_n2966_bF_buf50), .Y(u2_root_133__FF_INPUT) );
  AND2X2 AND2X2_9533 ( .A(u2__abc_44228_n3062_bF_buf66), .B(sqrto_133_), .Y(u2__abc_44228_n19371) );
  AND2X2 AND2X2_9534 ( .A(u2__abc_44228_n19361), .B(sqrto_132_), .Y(u2__abc_44228_n19373) );
  AND2X2 AND2X2_9535 ( .A(u2__abc_44228_n19374), .B(u2__abc_44228_n19372), .Y(u2__abc_44228_n19375) );
  AND2X2 AND2X2_9536 ( .A(u2__abc_44228_n2983_bF_buf66), .B(u2__abc_44228_n5197), .Y(u2__abc_44228_n19377) );
  AND2X2 AND2X2_9537 ( .A(u2__abc_44228_n19378), .B(u2__abc_44228_n2972_bF_buf54), .Y(u2__abc_44228_n19379) );
  AND2X2 AND2X2_9538 ( .A(u2__abc_44228_n19376), .B(u2__abc_44228_n19379), .Y(u2__abc_44228_n19380) );
  AND2X2 AND2X2_9539 ( .A(u2__abc_44228_n19381), .B(u2__abc_44228_n2966_bF_buf49), .Y(u2_root_134__FF_INPUT) );
  AND2X2 AND2X2_954 ( .A(u2__abc_44228_n3783), .B(u2__abc_44228_n3902), .Y(u2__abc_44228_n3903_1) );
  AND2X2 AND2X2_9540 ( .A(u2__abc_44228_n3062_bF_buf65), .B(sqrto_134_), .Y(u2__abc_44228_n19383) );
  AND2X2 AND2X2_9541 ( .A(u2__abc_44228_n19373), .B(sqrto_133_), .Y(u2__abc_44228_n19385) );
  AND2X2 AND2X2_9542 ( .A(u2__abc_44228_n19386), .B(u2__abc_44228_n19384), .Y(u2__abc_44228_n19387) );
  AND2X2 AND2X2_9543 ( .A(u2__abc_44228_n2983_bF_buf64), .B(u2__abc_44228_n5174), .Y(u2__abc_44228_n19389) );
  AND2X2 AND2X2_9544 ( .A(u2__abc_44228_n19390), .B(u2__abc_44228_n2972_bF_buf53), .Y(u2__abc_44228_n19391) );
  AND2X2 AND2X2_9545 ( .A(u2__abc_44228_n19388), .B(u2__abc_44228_n19391), .Y(u2__abc_44228_n19392) );
  AND2X2 AND2X2_9546 ( .A(u2__abc_44228_n19393), .B(u2__abc_44228_n2966_bF_buf48), .Y(u2_root_135__FF_INPUT) );
  AND2X2 AND2X2_9547 ( .A(u2__abc_44228_n3062_bF_buf64), .B(sqrto_135_), .Y(u2__abc_44228_n19395) );
  AND2X2 AND2X2_9548 ( .A(u2__abc_44228_n19385), .B(sqrto_134_), .Y(u2__abc_44228_n19397) );
  AND2X2 AND2X2_9549 ( .A(u2__abc_44228_n19398), .B(u2__abc_44228_n19396), .Y(u2__abc_44228_n19399) );
  AND2X2 AND2X2_955 ( .A(u2__abc_44228_n3904), .B(u2_remHi_93_), .Y(u2__abc_44228_n3905) );
  AND2X2 AND2X2_9550 ( .A(u2__abc_44228_n2983_bF_buf62), .B(u2__abc_44228_n5167), .Y(u2__abc_44228_n19401) );
  AND2X2 AND2X2_9551 ( .A(u2__abc_44228_n19402), .B(u2__abc_44228_n2972_bF_buf52), .Y(u2__abc_44228_n19403) );
  AND2X2 AND2X2_9552 ( .A(u2__abc_44228_n19400), .B(u2__abc_44228_n19403), .Y(u2__abc_44228_n19404) );
  AND2X2 AND2X2_9553 ( .A(u2__abc_44228_n19405), .B(u2__abc_44228_n2966_bF_buf47), .Y(u2_root_136__FF_INPUT) );
  AND2X2 AND2X2_9554 ( .A(u2__abc_44228_n3062_bF_buf63), .B(sqrto_136_), .Y(u2__abc_44228_n19407) );
  AND2X2 AND2X2_9555 ( .A(u2__abc_44228_n19397), .B(sqrto_135_), .Y(u2__abc_44228_n19409) );
  AND2X2 AND2X2_9556 ( .A(u2__abc_44228_n19410), .B(u2__abc_44228_n19408), .Y(u2__abc_44228_n19411) );
  AND2X2 AND2X2_9557 ( .A(u2__abc_44228_n2983_bF_buf60), .B(u2__abc_44228_n5188), .Y(u2__abc_44228_n19413) );
  AND2X2 AND2X2_9558 ( .A(u2__abc_44228_n19414), .B(u2__abc_44228_n2972_bF_buf51), .Y(u2__abc_44228_n19415) );
  AND2X2 AND2X2_9559 ( .A(u2__abc_44228_n19412), .B(u2__abc_44228_n19415), .Y(u2__abc_44228_n19416) );
  AND2X2 AND2X2_956 ( .A(u2__abc_44228_n3907), .B(sqrto_93_), .Y(u2__abc_44228_n3908) );
  AND2X2 AND2X2_9560 ( .A(u2__abc_44228_n19417), .B(u2__abc_44228_n2966_bF_buf46), .Y(u2_root_137__FF_INPUT) );
  AND2X2 AND2X2_9561 ( .A(u2__abc_44228_n3062_bF_buf62), .B(sqrto_137_), .Y(u2__abc_44228_n19419) );
  AND2X2 AND2X2_9562 ( .A(u2__abc_44228_n19409), .B(sqrto_136_), .Y(u2__abc_44228_n19421) );
  AND2X2 AND2X2_9563 ( .A(u2__abc_44228_n19422), .B(u2__abc_44228_n19420), .Y(u2__abc_44228_n19423) );
  AND2X2 AND2X2_9564 ( .A(u2__abc_44228_n2983_bF_buf58), .B(u2__abc_44228_n5181), .Y(u2__abc_44228_n19425) );
  AND2X2 AND2X2_9565 ( .A(u2__abc_44228_n19426), .B(u2__abc_44228_n2972_bF_buf50), .Y(u2__abc_44228_n19427) );
  AND2X2 AND2X2_9566 ( .A(u2__abc_44228_n19424), .B(u2__abc_44228_n19427), .Y(u2__abc_44228_n19428) );
  AND2X2 AND2X2_9567 ( .A(u2__abc_44228_n19429), .B(u2__abc_44228_n2966_bF_buf45), .Y(u2_root_138__FF_INPUT) );
  AND2X2 AND2X2_9568 ( .A(u2__abc_44228_n3062_bF_buf61), .B(sqrto_138_), .Y(u2__abc_44228_n19431) );
  AND2X2 AND2X2_9569 ( .A(u2__abc_44228_n19421), .B(sqrto_137_), .Y(u2__abc_44228_n19433) );
  AND2X2 AND2X2_957 ( .A(u2__abc_44228_n3906), .B(u2__abc_44228_n3909), .Y(u2__abc_44228_n3910) );
  AND2X2 AND2X2_9570 ( .A(u2__abc_44228_n19434), .B(u2__abc_44228_n19432), .Y(u2__abc_44228_n19435) );
  AND2X2 AND2X2_9571 ( .A(u2__abc_44228_n2983_bF_buf56), .B(u2__abc_44228_n5159), .Y(u2__abc_44228_n19437) );
  AND2X2 AND2X2_9572 ( .A(u2__abc_44228_n19438), .B(u2__abc_44228_n2972_bF_buf49), .Y(u2__abc_44228_n19439) );
  AND2X2 AND2X2_9573 ( .A(u2__abc_44228_n19436), .B(u2__abc_44228_n19439), .Y(u2__abc_44228_n19440) );
  AND2X2 AND2X2_9574 ( .A(u2__abc_44228_n19441), .B(u2__abc_44228_n2966_bF_buf44), .Y(u2_root_139__FF_INPUT) );
  AND2X2 AND2X2_9575 ( .A(u2__abc_44228_n3062_bF_buf60), .B(sqrto_139_), .Y(u2__abc_44228_n19443) );
  AND2X2 AND2X2_9576 ( .A(u2__abc_44228_n19433), .B(sqrto_138_), .Y(u2__abc_44228_n19445) );
  AND2X2 AND2X2_9577 ( .A(u2__abc_44228_n19446), .B(u2__abc_44228_n19444), .Y(u2__abc_44228_n19447) );
  AND2X2 AND2X2_9578 ( .A(u2__abc_44228_n2983_bF_buf54), .B(u2__abc_44228_n5152), .Y(u2__abc_44228_n19449) );
  AND2X2 AND2X2_9579 ( .A(u2__abc_44228_n19450), .B(u2__abc_44228_n2972_bF_buf48), .Y(u2__abc_44228_n19451) );
  AND2X2 AND2X2_958 ( .A(u2__abc_44228_n3911), .B(u2_remHi_92_), .Y(u2__abc_44228_n3912_1) );
  AND2X2 AND2X2_9580 ( .A(u2__abc_44228_n19448), .B(u2__abc_44228_n19451), .Y(u2__abc_44228_n19452) );
  AND2X2 AND2X2_9581 ( .A(u2__abc_44228_n19453), .B(u2__abc_44228_n2966_bF_buf43), .Y(u2_root_140__FF_INPUT) );
  AND2X2 AND2X2_9582 ( .A(u2__abc_44228_n3062_bF_buf59), .B(sqrto_140_), .Y(u2__abc_44228_n19455) );
  AND2X2 AND2X2_9583 ( .A(u2__abc_44228_n19445), .B(sqrto_139_), .Y(u2__abc_44228_n19457) );
  AND2X2 AND2X2_9584 ( .A(u2__abc_44228_n19458), .B(u2__abc_44228_n19456), .Y(u2__abc_44228_n19459) );
  AND2X2 AND2X2_9585 ( .A(u2__abc_44228_n2983_bF_buf52), .B(u2__abc_44228_n5145), .Y(u2__abc_44228_n19461) );
  AND2X2 AND2X2_9586 ( .A(u2__abc_44228_n19462), .B(u2__abc_44228_n2972_bF_buf47), .Y(u2__abc_44228_n19463) );
  AND2X2 AND2X2_9587 ( .A(u2__abc_44228_n19460), .B(u2__abc_44228_n19463), .Y(u2__abc_44228_n19464) );
  AND2X2 AND2X2_9588 ( .A(u2__abc_44228_n19465), .B(u2__abc_44228_n2966_bF_buf42), .Y(u2_root_141__FF_INPUT) );
  AND2X2 AND2X2_9589 ( .A(u2__abc_44228_n3062_bF_buf58), .B(sqrto_141_), .Y(u2__abc_44228_n19467) );
  AND2X2 AND2X2_959 ( .A(u2__abc_44228_n3913), .B(sqrto_92_), .Y(u2__abc_44228_n3914) );
  AND2X2 AND2X2_9590 ( .A(u2__abc_44228_n19457), .B(sqrto_140_), .Y(u2__abc_44228_n19469) );
  AND2X2 AND2X2_9591 ( .A(u2__abc_44228_n19470), .B(u2__abc_44228_n19468), .Y(u2__abc_44228_n19471) );
  AND2X2 AND2X2_9592 ( .A(u2__abc_44228_n2983_bF_buf50), .B(u2__abc_44228_n5138), .Y(u2__abc_44228_n19473) );
  AND2X2 AND2X2_9593 ( .A(u2__abc_44228_n19474), .B(u2__abc_44228_n2972_bF_buf46), .Y(u2__abc_44228_n19475) );
  AND2X2 AND2X2_9594 ( .A(u2__abc_44228_n19472), .B(u2__abc_44228_n19475), .Y(u2__abc_44228_n19476) );
  AND2X2 AND2X2_9595 ( .A(u2__abc_44228_n19477), .B(u2__abc_44228_n2966_bF_buf41), .Y(u2_root_142__FF_INPUT) );
  AND2X2 AND2X2_9596 ( .A(u2__abc_44228_n3062_bF_buf57), .B(sqrto_142_), .Y(u2__abc_44228_n19479) );
  AND2X2 AND2X2_9597 ( .A(u2__abc_44228_n19469), .B(sqrto_141_), .Y(u2__abc_44228_n19481) );
  AND2X2 AND2X2_9598 ( .A(u2__abc_44228_n19482), .B(u2__abc_44228_n19480), .Y(u2__abc_44228_n19483) );
  AND2X2 AND2X2_9599 ( .A(u2__abc_44228_n2983_bF_buf48), .B(u2__abc_44228_n5128), .Y(u2__abc_44228_n19485) );
  AND2X2 AND2X2_96 ( .A(_abc_64468_n888), .B(_abc_64468_n887), .Y(_auto_iopadmap_cc_313_execute_65414_131_) );
  AND2X2 AND2X2_960 ( .A(u2__abc_44228_n3916), .B(u2__abc_44228_n3910), .Y(u2__abc_44228_n3917) );
  AND2X2 AND2X2_9600 ( .A(u2__abc_44228_n19486), .B(u2__abc_44228_n2972_bF_buf45), .Y(u2__abc_44228_n19487) );
  AND2X2 AND2X2_9601 ( .A(u2__abc_44228_n19484), .B(u2__abc_44228_n19487), .Y(u2__abc_44228_n19488) );
  AND2X2 AND2X2_9602 ( .A(u2__abc_44228_n19489), .B(u2__abc_44228_n2966_bF_buf40), .Y(u2_root_143__FF_INPUT) );
  AND2X2 AND2X2_9603 ( .A(u2__abc_44228_n3062_bF_buf56), .B(sqrto_143_), .Y(u2__abc_44228_n19491) );
  AND2X2 AND2X2_9604 ( .A(u2__abc_44228_n19481), .B(sqrto_142_), .Y(u2__abc_44228_n19493) );
  AND2X2 AND2X2_9605 ( .A(u2__abc_44228_n19494), .B(u2__abc_44228_n19492), .Y(u2__abc_44228_n19495) );
  AND2X2 AND2X2_9606 ( .A(u2__abc_44228_n2983_bF_buf46), .B(u2__abc_44228_n5121), .Y(u2__abc_44228_n19497) );
  AND2X2 AND2X2_9607 ( .A(u2__abc_44228_n19498), .B(u2__abc_44228_n2972_bF_buf44), .Y(u2__abc_44228_n19499) );
  AND2X2 AND2X2_9608 ( .A(u2__abc_44228_n19496), .B(u2__abc_44228_n19499), .Y(u2__abc_44228_n19500) );
  AND2X2 AND2X2_9609 ( .A(u2__abc_44228_n19501), .B(u2__abc_44228_n2966_bF_buf39), .Y(u2_root_144__FF_INPUT) );
  AND2X2 AND2X2_961 ( .A(u2__abc_44228_n3918), .B(u2_remHi_90_), .Y(u2__abc_44228_n3919) );
  AND2X2 AND2X2_9610 ( .A(u2__abc_44228_n3062_bF_buf55), .B(sqrto_144_), .Y(u2__abc_44228_n19503) );
  AND2X2 AND2X2_9611 ( .A(u2__abc_44228_n19493), .B(sqrto_143_), .Y(u2__abc_44228_n19505) );
  AND2X2 AND2X2_9612 ( .A(u2__abc_44228_n19506), .B(u2__abc_44228_n19504), .Y(u2__abc_44228_n19507) );
  AND2X2 AND2X2_9613 ( .A(u2__abc_44228_n2983_bF_buf44), .B(u2__abc_44228_n5114), .Y(u2__abc_44228_n19509) );
  AND2X2 AND2X2_9614 ( .A(u2__abc_44228_n19510), .B(u2__abc_44228_n2972_bF_buf43), .Y(u2__abc_44228_n19511) );
  AND2X2 AND2X2_9615 ( .A(u2__abc_44228_n19508), .B(u2__abc_44228_n19511), .Y(u2__abc_44228_n19512) );
  AND2X2 AND2X2_9616 ( .A(u2__abc_44228_n19513), .B(u2__abc_44228_n2966_bF_buf38), .Y(u2_root_145__FF_INPUT) );
  AND2X2 AND2X2_9617 ( .A(u2__abc_44228_n3062_bF_buf54), .B(sqrto_145_), .Y(u2__abc_44228_n19515) );
  AND2X2 AND2X2_9618 ( .A(u2__abc_44228_n19505), .B(sqrto_144_), .Y(u2__abc_44228_n19517) );
  AND2X2 AND2X2_9619 ( .A(u2__abc_44228_n19518), .B(u2__abc_44228_n19516), .Y(u2__abc_44228_n19519) );
  AND2X2 AND2X2_962 ( .A(u2__abc_44228_n3920), .B(sqrto_90_), .Y(u2__abc_44228_n3921_1) );
  AND2X2 AND2X2_9620 ( .A(u2__abc_44228_n2983_bF_buf42), .B(u2__abc_44228_n5107), .Y(u2__abc_44228_n19521) );
  AND2X2 AND2X2_9621 ( .A(u2__abc_44228_n19522), .B(u2__abc_44228_n2972_bF_buf42), .Y(u2__abc_44228_n19523) );
  AND2X2 AND2X2_9622 ( .A(u2__abc_44228_n19520), .B(u2__abc_44228_n19523), .Y(u2__abc_44228_n19524) );
  AND2X2 AND2X2_9623 ( .A(u2__abc_44228_n19525), .B(u2__abc_44228_n2966_bF_buf37), .Y(u2_root_146__FF_INPUT) );
  AND2X2 AND2X2_9624 ( .A(u2__abc_44228_n3062_bF_buf53), .B(sqrto_146_), .Y(u2__abc_44228_n19527) );
  AND2X2 AND2X2_9625 ( .A(u2__abc_44228_n19517), .B(sqrto_145_), .Y(u2__abc_44228_n19529) );
  AND2X2 AND2X2_9626 ( .A(u2__abc_44228_n19530), .B(u2__abc_44228_n19528), .Y(u2__abc_44228_n19531) );
  AND2X2 AND2X2_9627 ( .A(u2__abc_44228_n2983_bF_buf40), .B(u2__abc_44228_n5092), .Y(u2__abc_44228_n19533) );
  AND2X2 AND2X2_9628 ( .A(u2__abc_44228_n19534), .B(u2__abc_44228_n2972_bF_buf41), .Y(u2__abc_44228_n19535) );
  AND2X2 AND2X2_9629 ( .A(u2__abc_44228_n19532), .B(u2__abc_44228_n19535), .Y(u2__abc_44228_n19536) );
  AND2X2 AND2X2_963 ( .A(u2__abc_44228_n3924), .B(u2_remHi_91_), .Y(u2__abc_44228_n3925) );
  AND2X2 AND2X2_9630 ( .A(u2__abc_44228_n19537), .B(u2__abc_44228_n2966_bF_buf36), .Y(u2_root_147__FF_INPUT) );
  AND2X2 AND2X2_9631 ( .A(u2__abc_44228_n3062_bF_buf52), .B(sqrto_147_), .Y(u2__abc_44228_n19539) );
  AND2X2 AND2X2_9632 ( .A(u2__abc_44228_n19529), .B(sqrto_146_), .Y(u2__abc_44228_n19541) );
  AND2X2 AND2X2_9633 ( .A(u2__abc_44228_n19542), .B(u2__abc_44228_n19540), .Y(u2__abc_44228_n19543) );
  AND2X2 AND2X2_9634 ( .A(u2__abc_44228_n2983_bF_buf38), .B(u2__abc_44228_n5098), .Y(u2__abc_44228_n19545) );
  AND2X2 AND2X2_9635 ( .A(u2__abc_44228_n19546), .B(u2__abc_44228_n2972_bF_buf40), .Y(u2__abc_44228_n19547) );
  AND2X2 AND2X2_9636 ( .A(u2__abc_44228_n19544), .B(u2__abc_44228_n19547), .Y(u2__abc_44228_n19548) );
  AND2X2 AND2X2_9637 ( .A(u2__abc_44228_n19549), .B(u2__abc_44228_n2966_bF_buf35), .Y(u2_root_148__FF_INPUT) );
  AND2X2 AND2X2_9638 ( .A(u2__abc_44228_n3062_bF_buf51), .B(sqrto_148_), .Y(u2__abc_44228_n19551) );
  AND2X2 AND2X2_9639 ( .A(u2__abc_44228_n19541), .B(sqrto_147_), .Y(u2__abc_44228_n19553) );
  AND2X2 AND2X2_964 ( .A(u2__abc_44228_n3927), .B(sqrto_91_), .Y(u2__abc_44228_n3928) );
  AND2X2 AND2X2_9640 ( .A(u2__abc_44228_n19554), .B(u2__abc_44228_n19552), .Y(u2__abc_44228_n19555) );
  AND2X2 AND2X2_9641 ( .A(u2__abc_44228_n2983_bF_buf36), .B(u2__abc_44228_n5085), .Y(u2__abc_44228_n19557) );
  AND2X2 AND2X2_9642 ( .A(u2__abc_44228_n19558), .B(u2__abc_44228_n2972_bF_buf39), .Y(u2__abc_44228_n19559) );
  AND2X2 AND2X2_9643 ( .A(u2__abc_44228_n19556), .B(u2__abc_44228_n19559), .Y(u2__abc_44228_n19560) );
  AND2X2 AND2X2_9644 ( .A(u2__abc_44228_n19561), .B(u2__abc_44228_n2966_bF_buf34), .Y(u2_root_149__FF_INPUT) );
  AND2X2 AND2X2_9645 ( .A(u2__abc_44228_n3062_bF_buf50), .B(sqrto_149_), .Y(u2__abc_44228_n19563) );
  AND2X2 AND2X2_9646 ( .A(u2__abc_44228_n19553), .B(sqrto_148_), .Y(u2__abc_44228_n19565) );
  AND2X2 AND2X2_9647 ( .A(u2__abc_44228_n19566), .B(u2__abc_44228_n19564), .Y(u2__abc_44228_n19567) );
  AND2X2 AND2X2_9648 ( .A(u2__abc_44228_n2983_bF_buf34), .B(u2__abc_44228_n5078), .Y(u2__abc_44228_n19569) );
  AND2X2 AND2X2_9649 ( .A(u2__abc_44228_n19570), .B(u2__abc_44228_n2972_bF_buf38), .Y(u2__abc_44228_n19571) );
  AND2X2 AND2X2_965 ( .A(u2__abc_44228_n3926), .B(u2__abc_44228_n3929), .Y(u2__abc_44228_n3930_1) );
  AND2X2 AND2X2_9650 ( .A(u2__abc_44228_n19568), .B(u2__abc_44228_n19571), .Y(u2__abc_44228_n19572) );
  AND2X2 AND2X2_9651 ( .A(u2__abc_44228_n19573), .B(u2__abc_44228_n2966_bF_buf33), .Y(u2_root_150__FF_INPUT) );
  AND2X2 AND2X2_9652 ( .A(u2__abc_44228_n3062_bF_buf49), .B(sqrto_150_), .Y(u2__abc_44228_n19575) );
  AND2X2 AND2X2_9653 ( .A(u2__abc_44228_n19565), .B(sqrto_149_), .Y(u2__abc_44228_n19577) );
  AND2X2 AND2X2_9654 ( .A(u2__abc_44228_n19578), .B(u2__abc_44228_n19576), .Y(u2__abc_44228_n19579) );
  AND2X2 AND2X2_9655 ( .A(u2__abc_44228_n2983_bF_buf32), .B(u2__abc_44228_n5062), .Y(u2__abc_44228_n19581) );
  AND2X2 AND2X2_9656 ( .A(u2__abc_44228_n19582), .B(u2__abc_44228_n2972_bF_buf37), .Y(u2__abc_44228_n19583) );
  AND2X2 AND2X2_9657 ( .A(u2__abc_44228_n19580), .B(u2__abc_44228_n19583), .Y(u2__abc_44228_n19584) );
  AND2X2 AND2X2_9658 ( .A(u2__abc_44228_n19585), .B(u2__abc_44228_n2966_bF_buf32), .Y(u2_root_151__FF_INPUT) );
  AND2X2 AND2X2_9659 ( .A(u2__abc_44228_n3062_bF_buf48), .B(sqrto_151_), .Y(u2__abc_44228_n19587) );
  AND2X2 AND2X2_966 ( .A(u2__abc_44228_n3923), .B(u2__abc_44228_n3930_1), .Y(u2__abc_44228_n3931) );
  AND2X2 AND2X2_9660 ( .A(u2__abc_44228_n19577), .B(sqrto_150_), .Y(u2__abc_44228_n19589) );
  AND2X2 AND2X2_9661 ( .A(u2__abc_44228_n19590), .B(u2__abc_44228_n19588), .Y(u2__abc_44228_n19591) );
  AND2X2 AND2X2_9662 ( .A(u2__abc_44228_n2983_bF_buf30), .B(u2__abc_44228_n5068), .Y(u2__abc_44228_n19593) );
  AND2X2 AND2X2_9663 ( .A(u2__abc_44228_n19594), .B(u2__abc_44228_n2972_bF_buf36), .Y(u2__abc_44228_n19595) );
  AND2X2 AND2X2_9664 ( .A(u2__abc_44228_n19592), .B(u2__abc_44228_n19595), .Y(u2__abc_44228_n19596) );
  AND2X2 AND2X2_9665 ( .A(u2__abc_44228_n19597), .B(u2__abc_44228_n2966_bF_buf31), .Y(u2_root_152__FF_INPUT) );
  AND2X2 AND2X2_9666 ( .A(u2__abc_44228_n3062_bF_buf47), .B(sqrto_152_), .Y(u2__abc_44228_n19599) );
  AND2X2 AND2X2_9667 ( .A(u2__abc_44228_n19589), .B(sqrto_151_), .Y(u2__abc_44228_n19601) );
  AND2X2 AND2X2_9668 ( .A(u2__abc_44228_n19602), .B(u2__abc_44228_n19600), .Y(u2__abc_44228_n19603) );
  AND2X2 AND2X2_9669 ( .A(u2__abc_44228_n2983_bF_buf28), .B(u2__abc_44228_n5055), .Y(u2__abc_44228_n19605) );
  AND2X2 AND2X2_967 ( .A(u2__abc_44228_n3917), .B(u2__abc_44228_n3931), .Y(u2__abc_44228_n3932) );
  AND2X2 AND2X2_9670 ( .A(u2__abc_44228_n19606), .B(u2__abc_44228_n2972_bF_buf35), .Y(u2__abc_44228_n19607) );
  AND2X2 AND2X2_9671 ( .A(u2__abc_44228_n19604), .B(u2__abc_44228_n19607), .Y(u2__abc_44228_n19608) );
  AND2X2 AND2X2_9672 ( .A(u2__abc_44228_n19609), .B(u2__abc_44228_n2966_bF_buf30), .Y(u2_root_153__FF_INPUT) );
  AND2X2 AND2X2_9673 ( .A(u2__abc_44228_n3062_bF_buf46), .B(sqrto_153_), .Y(u2__abc_44228_n19611) );
  AND2X2 AND2X2_9674 ( .A(u2__abc_44228_n19601), .B(sqrto_152_), .Y(u2__abc_44228_n19613) );
  AND2X2 AND2X2_9675 ( .A(u2__abc_44228_n19614), .B(u2__abc_44228_n19612), .Y(u2__abc_44228_n19615) );
  AND2X2 AND2X2_9676 ( .A(u2__abc_44228_n2983_bF_buf26), .B(u2__abc_44228_n5048), .Y(u2__abc_44228_n19617) );
  AND2X2 AND2X2_9677 ( .A(u2__abc_44228_n19618), .B(u2__abc_44228_n2972_bF_buf34), .Y(u2__abc_44228_n19619) );
  AND2X2 AND2X2_9678 ( .A(u2__abc_44228_n19616), .B(u2__abc_44228_n19619), .Y(u2__abc_44228_n19620) );
  AND2X2 AND2X2_9679 ( .A(u2__abc_44228_n19621), .B(u2__abc_44228_n2966_bF_buf29), .Y(u2_root_154__FF_INPUT) );
  AND2X2 AND2X2_968 ( .A(u2__abc_44228_n3933), .B(u2_remHi_89_), .Y(u2__abc_44228_n3934) );
  AND2X2 AND2X2_9680 ( .A(u2__abc_44228_n3062_bF_buf45), .B(sqrto_154_), .Y(u2__abc_44228_n19623) );
  AND2X2 AND2X2_9681 ( .A(u2__abc_44228_n19613), .B(sqrto_153_), .Y(u2__abc_44228_n19625) );
  AND2X2 AND2X2_9682 ( .A(u2__abc_44228_n19626), .B(u2__abc_44228_n19624), .Y(u2__abc_44228_n19627) );
  AND2X2 AND2X2_9683 ( .A(u2__abc_44228_n2983_bF_buf24), .B(u2__abc_44228_n5040), .Y(u2__abc_44228_n19629) );
  AND2X2 AND2X2_9684 ( .A(u2__abc_44228_n19630), .B(u2__abc_44228_n2972_bF_buf33), .Y(u2__abc_44228_n19631) );
  AND2X2 AND2X2_9685 ( .A(u2__abc_44228_n19628), .B(u2__abc_44228_n19631), .Y(u2__abc_44228_n19632) );
  AND2X2 AND2X2_9686 ( .A(u2__abc_44228_n19633), .B(u2__abc_44228_n2966_bF_buf28), .Y(u2_root_155__FF_INPUT) );
  AND2X2 AND2X2_9687 ( .A(u2__abc_44228_n3062_bF_buf44), .B(sqrto_155_), .Y(u2__abc_44228_n19635) );
  AND2X2 AND2X2_9688 ( .A(u2__abc_44228_n19625), .B(sqrto_154_), .Y(u2__abc_44228_n19637) );
  AND2X2 AND2X2_9689 ( .A(u2__abc_44228_n19638), .B(u2__abc_44228_n19636), .Y(u2__abc_44228_n19639) );
  AND2X2 AND2X2_969 ( .A(u2__abc_44228_n3936), .B(sqrto_89_), .Y(u2__abc_44228_n3937) );
  AND2X2 AND2X2_9690 ( .A(u2__abc_44228_n2983_bF_buf22), .B(u2__abc_44228_n5033), .Y(u2__abc_44228_n19641) );
  AND2X2 AND2X2_9691 ( .A(u2__abc_44228_n19642), .B(u2__abc_44228_n2972_bF_buf32), .Y(u2__abc_44228_n19643) );
  AND2X2 AND2X2_9692 ( .A(u2__abc_44228_n19640), .B(u2__abc_44228_n19643), .Y(u2__abc_44228_n19644) );
  AND2X2 AND2X2_9693 ( .A(u2__abc_44228_n19645), .B(u2__abc_44228_n2966_bF_buf27), .Y(u2_root_156__FF_INPUT) );
  AND2X2 AND2X2_9694 ( .A(u2__abc_44228_n3062_bF_buf43), .B(sqrto_156_), .Y(u2__abc_44228_n19647) );
  AND2X2 AND2X2_9695 ( .A(u2__abc_44228_n19637), .B(sqrto_155_), .Y(u2__abc_44228_n19649) );
  AND2X2 AND2X2_9696 ( .A(u2__abc_44228_n19650), .B(u2__abc_44228_n19648), .Y(u2__abc_44228_n19651) );
  AND2X2 AND2X2_9697 ( .A(u2__abc_44228_n2983_bF_buf20), .B(u2__abc_44228_n5026), .Y(u2__abc_44228_n19653) );
  AND2X2 AND2X2_9698 ( .A(u2__abc_44228_n19654), .B(u2__abc_44228_n2972_bF_buf31), .Y(u2__abc_44228_n19655) );
  AND2X2 AND2X2_9699 ( .A(u2__abc_44228_n19652), .B(u2__abc_44228_n19655), .Y(u2__abc_44228_n19656) );
  AND2X2 AND2X2_97 ( .A(_abc_64468_n891), .B(_abc_64468_n890), .Y(_auto_iopadmap_cc_313_execute_65414_132_) );
  AND2X2 AND2X2_970 ( .A(u2__abc_44228_n3935), .B(u2__abc_44228_n3938), .Y(u2__abc_44228_n3939) );
  AND2X2 AND2X2_9700 ( .A(u2__abc_44228_n19657), .B(u2__abc_44228_n2966_bF_buf26), .Y(u2_root_157__FF_INPUT) );
  AND2X2 AND2X2_9701 ( .A(u2__abc_44228_n3062_bF_buf42), .B(sqrto_157_), .Y(u2__abc_44228_n19659) );
  AND2X2 AND2X2_9702 ( .A(u2__abc_44228_n19649), .B(sqrto_156_), .Y(u2__abc_44228_n19661) );
  AND2X2 AND2X2_9703 ( .A(u2__abc_44228_n19662), .B(u2__abc_44228_n19660), .Y(u2__abc_44228_n19663) );
  AND2X2 AND2X2_9704 ( .A(u2__abc_44228_n2983_bF_buf18), .B(u2__abc_44228_n5019), .Y(u2__abc_44228_n19665) );
  AND2X2 AND2X2_9705 ( .A(u2__abc_44228_n19666), .B(u2__abc_44228_n2972_bF_buf30), .Y(u2__abc_44228_n19667) );
  AND2X2 AND2X2_9706 ( .A(u2__abc_44228_n19664), .B(u2__abc_44228_n19667), .Y(u2__abc_44228_n19668) );
  AND2X2 AND2X2_9707 ( .A(u2__abc_44228_n19669), .B(u2__abc_44228_n2966_bF_buf25), .Y(u2_root_158__FF_INPUT) );
  AND2X2 AND2X2_9708 ( .A(u2__abc_44228_n3062_bF_buf41), .B(sqrto_158_), .Y(u2__abc_44228_n19671) );
  AND2X2 AND2X2_9709 ( .A(u2__abc_44228_n19661), .B(sqrto_157_), .Y(u2__abc_44228_n19673) );
  AND2X2 AND2X2_971 ( .A(u2__abc_44228_n3940_1), .B(u2_remHi_88_), .Y(u2__abc_44228_n3941) );
  AND2X2 AND2X2_9710 ( .A(u2__abc_44228_n19674), .B(u2__abc_44228_n19672), .Y(u2__abc_44228_n19675) );
  AND2X2 AND2X2_9711 ( .A(u2__abc_44228_n2983_bF_buf16), .B(u2__abc_44228_n5001), .Y(u2__abc_44228_n19677) );
  AND2X2 AND2X2_9712 ( .A(u2__abc_44228_n19678), .B(u2__abc_44228_n2972_bF_buf29), .Y(u2__abc_44228_n19679) );
  AND2X2 AND2X2_9713 ( .A(u2__abc_44228_n19676), .B(u2__abc_44228_n19679), .Y(u2__abc_44228_n19680) );
  AND2X2 AND2X2_9714 ( .A(u2__abc_44228_n19681), .B(u2__abc_44228_n2966_bF_buf24), .Y(u2_root_159__FF_INPUT) );
  AND2X2 AND2X2_9715 ( .A(u2__abc_44228_n3062_bF_buf40), .B(sqrto_159_), .Y(u2__abc_44228_n19683) );
  AND2X2 AND2X2_9716 ( .A(u2__abc_44228_n19673), .B(sqrto_158_), .Y(u2__abc_44228_n19685) );
  AND2X2 AND2X2_9717 ( .A(u2__abc_44228_n19686), .B(u2__abc_44228_n19684), .Y(u2__abc_44228_n19687) );
  AND2X2 AND2X2_9718 ( .A(u2__abc_44228_n2983_bF_buf14), .B(u2__abc_44228_n5007), .Y(u2__abc_44228_n19689) );
  AND2X2 AND2X2_9719 ( .A(u2__abc_44228_n19690), .B(u2__abc_44228_n2972_bF_buf28), .Y(u2__abc_44228_n19691) );
  AND2X2 AND2X2_972 ( .A(u2__abc_44228_n3942), .B(sqrto_88_), .Y(u2__abc_44228_n3943) );
  AND2X2 AND2X2_9720 ( .A(u2__abc_44228_n19688), .B(u2__abc_44228_n19691), .Y(u2__abc_44228_n19692) );
  AND2X2 AND2X2_9721 ( .A(u2__abc_44228_n19693), .B(u2__abc_44228_n2966_bF_buf23), .Y(u2_root_160__FF_INPUT) );
  AND2X2 AND2X2_9722 ( .A(u2__abc_44228_n3062_bF_buf39), .B(sqrto_160_), .Y(u2__abc_44228_n19695) );
  AND2X2 AND2X2_9723 ( .A(u2__abc_44228_n19685), .B(sqrto_159_), .Y(u2__abc_44228_n19697) );
  AND2X2 AND2X2_9724 ( .A(u2__abc_44228_n19698), .B(u2__abc_44228_n19696), .Y(u2__abc_44228_n19699) );
  AND2X2 AND2X2_9725 ( .A(u2__abc_44228_n2983_bF_buf12), .B(u2__abc_44228_n4994), .Y(u2__abc_44228_n19701) );
  AND2X2 AND2X2_9726 ( .A(u2__abc_44228_n19702), .B(u2__abc_44228_n2972_bF_buf27), .Y(u2__abc_44228_n19703) );
  AND2X2 AND2X2_9727 ( .A(u2__abc_44228_n19700), .B(u2__abc_44228_n19703), .Y(u2__abc_44228_n19704) );
  AND2X2 AND2X2_9728 ( .A(u2__abc_44228_n19705), .B(u2__abc_44228_n2966_bF_buf22), .Y(u2_root_161__FF_INPUT) );
  AND2X2 AND2X2_9729 ( .A(u2__abc_44228_n3062_bF_buf38), .B(sqrto_161_), .Y(u2__abc_44228_n19707) );
  AND2X2 AND2X2_973 ( .A(u2__abc_44228_n3945), .B(u2__abc_44228_n3939), .Y(u2__abc_44228_n3946) );
  AND2X2 AND2X2_9730 ( .A(u2__abc_44228_n19697), .B(sqrto_160_), .Y(u2__abc_44228_n19709) );
  AND2X2 AND2X2_9731 ( .A(u2__abc_44228_n19710), .B(u2__abc_44228_n19708), .Y(u2__abc_44228_n19711) );
  AND2X2 AND2X2_9732 ( .A(u2__abc_44228_n2983_bF_buf10), .B(u2__abc_44228_n4987), .Y(u2__abc_44228_n19713) );
  AND2X2 AND2X2_9733 ( .A(u2__abc_44228_n19714), .B(u2__abc_44228_n2972_bF_buf26), .Y(u2__abc_44228_n19715) );
  AND2X2 AND2X2_9734 ( .A(u2__abc_44228_n19712), .B(u2__abc_44228_n19715), .Y(u2__abc_44228_n19716) );
  AND2X2 AND2X2_9735 ( .A(u2__abc_44228_n19717), .B(u2__abc_44228_n2966_bF_buf21), .Y(u2_root_162__FF_INPUT) );
  AND2X2 AND2X2_9736 ( .A(u2__abc_44228_n3062_bF_buf37), .B(sqrto_162_), .Y(u2__abc_44228_n19719) );
  AND2X2 AND2X2_9737 ( .A(u2__abc_44228_n19709), .B(sqrto_161_), .Y(u2__abc_44228_n19721) );
  AND2X2 AND2X2_9738 ( .A(u2__abc_44228_n19722), .B(u2__abc_44228_n19720), .Y(u2__abc_44228_n19723) );
  AND2X2 AND2X2_9739 ( .A(u2__abc_44228_n2983_bF_buf8), .B(u2__abc_44228_n4972), .Y(u2__abc_44228_n19725) );
  AND2X2 AND2X2_974 ( .A(u2__abc_44228_n3947), .B(u2_remHi_86_), .Y(u2__abc_44228_n3948) );
  AND2X2 AND2X2_9740 ( .A(u2__abc_44228_n19726), .B(u2__abc_44228_n2972_bF_buf25), .Y(u2__abc_44228_n19727) );
  AND2X2 AND2X2_9741 ( .A(u2__abc_44228_n19724), .B(u2__abc_44228_n19727), .Y(u2__abc_44228_n19728) );
  AND2X2 AND2X2_9742 ( .A(u2__abc_44228_n19729), .B(u2__abc_44228_n2966_bF_buf20), .Y(u2_root_163__FF_INPUT) );
  AND2X2 AND2X2_9743 ( .A(u2__abc_44228_n3062_bF_buf36), .B(sqrto_163_), .Y(u2__abc_44228_n19731) );
  AND2X2 AND2X2_9744 ( .A(u2__abc_44228_n19721), .B(sqrto_162_), .Y(u2__abc_44228_n19733) );
  AND2X2 AND2X2_9745 ( .A(u2__abc_44228_n19734), .B(u2__abc_44228_n19732), .Y(u2__abc_44228_n19735) );
  AND2X2 AND2X2_9746 ( .A(u2__abc_44228_n2983_bF_buf6), .B(u2__abc_44228_n4978), .Y(u2__abc_44228_n19737) );
  AND2X2 AND2X2_9747 ( .A(u2__abc_44228_n19738), .B(u2__abc_44228_n2972_bF_buf24), .Y(u2__abc_44228_n19739) );
  AND2X2 AND2X2_9748 ( .A(u2__abc_44228_n19736), .B(u2__abc_44228_n19739), .Y(u2__abc_44228_n19740) );
  AND2X2 AND2X2_9749 ( .A(u2__abc_44228_n19741), .B(u2__abc_44228_n2966_bF_buf19), .Y(u2_root_164__FF_INPUT) );
  AND2X2 AND2X2_975 ( .A(u2__abc_44228_n3949_1), .B(sqrto_86_), .Y(u2__abc_44228_n3950) );
  AND2X2 AND2X2_9750 ( .A(u2__abc_44228_n3062_bF_buf35), .B(sqrto_164_), .Y(u2__abc_44228_n19743) );
  AND2X2 AND2X2_9751 ( .A(u2__abc_44228_n19733), .B(sqrto_163_), .Y(u2__abc_44228_n19745) );
  AND2X2 AND2X2_9752 ( .A(u2__abc_44228_n19746), .B(u2__abc_44228_n19744), .Y(u2__abc_44228_n19747) );
  AND2X2 AND2X2_9753 ( .A(u2__abc_44228_n2983_bF_buf4), .B(u2__abc_44228_n4965), .Y(u2__abc_44228_n19749) );
  AND2X2 AND2X2_9754 ( .A(u2__abc_44228_n19750), .B(u2__abc_44228_n2972_bF_buf23), .Y(u2__abc_44228_n19751) );
  AND2X2 AND2X2_9755 ( .A(u2__abc_44228_n19748), .B(u2__abc_44228_n19751), .Y(u2__abc_44228_n19752) );
  AND2X2 AND2X2_9756 ( .A(u2__abc_44228_n19753), .B(u2__abc_44228_n2966_bF_buf18), .Y(u2_root_165__FF_INPUT) );
  AND2X2 AND2X2_9757 ( .A(u2__abc_44228_n3062_bF_buf34), .B(sqrto_165_), .Y(u2__abc_44228_n19755) );
  AND2X2 AND2X2_9758 ( .A(u2__abc_44228_n19745), .B(sqrto_164_), .Y(u2__abc_44228_n19757) );
  AND2X2 AND2X2_9759 ( .A(u2__abc_44228_n19758), .B(u2__abc_44228_n19756), .Y(u2__abc_44228_n19759) );
  AND2X2 AND2X2_976 ( .A(u2__abc_44228_n3953), .B(u2_remHi_87_), .Y(u2__abc_44228_n3954) );
  AND2X2 AND2X2_9760 ( .A(u2__abc_44228_n2983_bF_buf2), .B(u2__abc_44228_n4958), .Y(u2__abc_44228_n19761) );
  AND2X2 AND2X2_9761 ( .A(u2__abc_44228_n19762), .B(u2__abc_44228_n2972_bF_buf22), .Y(u2__abc_44228_n19763) );
  AND2X2 AND2X2_9762 ( .A(u2__abc_44228_n19760), .B(u2__abc_44228_n19763), .Y(u2__abc_44228_n19764) );
  AND2X2 AND2X2_9763 ( .A(u2__abc_44228_n19765), .B(u2__abc_44228_n2966_bF_buf17), .Y(u2_root_166__FF_INPUT) );
  AND2X2 AND2X2_9764 ( .A(u2__abc_44228_n3062_bF_buf33), .B(sqrto_166_), .Y(u2__abc_44228_n19767) );
  AND2X2 AND2X2_9765 ( .A(u2__abc_44228_n19757), .B(sqrto_165_), .Y(u2__abc_44228_n19769) );
  AND2X2 AND2X2_9766 ( .A(u2__abc_44228_n19770), .B(u2__abc_44228_n19768), .Y(u2__abc_44228_n19771) );
  AND2X2 AND2X2_9767 ( .A(u2__abc_44228_n2983_bF_buf0), .B(u2__abc_44228_n4942), .Y(u2__abc_44228_n19773) );
  AND2X2 AND2X2_9768 ( .A(u2__abc_44228_n19774), .B(u2__abc_44228_n2972_bF_buf21), .Y(u2__abc_44228_n19775) );
  AND2X2 AND2X2_9769 ( .A(u2__abc_44228_n19772), .B(u2__abc_44228_n19775), .Y(u2__abc_44228_n19776) );
  AND2X2 AND2X2_977 ( .A(u2__abc_44228_n3956), .B(sqrto_87_), .Y(u2__abc_44228_n3957) );
  AND2X2 AND2X2_9770 ( .A(u2__abc_44228_n19777), .B(u2__abc_44228_n2966_bF_buf16), .Y(u2_root_167__FF_INPUT) );
  AND2X2 AND2X2_9771 ( .A(u2__abc_44228_n3062_bF_buf32), .B(sqrto_167_), .Y(u2__abc_44228_n19779) );
  AND2X2 AND2X2_9772 ( .A(u2__abc_44228_n19769), .B(sqrto_166_), .Y(u2__abc_44228_n19781) );
  AND2X2 AND2X2_9773 ( .A(u2__abc_44228_n19782), .B(u2__abc_44228_n19780), .Y(u2__abc_44228_n19783) );
  AND2X2 AND2X2_9774 ( .A(u2__abc_44228_n2983_bF_buf140), .B(u2__abc_44228_n4948_1), .Y(u2__abc_44228_n19785) );
  AND2X2 AND2X2_9775 ( .A(u2__abc_44228_n19786), .B(u2__abc_44228_n2972_bF_buf20), .Y(u2__abc_44228_n19787) );
  AND2X2 AND2X2_9776 ( .A(u2__abc_44228_n19784), .B(u2__abc_44228_n19787), .Y(u2__abc_44228_n19788) );
  AND2X2 AND2X2_9777 ( .A(u2__abc_44228_n19789), .B(u2__abc_44228_n2966_bF_buf15), .Y(u2_root_168__FF_INPUT) );
  AND2X2 AND2X2_9778 ( .A(u2__abc_44228_n3062_bF_buf31), .B(sqrto_168_), .Y(u2__abc_44228_n19791) );
  AND2X2 AND2X2_9779 ( .A(u2__abc_44228_n19781), .B(sqrto_167_), .Y(u2__abc_44228_n19793) );
  AND2X2 AND2X2_978 ( .A(u2__abc_44228_n3955), .B(u2__abc_44228_n3958_1), .Y(u2__abc_44228_n3959) );
  AND2X2 AND2X2_9780 ( .A(u2__abc_44228_n19794), .B(u2__abc_44228_n19792), .Y(u2__abc_44228_n19795) );
  AND2X2 AND2X2_9781 ( .A(u2__abc_44228_n2983_bF_buf138), .B(u2__abc_44228_n4935), .Y(u2__abc_44228_n19797) );
  AND2X2 AND2X2_9782 ( .A(u2__abc_44228_n19798), .B(u2__abc_44228_n2972_bF_buf19), .Y(u2__abc_44228_n19799) );
  AND2X2 AND2X2_9783 ( .A(u2__abc_44228_n19796), .B(u2__abc_44228_n19799), .Y(u2__abc_44228_n19800) );
  AND2X2 AND2X2_9784 ( .A(u2__abc_44228_n19801), .B(u2__abc_44228_n2966_bF_buf14), .Y(u2_root_169__FF_INPUT) );
  AND2X2 AND2X2_9785 ( .A(u2__abc_44228_n3062_bF_buf30), .B(sqrto_169_), .Y(u2__abc_44228_n19803) );
  AND2X2 AND2X2_9786 ( .A(u2__abc_44228_n19793), .B(sqrto_168_), .Y(u2__abc_44228_n19805) );
  AND2X2 AND2X2_9787 ( .A(u2__abc_44228_n19806), .B(u2__abc_44228_n19804), .Y(u2__abc_44228_n19807) );
  AND2X2 AND2X2_9788 ( .A(u2__abc_44228_n2983_bF_buf136), .B(u2__abc_44228_n4928), .Y(u2__abc_44228_n19809) );
  AND2X2 AND2X2_9789 ( .A(u2__abc_44228_n19810), .B(u2__abc_44228_n2972_bF_buf18), .Y(u2__abc_44228_n19811) );
  AND2X2 AND2X2_979 ( .A(u2__abc_44228_n3952), .B(u2__abc_44228_n3959), .Y(u2__abc_44228_n3960) );
  AND2X2 AND2X2_9790 ( .A(u2__abc_44228_n19808), .B(u2__abc_44228_n19811), .Y(u2__abc_44228_n19812) );
  AND2X2 AND2X2_9791 ( .A(u2__abc_44228_n19813), .B(u2__abc_44228_n2966_bF_buf13), .Y(u2_root_170__FF_INPUT) );
  AND2X2 AND2X2_9792 ( .A(u2__abc_44228_n3062_bF_buf29), .B(sqrto_170_), .Y(u2__abc_44228_n19815) );
  AND2X2 AND2X2_9793 ( .A(u2__abc_44228_n19805), .B(sqrto_169_), .Y(u2__abc_44228_n19817) );
  AND2X2 AND2X2_9794 ( .A(u2__abc_44228_n19818), .B(u2__abc_44228_n19816), .Y(u2__abc_44228_n19819) );
  AND2X2 AND2X2_9795 ( .A(u2__abc_44228_n2983_bF_buf134), .B(u2__abc_44228_n4913), .Y(u2__abc_44228_n19821) );
  AND2X2 AND2X2_9796 ( .A(u2__abc_44228_n19822), .B(u2__abc_44228_n2972_bF_buf17), .Y(u2__abc_44228_n19823) );
  AND2X2 AND2X2_9797 ( .A(u2__abc_44228_n19820), .B(u2__abc_44228_n19823), .Y(u2__abc_44228_n19824) );
  AND2X2 AND2X2_9798 ( .A(u2__abc_44228_n19825), .B(u2__abc_44228_n2966_bF_buf12), .Y(u2_root_171__FF_INPUT) );
  AND2X2 AND2X2_9799 ( .A(u2__abc_44228_n3062_bF_buf28), .B(sqrto_171_), .Y(u2__abc_44228_n19827) );
  AND2X2 AND2X2_98 ( .A(_abc_64468_n894), .B(_abc_64468_n893), .Y(_auto_iopadmap_cc_313_execute_65414_133_) );
  AND2X2 AND2X2_980 ( .A(u2__abc_44228_n3946), .B(u2__abc_44228_n3960), .Y(u2__abc_44228_n3961) );
  AND2X2 AND2X2_9800 ( .A(u2__abc_44228_n19817), .B(sqrto_170_), .Y(u2__abc_44228_n19829) );
  AND2X2 AND2X2_9801 ( .A(u2__abc_44228_n19830), .B(u2__abc_44228_n19828), .Y(u2__abc_44228_n19831) );
  AND2X2 AND2X2_9802 ( .A(u2__abc_44228_n2983_bF_buf132), .B(u2__abc_44228_n4919), .Y(u2__abc_44228_n19833) );
  AND2X2 AND2X2_9803 ( .A(u2__abc_44228_n19834), .B(u2__abc_44228_n2972_bF_buf16), .Y(u2__abc_44228_n19835) );
  AND2X2 AND2X2_9804 ( .A(u2__abc_44228_n19832), .B(u2__abc_44228_n19835), .Y(u2__abc_44228_n19836) );
  AND2X2 AND2X2_9805 ( .A(u2__abc_44228_n19837), .B(u2__abc_44228_n2966_bF_buf11), .Y(u2_root_172__FF_INPUT) );
  AND2X2 AND2X2_9806 ( .A(u2__abc_44228_n3062_bF_buf27), .B(sqrto_172_), .Y(u2__abc_44228_n19839) );
  AND2X2 AND2X2_9807 ( .A(u2__abc_44228_n19829), .B(sqrto_171_), .Y(u2__abc_44228_n19841) );
  AND2X2 AND2X2_9808 ( .A(u2__abc_44228_n19842), .B(u2__abc_44228_n19840), .Y(u2__abc_44228_n19843) );
  AND2X2 AND2X2_9809 ( .A(u2__abc_44228_n2983_bF_buf130), .B(u2__abc_44228_n4906), .Y(u2__abc_44228_n19845) );
  AND2X2 AND2X2_981 ( .A(u2__abc_44228_n3932), .B(u2__abc_44228_n3961), .Y(u2__abc_44228_n3962) );
  AND2X2 AND2X2_9810 ( .A(u2__abc_44228_n19846), .B(u2__abc_44228_n2972_bF_buf15), .Y(u2__abc_44228_n19847) );
  AND2X2 AND2X2_9811 ( .A(u2__abc_44228_n19844), .B(u2__abc_44228_n19847), .Y(u2__abc_44228_n19848) );
  AND2X2 AND2X2_9812 ( .A(u2__abc_44228_n19849), .B(u2__abc_44228_n2966_bF_buf10), .Y(u2_root_173__FF_INPUT) );
  AND2X2 AND2X2_9813 ( .A(u2__abc_44228_n3062_bF_buf26), .B(sqrto_173_), .Y(u2__abc_44228_n19851) );
  AND2X2 AND2X2_9814 ( .A(u2__abc_44228_n19841), .B(sqrto_172_), .Y(u2__abc_44228_n19853) );
  AND2X2 AND2X2_9815 ( .A(u2__abc_44228_n19854), .B(u2__abc_44228_n19852), .Y(u2__abc_44228_n19855) );
  AND2X2 AND2X2_9816 ( .A(u2__abc_44228_n2983_bF_buf128), .B(u2__abc_44228_n4899), .Y(u2__abc_44228_n19857) );
  AND2X2 AND2X2_9817 ( .A(u2__abc_44228_n19858), .B(u2__abc_44228_n2972_bF_buf14), .Y(u2__abc_44228_n19859) );
  AND2X2 AND2X2_9818 ( .A(u2__abc_44228_n19856), .B(u2__abc_44228_n19859), .Y(u2__abc_44228_n19860) );
  AND2X2 AND2X2_9819 ( .A(u2__abc_44228_n19861), .B(u2__abc_44228_n2966_bF_buf9), .Y(u2_root_174__FF_INPUT) );
  AND2X2 AND2X2_982 ( .A(u2__abc_44228_n3963), .B(u2_remHi_85_), .Y(u2__abc_44228_n3964) );
  AND2X2 AND2X2_9820 ( .A(u2__abc_44228_n3062_bF_buf25), .B(sqrto_174_), .Y(u2__abc_44228_n19863) );
  AND2X2 AND2X2_9821 ( .A(u2__abc_44228_n19853), .B(sqrto_173_), .Y(u2__abc_44228_n19865) );
  AND2X2 AND2X2_9822 ( .A(u2__abc_44228_n19866), .B(u2__abc_44228_n19864), .Y(u2__abc_44228_n19867) );
  AND2X2 AND2X2_9823 ( .A(u2__abc_44228_n2983_bF_buf126), .B(u2__abc_44228_n4889), .Y(u2__abc_44228_n19869) );
  AND2X2 AND2X2_9824 ( .A(u2__abc_44228_n19870), .B(u2__abc_44228_n2972_bF_buf13), .Y(u2__abc_44228_n19871) );
  AND2X2 AND2X2_9825 ( .A(u2__abc_44228_n19868), .B(u2__abc_44228_n19871), .Y(u2__abc_44228_n19872) );
  AND2X2 AND2X2_9826 ( .A(u2__abc_44228_n19873), .B(u2__abc_44228_n2966_bF_buf8), .Y(u2_root_175__FF_INPUT) );
  AND2X2 AND2X2_9827 ( .A(u2__abc_44228_n3062_bF_buf24), .B(sqrto_175_), .Y(u2__abc_44228_n19875) );
  AND2X2 AND2X2_9828 ( .A(u2__abc_44228_n19865), .B(sqrto_174_), .Y(u2__abc_44228_n19877) );
  AND2X2 AND2X2_9829 ( .A(u2__abc_44228_n19878), .B(u2__abc_44228_n19876), .Y(u2__abc_44228_n19879) );
  AND2X2 AND2X2_983 ( .A(u2__abc_44228_n3966), .B(sqrto_85_), .Y(u2__abc_44228_n3967_1) );
  AND2X2 AND2X2_9830 ( .A(u2__abc_44228_n2983_bF_buf124), .B(u2__abc_44228_n4882_1), .Y(u2__abc_44228_n19881) );
  AND2X2 AND2X2_9831 ( .A(u2__abc_44228_n19882), .B(u2__abc_44228_n2972_bF_buf12), .Y(u2__abc_44228_n19883) );
  AND2X2 AND2X2_9832 ( .A(u2__abc_44228_n19880), .B(u2__abc_44228_n19883), .Y(u2__abc_44228_n19884) );
  AND2X2 AND2X2_9833 ( .A(u2__abc_44228_n19885), .B(u2__abc_44228_n2966_bF_buf7), .Y(u2_root_176__FF_INPUT) );
  AND2X2 AND2X2_9834 ( .A(u2__abc_44228_n3062_bF_buf23), .B(sqrto_176_), .Y(u2__abc_44228_n19887) );
  AND2X2 AND2X2_9835 ( .A(u2__abc_44228_n19877), .B(sqrto_175_), .Y(u2__abc_44228_n19889) );
  AND2X2 AND2X2_9836 ( .A(u2__abc_44228_n19890), .B(u2__abc_44228_n19888), .Y(u2__abc_44228_n19891) );
  AND2X2 AND2X2_9837 ( .A(u2__abc_44228_n2983_bF_buf122), .B(u2__abc_44228_n4875), .Y(u2__abc_44228_n19893) );
  AND2X2 AND2X2_9838 ( .A(u2__abc_44228_n19894), .B(u2__abc_44228_n2972_bF_buf11), .Y(u2__abc_44228_n19895) );
  AND2X2 AND2X2_9839 ( .A(u2__abc_44228_n19892), .B(u2__abc_44228_n19895), .Y(u2__abc_44228_n19896) );
  AND2X2 AND2X2_984 ( .A(u2__abc_44228_n3965), .B(u2__abc_44228_n3968), .Y(u2__abc_44228_n3969) );
  AND2X2 AND2X2_9840 ( .A(u2__abc_44228_n19897), .B(u2__abc_44228_n2966_bF_buf6), .Y(u2_root_177__FF_INPUT) );
  AND2X2 AND2X2_9841 ( .A(u2__abc_44228_n3062_bF_buf22), .B(sqrto_177_), .Y(u2__abc_44228_n19899) );
  AND2X2 AND2X2_9842 ( .A(u2__abc_44228_n19889), .B(sqrto_176_), .Y(u2__abc_44228_n19901) );
  AND2X2 AND2X2_9843 ( .A(u2__abc_44228_n19902), .B(u2__abc_44228_n19900), .Y(u2__abc_44228_n19903) );
  AND2X2 AND2X2_9844 ( .A(u2__abc_44228_n2983_bF_buf120), .B(u2__abc_44228_n4868), .Y(u2__abc_44228_n19905) );
  AND2X2 AND2X2_9845 ( .A(u2__abc_44228_n19906), .B(u2__abc_44228_n2972_bF_buf10), .Y(u2__abc_44228_n19907) );
  AND2X2 AND2X2_9846 ( .A(u2__abc_44228_n19904), .B(u2__abc_44228_n19907), .Y(u2__abc_44228_n19908) );
  AND2X2 AND2X2_9847 ( .A(u2__abc_44228_n19909), .B(u2__abc_44228_n2966_bF_buf5), .Y(u2_root_178__FF_INPUT) );
  AND2X2 AND2X2_9848 ( .A(u2__abc_44228_n3062_bF_buf21), .B(sqrto_178_), .Y(u2__abc_44228_n19911) );
  AND2X2 AND2X2_9849 ( .A(u2__abc_44228_n19901), .B(sqrto_177_), .Y(u2__abc_44228_n19913) );
  AND2X2 AND2X2_985 ( .A(u2__abc_44228_n3970), .B(u2_remHi_84_), .Y(u2__abc_44228_n3971) );
  AND2X2 AND2X2_9850 ( .A(u2__abc_44228_n19914), .B(u2__abc_44228_n19912), .Y(u2__abc_44228_n19915) );
  AND2X2 AND2X2_9851 ( .A(u2__abc_44228_n2983_bF_buf118), .B(u2__abc_44228_n4860), .Y(u2__abc_44228_n19917) );
  AND2X2 AND2X2_9852 ( .A(u2__abc_44228_n19918), .B(u2__abc_44228_n2972_bF_buf9), .Y(u2__abc_44228_n19919) );
  AND2X2 AND2X2_9853 ( .A(u2__abc_44228_n19916), .B(u2__abc_44228_n19919), .Y(u2__abc_44228_n19920) );
  AND2X2 AND2X2_9854 ( .A(u2__abc_44228_n19921), .B(u2__abc_44228_n2966_bF_buf4), .Y(u2_root_179__FF_INPUT) );
  AND2X2 AND2X2_9855 ( .A(u2__abc_44228_n3062_bF_buf20), .B(sqrto_179_), .Y(u2__abc_44228_n19923) );
  AND2X2 AND2X2_9856 ( .A(u2__abc_44228_n19913), .B(sqrto_178_), .Y(u2__abc_44228_n19925) );
  AND2X2 AND2X2_9857 ( .A(u2__abc_44228_n19926), .B(u2__abc_44228_n19924), .Y(u2__abc_44228_n19927) );
  AND2X2 AND2X2_9858 ( .A(u2__abc_44228_n2983_bF_buf116), .B(u2__abc_44228_n4853), .Y(u2__abc_44228_n19929) );
  AND2X2 AND2X2_9859 ( .A(u2__abc_44228_n19930), .B(u2__abc_44228_n2972_bF_buf8), .Y(u2__abc_44228_n19931) );
  AND2X2 AND2X2_986 ( .A(u2__abc_44228_n3972), .B(sqrto_84_), .Y(u2__abc_44228_n3973) );
  AND2X2 AND2X2_9860 ( .A(u2__abc_44228_n19928), .B(u2__abc_44228_n19931), .Y(u2__abc_44228_n19932) );
  AND2X2 AND2X2_9861 ( .A(u2__abc_44228_n19933), .B(u2__abc_44228_n2966_bF_buf3), .Y(u2_root_180__FF_INPUT) );
  AND2X2 AND2X2_9862 ( .A(u2__abc_44228_n3062_bF_buf19), .B(sqrto_180_), .Y(u2__abc_44228_n19935) );
  AND2X2 AND2X2_9863 ( .A(u2__abc_44228_n19925), .B(sqrto_179_), .Y(u2__abc_44228_n19937) );
  AND2X2 AND2X2_9864 ( .A(u2__abc_44228_n19938), .B(u2__abc_44228_n19936), .Y(u2__abc_44228_n19939) );
  AND2X2 AND2X2_9865 ( .A(u2__abc_44228_n2983_bF_buf114), .B(u2__abc_44228_n4846_1), .Y(u2__abc_44228_n19941) );
  AND2X2 AND2X2_9866 ( .A(u2__abc_44228_n19942), .B(u2__abc_44228_n2972_bF_buf7), .Y(u2__abc_44228_n19943) );
  AND2X2 AND2X2_9867 ( .A(u2__abc_44228_n19940), .B(u2__abc_44228_n19943), .Y(u2__abc_44228_n19944) );
  AND2X2 AND2X2_9868 ( .A(u2__abc_44228_n19945), .B(u2__abc_44228_n2966_bF_buf2), .Y(u2_root_181__FF_INPUT) );
  AND2X2 AND2X2_9869 ( .A(u2__abc_44228_n3062_bF_buf18), .B(sqrto_181_), .Y(u2__abc_44228_n19947) );
  AND2X2 AND2X2_987 ( .A(u2__abc_44228_n3975), .B(u2__abc_44228_n3969), .Y(u2__abc_44228_n3976_1) );
  AND2X2 AND2X2_9870 ( .A(u2__abc_44228_n19937), .B(sqrto_180_), .Y(u2__abc_44228_n19949) );
  AND2X2 AND2X2_9871 ( .A(u2__abc_44228_n19950), .B(u2__abc_44228_n19948), .Y(u2__abc_44228_n19951) );
  AND2X2 AND2X2_9872 ( .A(u2__abc_44228_n2983_bF_buf112), .B(u2__abc_44228_n4839), .Y(u2__abc_44228_n19953) );
  AND2X2 AND2X2_9873 ( .A(u2__abc_44228_n19954), .B(u2__abc_44228_n2972_bF_buf6), .Y(u2__abc_44228_n19955) );
  AND2X2 AND2X2_9874 ( .A(u2__abc_44228_n19952), .B(u2__abc_44228_n19955), .Y(u2__abc_44228_n19956) );
  AND2X2 AND2X2_9875 ( .A(u2__abc_44228_n19957), .B(u2__abc_44228_n2966_bF_buf1), .Y(u2_root_182__FF_INPUT) );
  AND2X2 AND2X2_9876 ( .A(u2__abc_44228_n3062_bF_buf17), .B(sqrto_182_), .Y(u2__abc_44228_n19959) );
  AND2X2 AND2X2_9877 ( .A(u2__abc_44228_n19949), .B(sqrto_181_), .Y(u2__abc_44228_n19961) );
  AND2X2 AND2X2_9878 ( .A(u2__abc_44228_n19962), .B(u2__abc_44228_n19960), .Y(u2__abc_44228_n19963) );
  AND2X2 AND2X2_9879 ( .A(u2__abc_44228_n2983_bF_buf110), .B(u2__abc_44228_n4816), .Y(u2__abc_44228_n19965) );
  AND2X2 AND2X2_988 ( .A(u2__abc_44228_n3977), .B(u2_remHi_82_), .Y(u2__abc_44228_n3978) );
  AND2X2 AND2X2_9880 ( .A(u2__abc_44228_n19966), .B(u2__abc_44228_n2972_bF_buf5), .Y(u2__abc_44228_n19967) );
  AND2X2 AND2X2_9881 ( .A(u2__abc_44228_n19964), .B(u2__abc_44228_n19967), .Y(u2__abc_44228_n19968) );
  AND2X2 AND2X2_9882 ( .A(u2__abc_44228_n19969), .B(u2__abc_44228_n2966_bF_buf0), .Y(u2_root_183__FF_INPUT) );
  AND2X2 AND2X2_9883 ( .A(u2__abc_44228_n3062_bF_buf16), .B(sqrto_183_), .Y(u2__abc_44228_n19971) );
  AND2X2 AND2X2_9884 ( .A(u2__abc_44228_n19961), .B(sqrto_182_), .Y(u2__abc_44228_n19973) );
  AND2X2 AND2X2_9885 ( .A(u2__abc_44228_n19974), .B(u2__abc_44228_n19972), .Y(u2__abc_44228_n19975) );
  AND2X2 AND2X2_9886 ( .A(u2__abc_44228_n2983_bF_buf108), .B(u2__abc_44228_n4809_1), .Y(u2__abc_44228_n19977) );
  AND2X2 AND2X2_9887 ( .A(u2__abc_44228_n19978), .B(u2__abc_44228_n2972_bF_buf4), .Y(u2__abc_44228_n19979) );
  AND2X2 AND2X2_9888 ( .A(u2__abc_44228_n19976), .B(u2__abc_44228_n19979), .Y(u2__abc_44228_n19980) );
  AND2X2 AND2X2_9889 ( .A(u2__abc_44228_n19981), .B(u2__abc_44228_n2966_bF_buf107), .Y(u2_root_184__FF_INPUT) );
  AND2X2 AND2X2_989 ( .A(u2__abc_44228_n3979), .B(sqrto_82_), .Y(u2__abc_44228_n3980) );
  AND2X2 AND2X2_9890 ( .A(u2__abc_44228_n3062_bF_buf15), .B(sqrto_184_), .Y(u2__abc_44228_n19983) );
  AND2X2 AND2X2_9891 ( .A(u2__abc_44228_n19973), .B(sqrto_183_), .Y(u2__abc_44228_n19985) );
  AND2X2 AND2X2_9892 ( .A(u2__abc_44228_n19986), .B(u2__abc_44228_n19984), .Y(u2__abc_44228_n19987) );
  AND2X2 AND2X2_9893 ( .A(u2__abc_44228_n2983_bF_buf106), .B(u2__abc_44228_n4830), .Y(u2__abc_44228_n19989) );
  AND2X2 AND2X2_9894 ( .A(u2__abc_44228_n19990), .B(u2__abc_44228_n2972_bF_buf3), .Y(u2__abc_44228_n19991) );
  AND2X2 AND2X2_9895 ( .A(u2__abc_44228_n19988), .B(u2__abc_44228_n19991), .Y(u2__abc_44228_n19992) );
  AND2X2 AND2X2_9896 ( .A(u2__abc_44228_n19993), .B(u2__abc_44228_n2966_bF_buf106), .Y(u2_root_185__FF_INPUT) );
  AND2X2 AND2X2_9897 ( .A(u2__abc_44228_n3062_bF_buf14), .B(sqrto_185_), .Y(u2__abc_44228_n19995) );
  AND2X2 AND2X2_9898 ( .A(u2__abc_44228_n19985), .B(sqrto_184_), .Y(u2__abc_44228_n19997) );
  AND2X2 AND2X2_9899 ( .A(u2__abc_44228_n19998), .B(u2__abc_44228_n19996), .Y(u2__abc_44228_n19999) );
  AND2X2 AND2X2_99 ( .A(_abc_64468_n897), .B(_abc_64468_n896), .Y(_auto_iopadmap_cc_313_execute_65414_134_) );
  AND2X2 AND2X2_990 ( .A(u2__abc_44228_n3983), .B(u2_remHi_83_), .Y(u2__abc_44228_n3984) );
  AND2X2 AND2X2_9900 ( .A(u2__abc_44228_n2983_bF_buf104), .B(u2__abc_44228_n4823), .Y(u2__abc_44228_n20001) );
  AND2X2 AND2X2_9901 ( .A(u2__abc_44228_n20002), .B(u2__abc_44228_n2972_bF_buf2), .Y(u2__abc_44228_n20003) );
  AND2X2 AND2X2_9902 ( .A(u2__abc_44228_n20000), .B(u2__abc_44228_n20003), .Y(u2__abc_44228_n20004) );
  AND2X2 AND2X2_9903 ( .A(u2__abc_44228_n20005), .B(u2__abc_44228_n2966_bF_buf105), .Y(u2_root_186__FF_INPUT) );
  AND2X2 AND2X2_9904 ( .A(u2__abc_44228_n3062_bF_buf13), .B(sqrto_186_), .Y(u2__abc_44228_n20007) );
  AND2X2 AND2X2_9905 ( .A(u2__abc_44228_n19997), .B(sqrto_185_), .Y(u2__abc_44228_n20009) );
  AND2X2 AND2X2_9906 ( .A(u2__abc_44228_n20010), .B(u2__abc_44228_n20008), .Y(u2__abc_44228_n20011) );
  AND2X2 AND2X2_9907 ( .A(u2__abc_44228_n2983_bF_buf102), .B(u2__abc_44228_n4801), .Y(u2__abc_44228_n20013) );
  AND2X2 AND2X2_9908 ( .A(u2__abc_44228_n20014), .B(u2__abc_44228_n2972_bF_buf1), .Y(u2__abc_44228_n20015) );
  AND2X2 AND2X2_9909 ( .A(u2__abc_44228_n20012), .B(u2__abc_44228_n20015), .Y(u2__abc_44228_n20016) );
  AND2X2 AND2X2_991 ( .A(u2__abc_44228_n3986_1), .B(sqrto_83_), .Y(u2__abc_44228_n3987) );
  AND2X2 AND2X2_9910 ( .A(u2__abc_44228_n20017), .B(u2__abc_44228_n2966_bF_buf104), .Y(u2_root_187__FF_INPUT) );
  AND2X2 AND2X2_9911 ( .A(u2__abc_44228_n3062_bF_buf12), .B(sqrto_187_), .Y(u2__abc_44228_n20019) );
  AND2X2 AND2X2_9912 ( .A(u2__abc_44228_n20009), .B(sqrto_186_), .Y(u2__abc_44228_n20021) );
  AND2X2 AND2X2_9913 ( .A(u2__abc_44228_n20022), .B(u2__abc_44228_n20020), .Y(u2__abc_44228_n20023) );
  AND2X2 AND2X2_9914 ( .A(u2__abc_44228_n2983_bF_buf100), .B(u2__abc_44228_n4794), .Y(u2__abc_44228_n20025) );
  AND2X2 AND2X2_9915 ( .A(u2__abc_44228_n20026), .B(u2__abc_44228_n2972_bF_buf0), .Y(u2__abc_44228_n20027) );
  AND2X2 AND2X2_9916 ( .A(u2__abc_44228_n20024), .B(u2__abc_44228_n20027), .Y(u2__abc_44228_n20028) );
  AND2X2 AND2X2_9917 ( .A(u2__abc_44228_n20029), .B(u2__abc_44228_n2966_bF_buf103), .Y(u2_root_188__FF_INPUT) );
  AND2X2 AND2X2_9918 ( .A(u2__abc_44228_n3062_bF_buf11), .B(sqrto_188_), .Y(u2__abc_44228_n20031) );
  AND2X2 AND2X2_9919 ( .A(u2__abc_44228_n20021), .B(sqrto_187_), .Y(u2__abc_44228_n20033) );
  AND2X2 AND2X2_992 ( .A(u2__abc_44228_n3985), .B(u2__abc_44228_n3988), .Y(u2__abc_44228_n3989) );
  AND2X2 AND2X2_9920 ( .A(u2__abc_44228_n20034), .B(u2__abc_44228_n20032), .Y(u2__abc_44228_n20035) );
  AND2X2 AND2X2_9921 ( .A(u2__abc_44228_n2983_bF_buf98), .B(u2__abc_44228_n4787), .Y(u2__abc_44228_n20037) );
  AND2X2 AND2X2_9922 ( .A(u2__abc_44228_n20038), .B(u2__abc_44228_n2972_bF_buf107), .Y(u2__abc_44228_n20039) );
  AND2X2 AND2X2_9923 ( .A(u2__abc_44228_n20036), .B(u2__abc_44228_n20039), .Y(u2__abc_44228_n20040) );
  AND2X2 AND2X2_9924 ( .A(u2__abc_44228_n20041), .B(u2__abc_44228_n2966_bF_buf102), .Y(u2_root_189__FF_INPUT) );
  AND2X2 AND2X2_9925 ( .A(u2__abc_44228_n3062_bF_buf10), .B(sqrto_189_), .Y(u2__abc_44228_n20043) );
  AND2X2 AND2X2_9926 ( .A(u2__abc_44228_n20033), .B(sqrto_188_), .Y(u2__abc_44228_n20045) );
  AND2X2 AND2X2_9927 ( .A(u2__abc_44228_n20046), .B(u2__abc_44228_n20044), .Y(u2__abc_44228_n20047) );
  AND2X2 AND2X2_9928 ( .A(u2__abc_44228_n2983_bF_buf96), .B(u2__abc_44228_n4780), .Y(u2__abc_44228_n20049) );
  AND2X2 AND2X2_9929 ( .A(u2__abc_44228_n20050), .B(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n20051) );
  AND2X2 AND2X2_993 ( .A(u2__abc_44228_n3982), .B(u2__abc_44228_n3989), .Y(u2__abc_44228_n3990) );
  AND2X2 AND2X2_9930 ( .A(u2__abc_44228_n20048), .B(u2__abc_44228_n20051), .Y(u2__abc_44228_n20052) );
  AND2X2 AND2X2_9931 ( .A(u2__abc_44228_n20053), .B(u2__abc_44228_n2966_bF_buf101), .Y(u2_root_190__FF_INPUT) );
  AND2X2 AND2X2_9932 ( .A(u2__abc_44228_n3062_bF_buf9), .B(sqrto_190_), .Y(u2__abc_44228_n20055) );
  AND2X2 AND2X2_9933 ( .A(u2__abc_44228_n20045), .B(sqrto_189_), .Y(u2__abc_44228_n20057) );
  AND2X2 AND2X2_9934 ( .A(u2__abc_44228_n20058), .B(u2__abc_44228_n20056), .Y(u2__abc_44228_n20059) );
  AND2X2 AND2X2_9935 ( .A(u2__abc_44228_n2983_bF_buf94), .B(u2__abc_44228_n4761), .Y(u2__abc_44228_n20061) );
  AND2X2 AND2X2_9936 ( .A(u2__abc_44228_n20062), .B(u2__abc_44228_n2972_bF_buf105), .Y(u2__abc_44228_n20063) );
  AND2X2 AND2X2_9937 ( .A(u2__abc_44228_n20060), .B(u2__abc_44228_n20063), .Y(u2__abc_44228_n20064) );
  AND2X2 AND2X2_9938 ( .A(u2__abc_44228_n20065), .B(u2__abc_44228_n2966_bF_buf100), .Y(u2_root_191__FF_INPUT) );
  AND2X2 AND2X2_9939 ( .A(u2__abc_44228_n3062_bF_buf8), .B(sqrto_191_), .Y(u2__abc_44228_n20067) );
  AND2X2 AND2X2_994 ( .A(u2__abc_44228_n3976_1), .B(u2__abc_44228_n3990), .Y(u2__abc_44228_n3991) );
  AND2X2 AND2X2_9940 ( .A(u2__abc_44228_n20057), .B(sqrto_190_), .Y(u2__abc_44228_n20069) );
  AND2X2 AND2X2_9941 ( .A(u2__abc_44228_n20070), .B(u2__abc_44228_n20068), .Y(u2__abc_44228_n20071) );
  AND2X2 AND2X2_9942 ( .A(u2__abc_44228_n2983_bF_buf92), .B(u2__abc_44228_n4767), .Y(u2__abc_44228_n20073) );
  AND2X2 AND2X2_9943 ( .A(u2__abc_44228_n20074), .B(u2__abc_44228_n2972_bF_buf104), .Y(u2__abc_44228_n20075) );
  AND2X2 AND2X2_9944 ( .A(u2__abc_44228_n20072), .B(u2__abc_44228_n20075), .Y(u2__abc_44228_n20076) );
  AND2X2 AND2X2_9945 ( .A(u2__abc_44228_n20077), .B(u2__abc_44228_n2966_bF_buf99), .Y(u2_root_192__FF_INPUT) );
  AND2X2 AND2X2_9946 ( .A(u2__abc_44228_n3062_bF_buf7), .B(sqrto_192_), .Y(u2__abc_44228_n20079) );
  AND2X2 AND2X2_9947 ( .A(u2__abc_44228_n20069), .B(sqrto_191_), .Y(u2__abc_44228_n20081) );
  AND2X2 AND2X2_9948 ( .A(u2__abc_44228_n20082), .B(u2__abc_44228_n20080), .Y(u2__abc_44228_n20083) );
  AND2X2 AND2X2_9949 ( .A(u2__abc_44228_n2983_bF_buf90), .B(u2__abc_44228_n4754), .Y(u2__abc_44228_n20085) );
  AND2X2 AND2X2_995 ( .A(u2__abc_44228_n3992), .B(u2_remHi_81_), .Y(u2__abc_44228_n3993) );
  AND2X2 AND2X2_9950 ( .A(u2__abc_44228_n20086), .B(u2__abc_44228_n2972_bF_buf103), .Y(u2__abc_44228_n20087) );
  AND2X2 AND2X2_9951 ( .A(u2__abc_44228_n20084), .B(u2__abc_44228_n20087), .Y(u2__abc_44228_n20088) );
  AND2X2 AND2X2_9952 ( .A(u2__abc_44228_n20089), .B(u2__abc_44228_n2966_bF_buf98), .Y(u2_root_193__FF_INPUT) );
  AND2X2 AND2X2_9953 ( .A(u2__abc_44228_n3062_bF_buf6), .B(sqrto_193_), .Y(u2__abc_44228_n20091) );
  AND2X2 AND2X2_9954 ( .A(u2__abc_44228_n20081), .B(sqrto_192_), .Y(u2__abc_44228_n20093) );
  AND2X2 AND2X2_9955 ( .A(u2__abc_44228_n20094), .B(u2__abc_44228_n20092), .Y(u2__abc_44228_n20095) );
  AND2X2 AND2X2_9956 ( .A(u2__abc_44228_n2983_bF_buf88), .B(u2__abc_44228_n4747), .Y(u2__abc_44228_n20097) );
  AND2X2 AND2X2_9957 ( .A(u2__abc_44228_n20098), .B(u2__abc_44228_n2972_bF_buf102), .Y(u2__abc_44228_n20099) );
  AND2X2 AND2X2_9958 ( .A(u2__abc_44228_n20096), .B(u2__abc_44228_n20099), .Y(u2__abc_44228_n20100) );
  AND2X2 AND2X2_9959 ( .A(u2__abc_44228_n20101), .B(u2__abc_44228_n2966_bF_buf97), .Y(u2_root_194__FF_INPUT) );
  AND2X2 AND2X2_996 ( .A(u2__abc_44228_n3995_1), .B(sqrto_81_), .Y(u2__abc_44228_n3996) );
  AND2X2 AND2X2_9960 ( .A(u2__abc_44228_n3062_bF_buf5), .B(sqrto_194_), .Y(u2__abc_44228_n20103) );
  AND2X2 AND2X2_9961 ( .A(u2__abc_44228_n20093), .B(sqrto_193_), .Y(u2__abc_44228_n20105) );
  AND2X2 AND2X2_9962 ( .A(u2__abc_44228_n20106), .B(u2__abc_44228_n20104), .Y(u2__abc_44228_n20107) );
  AND2X2 AND2X2_9963 ( .A(u2__abc_44228_n2983_bF_buf86), .B(u2__abc_44228_n4739), .Y(u2__abc_44228_n20109) );
  AND2X2 AND2X2_9964 ( .A(u2__abc_44228_n20110), .B(u2__abc_44228_n2972_bF_buf101), .Y(u2__abc_44228_n20111) );
  AND2X2 AND2X2_9965 ( .A(u2__abc_44228_n20108), .B(u2__abc_44228_n20111), .Y(u2__abc_44228_n20112) );
  AND2X2 AND2X2_9966 ( .A(u2__abc_44228_n20113), .B(u2__abc_44228_n2966_bF_buf96), .Y(u2_root_195__FF_INPUT) );
  AND2X2 AND2X2_9967 ( .A(u2__abc_44228_n3062_bF_buf4), .B(sqrto_195_), .Y(u2__abc_44228_n20115) );
  AND2X2 AND2X2_9968 ( .A(u2__abc_44228_n20105), .B(sqrto_194_), .Y(u2__abc_44228_n20117) );
  AND2X2 AND2X2_9969 ( .A(u2__abc_44228_n20118), .B(u2__abc_44228_n20116), .Y(u2__abc_44228_n20119) );
  AND2X2 AND2X2_997 ( .A(u2__abc_44228_n3994), .B(u2__abc_44228_n3997), .Y(u2__abc_44228_n3998) );
  AND2X2 AND2X2_9970 ( .A(u2__abc_44228_n2983_bF_buf84), .B(u2__abc_44228_n4732), .Y(u2__abc_44228_n20121) );
  AND2X2 AND2X2_9971 ( .A(u2__abc_44228_n20122), .B(u2__abc_44228_n2972_bF_buf100), .Y(u2__abc_44228_n20123) );
  AND2X2 AND2X2_9972 ( .A(u2__abc_44228_n20120), .B(u2__abc_44228_n20123), .Y(u2__abc_44228_n20124) );
  AND2X2 AND2X2_9973 ( .A(u2__abc_44228_n20125), .B(u2__abc_44228_n2966_bF_buf95), .Y(u2_root_196__FF_INPUT) );
  AND2X2 AND2X2_9974 ( .A(u2__abc_44228_n3062_bF_buf3), .B(sqrto_196_), .Y(u2__abc_44228_n20127) );
  AND2X2 AND2X2_9975 ( .A(u2__abc_44228_n20117), .B(sqrto_195_), .Y(u2__abc_44228_n20129) );
  AND2X2 AND2X2_9976 ( .A(u2__abc_44228_n20130), .B(u2__abc_44228_n20128), .Y(u2__abc_44228_n20131) );
  AND2X2 AND2X2_9977 ( .A(u2__abc_44228_n2983_bF_buf82), .B(u2__abc_44228_n4725), .Y(u2__abc_44228_n20133) );
  AND2X2 AND2X2_9978 ( .A(u2__abc_44228_n20134), .B(u2__abc_44228_n2972_bF_buf99), .Y(u2__abc_44228_n20135) );
  AND2X2 AND2X2_9979 ( .A(u2__abc_44228_n20132), .B(u2__abc_44228_n20135), .Y(u2__abc_44228_n20136) );
  AND2X2 AND2X2_998 ( .A(u2__abc_44228_n3999), .B(u2_remHi_80_), .Y(u2__abc_44228_n4000) );
  AND2X2 AND2X2_9980 ( .A(u2__abc_44228_n20137), .B(u2__abc_44228_n2966_bF_buf94), .Y(u2_root_197__FF_INPUT) );
  AND2X2 AND2X2_9981 ( .A(u2__abc_44228_n3062_bF_buf2), .B(sqrto_197_), .Y(u2__abc_44228_n20139) );
  AND2X2 AND2X2_9982 ( .A(u2__abc_44228_n20129), .B(sqrto_196_), .Y(u2__abc_44228_n20141) );
  AND2X2 AND2X2_9983 ( .A(u2__abc_44228_n20142), .B(u2__abc_44228_n20140), .Y(u2__abc_44228_n20143) );
  AND2X2 AND2X2_9984 ( .A(u2__abc_44228_n2983_bF_buf80), .B(u2__abc_44228_n4718), .Y(u2__abc_44228_n20145) );
  AND2X2 AND2X2_9985 ( .A(u2__abc_44228_n20146), .B(u2__abc_44228_n2972_bF_buf98), .Y(u2__abc_44228_n20147) );
  AND2X2 AND2X2_9986 ( .A(u2__abc_44228_n20144), .B(u2__abc_44228_n20147), .Y(u2__abc_44228_n20148) );
  AND2X2 AND2X2_9987 ( .A(u2__abc_44228_n20149), .B(u2__abc_44228_n2966_bF_buf93), .Y(u2_root_198__FF_INPUT) );
  AND2X2 AND2X2_9988 ( .A(u2__abc_44228_n3062_bF_buf1), .B(sqrto_198_), .Y(u2__abc_44228_n20151) );
  AND2X2 AND2X2_9989 ( .A(u2__abc_44228_n20141), .B(sqrto_197_), .Y(u2__abc_44228_n20153) );
  AND2X2 AND2X2_999 ( .A(u2__abc_44228_n4001), .B(sqrto_80_), .Y(u2__abc_44228_n4002) );
  AND2X2 AND2X2_9990 ( .A(u2__abc_44228_n20154), .B(u2__abc_44228_n20152), .Y(u2__abc_44228_n20155) );
  AND2X2 AND2X2_9991 ( .A(u2__abc_44228_n2983_bF_buf78), .B(u2__abc_44228_n4702), .Y(u2__abc_44228_n20157) );
  AND2X2 AND2X2_9992 ( .A(u2__abc_44228_n20158), .B(u2__abc_44228_n2972_bF_buf97), .Y(u2__abc_44228_n20159) );
  AND2X2 AND2X2_9993 ( .A(u2__abc_44228_n20156), .B(u2__abc_44228_n20159), .Y(u2__abc_44228_n20160) );
  AND2X2 AND2X2_9994 ( .A(u2__abc_44228_n20161), .B(u2__abc_44228_n2966_bF_buf92), .Y(u2_root_199__FF_INPUT) );
  AND2X2 AND2X2_9995 ( .A(u2__abc_44228_n3062_bF_buf0), .B(sqrto_199_), .Y(u2__abc_44228_n20163) );
  AND2X2 AND2X2_9996 ( .A(u2__abc_44228_n20153), .B(sqrto_198_), .Y(u2__abc_44228_n20165) );
  AND2X2 AND2X2_9997 ( .A(u2__abc_44228_n20166), .B(u2__abc_44228_n20164), .Y(u2__abc_44228_n20167) );
  AND2X2 AND2X2_9998 ( .A(u2__abc_44228_n2983_bF_buf76), .B(u2__abc_44228_n4708), .Y(u2__abc_44228_n20169) );
  AND2X2 AND2X2_9999 ( .A(u2__abc_44228_n20170), .B(u2__abc_44228_n2972_bF_buf96), .Y(u2__abc_44228_n20171) );
  BUFX2 BUFX2_1 ( .A(u2__abc_44228_n7548_1), .Y(u2__abc_44228_n7548_1_hier0_bF_buf6) );
  BUFX2 BUFX2_10 ( .A(clk), .Y(clk_hier0_bF_buf8) );
  BUFX2 BUFX2_100 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf2) );
  BUFX2 BUFX2_1000 ( .A(_auto_iopadmap_cc_313_execute_65414_89_), .Y(\o[89] ) );
  BUFX2 BUFX2_1001 ( .A(_auto_iopadmap_cc_313_execute_65414_90_), .Y(\o[90] ) );
  BUFX2 BUFX2_1002 ( .A(_auto_iopadmap_cc_313_execute_65414_91_), .Y(\o[91] ) );
  BUFX2 BUFX2_1003 ( .A(_auto_iopadmap_cc_313_execute_65414_92_), .Y(\o[92] ) );
  BUFX2 BUFX2_1004 ( .A(_auto_iopadmap_cc_313_execute_65414_93_), .Y(\o[93] ) );
  BUFX2 BUFX2_1005 ( .A(_auto_iopadmap_cc_313_execute_65414_94_), .Y(\o[94] ) );
  BUFX2 BUFX2_1006 ( .A(_auto_iopadmap_cc_313_execute_65414_95_), .Y(\o[95] ) );
  BUFX2 BUFX2_1007 ( .A(_auto_iopadmap_cc_313_execute_65414_96_), .Y(\o[96] ) );
  BUFX2 BUFX2_1008 ( .A(_auto_iopadmap_cc_313_execute_65414_97_), .Y(\o[97] ) );
  BUFX2 BUFX2_1009 ( .A(_auto_iopadmap_cc_313_execute_65414_98_), .Y(\o[98] ) );
  BUFX2 BUFX2_101 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf1) );
  BUFX2 BUFX2_1010 ( .A(_auto_iopadmap_cc_313_execute_65414_99_), .Y(\o[99] ) );
  BUFX2 BUFX2_1011 ( .A(_auto_iopadmap_cc_313_execute_65414_100_), .Y(\o[100] ) );
  BUFX2 BUFX2_1012 ( .A(_auto_iopadmap_cc_313_execute_65414_101_), .Y(\o[101] ) );
  BUFX2 BUFX2_1013 ( .A(_auto_iopadmap_cc_313_execute_65414_102_), .Y(\o[102] ) );
  BUFX2 BUFX2_1014 ( .A(_auto_iopadmap_cc_313_execute_65414_103_), .Y(\o[103] ) );
  BUFX2 BUFX2_1015 ( .A(_auto_iopadmap_cc_313_execute_65414_104_), .Y(\o[104] ) );
  BUFX2 BUFX2_1016 ( .A(_auto_iopadmap_cc_313_execute_65414_105_), .Y(\o[105] ) );
  BUFX2 BUFX2_1017 ( .A(_auto_iopadmap_cc_313_execute_65414_106_), .Y(\o[106] ) );
  BUFX2 BUFX2_1018 ( .A(_auto_iopadmap_cc_313_execute_65414_107_), .Y(\o[107] ) );
  BUFX2 BUFX2_1019 ( .A(_auto_iopadmap_cc_313_execute_65414_108_), .Y(\o[108] ) );
  BUFX2 BUFX2_102 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf0) );
  BUFX2 BUFX2_1020 ( .A(_auto_iopadmap_cc_313_execute_65414_109_), .Y(\o[109] ) );
  BUFX2 BUFX2_1021 ( .A(_auto_iopadmap_cc_313_execute_65414_110_), .Y(\o[110] ) );
  BUFX2 BUFX2_1022 ( .A(_auto_iopadmap_cc_313_execute_65414_111_), .Y(\o[111] ) );
  BUFX2 BUFX2_1023 ( .A(_auto_iopadmap_cc_313_execute_65414_112_), .Y(\o[112] ) );
  BUFX2 BUFX2_1024 ( .A(_auto_iopadmap_cc_313_execute_65414_113_), .Y(\o[113] ) );
  BUFX2 BUFX2_1025 ( .A(_auto_iopadmap_cc_313_execute_65414_114_), .Y(\o[114] ) );
  BUFX2 BUFX2_1026 ( .A(_auto_iopadmap_cc_313_execute_65414_115_), .Y(\o[115] ) );
  BUFX2 BUFX2_1027 ( .A(_auto_iopadmap_cc_313_execute_65414_116_), .Y(\o[116] ) );
  BUFX2 BUFX2_1028 ( .A(_auto_iopadmap_cc_313_execute_65414_117_), .Y(\o[117] ) );
  BUFX2 BUFX2_1029 ( .A(_auto_iopadmap_cc_313_execute_65414_118_), .Y(\o[118] ) );
  BUFX2 BUFX2_103 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf57) );
  BUFX2 BUFX2_1030 ( .A(_auto_iopadmap_cc_313_execute_65414_119_), .Y(\o[119] ) );
  BUFX2 BUFX2_1031 ( .A(_auto_iopadmap_cc_313_execute_65414_120_), .Y(\o[120] ) );
  BUFX2 BUFX2_1032 ( .A(_auto_iopadmap_cc_313_execute_65414_121_), .Y(\o[121] ) );
  BUFX2 BUFX2_1033 ( .A(_auto_iopadmap_cc_313_execute_65414_122_), .Y(\o[122] ) );
  BUFX2 BUFX2_1034 ( .A(_auto_iopadmap_cc_313_execute_65414_123_), .Y(\o[123] ) );
  BUFX2 BUFX2_1035 ( .A(_auto_iopadmap_cc_313_execute_65414_124_), .Y(\o[124] ) );
  BUFX2 BUFX2_1036 ( .A(_auto_iopadmap_cc_313_execute_65414_125_), .Y(\o[125] ) );
  BUFX2 BUFX2_1037 ( .A(_auto_iopadmap_cc_313_execute_65414_126_), .Y(\o[126] ) );
  BUFX2 BUFX2_1038 ( .A(_auto_iopadmap_cc_313_execute_65414_127_), .Y(\o[127] ) );
  BUFX2 BUFX2_1039 ( .A(_auto_iopadmap_cc_313_execute_65414_128_), .Y(\o[128] ) );
  BUFX2 BUFX2_104 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf56) );
  BUFX2 BUFX2_1040 ( .A(_auto_iopadmap_cc_313_execute_65414_129_), .Y(\o[129] ) );
  BUFX2 BUFX2_1041 ( .A(_auto_iopadmap_cc_313_execute_65414_130_), .Y(\o[130] ) );
  BUFX2 BUFX2_1042 ( .A(_auto_iopadmap_cc_313_execute_65414_131_), .Y(\o[131] ) );
  BUFX2 BUFX2_1043 ( .A(_auto_iopadmap_cc_313_execute_65414_132_), .Y(\o[132] ) );
  BUFX2 BUFX2_1044 ( .A(_auto_iopadmap_cc_313_execute_65414_133_), .Y(\o[133] ) );
  BUFX2 BUFX2_1045 ( .A(_auto_iopadmap_cc_313_execute_65414_134_), .Y(\o[134] ) );
  BUFX2 BUFX2_1046 ( .A(_auto_iopadmap_cc_313_execute_65414_135_), .Y(\o[135] ) );
  BUFX2 BUFX2_1047 ( .A(_auto_iopadmap_cc_313_execute_65414_136_), .Y(\o[136] ) );
  BUFX2 BUFX2_1048 ( .A(_auto_iopadmap_cc_313_execute_65414_137_), .Y(\o[137] ) );
  BUFX2 BUFX2_1049 ( .A(_auto_iopadmap_cc_313_execute_65414_138_), .Y(\o[138] ) );
  BUFX2 BUFX2_105 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf4), .Y(u2__abc_44228_n7548_1_bF_buf55) );
  BUFX2 BUFX2_1050 ( .A(_auto_iopadmap_cc_313_execute_65414_139_), .Y(\o[139] ) );
  BUFX2 BUFX2_1051 ( .A(_auto_iopadmap_cc_313_execute_65414_140_), .Y(\o[140] ) );
  BUFX2 BUFX2_1052 ( .A(_auto_iopadmap_cc_313_execute_65414_141_), .Y(\o[141] ) );
  BUFX2 BUFX2_1053 ( .A(_auto_iopadmap_cc_313_execute_65414_142_), .Y(\o[142] ) );
  BUFX2 BUFX2_1054 ( .A(_auto_iopadmap_cc_313_execute_65414_143_), .Y(\o[143] ) );
  BUFX2 BUFX2_1055 ( .A(_auto_iopadmap_cc_313_execute_65414_144_), .Y(\o[144] ) );
  BUFX2 BUFX2_1056 ( .A(_auto_iopadmap_cc_313_execute_65414_145_), .Y(\o[145] ) );
  BUFX2 BUFX2_1057 ( .A(_auto_iopadmap_cc_313_execute_65414_146_), .Y(\o[146] ) );
  BUFX2 BUFX2_1058 ( .A(_auto_iopadmap_cc_313_execute_65414_147_), .Y(\o[147] ) );
  BUFX2 BUFX2_1059 ( .A(_auto_iopadmap_cc_313_execute_65414_148_), .Y(\o[148] ) );
  BUFX2 BUFX2_106 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf3), .Y(u2__abc_44228_n7548_1_bF_buf54) );
  BUFX2 BUFX2_1060 ( .A(_auto_iopadmap_cc_313_execute_65414_149_), .Y(\o[149] ) );
  BUFX2 BUFX2_1061 ( .A(_auto_iopadmap_cc_313_execute_65414_150_), .Y(\o[150] ) );
  BUFX2 BUFX2_1062 ( .A(_auto_iopadmap_cc_313_execute_65414_151_), .Y(\o[151] ) );
  BUFX2 BUFX2_1063 ( .A(_auto_iopadmap_cc_313_execute_65414_152_), .Y(\o[152] ) );
  BUFX2 BUFX2_1064 ( .A(_auto_iopadmap_cc_313_execute_65414_153_), .Y(\o[153] ) );
  BUFX2 BUFX2_1065 ( .A(_auto_iopadmap_cc_313_execute_65414_154_), .Y(\o[154] ) );
  BUFX2 BUFX2_1066 ( .A(_auto_iopadmap_cc_313_execute_65414_155_), .Y(\o[155] ) );
  BUFX2 BUFX2_1067 ( .A(_auto_iopadmap_cc_313_execute_65414_156_), .Y(\o[156] ) );
  BUFX2 BUFX2_1068 ( .A(_auto_iopadmap_cc_313_execute_65414_157_), .Y(\o[157] ) );
  BUFX2 BUFX2_1069 ( .A(_auto_iopadmap_cc_313_execute_65414_158_), .Y(\o[158] ) );
  BUFX2 BUFX2_107 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf2), .Y(u2__abc_44228_n7548_1_bF_buf53) );
  BUFX2 BUFX2_1070 ( .A(_auto_iopadmap_cc_313_execute_65414_159_), .Y(\o[159] ) );
  BUFX2 BUFX2_1071 ( .A(_auto_iopadmap_cc_313_execute_65414_160_), .Y(\o[160] ) );
  BUFX2 BUFX2_1072 ( .A(_auto_iopadmap_cc_313_execute_65414_161_), .Y(\o[161] ) );
  BUFX2 BUFX2_1073 ( .A(_auto_iopadmap_cc_313_execute_65414_162_), .Y(\o[162] ) );
  BUFX2 BUFX2_1074 ( .A(_auto_iopadmap_cc_313_execute_65414_163_), .Y(\o[163] ) );
  BUFX2 BUFX2_1075 ( .A(_auto_iopadmap_cc_313_execute_65414_164_), .Y(\o[164] ) );
  BUFX2 BUFX2_1076 ( .A(_auto_iopadmap_cc_313_execute_65414_165_), .Y(\o[165] ) );
  BUFX2 BUFX2_1077 ( .A(_auto_iopadmap_cc_313_execute_65414_166_), .Y(\o[166] ) );
  BUFX2 BUFX2_1078 ( .A(_auto_iopadmap_cc_313_execute_65414_167_), .Y(\o[167] ) );
  BUFX2 BUFX2_1079 ( .A(_auto_iopadmap_cc_313_execute_65414_168_), .Y(\o[168] ) );
  BUFX2 BUFX2_108 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf1), .Y(u2__abc_44228_n7548_1_bF_buf52) );
  BUFX2 BUFX2_1080 ( .A(_auto_iopadmap_cc_313_execute_65414_169_), .Y(\o[169] ) );
  BUFX2 BUFX2_1081 ( .A(_auto_iopadmap_cc_313_execute_65414_170_), .Y(\o[170] ) );
  BUFX2 BUFX2_1082 ( .A(_auto_iopadmap_cc_313_execute_65414_171_), .Y(\o[171] ) );
  BUFX2 BUFX2_1083 ( .A(_auto_iopadmap_cc_313_execute_65414_172_), .Y(\o[172] ) );
  BUFX2 BUFX2_1084 ( .A(_auto_iopadmap_cc_313_execute_65414_173_), .Y(\o[173] ) );
  BUFX2 BUFX2_1085 ( .A(_auto_iopadmap_cc_313_execute_65414_174_), .Y(\o[174] ) );
  BUFX2 BUFX2_1086 ( .A(_auto_iopadmap_cc_313_execute_65414_175_), .Y(\o[175] ) );
  BUFX2 BUFX2_1087 ( .A(_auto_iopadmap_cc_313_execute_65414_176_), .Y(\o[176] ) );
  BUFX2 BUFX2_1088 ( .A(_auto_iopadmap_cc_313_execute_65414_177_), .Y(\o[177] ) );
  BUFX2 BUFX2_1089 ( .A(_auto_iopadmap_cc_313_execute_65414_178_), .Y(\o[178] ) );
  BUFX2 BUFX2_109 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf0), .Y(u2__abc_44228_n7548_1_bF_buf51) );
  BUFX2 BUFX2_1090 ( .A(_auto_iopadmap_cc_313_execute_65414_179_), .Y(\o[179] ) );
  BUFX2 BUFX2_1091 ( .A(_auto_iopadmap_cc_313_execute_65414_180_), .Y(\o[180] ) );
  BUFX2 BUFX2_1092 ( .A(_auto_iopadmap_cc_313_execute_65414_181_), .Y(\o[181] ) );
  BUFX2 BUFX2_1093 ( .A(_auto_iopadmap_cc_313_execute_65414_182_), .Y(\o[182] ) );
  BUFX2 BUFX2_1094 ( .A(_auto_iopadmap_cc_313_execute_65414_183_), .Y(\o[183] ) );
  BUFX2 BUFX2_1095 ( .A(_auto_iopadmap_cc_313_execute_65414_184_), .Y(\o[184] ) );
  BUFX2 BUFX2_1096 ( .A(_auto_iopadmap_cc_313_execute_65414_185_), .Y(\o[185] ) );
  BUFX2 BUFX2_1097 ( .A(_auto_iopadmap_cc_313_execute_65414_186_), .Y(\o[186] ) );
  BUFX2 BUFX2_1098 ( .A(_auto_iopadmap_cc_313_execute_65414_187_), .Y(\o[187] ) );
  BUFX2 BUFX2_1099 ( .A(_auto_iopadmap_cc_313_execute_65414_188_), .Y(\o[188] ) );
  BUFX2 BUFX2_11 ( .A(clk), .Y(clk_hier0_bF_buf7) );
  BUFX2 BUFX2_110 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf50) );
  BUFX2 BUFX2_1100 ( .A(_auto_iopadmap_cc_313_execute_65414_189_), .Y(\o[189] ) );
  BUFX2 BUFX2_1101 ( .A(_auto_iopadmap_cc_313_execute_65414_190_), .Y(\o[190] ) );
  BUFX2 BUFX2_1102 ( .A(_auto_iopadmap_cc_313_execute_65414_191_), .Y(\o[191] ) );
  BUFX2 BUFX2_1103 ( .A(_auto_iopadmap_cc_313_execute_65414_192_), .Y(\o[192] ) );
  BUFX2 BUFX2_1104 ( .A(_auto_iopadmap_cc_313_execute_65414_193_), .Y(\o[193] ) );
  BUFX2 BUFX2_1105 ( .A(_auto_iopadmap_cc_313_execute_65414_194_), .Y(\o[194] ) );
  BUFX2 BUFX2_1106 ( .A(_auto_iopadmap_cc_313_execute_65414_195_), .Y(\o[195] ) );
  BUFX2 BUFX2_1107 ( .A(_auto_iopadmap_cc_313_execute_65414_196_), .Y(\o[196] ) );
  BUFX2 BUFX2_1108 ( .A(_auto_iopadmap_cc_313_execute_65414_197_), .Y(\o[197] ) );
  BUFX2 BUFX2_1109 ( .A(_auto_iopadmap_cc_313_execute_65414_198_), .Y(\o[198] ) );
  BUFX2 BUFX2_111 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf49) );
  BUFX2 BUFX2_1110 ( .A(_auto_iopadmap_cc_313_execute_65414_199_), .Y(\o[199] ) );
  BUFX2 BUFX2_1111 ( .A(_auto_iopadmap_cc_313_execute_65414_200_), .Y(\o[200] ) );
  BUFX2 BUFX2_1112 ( .A(_auto_iopadmap_cc_313_execute_65414_201_), .Y(\o[201] ) );
  BUFX2 BUFX2_1113 ( .A(_auto_iopadmap_cc_313_execute_65414_202_), .Y(\o[202] ) );
  BUFX2 BUFX2_1114 ( .A(_auto_iopadmap_cc_313_execute_65414_203_), .Y(\o[203] ) );
  BUFX2 BUFX2_1115 ( .A(_auto_iopadmap_cc_313_execute_65414_204_), .Y(\o[204] ) );
  BUFX2 BUFX2_1116 ( .A(_auto_iopadmap_cc_313_execute_65414_205_), .Y(\o[205] ) );
  BUFX2 BUFX2_1117 ( .A(_auto_iopadmap_cc_313_execute_65414_206_), .Y(\o[206] ) );
  BUFX2 BUFX2_1118 ( .A(_auto_iopadmap_cc_313_execute_65414_207_), .Y(\o[207] ) );
  BUFX2 BUFX2_1119 ( .A(_auto_iopadmap_cc_313_execute_65414_208_), .Y(\o[208] ) );
  BUFX2 BUFX2_112 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf4), .Y(u2__abc_44228_n7548_1_bF_buf48) );
  BUFX2 BUFX2_1120 ( .A(_auto_iopadmap_cc_313_execute_65414_209_), .Y(\o[209] ) );
  BUFX2 BUFX2_1121 ( .A(_auto_iopadmap_cc_313_execute_65414_210_), .Y(\o[210] ) );
  BUFX2 BUFX2_1122 ( .A(_auto_iopadmap_cc_313_execute_65414_211_), .Y(\o[211] ) );
  BUFX2 BUFX2_1123 ( .A(_auto_iopadmap_cc_313_execute_65414_212_), .Y(\o[212] ) );
  BUFX2 BUFX2_1124 ( .A(_auto_iopadmap_cc_313_execute_65414_213_), .Y(\o[213] ) );
  BUFX2 BUFX2_1125 ( .A(_auto_iopadmap_cc_313_execute_65414_214_), .Y(\o[214] ) );
  BUFX2 BUFX2_1126 ( .A(_auto_iopadmap_cc_313_execute_65414_215_), .Y(\o[215] ) );
  BUFX2 BUFX2_1127 ( .A(_auto_iopadmap_cc_313_execute_65414_216_), .Y(\o[216] ) );
  BUFX2 BUFX2_1128 ( .A(_auto_iopadmap_cc_313_execute_65414_217_), .Y(\o[217] ) );
  BUFX2 BUFX2_1129 ( .A(_auto_iopadmap_cc_313_execute_65414_218_), .Y(\o[218] ) );
  BUFX2 BUFX2_113 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf3), .Y(u2__abc_44228_n7548_1_bF_buf47) );
  BUFX2 BUFX2_1130 ( .A(_auto_iopadmap_cc_313_execute_65414_219_), .Y(\o[219] ) );
  BUFX2 BUFX2_1131 ( .A(_auto_iopadmap_cc_313_execute_65414_220_), .Y(\o[220] ) );
  BUFX2 BUFX2_1132 ( .A(_auto_iopadmap_cc_313_execute_65414_221_), .Y(\o[221] ) );
  BUFX2 BUFX2_1133 ( .A(_auto_iopadmap_cc_313_execute_65414_222_), .Y(\o[222] ) );
  BUFX2 BUFX2_1134 ( .A(_auto_iopadmap_cc_313_execute_65414_223_), .Y(\o[223] ) );
  BUFX2 BUFX2_1135 ( .A(_auto_iopadmap_cc_313_execute_65414_224_), .Y(\o[224] ) );
  BUFX2 BUFX2_1136 ( .A(_auto_iopadmap_cc_313_execute_65414_225_), .Y(\o[225] ) );
  BUFX2 BUFX2_1137 ( .A(_auto_iopadmap_cc_313_execute_65414_226_), .Y(\o[226] ) );
  BUFX2 BUFX2_1138 ( .A(_auto_iopadmap_cc_313_execute_65414_227_), .Y(\o[227] ) );
  BUFX2 BUFX2_1139 ( .A(_auto_iopadmap_cc_313_execute_65414_228_), .Y(\o[228] ) );
  BUFX2 BUFX2_114 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf2), .Y(u2__abc_44228_n7548_1_bF_buf46) );
  BUFX2 BUFX2_1140 ( .A(_auto_iopadmap_cc_313_execute_65414_229_), .Y(\o[229] ) );
  BUFX2 BUFX2_1141 ( .A(_auto_iopadmap_cc_313_execute_65414_230_), .Y(\o[230] ) );
  BUFX2 BUFX2_1142 ( .A(_auto_iopadmap_cc_313_execute_65414_231_), .Y(\o[231] ) );
  BUFX2 BUFX2_1143 ( .A(_auto_iopadmap_cc_313_execute_65414_232_), .Y(\o[232] ) );
  BUFX2 BUFX2_1144 ( .A(_auto_iopadmap_cc_313_execute_65414_233_), .Y(\o[233] ) );
  BUFX2 BUFX2_1145 ( .A(_auto_iopadmap_cc_313_execute_65414_234_), .Y(\o[234] ) );
  BUFX2 BUFX2_1146 ( .A(_auto_iopadmap_cc_313_execute_65414_235_), .Y(\o[235] ) );
  BUFX2 BUFX2_1147 ( .A(_auto_iopadmap_cc_313_execute_65414_236_), .Y(\o[236] ) );
  BUFX2 BUFX2_1148 ( .A(_auto_iopadmap_cc_313_execute_65414_237_), .Y(\o[237] ) );
  BUFX2 BUFX2_1149 ( .A(_auto_iopadmap_cc_313_execute_65414_238_), .Y(\o[238] ) );
  BUFX2 BUFX2_115 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf1), .Y(u2__abc_44228_n7548_1_bF_buf45) );
  BUFX2 BUFX2_1150 ( .A(_auto_iopadmap_cc_313_execute_65414_239_), .Y(\o[239] ) );
  BUFX2 BUFX2_1151 ( .A(_auto_iopadmap_cc_313_execute_65414_240_), .Y(\o[240] ) );
  BUFX2 BUFX2_1152 ( .A(_auto_iopadmap_cc_313_execute_65414_241_), .Y(\o[241] ) );
  BUFX2 BUFX2_116 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf0), .Y(u2__abc_44228_n7548_1_bF_buf44) );
  BUFX2 BUFX2_117 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf43) );
  BUFX2 BUFX2_118 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf42) );
  BUFX2 BUFX2_119 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf4), .Y(u2__abc_44228_n7548_1_bF_buf41) );
  BUFX2 BUFX2_12 ( .A(clk), .Y(clk_hier0_bF_buf6) );
  BUFX2 BUFX2_120 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf3), .Y(u2__abc_44228_n7548_1_bF_buf40) );
  BUFX2 BUFX2_121 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf2), .Y(u2__abc_44228_n7548_1_bF_buf39) );
  BUFX2 BUFX2_122 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf1), .Y(u2__abc_44228_n7548_1_bF_buf38) );
  BUFX2 BUFX2_123 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf0), .Y(u2__abc_44228_n7548_1_bF_buf37) );
  BUFX2 BUFX2_124 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf36) );
  BUFX2 BUFX2_125 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf35) );
  BUFX2 BUFX2_126 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf4), .Y(u2__abc_44228_n7548_1_bF_buf34) );
  BUFX2 BUFX2_127 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf3), .Y(u2__abc_44228_n7548_1_bF_buf33) );
  BUFX2 BUFX2_128 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf2), .Y(u2__abc_44228_n7548_1_bF_buf32) );
  BUFX2 BUFX2_129 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf1), .Y(u2__abc_44228_n7548_1_bF_buf31) );
  BUFX2 BUFX2_13 ( .A(clk), .Y(clk_hier0_bF_buf5) );
  BUFX2 BUFX2_130 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf0), .Y(u2__abc_44228_n7548_1_bF_buf30) );
  BUFX2 BUFX2_131 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf29) );
  BUFX2 BUFX2_132 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf28) );
  BUFX2 BUFX2_133 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf4), .Y(u2__abc_44228_n7548_1_bF_buf27) );
  BUFX2 BUFX2_134 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf3), .Y(u2__abc_44228_n7548_1_bF_buf26) );
  BUFX2 BUFX2_135 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf2), .Y(u2__abc_44228_n7548_1_bF_buf25) );
  BUFX2 BUFX2_136 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf1), .Y(u2__abc_44228_n7548_1_bF_buf24) );
  BUFX2 BUFX2_137 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf0), .Y(u2__abc_44228_n7548_1_bF_buf23) );
  BUFX2 BUFX2_138 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf22) );
  BUFX2 BUFX2_139 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf21) );
  BUFX2 BUFX2_14 ( .A(clk), .Y(clk_hier0_bF_buf4) );
  BUFX2 BUFX2_140 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf4), .Y(u2__abc_44228_n7548_1_bF_buf20) );
  BUFX2 BUFX2_141 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf3), .Y(u2__abc_44228_n7548_1_bF_buf19) );
  BUFX2 BUFX2_142 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf2), .Y(u2__abc_44228_n7548_1_bF_buf18) );
  BUFX2 BUFX2_143 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf1), .Y(u2__abc_44228_n7548_1_bF_buf17) );
  BUFX2 BUFX2_144 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf0), .Y(u2__abc_44228_n7548_1_bF_buf16) );
  BUFX2 BUFX2_145 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf15) );
  BUFX2 BUFX2_146 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf14) );
  BUFX2 BUFX2_147 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf4), .Y(u2__abc_44228_n7548_1_bF_buf13) );
  BUFX2 BUFX2_148 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf3), .Y(u2__abc_44228_n7548_1_bF_buf12) );
  BUFX2 BUFX2_149 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf2), .Y(u2__abc_44228_n7548_1_bF_buf11) );
  BUFX2 BUFX2_15 ( .A(clk), .Y(clk_hier0_bF_buf3) );
  BUFX2 BUFX2_150 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf1), .Y(u2__abc_44228_n7548_1_bF_buf10) );
  BUFX2 BUFX2_151 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf0), .Y(u2__abc_44228_n7548_1_bF_buf9) );
  BUFX2 BUFX2_152 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf8) );
  BUFX2 BUFX2_153 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf7) );
  BUFX2 BUFX2_154 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf4), .Y(u2__abc_44228_n7548_1_bF_buf6) );
  BUFX2 BUFX2_155 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf3), .Y(u2__abc_44228_n7548_1_bF_buf5) );
  BUFX2 BUFX2_156 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf2), .Y(u2__abc_44228_n7548_1_bF_buf4) );
  BUFX2 BUFX2_157 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf1), .Y(u2__abc_44228_n7548_1_bF_buf3) );
  BUFX2 BUFX2_158 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf0), .Y(u2__abc_44228_n7548_1_bF_buf2) );
  BUFX2 BUFX2_159 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf6), .Y(u2__abc_44228_n7548_1_bF_buf1) );
  BUFX2 BUFX2_16 ( .A(clk), .Y(clk_hier0_bF_buf2) );
  BUFX2 BUFX2_160 ( .A(u2__abc_44228_n7548_1_hier0_bF_buf5), .Y(u2__abc_44228_n7548_1_bF_buf0) );
  BUFX2 BUFX2_161 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf121) );
  BUFX2 BUFX2_162 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf120) );
  BUFX2 BUFX2_163 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf119) );
  BUFX2 BUFX2_164 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf118) );
  BUFX2 BUFX2_165 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf117) );
  BUFX2 BUFX2_166 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf116) );
  BUFX2 BUFX2_167 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf115) );
  BUFX2 BUFX2_168 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf114) );
  BUFX2 BUFX2_169 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf113) );
  BUFX2 BUFX2_17 ( .A(clk), .Y(clk_hier0_bF_buf1) );
  BUFX2 BUFX2_170 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf112) );
  BUFX2 BUFX2_171 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf111) );
  BUFX2 BUFX2_172 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf110) );
  BUFX2 BUFX2_173 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf109) );
  BUFX2 BUFX2_174 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf108) );
  BUFX2 BUFX2_175 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf107) );
  BUFX2 BUFX2_176 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf106) );
  BUFX2 BUFX2_177 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf105) );
  BUFX2 BUFX2_178 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf104) );
  BUFX2 BUFX2_179 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf103) );
  BUFX2 BUFX2_18 ( .A(clk), .Y(clk_hier0_bF_buf0) );
  BUFX2 BUFX2_180 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf102) );
  BUFX2 BUFX2_181 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf101) );
  BUFX2 BUFX2_182 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf100) );
  BUFX2 BUFX2_183 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf99) );
  BUFX2 BUFX2_184 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf98) );
  BUFX2 BUFX2_185 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf97) );
  BUFX2 BUFX2_186 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf96) );
  BUFX2 BUFX2_187 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf95) );
  BUFX2 BUFX2_188 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf94) );
  BUFX2 BUFX2_189 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf93) );
  BUFX2 BUFX2_19 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf9) );
  BUFX2 BUFX2_190 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf92) );
  BUFX2 BUFX2_191 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf91) );
  BUFX2 BUFX2_192 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf90) );
  BUFX2 BUFX2_193 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf89) );
  BUFX2 BUFX2_194 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf88) );
  BUFX2 BUFX2_195 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf87) );
  BUFX2 BUFX2_196 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf86) );
  BUFX2 BUFX2_197 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf85) );
  BUFX2 BUFX2_198 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf84) );
  BUFX2 BUFX2_199 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf83) );
  BUFX2 BUFX2_2 ( .A(u2__abc_44228_n7548_1), .Y(u2__abc_44228_n7548_1_hier0_bF_buf5) );
  BUFX2 BUFX2_20 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf8) );
  BUFX2 BUFX2_200 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf82) );
  BUFX2 BUFX2_201 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf81) );
  BUFX2 BUFX2_202 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf80) );
  BUFX2 BUFX2_203 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf79) );
  BUFX2 BUFX2_204 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf78) );
  BUFX2 BUFX2_205 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf77) );
  BUFX2 BUFX2_206 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf76) );
  BUFX2 BUFX2_207 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf75) );
  BUFX2 BUFX2_208 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf74) );
  BUFX2 BUFX2_209 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf73) );
  BUFX2 BUFX2_21 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf7) );
  BUFX2 BUFX2_210 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf72) );
  BUFX2 BUFX2_211 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf71) );
  BUFX2 BUFX2_212 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf70) );
  BUFX2 BUFX2_213 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf69) );
  BUFX2 BUFX2_214 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf68) );
  BUFX2 BUFX2_215 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf67) );
  BUFX2 BUFX2_216 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf66) );
  BUFX2 BUFX2_217 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf65) );
  BUFX2 BUFX2_218 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf64) );
  BUFX2 BUFX2_219 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf63) );
  BUFX2 BUFX2_22 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf6) );
  BUFX2 BUFX2_220 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf62) );
  BUFX2 BUFX2_221 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf61) );
  BUFX2 BUFX2_222 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf60) );
  BUFX2 BUFX2_223 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf59) );
  BUFX2 BUFX2_224 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf58) );
  BUFX2 BUFX2_225 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf57) );
  BUFX2 BUFX2_226 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf56) );
  BUFX2 BUFX2_227 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf55) );
  BUFX2 BUFX2_228 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf54) );
  BUFX2 BUFX2_229 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf53) );
  BUFX2 BUFX2_23 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf5) );
  BUFX2 BUFX2_230 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf52) );
  BUFX2 BUFX2_231 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf51) );
  BUFX2 BUFX2_232 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf50) );
  BUFX2 BUFX2_233 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf49) );
  BUFX2 BUFX2_234 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf48) );
  BUFX2 BUFX2_235 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf47) );
  BUFX2 BUFX2_236 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf46) );
  BUFX2 BUFX2_237 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf45) );
  BUFX2 BUFX2_238 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf44) );
  BUFX2 BUFX2_239 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf43) );
  BUFX2 BUFX2_24 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf4) );
  BUFX2 BUFX2_240 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf42) );
  BUFX2 BUFX2_241 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf41) );
  BUFX2 BUFX2_242 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf40) );
  BUFX2 BUFX2_243 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf39) );
  BUFX2 BUFX2_244 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf38) );
  BUFX2 BUFX2_245 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf37) );
  BUFX2 BUFX2_246 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf36) );
  BUFX2 BUFX2_247 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf35) );
  BUFX2 BUFX2_248 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf34) );
  BUFX2 BUFX2_249 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf33) );
  BUFX2 BUFX2_25 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf3) );
  BUFX2 BUFX2_250 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf32) );
  BUFX2 BUFX2_251 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf31) );
  BUFX2 BUFX2_252 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf30) );
  BUFX2 BUFX2_253 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf29) );
  BUFX2 BUFX2_254 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf28) );
  BUFX2 BUFX2_255 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf27) );
  BUFX2 BUFX2_256 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf26) );
  BUFX2 BUFX2_257 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf25) );
  BUFX2 BUFX2_258 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf24) );
  BUFX2 BUFX2_259 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf23) );
  BUFX2 BUFX2_26 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf2) );
  BUFX2 BUFX2_260 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf22) );
  BUFX2 BUFX2_261 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf21) );
  BUFX2 BUFX2_262 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf20) );
  BUFX2 BUFX2_263 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf19) );
  BUFX2 BUFX2_264 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf18) );
  BUFX2 BUFX2_265 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf17) );
  BUFX2 BUFX2_266 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf16) );
  BUFX2 BUFX2_267 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf15) );
  BUFX2 BUFX2_268 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf14) );
  BUFX2 BUFX2_269 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf13) );
  BUFX2 BUFX2_27 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf1) );
  BUFX2 BUFX2_270 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf12) );
  BUFX2 BUFX2_271 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf11) );
  BUFX2 BUFX2_272 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf10) );
  BUFX2 BUFX2_273 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf9) );
  BUFX2 BUFX2_274 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf8) );
  BUFX2 BUFX2_275 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf7) );
  BUFX2 BUFX2_276 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf6) );
  BUFX2 BUFX2_277 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf5) );
  BUFX2 BUFX2_278 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf4) );
  BUFX2 BUFX2_279 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf3) );
  BUFX2 BUFX2_28 ( .A(u2__abc_44228_n2972), .Y(u2__abc_44228_n2972_hier0_bF_buf0) );
  BUFX2 BUFX2_280 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf2) );
  BUFX2 BUFX2_281 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf1) );
  BUFX2 BUFX2_282 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf0) );
  BUFX2 BUFX2_283 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf107) );
  BUFX2 BUFX2_284 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf106) );
  BUFX2 BUFX2_285 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf105) );
  BUFX2 BUFX2_286 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf104) );
  BUFX2 BUFX2_287 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf103) );
  BUFX2 BUFX2_288 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf102) );
  BUFX2 BUFX2_289 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf101) );
  BUFX2 BUFX2_29 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf8) );
  BUFX2 BUFX2_290 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf100) );
  BUFX2 BUFX2_291 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf99) );
  BUFX2 BUFX2_292 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf98) );
  BUFX2 BUFX2_293 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf97) );
  BUFX2 BUFX2_294 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf96) );
  BUFX2 BUFX2_295 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf95) );
  BUFX2 BUFX2_296 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf94) );
  BUFX2 BUFX2_297 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf93) );
  BUFX2 BUFX2_298 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf92) );
  BUFX2 BUFX2_299 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf91) );
  BUFX2 BUFX2_3 ( .A(u2__abc_44228_n7548_1), .Y(u2__abc_44228_n7548_1_hier0_bF_buf4) );
  BUFX2 BUFX2_30 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf7) );
  BUFX2 BUFX2_300 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf90) );
  BUFX2 BUFX2_301 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf89) );
  BUFX2 BUFX2_302 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf88) );
  BUFX2 BUFX2_303 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf87) );
  BUFX2 BUFX2_304 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf86) );
  BUFX2 BUFX2_305 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf85) );
  BUFX2 BUFX2_306 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf84) );
  BUFX2 BUFX2_307 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf83) );
  BUFX2 BUFX2_308 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf82) );
  BUFX2 BUFX2_309 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf81) );
  BUFX2 BUFX2_31 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf6) );
  BUFX2 BUFX2_310 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf80) );
  BUFX2 BUFX2_311 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf79) );
  BUFX2 BUFX2_312 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf78) );
  BUFX2 BUFX2_313 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf77) );
  BUFX2 BUFX2_314 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf76) );
  BUFX2 BUFX2_315 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf75) );
  BUFX2 BUFX2_316 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf74) );
  BUFX2 BUFX2_317 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf73) );
  BUFX2 BUFX2_318 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf72) );
  BUFX2 BUFX2_319 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf71) );
  BUFX2 BUFX2_32 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf5) );
  BUFX2 BUFX2_320 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf70) );
  BUFX2 BUFX2_321 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf69) );
  BUFX2 BUFX2_322 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf68) );
  BUFX2 BUFX2_323 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf67) );
  BUFX2 BUFX2_324 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf66) );
  BUFX2 BUFX2_325 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf65) );
  BUFX2 BUFX2_326 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf64) );
  BUFX2 BUFX2_327 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf63) );
  BUFX2 BUFX2_328 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf62) );
  BUFX2 BUFX2_329 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf61) );
  BUFX2 BUFX2_33 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf4) );
  BUFX2 BUFX2_330 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf60) );
  BUFX2 BUFX2_331 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf59) );
  BUFX2 BUFX2_332 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf58) );
  BUFX2 BUFX2_333 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf57) );
  BUFX2 BUFX2_334 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf56) );
  BUFX2 BUFX2_335 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf55) );
  BUFX2 BUFX2_336 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf54) );
  BUFX2 BUFX2_337 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf53) );
  BUFX2 BUFX2_338 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf52) );
  BUFX2 BUFX2_339 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf51) );
  BUFX2 BUFX2_34 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf3) );
  BUFX2 BUFX2_340 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf50) );
  BUFX2 BUFX2_341 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf49) );
  BUFX2 BUFX2_342 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf48) );
  BUFX2 BUFX2_343 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf47) );
  BUFX2 BUFX2_344 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf46) );
  BUFX2 BUFX2_345 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf45) );
  BUFX2 BUFX2_346 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf44) );
  BUFX2 BUFX2_347 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf43) );
  BUFX2 BUFX2_348 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf42) );
  BUFX2 BUFX2_349 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf41) );
  BUFX2 BUFX2_35 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf2) );
  BUFX2 BUFX2_350 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf40) );
  BUFX2 BUFX2_351 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf39) );
  BUFX2 BUFX2_352 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf38) );
  BUFX2 BUFX2_353 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf37) );
  BUFX2 BUFX2_354 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf36) );
  BUFX2 BUFX2_355 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf35) );
  BUFX2 BUFX2_356 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf34) );
  BUFX2 BUFX2_357 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf33) );
  BUFX2 BUFX2_358 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf32) );
  BUFX2 BUFX2_359 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf31) );
  BUFX2 BUFX2_36 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf1) );
  BUFX2 BUFX2_360 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf30) );
  BUFX2 BUFX2_361 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf29) );
  BUFX2 BUFX2_362 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf28) );
  BUFX2 BUFX2_363 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf27) );
  BUFX2 BUFX2_364 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf26) );
  BUFX2 BUFX2_365 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf25) );
  BUFX2 BUFX2_366 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf24) );
  BUFX2 BUFX2_367 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf23) );
  BUFX2 BUFX2_368 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf22) );
  BUFX2 BUFX2_369 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf21) );
  BUFX2 BUFX2_37 ( .A(u2__abc_44228_n3062), .Y(u2__abc_44228_n3062_hier0_bF_buf0) );
  BUFX2 BUFX2_370 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf20) );
  BUFX2 BUFX2_371 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf19) );
  BUFX2 BUFX2_372 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf18) );
  BUFX2 BUFX2_373 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf17) );
  BUFX2 BUFX2_374 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf16) );
  BUFX2 BUFX2_375 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf15) );
  BUFX2 BUFX2_376 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf14) );
  BUFX2 BUFX2_377 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf13) );
  BUFX2 BUFX2_378 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf12) );
  BUFX2 BUFX2_379 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf11) );
  BUFX2 BUFX2_38 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf9) );
  BUFX2 BUFX2_380 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf10) );
  BUFX2 BUFX2_381 ( .A(u2__abc_44228_n2972_hier0_bF_buf1), .Y(u2__abc_44228_n2972_bF_buf9) );
  BUFX2 BUFX2_382 ( .A(u2__abc_44228_n2972_hier0_bF_buf0), .Y(u2__abc_44228_n2972_bF_buf8) );
  BUFX2 BUFX2_383 ( .A(u2__abc_44228_n2972_hier0_bF_buf9), .Y(u2__abc_44228_n2972_bF_buf7) );
  BUFX2 BUFX2_384 ( .A(u2__abc_44228_n2972_hier0_bF_buf8), .Y(u2__abc_44228_n2972_bF_buf6) );
  BUFX2 BUFX2_385 ( .A(u2__abc_44228_n2972_hier0_bF_buf7), .Y(u2__abc_44228_n2972_bF_buf5) );
  BUFX2 BUFX2_386 ( .A(u2__abc_44228_n2972_hier0_bF_buf6), .Y(u2__abc_44228_n2972_bF_buf4) );
  BUFX2 BUFX2_387 ( .A(u2__abc_44228_n2972_hier0_bF_buf5), .Y(u2__abc_44228_n2972_bF_buf3) );
  BUFX2 BUFX2_388 ( .A(u2__abc_44228_n2972_hier0_bF_buf4), .Y(u2__abc_44228_n2972_bF_buf2) );
  BUFX2 BUFX2_389 ( .A(u2__abc_44228_n2972_hier0_bF_buf3), .Y(u2__abc_44228_n2972_bF_buf1) );
  BUFX2 BUFX2_39 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf8) );
  BUFX2 BUFX2_390 ( .A(u2__abc_44228_n2972_hier0_bF_buf2), .Y(u2__abc_44228_n2972_bF_buf0) );
  BUFX2 BUFX2_391 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf92) );
  BUFX2 BUFX2_392 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf91) );
  BUFX2 BUFX2_393 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf90) );
  BUFX2 BUFX2_394 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf89) );
  BUFX2 BUFX2_395 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf88) );
  BUFX2 BUFX2_396 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf87) );
  BUFX2 BUFX2_397 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf86) );
  BUFX2 BUFX2_398 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf85) );
  BUFX2 BUFX2_399 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf84) );
  BUFX2 BUFX2_4 ( .A(u2__abc_44228_n7548_1), .Y(u2__abc_44228_n7548_1_hier0_bF_buf3) );
  BUFX2 BUFX2_40 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf7) );
  BUFX2 BUFX2_400 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf83) );
  BUFX2 BUFX2_401 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf82) );
  BUFX2 BUFX2_402 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf81) );
  BUFX2 BUFX2_403 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf80) );
  BUFX2 BUFX2_404 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf79) );
  BUFX2 BUFX2_405 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf78) );
  BUFX2 BUFX2_406 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf77) );
  BUFX2 BUFX2_407 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf76) );
  BUFX2 BUFX2_408 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf75) );
  BUFX2 BUFX2_409 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf74) );
  BUFX2 BUFX2_41 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf6) );
  BUFX2 BUFX2_410 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf73) );
  BUFX2 BUFX2_411 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf72) );
  BUFX2 BUFX2_412 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf71) );
  BUFX2 BUFX2_413 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf70) );
  BUFX2 BUFX2_414 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf69) );
  BUFX2 BUFX2_415 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf68) );
  BUFX2 BUFX2_416 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf67) );
  BUFX2 BUFX2_417 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf66) );
  BUFX2 BUFX2_418 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf65) );
  BUFX2 BUFX2_419 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf64) );
  BUFX2 BUFX2_42 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf5) );
  BUFX2 BUFX2_420 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf63) );
  BUFX2 BUFX2_421 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf62) );
  BUFX2 BUFX2_422 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf61) );
  BUFX2 BUFX2_423 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf60) );
  BUFX2 BUFX2_424 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf59) );
  BUFX2 BUFX2_425 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf58) );
  BUFX2 BUFX2_426 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf57) );
  BUFX2 BUFX2_427 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf56) );
  BUFX2 BUFX2_428 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf55) );
  BUFX2 BUFX2_429 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf54) );
  BUFX2 BUFX2_43 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf4) );
  BUFX2 BUFX2_430 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf53) );
  BUFX2 BUFX2_431 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf52) );
  BUFX2 BUFX2_432 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf51) );
  BUFX2 BUFX2_433 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf50) );
  BUFX2 BUFX2_434 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf49) );
  BUFX2 BUFX2_435 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf48) );
  BUFX2 BUFX2_436 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf47) );
  BUFX2 BUFX2_437 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf46) );
  BUFX2 BUFX2_438 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf45) );
  BUFX2 BUFX2_439 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf44) );
  BUFX2 BUFX2_44 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf3) );
  BUFX2 BUFX2_440 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf43) );
  BUFX2 BUFX2_441 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf42) );
  BUFX2 BUFX2_442 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf41) );
  BUFX2 BUFX2_443 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf40) );
  BUFX2 BUFX2_444 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf39) );
  BUFX2 BUFX2_445 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf38) );
  BUFX2 BUFX2_446 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf37) );
  BUFX2 BUFX2_447 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf36) );
  BUFX2 BUFX2_448 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf35) );
  BUFX2 BUFX2_449 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf34) );
  BUFX2 BUFX2_45 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf2) );
  BUFX2 BUFX2_450 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf33) );
  BUFX2 BUFX2_451 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf32) );
  BUFX2 BUFX2_452 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf31) );
  BUFX2 BUFX2_453 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf30) );
  BUFX2 BUFX2_454 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf29) );
  BUFX2 BUFX2_455 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf28) );
  BUFX2 BUFX2_456 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf27) );
  BUFX2 BUFX2_457 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf26) );
  BUFX2 BUFX2_458 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf25) );
  BUFX2 BUFX2_459 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf24) );
  BUFX2 BUFX2_46 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf1) );
  BUFX2 BUFX2_460 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf23) );
  BUFX2 BUFX2_461 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf22) );
  BUFX2 BUFX2_462 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf21) );
  BUFX2 BUFX2_463 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf20) );
  BUFX2 BUFX2_464 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf19) );
  BUFX2 BUFX2_465 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf18) );
  BUFX2 BUFX2_466 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf17) );
  BUFX2 BUFX2_467 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf16) );
  BUFX2 BUFX2_468 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf15) );
  BUFX2 BUFX2_469 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf14) );
  BUFX2 BUFX2_47 ( .A(u2__abc_44228_n2966), .Y(u2__abc_44228_n2966_hier0_bF_buf0) );
  BUFX2 BUFX2_470 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf13) );
  BUFX2 BUFX2_471 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf12) );
  BUFX2 BUFX2_472 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf11) );
  BUFX2 BUFX2_473 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf10) );
  BUFX2 BUFX2_474 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf9) );
  BUFX2 BUFX2_475 ( .A(u2__abc_44228_n3062_hier0_bF_buf5), .Y(u2__abc_44228_n3062_bF_buf8) );
  BUFX2 BUFX2_476 ( .A(u2__abc_44228_n3062_hier0_bF_buf4), .Y(u2__abc_44228_n3062_bF_buf7) );
  BUFX2 BUFX2_477 ( .A(u2__abc_44228_n3062_hier0_bF_buf3), .Y(u2__abc_44228_n3062_bF_buf6) );
  BUFX2 BUFX2_478 ( .A(u2__abc_44228_n3062_hier0_bF_buf2), .Y(u2__abc_44228_n3062_bF_buf5) );
  BUFX2 BUFX2_479 ( .A(u2__abc_44228_n3062_hier0_bF_buf1), .Y(u2__abc_44228_n3062_bF_buf4) );
  BUFX2 BUFX2_48 ( .A(u2__abc_44228_n7547), .Y(u2__abc_44228_n7547_hier0_bF_buf6) );
  BUFX2 BUFX2_480 ( .A(u2__abc_44228_n3062_hier0_bF_buf0), .Y(u2__abc_44228_n3062_bF_buf3) );
  BUFX2 BUFX2_481 ( .A(u2__abc_44228_n3062_hier0_bF_buf8), .Y(u2__abc_44228_n3062_bF_buf2) );
  BUFX2 BUFX2_482 ( .A(u2__abc_44228_n3062_hier0_bF_buf7), .Y(u2__abc_44228_n3062_bF_buf1) );
  BUFX2 BUFX2_483 ( .A(u2__abc_44228_n3062_hier0_bF_buf6), .Y(u2__abc_44228_n3062_bF_buf0) );
  BUFX2 BUFX2_484 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf9) );
  BUFX2 BUFX2_485 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf8) );
  BUFX2 BUFX2_486 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf7) );
  BUFX2 BUFX2_487 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf6) );
  BUFX2 BUFX2_488 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf5) );
  BUFX2 BUFX2_489 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf4) );
  BUFX2 BUFX2_49 ( .A(u2__abc_44228_n7547), .Y(u2__abc_44228_n7547_hier0_bF_buf5) );
  BUFX2 BUFX2_490 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf3) );
  BUFX2 BUFX2_491 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf2) );
  BUFX2 BUFX2_492 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf1) );
  BUFX2 BUFX2_493 ( .A(u2__abc_44228_n8209), .Y(u2__abc_44228_n8209_bF_buf0) );
  BUFX2 BUFX2_494 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf9) );
  BUFX2 BUFX2_495 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf8) );
  BUFX2 BUFX2_496 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf7) );
  BUFX2 BUFX2_497 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf6) );
  BUFX2 BUFX2_498 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf5) );
  BUFX2 BUFX2_499 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf4) );
  BUFX2 BUFX2_5 ( .A(u2__abc_44228_n7548_1), .Y(u2__abc_44228_n7548_1_hier0_bF_buf2) );
  BUFX2 BUFX2_50 ( .A(u2__abc_44228_n7547), .Y(u2__abc_44228_n7547_hier0_bF_buf4) );
  BUFX2 BUFX2_500 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf3) );
  BUFX2 BUFX2_501 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf2) );
  BUFX2 BUFX2_502 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf1) );
  BUFX2 BUFX2_503 ( .A(_abc_64468_n1170), .Y(_abc_64468_n1170_bF_buf0) );
  BUFX2 BUFX2_504 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf14) );
  BUFX2 BUFX2_505 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf13) );
  BUFX2 BUFX2_506 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf12) );
  BUFX2 BUFX2_507 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf11) );
  BUFX2 BUFX2_508 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf10) );
  BUFX2 BUFX2_509 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf9) );
  BUFX2 BUFX2_51 ( .A(u2__abc_44228_n7547), .Y(u2__abc_44228_n7547_hier0_bF_buf3) );
  BUFX2 BUFX2_510 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf8) );
  BUFX2 BUFX2_511 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf7) );
  BUFX2 BUFX2_512 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf6) );
  BUFX2 BUFX2_513 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf5) );
  BUFX2 BUFX2_514 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf4) );
  BUFX2 BUFX2_515 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf3) );
  BUFX2 BUFX2_516 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf2) );
  BUFX2 BUFX2_517 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf1) );
  BUFX2 BUFX2_518 ( .A(u2__abc_44228_n15247), .Y(u2__abc_44228_n15247_bF_buf0) );
  BUFX2 BUFX2_519 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf107) );
  BUFX2 BUFX2_52 ( .A(u2__abc_44228_n7547), .Y(u2__abc_44228_n7547_hier0_bF_buf2) );
  BUFX2 BUFX2_520 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf106) );
  BUFX2 BUFX2_521 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf105) );
  BUFX2 BUFX2_522 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf104) );
  BUFX2 BUFX2_523 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf103) );
  BUFX2 BUFX2_524 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf102) );
  BUFX2 BUFX2_525 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf101) );
  BUFX2 BUFX2_526 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf100) );
  BUFX2 BUFX2_527 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf99) );
  BUFX2 BUFX2_528 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf98) );
  BUFX2 BUFX2_529 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf97) );
  BUFX2 BUFX2_53 ( .A(u2__abc_44228_n7547), .Y(u2__abc_44228_n7547_hier0_bF_buf1) );
  BUFX2 BUFX2_530 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf96) );
  BUFX2 BUFX2_531 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf95) );
  BUFX2 BUFX2_532 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf94) );
  BUFX2 BUFX2_533 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf93) );
  BUFX2 BUFX2_534 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf92) );
  BUFX2 BUFX2_535 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf91) );
  BUFX2 BUFX2_536 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf90) );
  BUFX2 BUFX2_537 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf89) );
  BUFX2 BUFX2_538 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf88) );
  BUFX2 BUFX2_539 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf87) );
  BUFX2 BUFX2_54 ( .A(u2__abc_44228_n7547), .Y(u2__abc_44228_n7547_hier0_bF_buf0) );
  BUFX2 BUFX2_540 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf86) );
  BUFX2 BUFX2_541 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf85) );
  BUFX2 BUFX2_542 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf84) );
  BUFX2 BUFX2_543 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf83) );
  BUFX2 BUFX2_544 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf82) );
  BUFX2 BUFX2_545 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf81) );
  BUFX2 BUFX2_546 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf80) );
  BUFX2 BUFX2_547 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf79) );
  BUFX2 BUFX2_548 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf78) );
  BUFX2 BUFX2_549 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf77) );
  BUFX2 BUFX2_55 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf10) );
  BUFX2 BUFX2_550 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf76) );
  BUFX2 BUFX2_551 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf75) );
  BUFX2 BUFX2_552 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf74) );
  BUFX2 BUFX2_553 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf73) );
  BUFX2 BUFX2_554 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf72) );
  BUFX2 BUFX2_555 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf71) );
  BUFX2 BUFX2_556 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf70) );
  BUFX2 BUFX2_557 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf69) );
  BUFX2 BUFX2_558 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf68) );
  BUFX2 BUFX2_559 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf67) );
  BUFX2 BUFX2_56 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf9) );
  BUFX2 BUFX2_560 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf66) );
  BUFX2 BUFX2_561 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf65) );
  BUFX2 BUFX2_562 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf64) );
  BUFX2 BUFX2_563 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf63) );
  BUFX2 BUFX2_564 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf62) );
  BUFX2 BUFX2_565 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf61) );
  BUFX2 BUFX2_566 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf60) );
  BUFX2 BUFX2_567 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf59) );
  BUFX2 BUFX2_568 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf58) );
  BUFX2 BUFX2_569 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf57) );
  BUFX2 BUFX2_57 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf8) );
  BUFX2 BUFX2_570 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf56) );
  BUFX2 BUFX2_571 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf55) );
  BUFX2 BUFX2_572 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf54) );
  BUFX2 BUFX2_573 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf53) );
  BUFX2 BUFX2_574 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf52) );
  BUFX2 BUFX2_575 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf51) );
  BUFX2 BUFX2_576 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf50) );
  BUFX2 BUFX2_577 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf49) );
  BUFX2 BUFX2_578 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf48) );
  BUFX2 BUFX2_579 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf47) );
  BUFX2 BUFX2_58 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf7) );
  BUFX2 BUFX2_580 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf46) );
  BUFX2 BUFX2_581 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf45) );
  BUFX2 BUFX2_582 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf44) );
  BUFX2 BUFX2_583 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf43) );
  BUFX2 BUFX2_584 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf42) );
  BUFX2 BUFX2_585 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf41) );
  BUFX2 BUFX2_586 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf40) );
  BUFX2 BUFX2_587 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf39) );
  BUFX2 BUFX2_588 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf38) );
  BUFX2 BUFX2_589 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf37) );
  BUFX2 BUFX2_59 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf6) );
  BUFX2 BUFX2_590 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf36) );
  BUFX2 BUFX2_591 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf35) );
  BUFX2 BUFX2_592 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf34) );
  BUFX2 BUFX2_593 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf33) );
  BUFX2 BUFX2_594 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf32) );
  BUFX2 BUFX2_595 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf31) );
  BUFX2 BUFX2_596 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf30) );
  BUFX2 BUFX2_597 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf29) );
  BUFX2 BUFX2_598 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf28) );
  BUFX2 BUFX2_599 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf27) );
  BUFX2 BUFX2_6 ( .A(u2__abc_44228_n7548_1), .Y(u2__abc_44228_n7548_1_hier0_bF_buf1) );
  BUFX2 BUFX2_60 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf5) );
  BUFX2 BUFX2_600 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf26) );
  BUFX2 BUFX2_601 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf25) );
  BUFX2 BUFX2_602 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf24) );
  BUFX2 BUFX2_603 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf23) );
  BUFX2 BUFX2_604 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf22) );
  BUFX2 BUFX2_605 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf21) );
  BUFX2 BUFX2_606 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf20) );
  BUFX2 BUFX2_607 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf19) );
  BUFX2 BUFX2_608 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf18) );
  BUFX2 BUFX2_609 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf17) );
  BUFX2 BUFX2_61 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf4) );
  BUFX2 BUFX2_610 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf16) );
  BUFX2 BUFX2_611 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf15) );
  BUFX2 BUFX2_612 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf14) );
  BUFX2 BUFX2_613 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf13) );
  BUFX2 BUFX2_614 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf12) );
  BUFX2 BUFX2_615 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf11) );
  BUFX2 BUFX2_616 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf10) );
  BUFX2 BUFX2_617 ( .A(u2__abc_44228_n2966_hier0_bF_buf1), .Y(u2__abc_44228_n2966_bF_buf9) );
  BUFX2 BUFX2_618 ( .A(u2__abc_44228_n2966_hier0_bF_buf0), .Y(u2__abc_44228_n2966_bF_buf8) );
  BUFX2 BUFX2_619 ( .A(u2__abc_44228_n2966_hier0_bF_buf9), .Y(u2__abc_44228_n2966_bF_buf7) );
  BUFX2 BUFX2_62 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf3) );
  BUFX2 BUFX2_620 ( .A(u2__abc_44228_n2966_hier0_bF_buf8), .Y(u2__abc_44228_n2966_bF_buf6) );
  BUFX2 BUFX2_621 ( .A(u2__abc_44228_n2966_hier0_bF_buf7), .Y(u2__abc_44228_n2966_bF_buf5) );
  BUFX2 BUFX2_622 ( .A(u2__abc_44228_n2966_hier0_bF_buf6), .Y(u2__abc_44228_n2966_bF_buf4) );
  BUFX2 BUFX2_623 ( .A(u2__abc_44228_n2966_hier0_bF_buf5), .Y(u2__abc_44228_n2966_bF_buf3) );
  BUFX2 BUFX2_624 ( .A(u2__abc_44228_n2966_hier0_bF_buf4), .Y(u2__abc_44228_n2966_bF_buf2) );
  BUFX2 BUFX2_625 ( .A(u2__abc_44228_n2966_hier0_bF_buf3), .Y(u2__abc_44228_n2966_bF_buf1) );
  BUFX2 BUFX2_626 ( .A(u2__abc_44228_n2966_hier0_bF_buf2), .Y(u2__abc_44228_n2966_bF_buf0) );
  BUFX2 BUFX2_627 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf57) );
  BUFX2 BUFX2_628 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf56) );
  BUFX2 BUFX2_629 ( .A(u2__abc_44228_n7547_hier0_bF_buf4), .Y(u2__abc_44228_n7547_bF_buf55) );
  BUFX2 BUFX2_63 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf2) );
  BUFX2 BUFX2_630 ( .A(u2__abc_44228_n7547_hier0_bF_buf3), .Y(u2__abc_44228_n7547_bF_buf54) );
  BUFX2 BUFX2_631 ( .A(u2__abc_44228_n7547_hier0_bF_buf2), .Y(u2__abc_44228_n7547_bF_buf53) );
  BUFX2 BUFX2_632 ( .A(u2__abc_44228_n7547_hier0_bF_buf1), .Y(u2__abc_44228_n7547_bF_buf52) );
  BUFX2 BUFX2_633 ( .A(u2__abc_44228_n7547_hier0_bF_buf0), .Y(u2__abc_44228_n7547_bF_buf51) );
  BUFX2 BUFX2_634 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf50) );
  BUFX2 BUFX2_635 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf49) );
  BUFX2 BUFX2_636 ( .A(u2__abc_44228_n7547_hier0_bF_buf4), .Y(u2__abc_44228_n7547_bF_buf48) );
  BUFX2 BUFX2_637 ( .A(u2__abc_44228_n7547_hier0_bF_buf3), .Y(u2__abc_44228_n7547_bF_buf47) );
  BUFX2 BUFX2_638 ( .A(u2__abc_44228_n7547_hier0_bF_buf2), .Y(u2__abc_44228_n7547_bF_buf46) );
  BUFX2 BUFX2_639 ( .A(u2__abc_44228_n7547_hier0_bF_buf1), .Y(u2__abc_44228_n7547_bF_buf45) );
  BUFX2 BUFX2_64 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf1) );
  BUFX2 BUFX2_640 ( .A(u2__abc_44228_n7547_hier0_bF_buf0), .Y(u2__abc_44228_n7547_bF_buf44) );
  BUFX2 BUFX2_641 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf43) );
  BUFX2 BUFX2_642 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf42) );
  BUFX2 BUFX2_643 ( .A(u2__abc_44228_n7547_hier0_bF_buf4), .Y(u2__abc_44228_n7547_bF_buf41) );
  BUFX2 BUFX2_644 ( .A(u2__abc_44228_n7547_hier0_bF_buf3), .Y(u2__abc_44228_n7547_bF_buf40) );
  BUFX2 BUFX2_645 ( .A(u2__abc_44228_n7547_hier0_bF_buf2), .Y(u2__abc_44228_n7547_bF_buf39) );
  BUFX2 BUFX2_646 ( .A(u2__abc_44228_n7547_hier0_bF_buf1), .Y(u2__abc_44228_n7547_bF_buf38) );
  BUFX2 BUFX2_647 ( .A(u2__abc_44228_n7547_hier0_bF_buf0), .Y(u2__abc_44228_n7547_bF_buf37) );
  BUFX2 BUFX2_648 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf36) );
  BUFX2 BUFX2_649 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf35) );
  BUFX2 BUFX2_65 ( .A(u2__abc_44228_n2983), .Y(u2__abc_44228_n2983_hier0_bF_buf0) );
  BUFX2 BUFX2_650 ( .A(u2__abc_44228_n7547_hier0_bF_buf4), .Y(u2__abc_44228_n7547_bF_buf34) );
  BUFX2 BUFX2_651 ( .A(u2__abc_44228_n7547_hier0_bF_buf3), .Y(u2__abc_44228_n7547_bF_buf33) );
  BUFX2 BUFX2_652 ( .A(u2__abc_44228_n7547_hier0_bF_buf2), .Y(u2__abc_44228_n7547_bF_buf32) );
  BUFX2 BUFX2_653 ( .A(u2__abc_44228_n7547_hier0_bF_buf1), .Y(u2__abc_44228_n7547_bF_buf31) );
  BUFX2 BUFX2_654 ( .A(u2__abc_44228_n7547_hier0_bF_buf0), .Y(u2__abc_44228_n7547_bF_buf30) );
  BUFX2 BUFX2_655 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf29) );
  BUFX2 BUFX2_656 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf28) );
  BUFX2 BUFX2_657 ( .A(u2__abc_44228_n7547_hier0_bF_buf4), .Y(u2__abc_44228_n7547_bF_buf27) );
  BUFX2 BUFX2_658 ( .A(u2__abc_44228_n7547_hier0_bF_buf3), .Y(u2__abc_44228_n7547_bF_buf26) );
  BUFX2 BUFX2_659 ( .A(u2__abc_44228_n7547_hier0_bF_buf2), .Y(u2__abc_44228_n7547_bF_buf25) );
  BUFX2 BUFX2_66 ( .A(u2__abc_44228_n15402), .Y(u2__abc_44228_n15402_bF_buf3) );
  BUFX2 BUFX2_660 ( .A(u2__abc_44228_n7547_hier0_bF_buf1), .Y(u2__abc_44228_n7547_bF_buf24) );
  BUFX2 BUFX2_661 ( .A(u2__abc_44228_n7547_hier0_bF_buf0), .Y(u2__abc_44228_n7547_bF_buf23) );
  BUFX2 BUFX2_662 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf22) );
  BUFX2 BUFX2_663 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf21) );
  BUFX2 BUFX2_664 ( .A(u2__abc_44228_n7547_hier0_bF_buf4), .Y(u2__abc_44228_n7547_bF_buf20) );
  BUFX2 BUFX2_665 ( .A(u2__abc_44228_n7547_hier0_bF_buf3), .Y(u2__abc_44228_n7547_bF_buf19) );
  BUFX2 BUFX2_666 ( .A(u2__abc_44228_n7547_hier0_bF_buf2), .Y(u2__abc_44228_n7547_bF_buf18) );
  BUFX2 BUFX2_667 ( .A(u2__abc_44228_n7547_hier0_bF_buf1), .Y(u2__abc_44228_n7547_bF_buf17) );
  BUFX2 BUFX2_668 ( .A(u2__abc_44228_n7547_hier0_bF_buf0), .Y(u2__abc_44228_n7547_bF_buf16) );
  BUFX2 BUFX2_669 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf15) );
  BUFX2 BUFX2_67 ( .A(u2__abc_44228_n15402), .Y(u2__abc_44228_n15402_bF_buf2) );
  BUFX2 BUFX2_670 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf14) );
  BUFX2 BUFX2_671 ( .A(u2__abc_44228_n7547_hier0_bF_buf4), .Y(u2__abc_44228_n7547_bF_buf13) );
  BUFX2 BUFX2_672 ( .A(u2__abc_44228_n7547_hier0_bF_buf3), .Y(u2__abc_44228_n7547_bF_buf12) );
  BUFX2 BUFX2_673 ( .A(u2__abc_44228_n7547_hier0_bF_buf2), .Y(u2__abc_44228_n7547_bF_buf11) );
  BUFX2 BUFX2_674 ( .A(u2__abc_44228_n7547_hier0_bF_buf1), .Y(u2__abc_44228_n7547_bF_buf10) );
  BUFX2 BUFX2_675 ( .A(u2__abc_44228_n7547_hier0_bF_buf0), .Y(u2__abc_44228_n7547_bF_buf9) );
  BUFX2 BUFX2_676 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf8) );
  BUFX2 BUFX2_677 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf7) );
  BUFX2 BUFX2_678 ( .A(u2__abc_44228_n7547_hier0_bF_buf4), .Y(u2__abc_44228_n7547_bF_buf6) );
  BUFX2 BUFX2_679 ( .A(u2__abc_44228_n7547_hier0_bF_buf3), .Y(u2__abc_44228_n7547_bF_buf5) );
  BUFX2 BUFX2_68 ( .A(u2__abc_44228_n15402), .Y(u2__abc_44228_n15402_bF_buf1) );
  BUFX2 BUFX2_680 ( .A(u2__abc_44228_n7547_hier0_bF_buf2), .Y(u2__abc_44228_n7547_bF_buf4) );
  BUFX2 BUFX2_681 ( .A(u2__abc_44228_n7547_hier0_bF_buf1), .Y(u2__abc_44228_n7547_bF_buf3) );
  BUFX2 BUFX2_682 ( .A(u2__abc_44228_n7547_hier0_bF_buf0), .Y(u2__abc_44228_n7547_bF_buf2) );
  BUFX2 BUFX2_683 ( .A(u2__abc_44228_n7547_hier0_bF_buf6), .Y(u2__abc_44228_n7547_bF_buf1) );
  BUFX2 BUFX2_684 ( .A(u2__abc_44228_n7547_hier0_bF_buf5), .Y(u2__abc_44228_n7547_bF_buf0) );
  BUFX2 BUFX2_685 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf13) );
  BUFX2 BUFX2_686 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf12) );
  BUFX2 BUFX2_687 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf11) );
  BUFX2 BUFX2_688 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf10) );
  BUFX2 BUFX2_689 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf9) );
  BUFX2 BUFX2_69 ( .A(u2__abc_44228_n15402), .Y(u2__abc_44228_n15402_bF_buf0) );
  BUFX2 BUFX2_690 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf8) );
  BUFX2 BUFX2_691 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf7) );
  BUFX2 BUFX2_692 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf6) );
  BUFX2 BUFX2_693 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf5) );
  BUFX2 BUFX2_694 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf4) );
  BUFX2 BUFX2_695 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf3) );
  BUFX2 BUFX2_696 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf2) );
  BUFX2 BUFX2_697 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf1) );
  BUFX2 BUFX2_698 ( .A(_abc_64468_n753), .Y(_abc_64468_n753_bF_buf0) );
  BUFX2 BUFX2_699 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf141) );
  BUFX2 BUFX2_7 ( .A(u2__abc_44228_n7548_1), .Y(u2__abc_44228_n7548_1_hier0_bF_buf0) );
  BUFX2 BUFX2_70 ( .A(u2__abc_44228_n15403), .Y(u2__abc_44228_n15403_bF_buf3) );
  BUFX2 BUFX2_700 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf140) );
  BUFX2 BUFX2_701 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf139) );
  BUFX2 BUFX2_702 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf138) );
  BUFX2 BUFX2_703 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf137) );
  BUFX2 BUFX2_704 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf136) );
  BUFX2 BUFX2_705 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf135) );
  BUFX2 BUFX2_706 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf134) );
  BUFX2 BUFX2_707 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf133) );
  BUFX2 BUFX2_708 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf132) );
  BUFX2 BUFX2_709 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf131) );
  BUFX2 BUFX2_71 ( .A(u2__abc_44228_n15403), .Y(u2__abc_44228_n15403_bF_buf2) );
  BUFX2 BUFX2_710 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf130) );
  BUFX2 BUFX2_711 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf129) );
  BUFX2 BUFX2_712 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf128) );
  BUFX2 BUFX2_713 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf127) );
  BUFX2 BUFX2_714 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf126) );
  BUFX2 BUFX2_715 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf125) );
  BUFX2 BUFX2_716 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf124) );
  BUFX2 BUFX2_717 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf123) );
  BUFX2 BUFX2_718 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf122) );
  BUFX2 BUFX2_719 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf121) );
  BUFX2 BUFX2_72 ( .A(u2__abc_44228_n15403), .Y(u2__abc_44228_n15403_bF_buf1) );
  BUFX2 BUFX2_720 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf120) );
  BUFX2 BUFX2_721 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf119) );
  BUFX2 BUFX2_722 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf118) );
  BUFX2 BUFX2_723 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf117) );
  BUFX2 BUFX2_724 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf116) );
  BUFX2 BUFX2_725 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf115) );
  BUFX2 BUFX2_726 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf114) );
  BUFX2 BUFX2_727 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf113) );
  BUFX2 BUFX2_728 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf112) );
  BUFX2 BUFX2_729 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf111) );
  BUFX2 BUFX2_73 ( .A(u2__abc_44228_n15403), .Y(u2__abc_44228_n15403_bF_buf0) );
  BUFX2 BUFX2_730 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf110) );
  BUFX2 BUFX2_731 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf109) );
  BUFX2 BUFX2_732 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf108) );
  BUFX2 BUFX2_733 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf107) );
  BUFX2 BUFX2_734 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf106) );
  BUFX2 BUFX2_735 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf105) );
  BUFX2 BUFX2_736 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf104) );
  BUFX2 BUFX2_737 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf103) );
  BUFX2 BUFX2_738 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf102) );
  BUFX2 BUFX2_739 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf101) );
  BUFX2 BUFX2_74 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf13) );
  BUFX2 BUFX2_740 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf100) );
  BUFX2 BUFX2_741 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf99) );
  BUFX2 BUFX2_742 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf98) );
  BUFX2 BUFX2_743 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf97) );
  BUFX2 BUFX2_744 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf96) );
  BUFX2 BUFX2_745 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf95) );
  BUFX2 BUFX2_746 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf94) );
  BUFX2 BUFX2_747 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf93) );
  BUFX2 BUFX2_748 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf92) );
  BUFX2 BUFX2_749 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf91) );
  BUFX2 BUFX2_75 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf12) );
  BUFX2 BUFX2_750 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf90) );
  BUFX2 BUFX2_751 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf89) );
  BUFX2 BUFX2_752 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf88) );
  BUFX2 BUFX2_753 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf87) );
  BUFX2 BUFX2_754 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf86) );
  BUFX2 BUFX2_755 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf85) );
  BUFX2 BUFX2_756 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf84) );
  BUFX2 BUFX2_757 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf83) );
  BUFX2 BUFX2_758 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf82) );
  BUFX2 BUFX2_759 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf81) );
  BUFX2 BUFX2_76 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf11) );
  BUFX2 BUFX2_760 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf80) );
  BUFX2 BUFX2_761 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf79) );
  BUFX2 BUFX2_762 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf78) );
  BUFX2 BUFX2_763 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf77) );
  BUFX2 BUFX2_764 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf76) );
  BUFX2 BUFX2_765 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf75) );
  BUFX2 BUFX2_766 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf74) );
  BUFX2 BUFX2_767 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf73) );
  BUFX2 BUFX2_768 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf72) );
  BUFX2 BUFX2_769 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf71) );
  BUFX2 BUFX2_77 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf10) );
  BUFX2 BUFX2_770 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf70) );
  BUFX2 BUFX2_771 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf69) );
  BUFX2 BUFX2_772 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf68) );
  BUFX2 BUFX2_773 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf67) );
  BUFX2 BUFX2_774 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf66) );
  BUFX2 BUFX2_775 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf65) );
  BUFX2 BUFX2_776 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf64) );
  BUFX2 BUFX2_777 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf63) );
  BUFX2 BUFX2_778 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf62) );
  BUFX2 BUFX2_779 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf61) );
  BUFX2 BUFX2_78 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf9) );
  BUFX2 BUFX2_780 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf60) );
  BUFX2 BUFX2_781 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf59) );
  BUFX2 BUFX2_782 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf58) );
  BUFX2 BUFX2_783 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf57) );
  BUFX2 BUFX2_784 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf56) );
  BUFX2 BUFX2_785 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf55) );
  BUFX2 BUFX2_786 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf54) );
  BUFX2 BUFX2_787 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf53) );
  BUFX2 BUFX2_788 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf52) );
  BUFX2 BUFX2_789 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf51) );
  BUFX2 BUFX2_79 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf8) );
  BUFX2 BUFX2_790 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf50) );
  BUFX2 BUFX2_791 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf49) );
  BUFX2 BUFX2_792 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf48) );
  BUFX2 BUFX2_793 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf47) );
  BUFX2 BUFX2_794 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf46) );
  BUFX2 BUFX2_795 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf45) );
  BUFX2 BUFX2_796 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf44) );
  BUFX2 BUFX2_797 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf43) );
  BUFX2 BUFX2_798 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf42) );
  BUFX2 BUFX2_799 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf41) );
  BUFX2 BUFX2_8 ( .A(clk), .Y(clk_hier0_bF_buf10) );
  BUFX2 BUFX2_80 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf7) );
  BUFX2 BUFX2_800 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf40) );
  BUFX2 BUFX2_801 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf39) );
  BUFX2 BUFX2_802 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf38) );
  BUFX2 BUFX2_803 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf37) );
  BUFX2 BUFX2_804 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf36) );
  BUFX2 BUFX2_805 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf35) );
  BUFX2 BUFX2_806 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf34) );
  BUFX2 BUFX2_807 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf33) );
  BUFX2 BUFX2_808 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf32) );
  BUFX2 BUFX2_809 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf31) );
  BUFX2 BUFX2_81 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf6) );
  BUFX2 BUFX2_810 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf30) );
  BUFX2 BUFX2_811 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf29) );
  BUFX2 BUFX2_812 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf28) );
  BUFX2 BUFX2_813 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf27) );
  BUFX2 BUFX2_814 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf26) );
  BUFX2 BUFX2_815 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf25) );
  BUFX2 BUFX2_816 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf24) );
  BUFX2 BUFX2_817 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf23) );
  BUFX2 BUFX2_818 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf22) );
  BUFX2 BUFX2_819 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf21) );
  BUFX2 BUFX2_82 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf5) );
  BUFX2 BUFX2_820 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf20) );
  BUFX2 BUFX2_821 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf19) );
  BUFX2 BUFX2_822 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf18) );
  BUFX2 BUFX2_823 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf17) );
  BUFX2 BUFX2_824 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf16) );
  BUFX2 BUFX2_825 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf15) );
  BUFX2 BUFX2_826 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf14) );
  BUFX2 BUFX2_827 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf13) );
  BUFX2 BUFX2_828 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf12) );
  BUFX2 BUFX2_829 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf11) );
  BUFX2 BUFX2_83 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf4) );
  BUFX2 BUFX2_830 ( .A(u2__abc_44228_n2983_hier0_bF_buf0), .Y(u2__abc_44228_n2983_bF_buf10) );
  BUFX2 BUFX2_831 ( .A(u2__abc_44228_n2983_hier0_bF_buf10), .Y(u2__abc_44228_n2983_bF_buf9) );
  BUFX2 BUFX2_832 ( .A(u2__abc_44228_n2983_hier0_bF_buf9), .Y(u2__abc_44228_n2983_bF_buf8) );
  BUFX2 BUFX2_833 ( .A(u2__abc_44228_n2983_hier0_bF_buf8), .Y(u2__abc_44228_n2983_bF_buf7) );
  BUFX2 BUFX2_834 ( .A(u2__abc_44228_n2983_hier0_bF_buf7), .Y(u2__abc_44228_n2983_bF_buf6) );
  BUFX2 BUFX2_835 ( .A(u2__abc_44228_n2983_hier0_bF_buf6), .Y(u2__abc_44228_n2983_bF_buf5) );
  BUFX2 BUFX2_836 ( .A(u2__abc_44228_n2983_hier0_bF_buf5), .Y(u2__abc_44228_n2983_bF_buf4) );
  BUFX2 BUFX2_837 ( .A(u2__abc_44228_n2983_hier0_bF_buf4), .Y(u2__abc_44228_n2983_bF_buf3) );
  BUFX2 BUFX2_838 ( .A(u2__abc_44228_n2983_hier0_bF_buf3), .Y(u2__abc_44228_n2983_bF_buf2) );
  BUFX2 BUFX2_839 ( .A(u2__abc_44228_n2983_hier0_bF_buf2), .Y(u2__abc_44228_n2983_bF_buf1) );
  BUFX2 BUFX2_84 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf3) );
  BUFX2 BUFX2_840 ( .A(u2__abc_44228_n2983_hier0_bF_buf1), .Y(u2__abc_44228_n2983_bF_buf0) );
  BUFX2 BUFX2_841 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf14) );
  BUFX2 BUFX2_842 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf13) );
  BUFX2 BUFX2_843 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf12) );
  BUFX2 BUFX2_844 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf11) );
  BUFX2 BUFX2_845 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf10) );
  BUFX2 BUFX2_846 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf9) );
  BUFX2 BUFX2_847 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf8) );
  BUFX2 BUFX2_848 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf7) );
  BUFX2 BUFX2_849 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf6) );
  BUFX2 BUFX2_85 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf2) );
  BUFX2 BUFX2_850 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf5) );
  BUFX2 BUFX2_851 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf4) );
  BUFX2 BUFX2_852 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf3) );
  BUFX2 BUFX2_853 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf2) );
  BUFX2 BUFX2_854 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf1) );
  BUFX2 BUFX2_855 ( .A(u2__abc_44228_n2984), .Y(u2__abc_44228_n2984_bF_buf0) );
  BUFX2 BUFX2_856 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf14) );
  BUFX2 BUFX2_857 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf13) );
  BUFX2 BUFX2_858 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf12) );
  BUFX2 BUFX2_859 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf11) );
  BUFX2 BUFX2_86 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf1) );
  BUFX2 BUFX2_860 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf10) );
  BUFX2 BUFX2_861 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf9) );
  BUFX2 BUFX2_862 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf8) );
  BUFX2 BUFX2_863 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf7) );
  BUFX2 BUFX2_864 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf6) );
  BUFX2 BUFX2_865 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf5) );
  BUFX2 BUFX2_866 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf4) );
  BUFX2 BUFX2_867 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf3) );
  BUFX2 BUFX2_868 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf2) );
  BUFX2 BUFX2_869 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf1) );
  BUFX2 BUFX2_87 ( .A(u2__abc_44228_n15405), .Y(u2__abc_44228_n15405_bF_buf0) );
  BUFX2 BUFX2_870 ( .A(u2__abc_44228_n2987), .Y(u2__abc_44228_n2987_bF_buf0) );
  BUFX2 BUFX2_871 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf13) );
  BUFX2 BUFX2_872 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf12) );
  BUFX2 BUFX2_873 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf11) );
  BUFX2 BUFX2_874 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf10) );
  BUFX2 BUFX2_875 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf9) );
  BUFX2 BUFX2_876 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf8) );
  BUFX2 BUFX2_877 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf7) );
  BUFX2 BUFX2_878 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf6) );
  BUFX2 BUFX2_879 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf5) );
  BUFX2 BUFX2_88 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf14) );
  BUFX2 BUFX2_880 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf4) );
  BUFX2 BUFX2_881 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf3) );
  BUFX2 BUFX2_882 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf2) );
  BUFX2 BUFX2_883 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf1) );
  BUFX2 BUFX2_884 ( .A(u2__abc_44228_n2988), .Y(u2__abc_44228_n2988_bF_buf0) );
  BUFX2 BUFX2_885 ( .A(u2__abc_44228_n2989), .Y(u2__abc_44228_n2989_bF_buf3) );
  BUFX2 BUFX2_886 ( .A(u2__abc_44228_n2989), .Y(u2__abc_44228_n2989_bF_buf2) );
  BUFX2 BUFX2_887 ( .A(u2__abc_44228_n2989), .Y(u2__abc_44228_n2989_bF_buf1) );
  BUFX2 BUFX2_888 ( .A(u2__abc_44228_n2989), .Y(u2__abc_44228_n2989_bF_buf0) );
  BUFX2 BUFX2_889 ( .A(\a[112] ), .Y(a_112_bF_buf9) );
  BUFX2 BUFX2_89 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf13) );
  BUFX2 BUFX2_890 ( .A(\a[112] ), .Y(a_112_bF_buf8) );
  BUFX2 BUFX2_891 ( .A(\a[112] ), .Y(a_112_bF_buf7) );
  BUFX2 BUFX2_892 ( .A(\a[112] ), .Y(a_112_bF_buf6) );
  BUFX2 BUFX2_893 ( .A(\a[112] ), .Y(a_112_bF_buf5) );
  BUFX2 BUFX2_894 ( .A(\a[112] ), .Y(a_112_bF_buf4) );
  BUFX2 BUFX2_895 ( .A(\a[112] ), .Y(a_112_bF_buf3) );
  BUFX2 BUFX2_896 ( .A(\a[112] ), .Y(a_112_bF_buf2) );
  BUFX2 BUFX2_897 ( .A(\a[112] ), .Y(a_112_bF_buf1) );
  BUFX2 BUFX2_898 ( .A(\a[112] ), .Y(a_112_bF_buf0) );
  BUFX2 BUFX2_899 ( .A(aNan), .Y(aNan_bF_buf10) );
  BUFX2 BUFX2_9 ( .A(clk), .Y(clk_hier0_bF_buf9) );
  BUFX2 BUFX2_90 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf12) );
  BUFX2 BUFX2_900 ( .A(aNan), .Y(aNan_bF_buf9) );
  BUFX2 BUFX2_901 ( .A(aNan), .Y(aNan_bF_buf8) );
  BUFX2 BUFX2_902 ( .A(aNan), .Y(aNan_bF_buf7) );
  BUFX2 BUFX2_903 ( .A(aNan), .Y(aNan_bF_buf6) );
  BUFX2 BUFX2_904 ( .A(aNan), .Y(aNan_bF_buf5) );
  BUFX2 BUFX2_905 ( .A(aNan), .Y(aNan_bF_buf4) );
  BUFX2 BUFX2_906 ( .A(aNan), .Y(aNan_bF_buf3) );
  BUFX2 BUFX2_907 ( .A(aNan), .Y(aNan_bF_buf2) );
  BUFX2 BUFX2_908 ( .A(aNan), .Y(aNan_bF_buf1) );
  BUFX2 BUFX2_909 ( .A(aNan), .Y(aNan_bF_buf0) );
  BUFX2 BUFX2_91 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf11) );
  BUFX2 BUFX2_910 ( .A(_auto_iopadmap_cc_313_execute_65412), .Y(done) );
  BUFX2 BUFX2_911 ( .A(1'b0), .Y(\o[0] ) );
  BUFX2 BUFX2_912 ( .A(1'b0), .Y(\o[1] ) );
  BUFX2 BUFX2_913 ( .A(1'b0), .Y(\o[2] ) );
  BUFX2 BUFX2_914 ( .A(1'b0), .Y(\o[3] ) );
  BUFX2 BUFX2_915 ( .A(1'b0), .Y(\o[4] ) );
  BUFX2 BUFX2_916 ( .A(1'b0), .Y(\o[5] ) );
  BUFX2 BUFX2_917 ( .A(1'b0), .Y(\o[6] ) );
  BUFX2 BUFX2_918 ( .A(1'b0), .Y(\o[7] ) );
  BUFX2 BUFX2_919 ( .A(1'b0), .Y(\o[8] ) );
  BUFX2 BUFX2_92 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf10) );
  BUFX2 BUFX2_920 ( .A(1'b0), .Y(\o[9] ) );
  BUFX2 BUFX2_921 ( .A(1'b0), .Y(\o[10] ) );
  BUFX2 BUFX2_922 ( .A(1'b0), .Y(\o[11] ) );
  BUFX2 BUFX2_923 ( .A(1'b0), .Y(\o[12] ) );
  BUFX2 BUFX2_924 ( .A(1'b0), .Y(\o[13] ) );
  BUFX2 BUFX2_925 ( .A(1'b0), .Y(\o[14] ) );
  BUFX2 BUFX2_926 ( .A(1'b0), .Y(\o[15] ) );
  BUFX2 BUFX2_927 ( .A(1'b0), .Y(\o[16] ) );
  BUFX2 BUFX2_928 ( .A(1'b0), .Y(\o[17] ) );
  BUFX2 BUFX2_929 ( .A(1'b0), .Y(\o[18] ) );
  BUFX2 BUFX2_93 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf9) );
  BUFX2 BUFX2_930 ( .A(1'b0), .Y(\o[19] ) );
  BUFX2 BUFX2_931 ( .A(1'b0), .Y(\o[20] ) );
  BUFX2 BUFX2_932 ( .A(1'b0), .Y(\o[21] ) );
  BUFX2 BUFX2_933 ( .A(1'b0), .Y(\o[22] ) );
  BUFX2 BUFX2_934 ( .A(1'b0), .Y(\o[23] ) );
  BUFX2 BUFX2_935 ( .A(1'b0), .Y(\o[24] ) );
  BUFX2 BUFX2_936 ( .A(1'b0), .Y(\o[25] ) );
  BUFX2 BUFX2_937 ( .A(1'b0), .Y(\o[26] ) );
  BUFX2 BUFX2_938 ( .A(1'b0), .Y(\o[27] ) );
  BUFX2 BUFX2_939 ( .A(1'b0), .Y(\o[28] ) );
  BUFX2 BUFX2_94 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf8) );
  BUFX2 BUFX2_940 ( .A(1'b0), .Y(\o[29] ) );
  BUFX2 BUFX2_941 ( .A(1'b0), .Y(\o[30] ) );
  BUFX2 BUFX2_942 ( .A(1'b0), .Y(\o[31] ) );
  BUFX2 BUFX2_943 ( .A(1'b0), .Y(\o[32] ) );
  BUFX2 BUFX2_944 ( .A(1'b0), .Y(\o[33] ) );
  BUFX2 BUFX2_945 ( .A(1'b0), .Y(\o[34] ) );
  BUFX2 BUFX2_946 ( .A(1'b0), .Y(\o[35] ) );
  BUFX2 BUFX2_947 ( .A(_auto_iopadmap_cc_313_execute_65414_36_), .Y(\o[36] ) );
  BUFX2 BUFX2_948 ( .A(_auto_iopadmap_cc_313_execute_65414_37_), .Y(\o[37] ) );
  BUFX2 BUFX2_949 ( .A(_auto_iopadmap_cc_313_execute_65414_38_), .Y(\o[38] ) );
  BUFX2 BUFX2_95 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf7) );
  BUFX2 BUFX2_950 ( .A(_auto_iopadmap_cc_313_execute_65414_39_), .Y(\o[39] ) );
  BUFX2 BUFX2_951 ( .A(_auto_iopadmap_cc_313_execute_65414_40_), .Y(\o[40] ) );
  BUFX2 BUFX2_952 ( .A(_auto_iopadmap_cc_313_execute_65414_41_), .Y(\o[41] ) );
  BUFX2 BUFX2_953 ( .A(_auto_iopadmap_cc_313_execute_65414_42_), .Y(\o[42] ) );
  BUFX2 BUFX2_954 ( .A(_auto_iopadmap_cc_313_execute_65414_43_), .Y(\o[43] ) );
  BUFX2 BUFX2_955 ( .A(_auto_iopadmap_cc_313_execute_65414_44_), .Y(\o[44] ) );
  BUFX2 BUFX2_956 ( .A(_auto_iopadmap_cc_313_execute_65414_45_), .Y(\o[45] ) );
  BUFX2 BUFX2_957 ( .A(_auto_iopadmap_cc_313_execute_65414_46_), .Y(\o[46] ) );
  BUFX2 BUFX2_958 ( .A(_auto_iopadmap_cc_313_execute_65414_47_), .Y(\o[47] ) );
  BUFX2 BUFX2_959 ( .A(_auto_iopadmap_cc_313_execute_65414_48_), .Y(\o[48] ) );
  BUFX2 BUFX2_96 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf6) );
  BUFX2 BUFX2_960 ( .A(_auto_iopadmap_cc_313_execute_65414_49_), .Y(\o[49] ) );
  BUFX2 BUFX2_961 ( .A(_auto_iopadmap_cc_313_execute_65414_50_), .Y(\o[50] ) );
  BUFX2 BUFX2_962 ( .A(_auto_iopadmap_cc_313_execute_65414_51_), .Y(\o[51] ) );
  BUFX2 BUFX2_963 ( .A(_auto_iopadmap_cc_313_execute_65414_52_), .Y(\o[52] ) );
  BUFX2 BUFX2_964 ( .A(_auto_iopadmap_cc_313_execute_65414_53_), .Y(\o[53] ) );
  BUFX2 BUFX2_965 ( .A(_auto_iopadmap_cc_313_execute_65414_54_), .Y(\o[54] ) );
  BUFX2 BUFX2_966 ( .A(_auto_iopadmap_cc_313_execute_65414_55_), .Y(\o[55] ) );
  BUFX2 BUFX2_967 ( .A(_auto_iopadmap_cc_313_execute_65414_56_), .Y(\o[56] ) );
  BUFX2 BUFX2_968 ( .A(_auto_iopadmap_cc_313_execute_65414_57_), .Y(\o[57] ) );
  BUFX2 BUFX2_969 ( .A(_auto_iopadmap_cc_313_execute_65414_58_), .Y(\o[58] ) );
  BUFX2 BUFX2_97 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf5) );
  BUFX2 BUFX2_970 ( .A(_auto_iopadmap_cc_313_execute_65414_59_), .Y(\o[59] ) );
  BUFX2 BUFX2_971 ( .A(_auto_iopadmap_cc_313_execute_65414_60_), .Y(\o[60] ) );
  BUFX2 BUFX2_972 ( .A(_auto_iopadmap_cc_313_execute_65414_61_), .Y(\o[61] ) );
  BUFX2 BUFX2_973 ( .A(_auto_iopadmap_cc_313_execute_65414_62_), .Y(\o[62] ) );
  BUFX2 BUFX2_974 ( .A(_auto_iopadmap_cc_313_execute_65414_63_), .Y(\o[63] ) );
  BUFX2 BUFX2_975 ( .A(_auto_iopadmap_cc_313_execute_65414_64_), .Y(\o[64] ) );
  BUFX2 BUFX2_976 ( .A(_auto_iopadmap_cc_313_execute_65414_65_), .Y(\o[65] ) );
  BUFX2 BUFX2_977 ( .A(_auto_iopadmap_cc_313_execute_65414_66_), .Y(\o[66] ) );
  BUFX2 BUFX2_978 ( .A(_auto_iopadmap_cc_313_execute_65414_67_), .Y(\o[67] ) );
  BUFX2 BUFX2_979 ( .A(_auto_iopadmap_cc_313_execute_65414_68_), .Y(\o[68] ) );
  BUFX2 BUFX2_98 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf4) );
  BUFX2 BUFX2_980 ( .A(_auto_iopadmap_cc_313_execute_65414_69_), .Y(\o[69] ) );
  BUFX2 BUFX2_981 ( .A(_auto_iopadmap_cc_313_execute_65414_70_), .Y(\o[70] ) );
  BUFX2 BUFX2_982 ( .A(_auto_iopadmap_cc_313_execute_65414_71_), .Y(\o[71] ) );
  BUFX2 BUFX2_983 ( .A(_auto_iopadmap_cc_313_execute_65414_72_), .Y(\o[72] ) );
  BUFX2 BUFX2_984 ( .A(_auto_iopadmap_cc_313_execute_65414_73_), .Y(\o[73] ) );
  BUFX2 BUFX2_985 ( .A(_auto_iopadmap_cc_313_execute_65414_74_), .Y(\o[74] ) );
  BUFX2 BUFX2_986 ( .A(_auto_iopadmap_cc_313_execute_65414_75_), .Y(\o[75] ) );
  BUFX2 BUFX2_987 ( .A(_auto_iopadmap_cc_313_execute_65414_76_), .Y(\o[76] ) );
  BUFX2 BUFX2_988 ( .A(_auto_iopadmap_cc_313_execute_65414_77_), .Y(\o[77] ) );
  BUFX2 BUFX2_989 ( .A(_auto_iopadmap_cc_313_execute_65414_78_), .Y(\o[78] ) );
  BUFX2 BUFX2_99 ( .A(u2__abc_44228_n15408), .Y(u2__abc_44228_n15408_bF_buf3) );
  BUFX2 BUFX2_990 ( .A(_auto_iopadmap_cc_313_execute_65414_79_), .Y(\o[79] ) );
  BUFX2 BUFX2_991 ( .A(_auto_iopadmap_cc_313_execute_65414_80_), .Y(\o[80] ) );
  BUFX2 BUFX2_992 ( .A(_auto_iopadmap_cc_313_execute_65414_81_), .Y(\o[81] ) );
  BUFX2 BUFX2_993 ( .A(_auto_iopadmap_cc_313_execute_65414_82_), .Y(\o[82] ) );
  BUFX2 BUFX2_994 ( .A(_auto_iopadmap_cc_313_execute_65414_83_), .Y(\o[83] ) );
  BUFX2 BUFX2_995 ( .A(_auto_iopadmap_cc_313_execute_65414_84_), .Y(\o[84] ) );
  BUFX2 BUFX2_996 ( .A(_auto_iopadmap_cc_313_execute_65414_85_), .Y(\o[85] ) );
  BUFX2 BUFX2_997 ( .A(_auto_iopadmap_cc_313_execute_65414_86_), .Y(\o[86] ) );
  BUFX2 BUFX2_998 ( .A(_auto_iopadmap_cc_313_execute_65414_87_), .Y(\o[87] ) );
  BUFX2 BUFX2_999 ( .A(_auto_iopadmap_cc_313_execute_65414_88_), .Y(\o[88] ) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf121), .D(u2__abc_29664_n1191), .Q(u2_state_0_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf112), .D(u2_root_6__FF_INPUT), .Q(sqrto_5_) );
  DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf22), .D(u2_root_96__FF_INPUT), .Q(sqrto_95_) );
  DFFPOSX1 DFFPOSX1_1000 ( .CLK(clk_bF_buf98), .D(u2_remHi_93__FF_INPUT), .Q(u2_remHi_93_) );
  DFFPOSX1 DFFPOSX1_1001 ( .CLK(clk_bF_buf97), .D(u2_remHi_94__FF_INPUT), .Q(u2_remHi_94_) );
  DFFPOSX1 DFFPOSX1_1002 ( .CLK(clk_bF_buf96), .D(u2_remHi_95__FF_INPUT), .Q(u2_remHi_95_) );
  DFFPOSX1 DFFPOSX1_1003 ( .CLK(clk_bF_buf95), .D(u2_remHi_96__FF_INPUT), .Q(u2_remHi_96_) );
  DFFPOSX1 DFFPOSX1_1004 ( .CLK(clk_bF_buf94), .D(u2_remHi_97__FF_INPUT), .Q(u2_remHi_97_) );
  DFFPOSX1 DFFPOSX1_1005 ( .CLK(clk_bF_buf93), .D(u2_remHi_98__FF_INPUT), .Q(u2_remHi_98_) );
  DFFPOSX1 DFFPOSX1_1006 ( .CLK(clk_bF_buf92), .D(u2_remHi_99__FF_INPUT), .Q(u2_remHi_99_) );
  DFFPOSX1 DFFPOSX1_1007 ( .CLK(clk_bF_buf91), .D(u2_remHi_100__FF_INPUT), .Q(u2_remHi_100_) );
  DFFPOSX1 DFFPOSX1_1008 ( .CLK(clk_bF_buf90), .D(u2_remHi_101__FF_INPUT), .Q(u2_remHi_101_) );
  DFFPOSX1 DFFPOSX1_1009 ( .CLK(clk_bF_buf89), .D(u2_remHi_102__FF_INPUT), .Q(u2_remHi_102_) );
  DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf21), .D(u2_root_97__FF_INPUT), .Q(sqrto_96_) );
  DFFPOSX1 DFFPOSX1_1010 ( .CLK(clk_bF_buf88), .D(u2_remHi_103__FF_INPUT), .Q(u2_remHi_103_) );
  DFFPOSX1 DFFPOSX1_1011 ( .CLK(clk_bF_buf87), .D(u2_remHi_104__FF_INPUT), .Q(u2_remHi_104_) );
  DFFPOSX1 DFFPOSX1_1012 ( .CLK(clk_bF_buf86), .D(u2_remHi_105__FF_INPUT), .Q(u2_remHi_105_) );
  DFFPOSX1 DFFPOSX1_1013 ( .CLK(clk_bF_buf85), .D(u2_remHi_106__FF_INPUT), .Q(u2_remHi_106_) );
  DFFPOSX1 DFFPOSX1_1014 ( .CLK(clk_bF_buf84), .D(u2_remHi_107__FF_INPUT), .Q(u2_remHi_107_) );
  DFFPOSX1 DFFPOSX1_1015 ( .CLK(clk_bF_buf83), .D(u2_remHi_108__FF_INPUT), .Q(u2_remHi_108_) );
  DFFPOSX1 DFFPOSX1_1016 ( .CLK(clk_bF_buf82), .D(u2_remHi_109__FF_INPUT), .Q(u2_remHi_109_) );
  DFFPOSX1 DFFPOSX1_1017 ( .CLK(clk_bF_buf81), .D(u2_remHi_110__FF_INPUT), .Q(u2_remHi_110_) );
  DFFPOSX1 DFFPOSX1_1018 ( .CLK(clk_bF_buf80), .D(u2_remHi_111__FF_INPUT), .Q(u2_remHi_111_) );
  DFFPOSX1 DFFPOSX1_1019 ( .CLK(clk_bF_buf79), .D(u2_remHi_112__FF_INPUT), .Q(u2_remHi_112_) );
  DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf20), .D(u2_root_98__FF_INPUT), .Q(sqrto_97_) );
  DFFPOSX1 DFFPOSX1_1020 ( .CLK(clk_bF_buf78), .D(u2_remHi_113__FF_INPUT), .Q(u2_remHi_113_) );
  DFFPOSX1 DFFPOSX1_1021 ( .CLK(clk_bF_buf77), .D(u2_remHi_114__FF_INPUT), .Q(u2_remHi_114_) );
  DFFPOSX1 DFFPOSX1_1022 ( .CLK(clk_bF_buf76), .D(u2_remHi_115__FF_INPUT), .Q(u2_remHi_115_) );
  DFFPOSX1 DFFPOSX1_1023 ( .CLK(clk_bF_buf75), .D(u2_remHi_116__FF_INPUT), .Q(u2_remHi_116_) );
  DFFPOSX1 DFFPOSX1_1024 ( .CLK(clk_bF_buf74), .D(u2_remHi_117__FF_INPUT), .Q(u2_remHi_117_) );
  DFFPOSX1 DFFPOSX1_1025 ( .CLK(clk_bF_buf73), .D(u2_remHi_118__FF_INPUT), .Q(u2_remHi_118_) );
  DFFPOSX1 DFFPOSX1_1026 ( .CLK(clk_bF_buf72), .D(u2_remHi_119__FF_INPUT), .Q(u2_remHi_119_) );
  DFFPOSX1 DFFPOSX1_1027 ( .CLK(clk_bF_buf71), .D(u2_remHi_120__FF_INPUT), .Q(u2_remHi_120_) );
  DFFPOSX1 DFFPOSX1_1028 ( .CLK(clk_bF_buf70), .D(u2_remHi_121__FF_INPUT), .Q(u2_remHi_121_) );
  DFFPOSX1 DFFPOSX1_1029 ( .CLK(clk_bF_buf69), .D(u2_remHi_122__FF_INPUT), .Q(u2_remHi_122_) );
  DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf19), .D(u2_root_99__FF_INPUT), .Q(sqrto_98_) );
  DFFPOSX1 DFFPOSX1_1030 ( .CLK(clk_bF_buf68), .D(u2_remHi_123__FF_INPUT), .Q(u2_remHi_123_) );
  DFFPOSX1 DFFPOSX1_1031 ( .CLK(clk_bF_buf67), .D(u2_remHi_124__FF_INPUT), .Q(u2_remHi_124_) );
  DFFPOSX1 DFFPOSX1_1032 ( .CLK(clk_bF_buf66), .D(u2_remHi_125__FF_INPUT), .Q(u2_remHi_125_) );
  DFFPOSX1 DFFPOSX1_1033 ( .CLK(clk_bF_buf65), .D(u2_remHi_126__FF_INPUT), .Q(u2_remHi_126_) );
  DFFPOSX1 DFFPOSX1_1034 ( .CLK(clk_bF_buf64), .D(u2_remHi_127__FF_INPUT), .Q(u2_remHi_127_) );
  DFFPOSX1 DFFPOSX1_1035 ( .CLK(clk_bF_buf63), .D(u2_remHi_128__FF_INPUT), .Q(u2_remHi_128_) );
  DFFPOSX1 DFFPOSX1_1036 ( .CLK(clk_bF_buf62), .D(u2_remHi_129__FF_INPUT), .Q(u2_remHi_129_) );
  DFFPOSX1 DFFPOSX1_1037 ( .CLK(clk_bF_buf61), .D(u2_remHi_130__FF_INPUT), .Q(u2_remHi_130_) );
  DFFPOSX1 DFFPOSX1_1038 ( .CLK(clk_bF_buf60), .D(u2_remHi_131__FF_INPUT), .Q(u2_remHi_131_) );
  DFFPOSX1 DFFPOSX1_1039 ( .CLK(clk_bF_buf59), .D(u2_remHi_132__FF_INPUT), .Q(u2_remHi_132_) );
  DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf18), .D(u2_root_100__FF_INPUT), .Q(sqrto_99_) );
  DFFPOSX1 DFFPOSX1_1040 ( .CLK(clk_bF_buf58), .D(u2_remHi_133__FF_INPUT), .Q(u2_remHi_133_) );
  DFFPOSX1 DFFPOSX1_1041 ( .CLK(clk_bF_buf57), .D(u2_remHi_134__FF_INPUT), .Q(u2_remHi_134_) );
  DFFPOSX1 DFFPOSX1_1042 ( .CLK(clk_bF_buf56), .D(u2_remHi_135__FF_INPUT), .Q(u2_remHi_135_) );
  DFFPOSX1 DFFPOSX1_1043 ( .CLK(clk_bF_buf55), .D(u2_remHi_136__FF_INPUT), .Q(u2_remHi_136_) );
  DFFPOSX1 DFFPOSX1_1044 ( .CLK(clk_bF_buf54), .D(u2_remHi_137__FF_INPUT), .Q(u2_remHi_137_) );
  DFFPOSX1 DFFPOSX1_1045 ( .CLK(clk_bF_buf53), .D(u2_remHi_138__FF_INPUT), .Q(u2_remHi_138_) );
  DFFPOSX1 DFFPOSX1_1046 ( .CLK(clk_bF_buf52), .D(u2_remHi_139__FF_INPUT), .Q(u2_remHi_139_) );
  DFFPOSX1 DFFPOSX1_1047 ( .CLK(clk_bF_buf51), .D(u2_remHi_140__FF_INPUT), .Q(u2_remHi_140_) );
  DFFPOSX1 DFFPOSX1_1048 ( .CLK(clk_bF_buf50), .D(u2_remHi_141__FF_INPUT), .Q(u2_remHi_141_) );
  DFFPOSX1 DFFPOSX1_1049 ( .CLK(clk_bF_buf49), .D(u2_remHi_142__FF_INPUT), .Q(u2_remHi_142_) );
  DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf17), .D(u2_root_101__FF_INPUT), .Q(sqrto_100_) );
  DFFPOSX1 DFFPOSX1_1050 ( .CLK(clk_bF_buf48), .D(u2_remHi_143__FF_INPUT), .Q(u2_remHi_143_) );
  DFFPOSX1 DFFPOSX1_1051 ( .CLK(clk_bF_buf47), .D(u2_remHi_144__FF_INPUT), .Q(u2_remHi_144_) );
  DFFPOSX1 DFFPOSX1_1052 ( .CLK(clk_bF_buf46), .D(u2_remHi_145__FF_INPUT), .Q(u2_remHi_145_) );
  DFFPOSX1 DFFPOSX1_1053 ( .CLK(clk_bF_buf45), .D(u2_remHi_146__FF_INPUT), .Q(u2_remHi_146_) );
  DFFPOSX1 DFFPOSX1_1054 ( .CLK(clk_bF_buf44), .D(u2_remHi_147__FF_INPUT), .Q(u2_remHi_147_) );
  DFFPOSX1 DFFPOSX1_1055 ( .CLK(clk_bF_buf43), .D(u2_remHi_148__FF_INPUT), .Q(u2_remHi_148_) );
  DFFPOSX1 DFFPOSX1_1056 ( .CLK(clk_bF_buf42), .D(u2_remHi_149__FF_INPUT), .Q(u2_remHi_149_) );
  DFFPOSX1 DFFPOSX1_1057 ( .CLK(clk_bF_buf41), .D(u2_remHi_150__FF_INPUT), .Q(u2_remHi_150_) );
  DFFPOSX1 DFFPOSX1_1058 ( .CLK(clk_bF_buf40), .D(u2_remHi_151__FF_INPUT), .Q(u2_remHi_151_) );
  DFFPOSX1 DFFPOSX1_1059 ( .CLK(clk_bF_buf39), .D(u2_remHi_152__FF_INPUT), .Q(u2_remHi_152_) );
  DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf16), .D(u2_root_102__FF_INPUT), .Q(sqrto_101_) );
  DFFPOSX1 DFFPOSX1_1060 ( .CLK(clk_bF_buf38), .D(u2_remHi_153__FF_INPUT), .Q(u2_remHi_153_) );
  DFFPOSX1 DFFPOSX1_1061 ( .CLK(clk_bF_buf37), .D(u2_remHi_154__FF_INPUT), .Q(u2_remHi_154_) );
  DFFPOSX1 DFFPOSX1_1062 ( .CLK(clk_bF_buf36), .D(u2_remHi_155__FF_INPUT), .Q(u2_remHi_155_) );
  DFFPOSX1 DFFPOSX1_1063 ( .CLK(clk_bF_buf35), .D(u2_remHi_156__FF_INPUT), .Q(u2_remHi_156_) );
  DFFPOSX1 DFFPOSX1_1064 ( .CLK(clk_bF_buf34), .D(u2_remHi_157__FF_INPUT), .Q(u2_remHi_157_) );
  DFFPOSX1 DFFPOSX1_1065 ( .CLK(clk_bF_buf33), .D(u2_remHi_158__FF_INPUT), .Q(u2_remHi_158_) );
  DFFPOSX1 DFFPOSX1_1066 ( .CLK(clk_bF_buf32), .D(u2_remHi_159__FF_INPUT), .Q(u2_remHi_159_) );
  DFFPOSX1 DFFPOSX1_1067 ( .CLK(clk_bF_buf31), .D(u2_remHi_160__FF_INPUT), .Q(u2_remHi_160_) );
  DFFPOSX1 DFFPOSX1_1068 ( .CLK(clk_bF_buf30), .D(u2_remHi_161__FF_INPUT), .Q(u2_remHi_161_) );
  DFFPOSX1 DFFPOSX1_1069 ( .CLK(clk_bF_buf29), .D(u2_remHi_162__FF_INPUT), .Q(u2_remHi_162_) );
  DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf15), .D(u2_root_103__FF_INPUT), .Q(sqrto_102_) );
  DFFPOSX1 DFFPOSX1_1070 ( .CLK(clk_bF_buf28), .D(u2_remHi_163__FF_INPUT), .Q(u2_remHi_163_) );
  DFFPOSX1 DFFPOSX1_1071 ( .CLK(clk_bF_buf27), .D(u2_remHi_164__FF_INPUT), .Q(u2_remHi_164_) );
  DFFPOSX1 DFFPOSX1_1072 ( .CLK(clk_bF_buf26), .D(u2_remHi_165__FF_INPUT), .Q(u2_remHi_165_) );
  DFFPOSX1 DFFPOSX1_1073 ( .CLK(clk_bF_buf25), .D(u2_remHi_166__FF_INPUT), .Q(u2_remHi_166_) );
  DFFPOSX1 DFFPOSX1_1074 ( .CLK(clk_bF_buf24), .D(u2_remHi_167__FF_INPUT), .Q(u2_remHi_167_) );
  DFFPOSX1 DFFPOSX1_1075 ( .CLK(clk_bF_buf23), .D(u2_remHi_168__FF_INPUT), .Q(u2_remHi_168_) );
  DFFPOSX1 DFFPOSX1_1076 ( .CLK(clk_bF_buf22), .D(u2_remHi_169__FF_INPUT), .Q(u2_remHi_169_) );
  DFFPOSX1 DFFPOSX1_1077 ( .CLK(clk_bF_buf21), .D(u2_remHi_170__FF_INPUT), .Q(u2_remHi_170_) );
  DFFPOSX1 DFFPOSX1_1078 ( .CLK(clk_bF_buf20), .D(u2_remHi_171__FF_INPUT), .Q(u2_remHi_171_) );
  DFFPOSX1 DFFPOSX1_1079 ( .CLK(clk_bF_buf19), .D(u2_remHi_172__FF_INPUT), .Q(u2_remHi_172_) );
  DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf14), .D(u2_root_104__FF_INPUT), .Q(sqrto_103_) );
  DFFPOSX1 DFFPOSX1_1080 ( .CLK(clk_bF_buf18), .D(u2_remHi_173__FF_INPUT), .Q(u2_remHi_173_) );
  DFFPOSX1 DFFPOSX1_1081 ( .CLK(clk_bF_buf17), .D(u2_remHi_174__FF_INPUT), .Q(u2_remHi_174_) );
  DFFPOSX1 DFFPOSX1_1082 ( .CLK(clk_bF_buf16), .D(u2_remHi_175__FF_INPUT), .Q(u2_remHi_175_) );
  DFFPOSX1 DFFPOSX1_1083 ( .CLK(clk_bF_buf15), .D(u2_remHi_176__FF_INPUT), .Q(u2_remHi_176_) );
  DFFPOSX1 DFFPOSX1_1084 ( .CLK(clk_bF_buf14), .D(u2_remHi_177__FF_INPUT), .Q(u2_remHi_177_) );
  DFFPOSX1 DFFPOSX1_1085 ( .CLK(clk_bF_buf13), .D(u2_remHi_178__FF_INPUT), .Q(u2_remHi_178_) );
  DFFPOSX1 DFFPOSX1_1086 ( .CLK(clk_bF_buf12), .D(u2_remHi_179__FF_INPUT), .Q(u2_remHi_179_) );
  DFFPOSX1 DFFPOSX1_1087 ( .CLK(clk_bF_buf11), .D(u2_remHi_180__FF_INPUT), .Q(u2_remHi_180_) );
  DFFPOSX1 DFFPOSX1_1088 ( .CLK(clk_bF_buf10), .D(u2_remHi_181__FF_INPUT), .Q(u2_remHi_181_) );
  DFFPOSX1 DFFPOSX1_1089 ( .CLK(clk_bF_buf9), .D(u2_remHi_182__FF_INPUT), .Q(u2_remHi_182_) );
  DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf13), .D(u2_root_105__FF_INPUT), .Q(sqrto_104_) );
  DFFPOSX1 DFFPOSX1_1090 ( .CLK(clk_bF_buf8), .D(u2_remHi_183__FF_INPUT), .Q(u2_remHi_183_) );
  DFFPOSX1 DFFPOSX1_1091 ( .CLK(clk_bF_buf7), .D(u2_remHi_184__FF_INPUT), .Q(u2_remHi_184_) );
  DFFPOSX1 DFFPOSX1_1092 ( .CLK(clk_bF_buf6), .D(u2_remHi_185__FF_INPUT), .Q(u2_remHi_185_) );
  DFFPOSX1 DFFPOSX1_1093 ( .CLK(clk_bF_buf5), .D(u2_remHi_186__FF_INPUT), .Q(u2_remHi_186_) );
  DFFPOSX1 DFFPOSX1_1094 ( .CLK(clk_bF_buf4), .D(u2_remHi_187__FF_INPUT), .Q(u2_remHi_187_) );
  DFFPOSX1 DFFPOSX1_1095 ( .CLK(clk_bF_buf3), .D(u2_remHi_188__FF_INPUT), .Q(u2_remHi_188_) );
  DFFPOSX1 DFFPOSX1_1096 ( .CLK(clk_bF_buf2), .D(u2_remHi_189__FF_INPUT), .Q(u2_remHi_189_) );
  DFFPOSX1 DFFPOSX1_1097 ( .CLK(clk_bF_buf1), .D(u2_remHi_190__FF_INPUT), .Q(u2_remHi_190_) );
  DFFPOSX1 DFFPOSX1_1098 ( .CLK(clk_bF_buf0), .D(u2_remHi_191__FF_INPUT), .Q(u2_remHi_191_) );
  DFFPOSX1 DFFPOSX1_1099 ( .CLK(clk_bF_buf121), .D(u2_remHi_192__FF_INPUT), .Q(u2_remHi_192_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf111), .D(u2_root_7__FF_INPUT), .Q(sqrto_6_) );
  DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf12), .D(u2_root_106__FF_INPUT), .Q(sqrto_105_) );
  DFFPOSX1 DFFPOSX1_1100 ( .CLK(clk_bF_buf120), .D(u2_remHi_193__FF_INPUT), .Q(u2_remHi_193_) );
  DFFPOSX1 DFFPOSX1_1101 ( .CLK(clk_bF_buf119), .D(u2_remHi_194__FF_INPUT), .Q(u2_remHi_194_) );
  DFFPOSX1 DFFPOSX1_1102 ( .CLK(clk_bF_buf118), .D(u2_remHi_195__FF_INPUT), .Q(u2_remHi_195_) );
  DFFPOSX1 DFFPOSX1_1103 ( .CLK(clk_bF_buf117), .D(u2_remHi_196__FF_INPUT), .Q(u2_remHi_196_) );
  DFFPOSX1 DFFPOSX1_1104 ( .CLK(clk_bF_buf116), .D(u2_remHi_197__FF_INPUT), .Q(u2_remHi_197_) );
  DFFPOSX1 DFFPOSX1_1105 ( .CLK(clk_bF_buf115), .D(u2_remHi_198__FF_INPUT), .Q(u2_remHi_198_) );
  DFFPOSX1 DFFPOSX1_1106 ( .CLK(clk_bF_buf114), .D(u2_remHi_199__FF_INPUT), .Q(u2_remHi_199_) );
  DFFPOSX1 DFFPOSX1_1107 ( .CLK(clk_bF_buf113), .D(u2_remHi_200__FF_INPUT), .Q(u2_remHi_200_) );
  DFFPOSX1 DFFPOSX1_1108 ( .CLK(clk_bF_buf112), .D(u2_remHi_201__FF_INPUT), .Q(u2_remHi_201_) );
  DFFPOSX1 DFFPOSX1_1109 ( .CLK(clk_bF_buf111), .D(u2_remHi_202__FF_INPUT), .Q(u2_remHi_202_) );
  DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf11), .D(u2_root_107__FF_INPUT), .Q(sqrto_106_) );
  DFFPOSX1 DFFPOSX1_1110 ( .CLK(clk_bF_buf110), .D(u2_remHi_203__FF_INPUT), .Q(u2_remHi_203_) );
  DFFPOSX1 DFFPOSX1_1111 ( .CLK(clk_bF_buf109), .D(u2_remHi_204__FF_INPUT), .Q(u2_remHi_204_) );
  DFFPOSX1 DFFPOSX1_1112 ( .CLK(clk_bF_buf108), .D(u2_remHi_205__FF_INPUT), .Q(u2_remHi_205_) );
  DFFPOSX1 DFFPOSX1_1113 ( .CLK(clk_bF_buf107), .D(u2_remHi_206__FF_INPUT), .Q(u2_remHi_206_) );
  DFFPOSX1 DFFPOSX1_1114 ( .CLK(clk_bF_buf106), .D(u2_remHi_207__FF_INPUT), .Q(u2_remHi_207_) );
  DFFPOSX1 DFFPOSX1_1115 ( .CLK(clk_bF_buf105), .D(u2_remHi_208__FF_INPUT), .Q(u2_remHi_208_) );
  DFFPOSX1 DFFPOSX1_1116 ( .CLK(clk_bF_buf104), .D(u2_remHi_209__FF_INPUT), .Q(u2_remHi_209_) );
  DFFPOSX1 DFFPOSX1_1117 ( .CLK(clk_bF_buf103), .D(u2_remHi_210__FF_INPUT), .Q(u2_remHi_210_) );
  DFFPOSX1 DFFPOSX1_1118 ( .CLK(clk_bF_buf102), .D(u2_remHi_211__FF_INPUT), .Q(u2_remHi_211_) );
  DFFPOSX1 DFFPOSX1_1119 ( .CLK(clk_bF_buf101), .D(u2_remHi_212__FF_INPUT), .Q(u2_remHi_212_) );
  DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf10), .D(u2_root_108__FF_INPUT), .Q(sqrto_107_) );
  DFFPOSX1 DFFPOSX1_1120 ( .CLK(clk_bF_buf100), .D(u2_remHi_213__FF_INPUT), .Q(u2_remHi_213_) );
  DFFPOSX1 DFFPOSX1_1121 ( .CLK(clk_bF_buf99), .D(u2_remHi_214__FF_INPUT), .Q(u2_remHi_214_) );
  DFFPOSX1 DFFPOSX1_1122 ( .CLK(clk_bF_buf98), .D(u2_remHi_215__FF_INPUT), .Q(u2_remHi_215_) );
  DFFPOSX1 DFFPOSX1_1123 ( .CLK(clk_bF_buf97), .D(u2_remHi_216__FF_INPUT), .Q(u2_remHi_216_) );
  DFFPOSX1 DFFPOSX1_1124 ( .CLK(clk_bF_buf96), .D(u2_remHi_217__FF_INPUT), .Q(u2_remHi_217_) );
  DFFPOSX1 DFFPOSX1_1125 ( .CLK(clk_bF_buf95), .D(u2_remHi_218__FF_INPUT), .Q(u2_remHi_218_) );
  DFFPOSX1 DFFPOSX1_1126 ( .CLK(clk_bF_buf94), .D(u2_remHi_219__FF_INPUT), .Q(u2_remHi_219_) );
  DFFPOSX1 DFFPOSX1_1127 ( .CLK(clk_bF_buf93), .D(u2_remHi_220__FF_INPUT), .Q(u2_remHi_220_) );
  DFFPOSX1 DFFPOSX1_1128 ( .CLK(clk_bF_buf92), .D(u2_remHi_221__FF_INPUT), .Q(u2_remHi_221_) );
  DFFPOSX1 DFFPOSX1_1129 ( .CLK(clk_bF_buf91), .D(u2_remHi_222__FF_INPUT), .Q(u2_remHi_222_) );
  DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf9), .D(u2_root_109__FF_INPUT), .Q(sqrto_108_) );
  DFFPOSX1 DFFPOSX1_1130 ( .CLK(clk_bF_buf90), .D(u2_remHi_223__FF_INPUT), .Q(u2_remHi_223_) );
  DFFPOSX1 DFFPOSX1_1131 ( .CLK(clk_bF_buf89), .D(u2_remHi_224__FF_INPUT), .Q(u2_remHi_224_) );
  DFFPOSX1 DFFPOSX1_1132 ( .CLK(clk_bF_buf88), .D(u2_remHi_225__FF_INPUT), .Q(u2_remHi_225_) );
  DFFPOSX1 DFFPOSX1_1133 ( .CLK(clk_bF_buf87), .D(u2_remHi_226__FF_INPUT), .Q(u2_remHi_226_) );
  DFFPOSX1 DFFPOSX1_1134 ( .CLK(clk_bF_buf86), .D(u2_remHi_227__FF_INPUT), .Q(u2_remHi_227_) );
  DFFPOSX1 DFFPOSX1_1135 ( .CLK(clk_bF_buf85), .D(u2_remHi_228__FF_INPUT), .Q(u2_remHi_228_) );
  DFFPOSX1 DFFPOSX1_1136 ( .CLK(clk_bF_buf84), .D(u2_remHi_229__FF_INPUT), .Q(u2_remHi_229_) );
  DFFPOSX1 DFFPOSX1_1137 ( .CLK(clk_bF_buf83), .D(u2_remHi_230__FF_INPUT), .Q(u2_remHi_230_) );
  DFFPOSX1 DFFPOSX1_1138 ( .CLK(clk_bF_buf82), .D(u2_remHi_231__FF_INPUT), .Q(u2_remHi_231_) );
  DFFPOSX1 DFFPOSX1_1139 ( .CLK(clk_bF_buf81), .D(u2_remHi_232__FF_INPUT), .Q(u2_remHi_232_) );
  DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf8), .D(u2_root_110__FF_INPUT), .Q(sqrto_109_) );
  DFFPOSX1 DFFPOSX1_1140 ( .CLK(clk_bF_buf80), .D(u2_remHi_233__FF_INPUT), .Q(u2_remHi_233_) );
  DFFPOSX1 DFFPOSX1_1141 ( .CLK(clk_bF_buf79), .D(u2_remHi_234__FF_INPUT), .Q(u2_remHi_234_) );
  DFFPOSX1 DFFPOSX1_1142 ( .CLK(clk_bF_buf78), .D(u2_remHi_235__FF_INPUT), .Q(u2_remHi_235_) );
  DFFPOSX1 DFFPOSX1_1143 ( .CLK(clk_bF_buf77), .D(u2_remHi_236__FF_INPUT), .Q(u2_remHi_236_) );
  DFFPOSX1 DFFPOSX1_1144 ( .CLK(clk_bF_buf76), .D(u2_remHi_237__FF_INPUT), .Q(u2_remHi_237_) );
  DFFPOSX1 DFFPOSX1_1145 ( .CLK(clk_bF_buf75), .D(u2_remHi_238__FF_INPUT), .Q(u2_remHi_238_) );
  DFFPOSX1 DFFPOSX1_1146 ( .CLK(clk_bF_buf74), .D(u2_remHi_239__FF_INPUT), .Q(u2_remHi_239_) );
  DFFPOSX1 DFFPOSX1_1147 ( .CLK(clk_bF_buf73), .D(u2_remHi_240__FF_INPUT), .Q(u2_remHi_240_) );
  DFFPOSX1 DFFPOSX1_1148 ( .CLK(clk_bF_buf72), .D(u2_remHi_241__FF_INPUT), .Q(u2_remHi_241_) );
  DFFPOSX1 DFFPOSX1_1149 ( .CLK(clk_bF_buf71), .D(u2_remHi_242__FF_INPUT), .Q(u2_remHi_242_) );
  DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf7), .D(u2_root_111__FF_INPUT), .Q(sqrto_110_) );
  DFFPOSX1 DFFPOSX1_1150 ( .CLK(clk_bF_buf70), .D(u2_remHi_243__FF_INPUT), .Q(u2_remHi_243_) );
  DFFPOSX1 DFFPOSX1_1151 ( .CLK(clk_bF_buf69), .D(u2_remHi_244__FF_INPUT), .Q(u2_remHi_244_) );
  DFFPOSX1 DFFPOSX1_1152 ( .CLK(clk_bF_buf68), .D(u2_remHi_245__FF_INPUT), .Q(u2_remHi_245_) );
  DFFPOSX1 DFFPOSX1_1153 ( .CLK(clk_bF_buf67), .D(u2_remHi_246__FF_INPUT), .Q(u2_remHi_246_) );
  DFFPOSX1 DFFPOSX1_1154 ( .CLK(clk_bF_buf66), .D(u2_remHi_247__FF_INPUT), .Q(u2_remHi_247_) );
  DFFPOSX1 DFFPOSX1_1155 ( .CLK(clk_bF_buf65), .D(u2_remHi_248__FF_INPUT), .Q(u2_remHi_248_) );
  DFFPOSX1 DFFPOSX1_1156 ( .CLK(clk_bF_buf64), .D(u2_remHi_249__FF_INPUT), .Q(u2_remHi_249_) );
  DFFPOSX1 DFFPOSX1_1157 ( .CLK(clk_bF_buf63), .D(u2_remHi_250__FF_INPUT), .Q(u2_remHi_250_) );
  DFFPOSX1 DFFPOSX1_1158 ( .CLK(clk_bF_buf62), .D(u2_remHi_251__FF_INPUT), .Q(u2_remHi_251_) );
  DFFPOSX1 DFFPOSX1_1159 ( .CLK(clk_bF_buf61), .D(u2_remHi_252__FF_INPUT), .Q(u2_remHi_252_) );
  DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf6), .D(u2_root_112__FF_INPUT), .Q(sqrto_111_) );
  DFFPOSX1 DFFPOSX1_1160 ( .CLK(clk_bF_buf60), .D(u2_remHi_253__FF_INPUT), .Q(u2_remHi_253_) );
  DFFPOSX1 DFFPOSX1_1161 ( .CLK(clk_bF_buf59), .D(u2_remHi_254__FF_INPUT), .Q(u2_remHi_254_) );
  DFFPOSX1 DFFPOSX1_1162 ( .CLK(clk_bF_buf58), .D(u2_remHi_255__FF_INPUT), .Q(u2_remHi_255_) );
  DFFPOSX1 DFFPOSX1_1163 ( .CLK(clk_bF_buf57), .D(u2_remHi_256__FF_INPUT), .Q(u2_remHi_256_) );
  DFFPOSX1 DFFPOSX1_1164 ( .CLK(clk_bF_buf56), .D(u2_remHi_257__FF_INPUT), .Q(u2_remHi_257_) );
  DFFPOSX1 DFFPOSX1_1165 ( .CLK(clk_bF_buf55), .D(u2_remHi_258__FF_INPUT), .Q(u2_remHi_258_) );
  DFFPOSX1 DFFPOSX1_1166 ( .CLK(clk_bF_buf54), .D(u2_remHi_259__FF_INPUT), .Q(u2_remHi_259_) );
  DFFPOSX1 DFFPOSX1_1167 ( .CLK(clk_bF_buf53), .D(u2_remHi_260__FF_INPUT), .Q(u2_remHi_260_) );
  DFFPOSX1 DFFPOSX1_1168 ( .CLK(clk_bF_buf52), .D(u2_remHi_261__FF_INPUT), .Q(u2_remHi_261_) );
  DFFPOSX1 DFFPOSX1_1169 ( .CLK(clk_bF_buf51), .D(u2_remHi_262__FF_INPUT), .Q(u2_remHi_262_) );
  DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf5), .D(u2_root_113__FF_INPUT), .Q(sqrto_112_) );
  DFFPOSX1 DFFPOSX1_1170 ( .CLK(clk_bF_buf50), .D(u2_remHi_263__FF_INPUT), .Q(u2_remHi_263_) );
  DFFPOSX1 DFFPOSX1_1171 ( .CLK(clk_bF_buf49), .D(u2_remHi_264__FF_INPUT), .Q(u2_remHi_264_) );
  DFFPOSX1 DFFPOSX1_1172 ( .CLK(clk_bF_buf48), .D(u2_remHi_265__FF_INPUT), .Q(u2_remHi_265_) );
  DFFPOSX1 DFFPOSX1_1173 ( .CLK(clk_bF_buf47), .D(u2_remHi_266__FF_INPUT), .Q(u2_remHi_266_) );
  DFFPOSX1 DFFPOSX1_1174 ( .CLK(clk_bF_buf46), .D(u2_remHi_267__FF_INPUT), .Q(u2_remHi_267_) );
  DFFPOSX1 DFFPOSX1_1175 ( .CLK(clk_bF_buf45), .D(u2_remHi_268__FF_INPUT), .Q(u2_remHi_268_) );
  DFFPOSX1 DFFPOSX1_1176 ( .CLK(clk_bF_buf44), .D(u2_remHi_269__FF_INPUT), .Q(u2_remHi_269_) );
  DFFPOSX1 DFFPOSX1_1177 ( .CLK(clk_bF_buf43), .D(u2_remHi_270__FF_INPUT), .Q(u2_remHi_270_) );
  DFFPOSX1 DFFPOSX1_1178 ( .CLK(clk_bF_buf42), .D(u2_remHi_271__FF_INPUT), .Q(u2_remHi_271_) );
  DFFPOSX1 DFFPOSX1_1179 ( .CLK(clk_bF_buf41), .D(u2_remHi_272__FF_INPUT), .Q(u2_remHi_272_) );
  DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf4), .D(u2_root_114__FF_INPUT), .Q(sqrto_113_) );
  DFFPOSX1 DFFPOSX1_1180 ( .CLK(clk_bF_buf40), .D(u2_remHi_273__FF_INPUT), .Q(u2_remHi_273_) );
  DFFPOSX1 DFFPOSX1_1181 ( .CLK(clk_bF_buf39), .D(u2_remHi_274__FF_INPUT), .Q(u2_remHi_274_) );
  DFFPOSX1 DFFPOSX1_1182 ( .CLK(clk_bF_buf38), .D(u2_remHi_275__FF_INPUT), .Q(u2_remHi_275_) );
  DFFPOSX1 DFFPOSX1_1183 ( .CLK(clk_bF_buf37), .D(u2_remHi_276__FF_INPUT), .Q(u2_remHi_276_) );
  DFFPOSX1 DFFPOSX1_1184 ( .CLK(clk_bF_buf36), .D(u2_remHi_277__FF_INPUT), .Q(u2_remHi_277_) );
  DFFPOSX1 DFFPOSX1_1185 ( .CLK(clk_bF_buf35), .D(u2_remHi_278__FF_INPUT), .Q(u2_remHi_278_) );
  DFFPOSX1 DFFPOSX1_1186 ( .CLK(clk_bF_buf34), .D(u2_remHi_279__FF_INPUT), .Q(u2_remHi_279_) );
  DFFPOSX1 DFFPOSX1_1187 ( .CLK(clk_bF_buf33), .D(u2_remHi_280__FF_INPUT), .Q(u2_remHi_280_) );
  DFFPOSX1 DFFPOSX1_1188 ( .CLK(clk_bF_buf32), .D(u2_remHi_281__FF_INPUT), .Q(u2_remHi_281_) );
  DFFPOSX1 DFFPOSX1_1189 ( .CLK(clk_bF_buf31), .D(u2_remHi_282__FF_INPUT), .Q(u2_remHi_282_) );
  DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf3), .D(u2_root_115__FF_INPUT), .Q(sqrto_114_) );
  DFFPOSX1 DFFPOSX1_1190 ( .CLK(clk_bF_buf30), .D(u2_remHi_283__FF_INPUT), .Q(u2_remHi_283_) );
  DFFPOSX1 DFFPOSX1_1191 ( .CLK(clk_bF_buf29), .D(u2_remHi_284__FF_INPUT), .Q(u2_remHi_284_) );
  DFFPOSX1 DFFPOSX1_1192 ( .CLK(clk_bF_buf28), .D(u2_remHi_285__FF_INPUT), .Q(u2_remHi_285_) );
  DFFPOSX1 DFFPOSX1_1193 ( .CLK(clk_bF_buf27), .D(u2_remHi_286__FF_INPUT), .Q(u2_remHi_286_) );
  DFFPOSX1 DFFPOSX1_1194 ( .CLK(clk_bF_buf26), .D(u2_remHi_287__FF_INPUT), .Q(u2_remHi_287_) );
  DFFPOSX1 DFFPOSX1_1195 ( .CLK(clk_bF_buf25), .D(u2_remHi_288__FF_INPUT), .Q(u2_remHi_288_) );
  DFFPOSX1 DFFPOSX1_1196 ( .CLK(clk_bF_buf24), .D(u2_remHi_289__FF_INPUT), .Q(u2_remHi_289_) );
  DFFPOSX1 DFFPOSX1_1197 ( .CLK(clk_bF_buf23), .D(u2_remHi_290__FF_INPUT), .Q(u2_remHi_290_) );
  DFFPOSX1 DFFPOSX1_1198 ( .CLK(clk_bF_buf22), .D(u2_remHi_291__FF_INPUT), .Q(u2_remHi_291_) );
  DFFPOSX1 DFFPOSX1_1199 ( .CLK(clk_bF_buf21), .D(u2_remHi_292__FF_INPUT), .Q(u2_remHi_292_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf110), .D(u2_root_8__FF_INPUT), .Q(sqrto_7_) );
  DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf2), .D(u2_root_116__FF_INPUT), .Q(sqrto_115_) );
  DFFPOSX1 DFFPOSX1_1200 ( .CLK(clk_bF_buf20), .D(u2_remHi_293__FF_INPUT), .Q(u2_remHi_293_) );
  DFFPOSX1 DFFPOSX1_1201 ( .CLK(clk_bF_buf19), .D(u2_remHi_294__FF_INPUT), .Q(u2_remHi_294_) );
  DFFPOSX1 DFFPOSX1_1202 ( .CLK(clk_bF_buf18), .D(u2_remHi_295__FF_INPUT), .Q(u2_remHi_295_) );
  DFFPOSX1 DFFPOSX1_1203 ( .CLK(clk_bF_buf17), .D(u2_remHi_296__FF_INPUT), .Q(u2_remHi_296_) );
  DFFPOSX1 DFFPOSX1_1204 ( .CLK(clk_bF_buf16), .D(u2_remHi_297__FF_INPUT), .Q(u2_remHi_297_) );
  DFFPOSX1 DFFPOSX1_1205 ( .CLK(clk_bF_buf15), .D(u2_remHi_298__FF_INPUT), .Q(u2_remHi_298_) );
  DFFPOSX1 DFFPOSX1_1206 ( .CLK(clk_bF_buf14), .D(u2_remHi_299__FF_INPUT), .Q(u2_remHi_299_) );
  DFFPOSX1 DFFPOSX1_1207 ( .CLK(clk_bF_buf13), .D(u2_remHi_300__FF_INPUT), .Q(u2_remHi_300_) );
  DFFPOSX1 DFFPOSX1_1208 ( .CLK(clk_bF_buf12), .D(u2_remHi_301__FF_INPUT), .Q(u2_remHi_301_) );
  DFFPOSX1 DFFPOSX1_1209 ( .CLK(clk_bF_buf11), .D(u2_remHi_302__FF_INPUT), .Q(u2_remHi_302_) );
  DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf1), .D(u2_root_117__FF_INPUT), .Q(sqrto_116_) );
  DFFPOSX1 DFFPOSX1_1210 ( .CLK(clk_bF_buf10), .D(u2_remHi_303__FF_INPUT), .Q(u2_remHi_303_) );
  DFFPOSX1 DFFPOSX1_1211 ( .CLK(clk_bF_buf9), .D(u2_remHi_304__FF_INPUT), .Q(u2_remHi_304_) );
  DFFPOSX1 DFFPOSX1_1212 ( .CLK(clk_bF_buf8), .D(u2_remHi_305__FF_INPUT), .Q(u2_remHi_305_) );
  DFFPOSX1 DFFPOSX1_1213 ( .CLK(clk_bF_buf7), .D(u2_remHi_306__FF_INPUT), .Q(u2_remHi_306_) );
  DFFPOSX1 DFFPOSX1_1214 ( .CLK(clk_bF_buf6), .D(u2_remHi_307__FF_INPUT), .Q(u2_remHi_307_) );
  DFFPOSX1 DFFPOSX1_1215 ( .CLK(clk_bF_buf5), .D(u2_remHi_308__FF_INPUT), .Q(u2_remHi_308_) );
  DFFPOSX1 DFFPOSX1_1216 ( .CLK(clk_bF_buf4), .D(u2_remHi_309__FF_INPUT), .Q(u2_remHi_309_) );
  DFFPOSX1 DFFPOSX1_1217 ( .CLK(clk_bF_buf3), .D(u2_remHi_310__FF_INPUT), .Q(u2_remHi_310_) );
  DFFPOSX1 DFFPOSX1_1218 ( .CLK(clk_bF_buf2), .D(u2_remHi_311__FF_INPUT), .Q(u2_remHi_311_) );
  DFFPOSX1 DFFPOSX1_1219 ( .CLK(clk_bF_buf1), .D(u2_remHi_312__FF_INPUT), .Q(u2_remHi_312_) );
  DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf0), .D(u2_root_118__FF_INPUT), .Q(sqrto_117_) );
  DFFPOSX1 DFFPOSX1_1220 ( .CLK(clk_bF_buf0), .D(u2_remHi_313__FF_INPUT), .Q(u2_remHi_313_) );
  DFFPOSX1 DFFPOSX1_1221 ( .CLK(clk_bF_buf121), .D(u2_remHi_314__FF_INPUT), .Q(u2_remHi_314_) );
  DFFPOSX1 DFFPOSX1_1222 ( .CLK(clk_bF_buf120), .D(u2_remHi_315__FF_INPUT), .Q(u2_remHi_315_) );
  DFFPOSX1 DFFPOSX1_1223 ( .CLK(clk_bF_buf119), .D(u2_remHi_316__FF_INPUT), .Q(u2_remHi_316_) );
  DFFPOSX1 DFFPOSX1_1224 ( .CLK(clk_bF_buf118), .D(u2_remHi_317__FF_INPUT), .Q(u2_remHi_317_) );
  DFFPOSX1 DFFPOSX1_1225 ( .CLK(clk_bF_buf117), .D(u2_remHi_318__FF_INPUT), .Q(u2_remHi_318_) );
  DFFPOSX1 DFFPOSX1_1226 ( .CLK(clk_bF_buf116), .D(u2_remHi_319__FF_INPUT), .Q(u2_remHi_319_) );
  DFFPOSX1 DFFPOSX1_1227 ( .CLK(clk_bF_buf115), .D(u2_remHi_320__FF_INPUT), .Q(u2_remHi_320_) );
  DFFPOSX1 DFFPOSX1_1228 ( .CLK(clk_bF_buf114), .D(u2_remHi_321__FF_INPUT), .Q(u2_remHi_321_) );
  DFFPOSX1 DFFPOSX1_1229 ( .CLK(clk_bF_buf113), .D(u2_remHi_322__FF_INPUT), .Q(u2_remHi_322_) );
  DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf121), .D(u2_root_119__FF_INPUT), .Q(sqrto_118_) );
  DFFPOSX1 DFFPOSX1_1230 ( .CLK(clk_bF_buf112), .D(u2_remHi_323__FF_INPUT), .Q(u2_remHi_323_) );
  DFFPOSX1 DFFPOSX1_1231 ( .CLK(clk_bF_buf111), .D(u2_remHi_324__FF_INPUT), .Q(u2_remHi_324_) );
  DFFPOSX1 DFFPOSX1_1232 ( .CLK(clk_bF_buf110), .D(u2_remHi_325__FF_INPUT), .Q(u2_remHi_325_) );
  DFFPOSX1 DFFPOSX1_1233 ( .CLK(clk_bF_buf109), .D(u2_remHi_326__FF_INPUT), .Q(u2_remHi_326_) );
  DFFPOSX1 DFFPOSX1_1234 ( .CLK(clk_bF_buf108), .D(u2_remHi_327__FF_INPUT), .Q(u2_remHi_327_) );
  DFFPOSX1 DFFPOSX1_1235 ( .CLK(clk_bF_buf107), .D(u2_remHi_328__FF_INPUT), .Q(u2_remHi_328_) );
  DFFPOSX1 DFFPOSX1_1236 ( .CLK(clk_bF_buf106), .D(u2_remHi_329__FF_INPUT), .Q(u2_remHi_329_) );
  DFFPOSX1 DFFPOSX1_1237 ( .CLK(clk_bF_buf105), .D(u2_remHi_330__FF_INPUT), .Q(u2_remHi_330_) );
  DFFPOSX1 DFFPOSX1_1238 ( .CLK(clk_bF_buf104), .D(u2_remHi_331__FF_INPUT), .Q(u2_remHi_331_) );
  DFFPOSX1 DFFPOSX1_1239 ( .CLK(clk_bF_buf103), .D(u2_remHi_332__FF_INPUT), .Q(u2_remHi_332_) );
  DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf120), .D(u2_root_120__FF_INPUT), .Q(sqrto_119_) );
  DFFPOSX1 DFFPOSX1_1240 ( .CLK(clk_bF_buf102), .D(u2_remHi_333__FF_INPUT), .Q(u2_remHi_333_) );
  DFFPOSX1 DFFPOSX1_1241 ( .CLK(clk_bF_buf101), .D(u2_remHi_334__FF_INPUT), .Q(u2_remHi_334_) );
  DFFPOSX1 DFFPOSX1_1242 ( .CLK(clk_bF_buf100), .D(u2_remHi_335__FF_INPUT), .Q(u2_remHi_335_) );
  DFFPOSX1 DFFPOSX1_1243 ( .CLK(clk_bF_buf99), .D(u2_remHi_336__FF_INPUT), .Q(u2_remHi_336_) );
  DFFPOSX1 DFFPOSX1_1244 ( .CLK(clk_bF_buf98), .D(u2_remHi_337__FF_INPUT), .Q(u2_remHi_337_) );
  DFFPOSX1 DFFPOSX1_1245 ( .CLK(clk_bF_buf97), .D(u2_remHi_338__FF_INPUT), .Q(u2_remHi_338_) );
  DFFPOSX1 DFFPOSX1_1246 ( .CLK(clk_bF_buf96), .D(u2_remHi_339__FF_INPUT), .Q(u2_remHi_339_) );
  DFFPOSX1 DFFPOSX1_1247 ( .CLK(clk_bF_buf95), .D(u2_remHi_340__FF_INPUT), .Q(u2_remHi_340_) );
  DFFPOSX1 DFFPOSX1_1248 ( .CLK(clk_bF_buf94), .D(u2_remHi_341__FF_INPUT), .Q(u2_remHi_341_) );
  DFFPOSX1 DFFPOSX1_1249 ( .CLK(clk_bF_buf93), .D(u2_remHi_342__FF_INPUT), .Q(u2_remHi_342_) );
  DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf119), .D(u2_root_121__FF_INPUT), .Q(sqrto_120_) );
  DFFPOSX1 DFFPOSX1_1250 ( .CLK(clk_bF_buf92), .D(u2_remHi_343__FF_INPUT), .Q(u2_remHi_343_) );
  DFFPOSX1 DFFPOSX1_1251 ( .CLK(clk_bF_buf91), .D(u2_remHi_344__FF_INPUT), .Q(u2_remHi_344_) );
  DFFPOSX1 DFFPOSX1_1252 ( .CLK(clk_bF_buf90), .D(u2_remHi_345__FF_INPUT), .Q(u2_remHi_345_) );
  DFFPOSX1 DFFPOSX1_1253 ( .CLK(clk_bF_buf89), .D(u2_remHi_346__FF_INPUT), .Q(u2_remHi_346_) );
  DFFPOSX1 DFFPOSX1_1254 ( .CLK(clk_bF_buf88), .D(u2_remHi_347__FF_INPUT), .Q(u2_remHi_347_) );
  DFFPOSX1 DFFPOSX1_1255 ( .CLK(clk_bF_buf87), .D(u2_remHi_348__FF_INPUT), .Q(u2_remHi_348_) );
  DFFPOSX1 DFFPOSX1_1256 ( .CLK(clk_bF_buf86), .D(u2_remHi_349__FF_INPUT), .Q(u2_remHi_349_) );
  DFFPOSX1 DFFPOSX1_1257 ( .CLK(clk_bF_buf85), .D(u2_remHi_350__FF_INPUT), .Q(u2_remHi_350_) );
  DFFPOSX1 DFFPOSX1_1258 ( .CLK(clk_bF_buf84), .D(u2_remHi_351__FF_INPUT), .Q(u2_remHi_351_) );
  DFFPOSX1 DFFPOSX1_1259 ( .CLK(clk_bF_buf83), .D(u2_remHi_352__FF_INPUT), .Q(u2_remHi_352_) );
  DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf118), .D(u2_root_122__FF_INPUT), .Q(sqrto_121_) );
  DFFPOSX1 DFFPOSX1_1260 ( .CLK(clk_bF_buf82), .D(u2_remHi_353__FF_INPUT), .Q(u2_remHi_353_) );
  DFFPOSX1 DFFPOSX1_1261 ( .CLK(clk_bF_buf81), .D(u2_remHi_354__FF_INPUT), .Q(u2_remHi_354_) );
  DFFPOSX1 DFFPOSX1_1262 ( .CLK(clk_bF_buf80), .D(u2_remHi_355__FF_INPUT), .Q(u2_remHi_355_) );
  DFFPOSX1 DFFPOSX1_1263 ( .CLK(clk_bF_buf79), .D(u2_remHi_356__FF_INPUT), .Q(u2_remHi_356_) );
  DFFPOSX1 DFFPOSX1_1264 ( .CLK(clk_bF_buf78), .D(u2_remHi_357__FF_INPUT), .Q(u2_remHi_357_) );
  DFFPOSX1 DFFPOSX1_1265 ( .CLK(clk_bF_buf77), .D(u2_remHi_358__FF_INPUT), .Q(u2_remHi_358_) );
  DFFPOSX1 DFFPOSX1_1266 ( .CLK(clk_bF_buf76), .D(u2_remHi_359__FF_INPUT), .Q(u2_remHi_359_) );
  DFFPOSX1 DFFPOSX1_1267 ( .CLK(clk_bF_buf75), .D(u2_remHi_360__FF_INPUT), .Q(u2_remHi_360_) );
  DFFPOSX1 DFFPOSX1_1268 ( .CLK(clk_bF_buf74), .D(u2_remHi_361__FF_INPUT), .Q(u2_remHi_361_) );
  DFFPOSX1 DFFPOSX1_1269 ( .CLK(clk_bF_buf73), .D(u2_remHi_362__FF_INPUT), .Q(u2_remHi_362_) );
  DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf117), .D(u2_root_123__FF_INPUT), .Q(sqrto_122_) );
  DFFPOSX1 DFFPOSX1_1270 ( .CLK(clk_bF_buf72), .D(u2_remHi_363__FF_INPUT), .Q(u2_remHi_363_) );
  DFFPOSX1 DFFPOSX1_1271 ( .CLK(clk_bF_buf71), .D(u2_remHi_364__FF_INPUT), .Q(u2_remHi_364_) );
  DFFPOSX1 DFFPOSX1_1272 ( .CLK(clk_bF_buf70), .D(u2_remHi_365__FF_INPUT), .Q(u2_remHi_365_) );
  DFFPOSX1 DFFPOSX1_1273 ( .CLK(clk_bF_buf69), .D(u2_remHi_366__FF_INPUT), .Q(u2_remHi_366_) );
  DFFPOSX1 DFFPOSX1_1274 ( .CLK(clk_bF_buf68), .D(u2_remHi_367__FF_INPUT), .Q(u2_remHi_367_) );
  DFFPOSX1 DFFPOSX1_1275 ( .CLK(clk_bF_buf67), .D(u2_remHi_368__FF_INPUT), .Q(u2_remHi_368_) );
  DFFPOSX1 DFFPOSX1_1276 ( .CLK(clk_bF_buf66), .D(u2_remHi_369__FF_INPUT), .Q(u2_remHi_369_) );
  DFFPOSX1 DFFPOSX1_1277 ( .CLK(clk_bF_buf65), .D(u2_remHi_370__FF_INPUT), .Q(u2_remHi_370_) );
  DFFPOSX1 DFFPOSX1_1278 ( .CLK(clk_bF_buf64), .D(u2_remHi_371__FF_INPUT), .Q(u2_remHi_371_) );
  DFFPOSX1 DFFPOSX1_1279 ( .CLK(clk_bF_buf63), .D(u2_remHi_372__FF_INPUT), .Q(u2_remHi_372_) );
  DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf116), .D(u2_root_124__FF_INPUT), .Q(sqrto_123_) );
  DFFPOSX1 DFFPOSX1_1280 ( .CLK(clk_bF_buf62), .D(u2_remHi_373__FF_INPUT), .Q(u2_remHi_373_) );
  DFFPOSX1 DFFPOSX1_1281 ( .CLK(clk_bF_buf61), .D(u2_remHi_374__FF_INPUT), .Q(u2_remHi_374_) );
  DFFPOSX1 DFFPOSX1_1282 ( .CLK(clk_bF_buf60), .D(u2_remHi_375__FF_INPUT), .Q(u2_remHi_375_) );
  DFFPOSX1 DFFPOSX1_1283 ( .CLK(clk_bF_buf59), .D(u2_remHi_376__FF_INPUT), .Q(u2_remHi_376_) );
  DFFPOSX1 DFFPOSX1_1284 ( .CLK(clk_bF_buf58), .D(u2_remHi_377__FF_INPUT), .Q(u2_remHi_377_) );
  DFFPOSX1 DFFPOSX1_1285 ( .CLK(clk_bF_buf57), .D(u2_remHi_378__FF_INPUT), .Q(u2_remHi_378_) );
  DFFPOSX1 DFFPOSX1_1286 ( .CLK(clk_bF_buf56), .D(u2_remHi_379__FF_INPUT), .Q(u2_remHi_379_) );
  DFFPOSX1 DFFPOSX1_1287 ( .CLK(clk_bF_buf55), .D(u2_remHi_380__FF_INPUT), .Q(u2_remHi_380_) );
  DFFPOSX1 DFFPOSX1_1288 ( .CLK(clk_bF_buf54), .D(u2_remHi_381__FF_INPUT), .Q(u2_remHi_381_) );
  DFFPOSX1 DFFPOSX1_1289 ( .CLK(clk_bF_buf53), .D(u2_remHi_382__FF_INPUT), .Q(u2_remHi_382_) );
  DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf115), .D(u2_root_125__FF_INPUT), .Q(sqrto_124_) );
  DFFPOSX1 DFFPOSX1_1290 ( .CLK(clk_bF_buf52), .D(u2_remHi_383__FF_INPUT), .Q(u2_remHi_383_) );
  DFFPOSX1 DFFPOSX1_1291 ( .CLK(clk_bF_buf51), .D(u2_remHi_384__FF_INPUT), .Q(u2_remHi_384_) );
  DFFPOSX1 DFFPOSX1_1292 ( .CLK(clk_bF_buf50), .D(u2_remHi_385__FF_INPUT), .Q(u2_remHi_385_) );
  DFFPOSX1 DFFPOSX1_1293 ( .CLK(clk_bF_buf49), .D(u2_remHi_386__FF_INPUT), .Q(u2_remHi_386_) );
  DFFPOSX1 DFFPOSX1_1294 ( .CLK(clk_bF_buf48), .D(u2_remHi_387__FF_INPUT), .Q(u2_remHi_387_) );
  DFFPOSX1 DFFPOSX1_1295 ( .CLK(clk_bF_buf47), .D(u2_remHi_388__FF_INPUT), .Q(u2_remHi_388_) );
  DFFPOSX1 DFFPOSX1_1296 ( .CLK(clk_bF_buf46), .D(u2_remHi_389__FF_INPUT), .Q(u2_remHi_389_) );
  DFFPOSX1 DFFPOSX1_1297 ( .CLK(clk_bF_buf45), .D(u2_remHi_390__FF_INPUT), .Q(u2_remHi_390_) );
  DFFPOSX1 DFFPOSX1_1298 ( .CLK(clk_bF_buf44), .D(u2_remHi_391__FF_INPUT), .Q(u2_remHi_391_) );
  DFFPOSX1 DFFPOSX1_1299 ( .CLK(clk_bF_buf43), .D(u2_remHi_392__FF_INPUT), .Q(u2_remHi_392_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf109), .D(u2_root_9__FF_INPUT), .Q(sqrto_8_) );
  DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf114), .D(u2_root_126__FF_INPUT), .Q(sqrto_125_) );
  DFFPOSX1 DFFPOSX1_1300 ( .CLK(clk_bF_buf42), .D(u2_remHi_393__FF_INPUT), .Q(u2_remHi_393_) );
  DFFPOSX1 DFFPOSX1_1301 ( .CLK(clk_bF_buf41), .D(u2_remHi_394__FF_INPUT), .Q(u2_remHi_394_) );
  DFFPOSX1 DFFPOSX1_1302 ( .CLK(clk_bF_buf40), .D(u2_remHi_395__FF_INPUT), .Q(u2_remHi_395_) );
  DFFPOSX1 DFFPOSX1_1303 ( .CLK(clk_bF_buf39), .D(u2_remHi_396__FF_INPUT), .Q(u2_remHi_396_) );
  DFFPOSX1 DFFPOSX1_1304 ( .CLK(clk_bF_buf38), .D(u2_remHi_397__FF_INPUT), .Q(u2_remHi_397_) );
  DFFPOSX1 DFFPOSX1_1305 ( .CLK(clk_bF_buf37), .D(u2_remHi_398__FF_INPUT), .Q(u2_remHi_398_) );
  DFFPOSX1 DFFPOSX1_1306 ( .CLK(clk_bF_buf36), .D(u2_remHi_399__FF_INPUT), .Q(u2_remHi_399_) );
  DFFPOSX1 DFFPOSX1_1307 ( .CLK(clk_bF_buf35), .D(u2_remHi_400__FF_INPUT), .Q(u2_remHi_400_) );
  DFFPOSX1 DFFPOSX1_1308 ( .CLK(clk_bF_buf34), .D(u2_remHi_401__FF_INPUT), .Q(u2_remHi_401_) );
  DFFPOSX1 DFFPOSX1_1309 ( .CLK(clk_bF_buf33), .D(u2_remHi_402__FF_INPUT), .Q(u2_remHi_402_) );
  DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf113), .D(u2_root_127__FF_INPUT), .Q(sqrto_126_) );
  DFFPOSX1 DFFPOSX1_1310 ( .CLK(clk_bF_buf32), .D(u2_remHi_403__FF_INPUT), .Q(u2_remHi_403_) );
  DFFPOSX1 DFFPOSX1_1311 ( .CLK(clk_bF_buf31), .D(u2_remHi_404__FF_INPUT), .Q(u2_remHi_404_) );
  DFFPOSX1 DFFPOSX1_1312 ( .CLK(clk_bF_buf30), .D(u2_remHi_405__FF_INPUT), .Q(u2_remHi_405_) );
  DFFPOSX1 DFFPOSX1_1313 ( .CLK(clk_bF_buf29), .D(u2_remHi_406__FF_INPUT), .Q(u2_remHi_406_) );
  DFFPOSX1 DFFPOSX1_1314 ( .CLK(clk_bF_buf28), .D(u2_remHi_407__FF_INPUT), .Q(u2_remHi_407_) );
  DFFPOSX1 DFFPOSX1_1315 ( .CLK(clk_bF_buf27), .D(u2_remHi_408__FF_INPUT), .Q(u2_remHi_408_) );
  DFFPOSX1 DFFPOSX1_1316 ( .CLK(clk_bF_buf26), .D(u2_remHi_409__FF_INPUT), .Q(u2_remHi_409_) );
  DFFPOSX1 DFFPOSX1_1317 ( .CLK(clk_bF_buf25), .D(u2_remHi_410__FF_INPUT), .Q(u2_remHi_410_) );
  DFFPOSX1 DFFPOSX1_1318 ( .CLK(clk_bF_buf24), .D(u2_remHi_411__FF_INPUT), .Q(u2_remHi_411_) );
  DFFPOSX1 DFFPOSX1_1319 ( .CLK(clk_bF_buf23), .D(u2_remHi_412__FF_INPUT), .Q(u2_remHi_412_) );
  DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf112), .D(u2_root_128__FF_INPUT), .Q(sqrto_127_) );
  DFFPOSX1 DFFPOSX1_1320 ( .CLK(clk_bF_buf22), .D(u2_remHi_413__FF_INPUT), .Q(u2_remHi_413_) );
  DFFPOSX1 DFFPOSX1_1321 ( .CLK(clk_bF_buf21), .D(u2_remHi_414__FF_INPUT), .Q(u2_remHi_414_) );
  DFFPOSX1 DFFPOSX1_1322 ( .CLK(clk_bF_buf20), .D(u2_remHi_415__FF_INPUT), .Q(u2_remHi_415_) );
  DFFPOSX1 DFFPOSX1_1323 ( .CLK(clk_bF_buf19), .D(u2_remHi_416__FF_INPUT), .Q(u2_remHi_416_) );
  DFFPOSX1 DFFPOSX1_1324 ( .CLK(clk_bF_buf18), .D(u2_remHi_417__FF_INPUT), .Q(u2_remHi_417_) );
  DFFPOSX1 DFFPOSX1_1325 ( .CLK(clk_bF_buf17), .D(u2_remHi_418__FF_INPUT), .Q(u2_remHi_418_) );
  DFFPOSX1 DFFPOSX1_1326 ( .CLK(clk_bF_buf16), .D(u2_remHi_419__FF_INPUT), .Q(u2_remHi_419_) );
  DFFPOSX1 DFFPOSX1_1327 ( .CLK(clk_bF_buf15), .D(u2_remHi_420__FF_INPUT), .Q(u2_remHi_420_) );
  DFFPOSX1 DFFPOSX1_1328 ( .CLK(clk_bF_buf14), .D(u2_remHi_421__FF_INPUT), .Q(u2_remHi_421_) );
  DFFPOSX1 DFFPOSX1_1329 ( .CLK(clk_bF_buf13), .D(u2_remHi_422__FF_INPUT), .Q(u2_remHi_422_) );
  DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf111), .D(u2_root_129__FF_INPUT), .Q(sqrto_128_) );
  DFFPOSX1 DFFPOSX1_1330 ( .CLK(clk_bF_buf12), .D(u2_remHi_423__FF_INPUT), .Q(u2_remHi_423_) );
  DFFPOSX1 DFFPOSX1_1331 ( .CLK(clk_bF_buf11), .D(u2_remHi_424__FF_INPUT), .Q(u2_remHi_424_) );
  DFFPOSX1 DFFPOSX1_1332 ( .CLK(clk_bF_buf10), .D(u2_remHi_425__FF_INPUT), .Q(u2_remHi_425_) );
  DFFPOSX1 DFFPOSX1_1333 ( .CLK(clk_bF_buf9), .D(u2_remHi_426__FF_INPUT), .Q(u2_remHi_426_) );
  DFFPOSX1 DFFPOSX1_1334 ( .CLK(clk_bF_buf8), .D(u2_remHi_427__FF_INPUT), .Q(u2_remHi_427_) );
  DFFPOSX1 DFFPOSX1_1335 ( .CLK(clk_bF_buf7), .D(u2_remHi_428__FF_INPUT), .Q(u2_remHi_428_) );
  DFFPOSX1 DFFPOSX1_1336 ( .CLK(clk_bF_buf6), .D(u2_remHi_429__FF_INPUT), .Q(u2_remHi_429_) );
  DFFPOSX1 DFFPOSX1_1337 ( .CLK(clk_bF_buf5), .D(u2_remHi_430__FF_INPUT), .Q(u2_remHi_430_) );
  DFFPOSX1 DFFPOSX1_1338 ( .CLK(clk_bF_buf4), .D(u2_remHi_431__FF_INPUT), .Q(u2_remHi_431_) );
  DFFPOSX1 DFFPOSX1_1339 ( .CLK(clk_bF_buf3), .D(u2_remHi_432__FF_INPUT), .Q(u2_remHi_432_) );
  DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf110), .D(u2_root_130__FF_INPUT), .Q(sqrto_129_) );
  DFFPOSX1 DFFPOSX1_1340 ( .CLK(clk_bF_buf2), .D(u2_remHi_433__FF_INPUT), .Q(u2_remHi_433_) );
  DFFPOSX1 DFFPOSX1_1341 ( .CLK(clk_bF_buf1), .D(u2_remHi_434__FF_INPUT), .Q(u2_remHi_434_) );
  DFFPOSX1 DFFPOSX1_1342 ( .CLK(clk_bF_buf0), .D(u2_remHi_435__FF_INPUT), .Q(u2_remHi_435_) );
  DFFPOSX1 DFFPOSX1_1343 ( .CLK(clk_bF_buf121), .D(u2_remHi_436__FF_INPUT), .Q(u2_remHi_436_) );
  DFFPOSX1 DFFPOSX1_1344 ( .CLK(clk_bF_buf120), .D(u2_remHi_437__FF_INPUT), .Q(u2_remHi_437_) );
  DFFPOSX1 DFFPOSX1_1345 ( .CLK(clk_bF_buf119), .D(u2_remHi_438__FF_INPUT), .Q(u2_remHi_438_) );
  DFFPOSX1 DFFPOSX1_1346 ( .CLK(clk_bF_buf118), .D(u2_remHi_439__FF_INPUT), .Q(u2_remHi_439_) );
  DFFPOSX1 DFFPOSX1_1347 ( .CLK(clk_bF_buf117), .D(u2_remHi_440__FF_INPUT), .Q(u2_remHi_440_) );
  DFFPOSX1 DFFPOSX1_1348 ( .CLK(clk_bF_buf116), .D(u2_remHi_441__FF_INPUT), .Q(u2_remHi_441_) );
  DFFPOSX1 DFFPOSX1_1349 ( .CLK(clk_bF_buf115), .D(u2_remHi_442__FF_INPUT), .Q(u2_remHi_442_) );
  DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf109), .D(u2_root_131__FF_INPUT), .Q(sqrto_130_) );
  DFFPOSX1 DFFPOSX1_1350 ( .CLK(clk_bF_buf114), .D(u2_remHi_443__FF_INPUT), .Q(u2_remHi_443_) );
  DFFPOSX1 DFFPOSX1_1351 ( .CLK(clk_bF_buf113), .D(u2_remHi_444__FF_INPUT), .Q(u2_remHi_444_) );
  DFFPOSX1 DFFPOSX1_1352 ( .CLK(clk_bF_buf112), .D(u2_remHi_445__FF_INPUT), .Q(u2_remHi_445_) );
  DFFPOSX1 DFFPOSX1_1353 ( .CLK(clk_bF_buf111), .D(u2_remHi_446__FF_INPUT), .Q(u2_remHi_446_) );
  DFFPOSX1 DFFPOSX1_1354 ( .CLK(clk_bF_buf110), .D(u2_remHi_447__FF_INPUT), .Q(u2_remHi_447_) );
  DFFPOSX1 DFFPOSX1_1355 ( .CLK(clk_bF_buf109), .D(u2_remHi_448__FF_INPUT), .Q(u2_remHi_448_) );
  DFFPOSX1 DFFPOSX1_1356 ( .CLK(clk_bF_buf108), .D(u2_remHi_449__FF_INPUT), .Q(u2_remHi_449_) );
  DFFPOSX1 DFFPOSX1_1357 ( .CLK(clk_bF_buf107), .D(u2_cnt_0__FF_INPUT), .Q(u2_cnt_0_) );
  DFFPOSX1 DFFPOSX1_1358 ( .CLK(clk_bF_buf106), .D(u2_cnt_1__FF_INPUT), .Q(u2_cnt_1_) );
  DFFPOSX1 DFFPOSX1_1359 ( .CLK(clk_bF_buf105), .D(u2_cnt_2__FF_INPUT), .Q(u2_cnt_2_) );
  DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf108), .D(u2_root_132__FF_INPUT), .Q(sqrto_131_) );
  DFFPOSX1 DFFPOSX1_1360 ( .CLK(clk_bF_buf104), .D(u2_cnt_3__FF_INPUT), .Q(u2_cnt_3_) );
  DFFPOSX1 DFFPOSX1_1361 ( .CLK(clk_bF_buf103), .D(u2_cnt_4__FF_INPUT), .Q(u2_cnt_4_) );
  DFFPOSX1 DFFPOSX1_1362 ( .CLK(clk_bF_buf102), .D(u2_cnt_5__FF_INPUT), .Q(u2_cnt_5_) );
  DFFPOSX1 DFFPOSX1_1363 ( .CLK(clk_bF_buf101), .D(u2_cnt_6__FF_INPUT), .Q(u2_cnt_6_) );
  DFFPOSX1 DFFPOSX1_1364 ( .CLK(clk_bF_buf100), .D(u2_cnt_7__FF_INPUT), .Q(u2_cnt_7_) );
  DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf107), .D(u2_root_133__FF_INPUT), .Q(sqrto_132_) );
  DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf106), .D(u2_root_134__FF_INPUT), .Q(sqrto_133_) );
  DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf105), .D(u2_root_135__FF_INPUT), .Q(sqrto_134_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf108), .D(u2_root_10__FF_INPUT), .Q(sqrto_9_) );
  DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf104), .D(u2_root_136__FF_INPUT), .Q(sqrto_135_) );
  DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf103), .D(u2_root_137__FF_INPUT), .Q(sqrto_136_) );
  DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf102), .D(u2_root_138__FF_INPUT), .Q(sqrto_137_) );
  DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf101), .D(u2_root_139__FF_INPUT), .Q(sqrto_138_) );
  DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf100), .D(u2_root_140__FF_INPUT), .Q(sqrto_139_) );
  DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf99), .D(u2_root_141__FF_INPUT), .Q(sqrto_140_) );
  DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf98), .D(u2_root_142__FF_INPUT), .Q(sqrto_141_) );
  DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf97), .D(u2_root_143__FF_INPUT), .Q(sqrto_142_) );
  DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf96), .D(u2_root_144__FF_INPUT), .Q(sqrto_143_) );
  DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf95), .D(u2_root_145__FF_INPUT), .Q(sqrto_144_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf107), .D(u2_root_11__FF_INPUT), .Q(sqrto_10_) );
  DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf94), .D(u2_root_146__FF_INPUT), .Q(sqrto_145_) );
  DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf93), .D(u2_root_147__FF_INPUT), .Q(sqrto_146_) );
  DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf92), .D(u2_root_148__FF_INPUT), .Q(sqrto_147_) );
  DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf91), .D(u2_root_149__FF_INPUT), .Q(sqrto_148_) );
  DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf90), .D(u2_root_150__FF_INPUT), .Q(sqrto_149_) );
  DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf89), .D(u2_root_151__FF_INPUT), .Q(sqrto_150_) );
  DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf88), .D(u2_root_152__FF_INPUT), .Q(sqrto_151_) );
  DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf87), .D(u2_root_153__FF_INPUT), .Q(sqrto_152_) );
  DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf86), .D(u2_root_154__FF_INPUT), .Q(sqrto_153_) );
  DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf85), .D(u2_root_155__FF_INPUT), .Q(sqrto_154_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf106), .D(u2_root_12__FF_INPUT), .Q(sqrto_11_) );
  DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf84), .D(u2_root_156__FF_INPUT), .Q(sqrto_155_) );
  DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf83), .D(u2_root_157__FF_INPUT), .Q(sqrto_156_) );
  DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf82), .D(u2_root_158__FF_INPUT), .Q(sqrto_157_) );
  DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf81), .D(u2_root_159__FF_INPUT), .Q(sqrto_158_) );
  DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf80), .D(u2_root_160__FF_INPUT), .Q(sqrto_159_) );
  DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf79), .D(u2_root_161__FF_INPUT), .Q(sqrto_160_) );
  DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf78), .D(u2_root_162__FF_INPUT), .Q(sqrto_161_) );
  DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf77), .D(u2_root_163__FF_INPUT), .Q(sqrto_162_) );
  DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf76), .D(u2_root_164__FF_INPUT), .Q(sqrto_163_) );
  DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf75), .D(u2_root_165__FF_INPUT), .Q(sqrto_164_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf105), .D(u2_root_13__FF_INPUT), .Q(sqrto_12_) );
  DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf74), .D(u2_root_166__FF_INPUT), .Q(sqrto_165_) );
  DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf73), .D(u2_root_167__FF_INPUT), .Q(sqrto_166_) );
  DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf72), .D(u2_root_168__FF_INPUT), .Q(sqrto_167_) );
  DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf71), .D(u2_root_169__FF_INPUT), .Q(sqrto_168_) );
  DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf70), .D(u2_root_170__FF_INPUT), .Q(sqrto_169_) );
  DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf69), .D(u2_root_171__FF_INPUT), .Q(sqrto_170_) );
  DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf68), .D(u2_root_172__FF_INPUT), .Q(sqrto_171_) );
  DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf67), .D(u2_root_173__FF_INPUT), .Q(sqrto_172_) );
  DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf66), .D(u2_root_174__FF_INPUT), .Q(sqrto_173_) );
  DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf65), .D(u2_root_175__FF_INPUT), .Q(sqrto_174_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf104), .D(u2_root_14__FF_INPUT), .Q(sqrto_13_) );
  DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf64), .D(u2_root_176__FF_INPUT), .Q(sqrto_175_) );
  DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf63), .D(u2_root_177__FF_INPUT), .Q(sqrto_176_) );
  DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf62), .D(u2_root_178__FF_INPUT), .Q(sqrto_177_) );
  DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf61), .D(u2_root_179__FF_INPUT), .Q(sqrto_178_) );
  DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf60), .D(u2_root_180__FF_INPUT), .Q(sqrto_179_) );
  DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf59), .D(u2_root_181__FF_INPUT), .Q(sqrto_180_) );
  DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf58), .D(u2_root_182__FF_INPUT), .Q(sqrto_181_) );
  DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf57), .D(u2_root_183__FF_INPUT), .Q(sqrto_182_) );
  DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf56), .D(u2_root_184__FF_INPUT), .Q(sqrto_183_) );
  DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf55), .D(u2_root_185__FF_INPUT), .Q(sqrto_184_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf103), .D(u2_root_15__FF_INPUT), .Q(sqrto_14_) );
  DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf54), .D(u2_root_186__FF_INPUT), .Q(sqrto_185_) );
  DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf53), .D(u2_root_187__FF_INPUT), .Q(sqrto_186_) );
  DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf52), .D(u2_root_188__FF_INPUT), .Q(sqrto_187_) );
  DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf51), .D(u2_root_189__FF_INPUT), .Q(sqrto_188_) );
  DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf50), .D(u2_root_190__FF_INPUT), .Q(sqrto_189_) );
  DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf49), .D(u2_root_191__FF_INPUT), .Q(sqrto_190_) );
  DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf48), .D(u2_root_192__FF_INPUT), .Q(sqrto_191_) );
  DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf47), .D(u2_root_193__FF_INPUT), .Q(sqrto_192_) );
  DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf46), .D(u2_root_194__FF_INPUT), .Q(sqrto_193_) );
  DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf45), .D(u2_root_195__FF_INPUT), .Q(sqrto_194_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf120), .D(u2__abc_29664_n3927), .Q(_auto_iopadmap_cc_313_execute_65412) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf102), .D(u2_root_16__FF_INPUT), .Q(sqrto_15_) );
  DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf44), .D(u2_root_196__FF_INPUT), .Q(sqrto_195_) );
  DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf43), .D(u2_root_197__FF_INPUT), .Q(sqrto_196_) );
  DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf42), .D(u2_root_198__FF_INPUT), .Q(sqrto_197_) );
  DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf41), .D(u2_root_199__FF_INPUT), .Q(sqrto_198_) );
  DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf40), .D(u2_root_200__FF_INPUT), .Q(sqrto_199_) );
  DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf39), .D(u2_root_201__FF_INPUT), .Q(sqrto_200_) );
  DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf38), .D(u2_root_202__FF_INPUT), .Q(sqrto_201_) );
  DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf37), .D(u2_root_203__FF_INPUT), .Q(sqrto_202_) );
  DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf36), .D(u2_root_204__FF_INPUT), .Q(sqrto_203_) );
  DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf35), .D(u2_root_205__FF_INPUT), .Q(sqrto_204_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf101), .D(u2_root_17__FF_INPUT), .Q(sqrto_16_) );
  DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf34), .D(u2_root_206__FF_INPUT), .Q(sqrto_205_) );
  DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf33), .D(u2_root_207__FF_INPUT), .Q(sqrto_206_) );
  DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf32), .D(u2_root_208__FF_INPUT), .Q(sqrto_207_) );
  DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf31), .D(u2_root_209__FF_INPUT), .Q(sqrto_208_) );
  DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf30), .D(u2_root_210__FF_INPUT), .Q(sqrto_209_) );
  DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf29), .D(u2_root_211__FF_INPUT), .Q(sqrto_210_) );
  DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf28), .D(u2_root_212__FF_INPUT), .Q(sqrto_211_) );
  DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf27), .D(u2_root_213__FF_INPUT), .Q(sqrto_212_) );
  DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf26), .D(u2_root_214__FF_INPUT), .Q(sqrto_213_) );
  DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf25), .D(u2_root_215__FF_INPUT), .Q(sqrto_214_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf100), .D(u2_root_18__FF_INPUT), .Q(sqrto_17_) );
  DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf24), .D(u2_root_216__FF_INPUT), .Q(sqrto_215_) );
  DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf23), .D(u2_root_217__FF_INPUT), .Q(sqrto_216_) );
  DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf22), .D(u2_root_218__FF_INPUT), .Q(sqrto_217_) );
  DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf21), .D(u2_root_219__FF_INPUT), .Q(sqrto_218_) );
  DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf20), .D(u2_root_220__FF_INPUT), .Q(sqrto_219_) );
  DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf19), .D(u2_root_221__FF_INPUT), .Q(sqrto_220_) );
  DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf18), .D(u2_root_222__FF_INPUT), .Q(sqrto_221_) );
  DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf17), .D(u2_root_223__FF_INPUT), .Q(sqrto_222_) );
  DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf16), .D(u2_root_224__FF_INPUT), .Q(sqrto_223_) );
  DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf15), .D(u2_root_225__FF_INPUT), .Q(sqrto_224_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf99), .D(u2_root_19__FF_INPUT), .Q(sqrto_18_) );
  DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf14), .D(u2_root_226__FF_INPUT), .Q(sqrto_225_) );
  DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf13), .D(u2_root_227__FF_INPUT), .Q(u2_o_226_) );
  DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf12), .D(u2_root_228__FF_INPUT), .Q(u2_o_227_) );
  DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf11), .D(u2_root_229__FF_INPUT), .Q(u2_o_228_) );
  DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf10), .D(u2_root_230__FF_INPUT), .Q(u2_o_229_) );
  DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf9), .D(u2_root_231__FF_INPUT), .Q(u2_o_230_) );
  DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf8), .D(u2_root_232__FF_INPUT), .Q(u2_o_231_) );
  DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf7), .D(u2_root_233__FF_INPUT), .Q(u2_o_232_) );
  DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf6), .D(u2_root_234__FF_INPUT), .Q(u2_o_233_) );
  DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf5), .D(u2_root_235__FF_INPUT), .Q(u2_o_234_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf98), .D(u2_root_20__FF_INPUT), .Q(sqrto_19_) );
  DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf4), .D(u2_root_236__FF_INPUT), .Q(u2_o_235_) );
  DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf3), .D(u2_root_237__FF_INPUT), .Q(u2_o_236_) );
  DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf2), .D(u2_root_238__FF_INPUT), .Q(u2_o_237_) );
  DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf1), .D(u2_root_239__FF_INPUT), .Q(u2_o_238_) );
  DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf0), .D(u2_root_240__FF_INPUT), .Q(u2_o_239_) );
  DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf121), .D(u2_root_241__FF_INPUT), .Q(u2_o_240_) );
  DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf120), .D(u2_root_242__FF_INPUT), .Q(u2_o_241_) );
  DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf119), .D(u2_root_243__FF_INPUT), .Q(u2_o_242_) );
  DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf118), .D(u2_root_244__FF_INPUT), .Q(u2_o_243_) );
  DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf117), .D(u2_root_245__FF_INPUT), .Q(u2_o_244_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf97), .D(u2_root_21__FF_INPUT), .Q(sqrto_20_) );
  DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf116), .D(u2_root_246__FF_INPUT), .Q(u2_o_245_) );
  DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf115), .D(u2_root_247__FF_INPUT), .Q(u2_o_246_) );
  DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf114), .D(u2_root_248__FF_INPUT), .Q(u2_o_247_) );
  DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf113), .D(u2_root_249__FF_INPUT), .Q(u2_o_248_) );
  DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf112), .D(u2_root_250__FF_INPUT), .Q(u2_o_249_) );
  DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf111), .D(u2_root_251__FF_INPUT), .Q(u2_o_250_) );
  DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf110), .D(u2_root_252__FF_INPUT), .Q(u2_o_251_) );
  DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf109), .D(u2_root_253__FF_INPUT), .Q(u2_o_252_) );
  DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf108), .D(u2_root_254__FF_INPUT), .Q(u2_o_253_) );
  DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf107), .D(u2_root_255__FF_INPUT), .Q(u2_o_254_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf96), .D(u2_root_22__FF_INPUT), .Q(sqrto_21_) );
  DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf106), .D(u2_root_256__FF_INPUT), .Q(u2_o_255_) );
  DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf105), .D(u2_root_257__FF_INPUT), .Q(u2_o_256_) );
  DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf104), .D(u2_root_258__FF_INPUT), .Q(u2_o_257_) );
  DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf103), .D(u2_root_259__FF_INPUT), .Q(u2_o_258_) );
  DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf102), .D(u2_root_260__FF_INPUT), .Q(u2_o_259_) );
  DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf101), .D(u2_root_261__FF_INPUT), .Q(u2_o_260_) );
  DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf100), .D(u2_root_262__FF_INPUT), .Q(u2_o_261_) );
  DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf99), .D(u2_root_263__FF_INPUT), .Q(u2_o_262_) );
  DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf98), .D(u2_root_264__FF_INPUT), .Q(u2_o_263_) );
  DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf97), .D(u2_root_265__FF_INPUT), .Q(u2_o_264_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf95), .D(u2_root_23__FF_INPUT), .Q(sqrto_22_) );
  DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf96), .D(u2_root_266__FF_INPUT), .Q(u2_o_265_) );
  DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf95), .D(u2_root_267__FF_INPUT), .Q(u2_o_266_) );
  DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf94), .D(u2_root_268__FF_INPUT), .Q(u2_o_267_) );
  DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf93), .D(u2_root_269__FF_INPUT), .Q(u2_o_268_) );
  DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf92), .D(u2_root_270__FF_INPUT), .Q(u2_o_269_) );
  DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf91), .D(u2_root_271__FF_INPUT), .Q(u2_o_270_) );
  DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf90), .D(u2_root_272__FF_INPUT), .Q(u2_o_271_) );
  DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf89), .D(u2_root_273__FF_INPUT), .Q(u2_o_272_) );
  DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf88), .D(u2_root_274__FF_INPUT), .Q(u2_o_273_) );
  DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf87), .D(u2_root_275__FF_INPUT), .Q(u2_o_274_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf94), .D(u2_root_24__FF_INPUT), .Q(sqrto_23_) );
  DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf86), .D(u2_root_276__FF_INPUT), .Q(u2_o_275_) );
  DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf85), .D(u2_root_277__FF_INPUT), .Q(u2_o_276_) );
  DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf84), .D(u2_root_278__FF_INPUT), .Q(u2_o_277_) );
  DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf83), .D(u2_root_279__FF_INPUT), .Q(u2_o_278_) );
  DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf82), .D(u2_root_280__FF_INPUT), .Q(u2_o_279_) );
  DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf81), .D(u2_root_281__FF_INPUT), .Q(u2_o_280_) );
  DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf80), .D(u2_root_282__FF_INPUT), .Q(u2_o_281_) );
  DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf79), .D(u2_root_283__FF_INPUT), .Q(u2_o_282_) );
  DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf78), .D(u2_root_284__FF_INPUT), .Q(u2_o_283_) );
  DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf77), .D(u2_root_285__FF_INPUT), .Q(u2_o_284_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf93), .D(u2_root_25__FF_INPUT), .Q(sqrto_24_) );
  DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf76), .D(u2_root_286__FF_INPUT), .Q(u2_o_285_) );
  DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf75), .D(u2_root_287__FF_INPUT), .Q(u2_o_286_) );
  DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf74), .D(u2_root_288__FF_INPUT), .Q(u2_o_287_) );
  DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf73), .D(u2_root_289__FF_INPUT), .Q(u2_o_288_) );
  DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf72), .D(u2_root_290__FF_INPUT), .Q(u2_o_289_) );
  DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf71), .D(u2_root_291__FF_INPUT), .Q(u2_o_290_) );
  DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf70), .D(u2_root_292__FF_INPUT), .Q(u2_o_291_) );
  DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf69), .D(u2_root_293__FF_INPUT), .Q(u2_o_292_) );
  DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf68), .D(u2_root_294__FF_INPUT), .Q(u2_o_293_) );
  DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf67), .D(u2_root_295__FF_INPUT), .Q(u2_o_294_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf119), .D(u2__abc_29664_n3922), .Q(u2_state_2_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf92), .D(u2_root_26__FF_INPUT), .Q(sqrto_25_) );
  DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf66), .D(u2_root_296__FF_INPUT), .Q(u2_o_295_) );
  DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf65), .D(u2_root_297__FF_INPUT), .Q(u2_o_296_) );
  DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf64), .D(u2_root_298__FF_INPUT), .Q(u2_o_297_) );
  DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf63), .D(u2_root_299__FF_INPUT), .Q(u2_o_298_) );
  DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf62), .D(u2_root_300__FF_INPUT), .Q(u2_o_299_) );
  DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf61), .D(u2_root_301__FF_INPUT), .Q(u2_o_300_) );
  DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf60), .D(u2_root_302__FF_INPUT), .Q(u2_o_301_) );
  DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf59), .D(u2_root_303__FF_INPUT), .Q(u2_o_302_) );
  DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf58), .D(u2_root_304__FF_INPUT), .Q(u2_o_303_) );
  DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf57), .D(u2_root_305__FF_INPUT), .Q(u2_o_304_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf91), .D(u2_root_27__FF_INPUT), .Q(sqrto_26_) );
  DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf56), .D(u2_root_306__FF_INPUT), .Q(u2_o_305_) );
  DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf55), .D(u2_root_307__FF_INPUT), .Q(u2_o_306_) );
  DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf54), .D(u2_root_308__FF_INPUT), .Q(u2_o_307_) );
  DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf53), .D(u2_root_309__FF_INPUT), .Q(u2_o_308_) );
  DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf52), .D(u2_root_310__FF_INPUT), .Q(u2_o_309_) );
  DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf51), .D(u2_root_311__FF_INPUT), .Q(u2_o_310_) );
  DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf50), .D(u2_root_312__FF_INPUT), .Q(u2_o_311_) );
  DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf49), .D(u2_root_313__FF_INPUT), .Q(u2_o_312_) );
  DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf48), .D(u2_root_314__FF_INPUT), .Q(u2_o_313_) );
  DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf47), .D(u2_root_315__FF_INPUT), .Q(u2_o_314_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf90), .D(u2_root_28__FF_INPUT), .Q(sqrto_27_) );
  DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf46), .D(u2_root_316__FF_INPUT), .Q(u2_o_315_) );
  DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf45), .D(u2_root_317__FF_INPUT), .Q(u2_o_316_) );
  DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf44), .D(u2_root_318__FF_INPUT), .Q(u2_o_317_) );
  DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf43), .D(u2_root_319__FF_INPUT), .Q(u2_o_318_) );
  DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf42), .D(u2_root_320__FF_INPUT), .Q(u2_o_319_) );
  DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf41), .D(u2_root_321__FF_INPUT), .Q(u2_o_320_) );
  DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf40), .D(u2_root_322__FF_INPUT), .Q(u2_o_321_) );
  DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf39), .D(u2_root_323__FF_INPUT), .Q(u2_o_322_) );
  DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf38), .D(u2_root_324__FF_INPUT), .Q(u2_o_323_) );
  DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf37), .D(u2_root_325__FF_INPUT), .Q(u2_o_324_) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf89), .D(u2_root_29__FF_INPUT), .Q(sqrto_28_) );
  DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf36), .D(u2_root_326__FF_INPUT), .Q(u2_o_325_) );
  DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf35), .D(u2_root_327__FF_INPUT), .Q(u2_o_326_) );
  DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf34), .D(u2_root_328__FF_INPUT), .Q(u2_o_327_) );
  DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf33), .D(u2_root_329__FF_INPUT), .Q(u2_o_328_) );
  DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf32), .D(u2_root_330__FF_INPUT), .Q(u2_o_329_) );
  DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf31), .D(u2_root_331__FF_INPUT), .Q(u2_o_330_) );
  DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf30), .D(u2_root_332__FF_INPUT), .Q(u2_o_331_) );
  DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf29), .D(u2_root_333__FF_INPUT), .Q(u2_o_332_) );
  DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf28), .D(u2_root_334__FF_INPUT), .Q(u2_o_333_) );
  DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf27), .D(u2_root_335__FF_INPUT), .Q(u2_o_334_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf88), .D(u2_root_30__FF_INPUT), .Q(sqrto_29_) );
  DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf26), .D(u2_root_336__FF_INPUT), .Q(u2_o_335_) );
  DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf25), .D(u2_root_337__FF_INPUT), .Q(u2_o_336_) );
  DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf24), .D(u2_root_338__FF_INPUT), .Q(u2_o_337_) );
  DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf23), .D(u2_root_339__FF_INPUT), .Q(u2_o_338_) );
  DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf22), .D(u2_root_340__FF_INPUT), .Q(u2_o_339_) );
  DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf21), .D(u2_root_341__FF_INPUT), .Q(u2_o_340_) );
  DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf20), .D(u2_root_342__FF_INPUT), .Q(u2_o_341_) );
  DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf19), .D(u2_root_343__FF_INPUT), .Q(u2_o_342_) );
  DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf18), .D(u2_root_344__FF_INPUT), .Q(u2_o_343_) );
  DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf17), .D(u2_root_345__FF_INPUT), .Q(u2_o_344_) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf87), .D(u2_root_31__FF_INPUT), .Q(sqrto_30_) );
  DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf16), .D(u2_root_346__FF_INPUT), .Q(u2_o_345_) );
  DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf15), .D(u2_root_347__FF_INPUT), .Q(u2_o_346_) );
  DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf14), .D(u2_root_348__FF_INPUT), .Q(u2_o_347_) );
  DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf13), .D(u2_root_349__FF_INPUT), .Q(u2_o_348_) );
  DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf12), .D(u2_root_350__FF_INPUT), .Q(u2_o_349_) );
  DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf11), .D(u2_root_351__FF_INPUT), .Q(u2_o_350_) );
  DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf10), .D(u2_root_352__FF_INPUT), .Q(u2_o_351_) );
  DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf9), .D(u2_root_353__FF_INPUT), .Q(u2_o_352_) );
  DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf8), .D(u2_root_354__FF_INPUT), .Q(u2_o_353_) );
  DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf7), .D(u2_root_355__FF_INPUT), .Q(u2_o_354_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf86), .D(u2_root_32__FF_INPUT), .Q(sqrto_31_) );
  DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf6), .D(u2_root_356__FF_INPUT), .Q(u2_o_355_) );
  DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf5), .D(u2_root_357__FF_INPUT), .Q(u2_o_356_) );
  DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf4), .D(u2_root_358__FF_INPUT), .Q(u2_o_357_) );
  DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf3), .D(u2_root_359__FF_INPUT), .Q(u2_o_358_) );
  DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf2), .D(u2_root_360__FF_INPUT), .Q(u2_o_359_) );
  DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf1), .D(u2_root_361__FF_INPUT), .Q(u2_o_360_) );
  DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf0), .D(u2_root_362__FF_INPUT), .Q(u2_o_361_) );
  DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf121), .D(u2_root_363__FF_INPUT), .Q(u2_o_362_) );
  DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf120), .D(u2_root_364__FF_INPUT), .Q(u2_o_363_) );
  DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf119), .D(u2_root_365__FF_INPUT), .Q(u2_o_364_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf85), .D(u2_root_33__FF_INPUT), .Q(sqrto_32_) );
  DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf118), .D(u2_root_366__FF_INPUT), .Q(u2_o_365_) );
  DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf117), .D(u2_root_367__FF_INPUT), .Q(u2_o_366_) );
  DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf116), .D(u2_root_368__FF_INPUT), .Q(u2_o_367_) );
  DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf115), .D(u2_root_369__FF_INPUT), .Q(u2_o_368_) );
  DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf114), .D(u2_root_370__FF_INPUT), .Q(u2_o_369_) );
  DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf113), .D(u2_root_371__FF_INPUT), .Q(u2_o_370_) );
  DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf112), .D(u2_root_372__FF_INPUT), .Q(u2_o_371_) );
  DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf111), .D(u2_root_373__FF_INPUT), .Q(u2_o_372_) );
  DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf110), .D(u2_root_374__FF_INPUT), .Q(u2_o_373_) );
  DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf109), .D(u2_root_375__FF_INPUT), .Q(u2_o_374_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf84), .D(u2_root_34__FF_INPUT), .Q(sqrto_33_) );
  DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf108), .D(u2_root_376__FF_INPUT), .Q(u2_o_375_) );
  DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf107), .D(u2_root_377__FF_INPUT), .Q(u2_o_376_) );
  DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf106), .D(u2_root_378__FF_INPUT), .Q(u2_o_377_) );
  DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf105), .D(u2_root_379__FF_INPUT), .Q(u2_o_378_) );
  DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf104), .D(u2_root_380__FF_INPUT), .Q(u2_o_379_) );
  DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf103), .D(u2_root_381__FF_INPUT), .Q(u2_o_380_) );
  DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf102), .D(u2_root_382__FF_INPUT), .Q(u2_o_381_) );
  DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf101), .D(u2_root_383__FF_INPUT), .Q(u2_o_382_) );
  DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf100), .D(u2_root_384__FF_INPUT), .Q(u2_o_383_) );
  DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf99), .D(u2_root_385__FF_INPUT), .Q(u2_o_384_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf83), .D(u2_root_35__FF_INPUT), .Q(sqrto_34_) );
  DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf98), .D(u2_root_386__FF_INPUT), .Q(u2_o_385_) );
  DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf97), .D(u2_root_387__FF_INPUT), .Q(u2_o_386_) );
  DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf96), .D(u2_root_388__FF_INPUT), .Q(u2_o_387_) );
  DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf95), .D(u2_root_389__FF_INPUT), .Q(u2_o_388_) );
  DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf94), .D(u2_root_390__FF_INPUT), .Q(u2_o_389_) );
  DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf93), .D(u2_root_391__FF_INPUT), .Q(u2_o_390_) );
  DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf92), .D(u2_root_392__FF_INPUT), .Q(u2_o_391_) );
  DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf91), .D(u2_root_393__FF_INPUT), .Q(u2_o_392_) );
  DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf90), .D(u2_root_394__FF_INPUT), .Q(u2_o_393_) );
  DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf89), .D(u2_root_395__FF_INPUT), .Q(u2_o_394_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf118), .D(u2_root_0__FF_INPUT), .Q(u2_root_0_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf82), .D(u2_root_36__FF_INPUT), .Q(sqrto_35_) );
  DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf88), .D(u2_root_396__FF_INPUT), .Q(u2_o_395_) );
  DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf87), .D(u2_root_397__FF_INPUT), .Q(u2_o_396_) );
  DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf86), .D(u2_root_398__FF_INPUT), .Q(u2_o_397_) );
  DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf85), .D(u2_root_399__FF_INPUT), .Q(u2_o_398_) );
  DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf84), .D(u2_root_400__FF_INPUT), .Q(u2_o_399_) );
  DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf83), .D(u2_root_401__FF_INPUT), .Q(u2_o_400_) );
  DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf82), .D(u2_root_402__FF_INPUT), .Q(u2_o_401_) );
  DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf81), .D(u2_root_403__FF_INPUT), .Q(u2_o_402_) );
  DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf80), .D(u2_root_404__FF_INPUT), .Q(u2_o_403_) );
  DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf79), .D(u2_root_405__FF_INPUT), .Q(u2_o_404_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf81), .D(u2_root_37__FF_INPUT), .Q(sqrto_36_) );
  DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf78), .D(u2_root_406__FF_INPUT), .Q(u2_o_405_) );
  DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf77), .D(u2_root_407__FF_INPUT), .Q(u2_o_406_) );
  DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf76), .D(u2_root_408__FF_INPUT), .Q(u2_o_407_) );
  DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf75), .D(u2_root_409__FF_INPUT), .Q(u2_o_408_) );
  DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf74), .D(u2_root_410__FF_INPUT), .Q(u2_o_409_) );
  DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf73), .D(u2_root_411__FF_INPUT), .Q(u2_o_410_) );
  DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf72), .D(u2_root_412__FF_INPUT), .Q(u2_o_411_) );
  DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf71), .D(u2_root_413__FF_INPUT), .Q(u2_o_412_) );
  DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf70), .D(u2_root_414__FF_INPUT), .Q(u2_o_413_) );
  DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf69), .D(u2_root_415__FF_INPUT), .Q(u2_o_414_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf80), .D(u2_root_38__FF_INPUT), .Q(sqrto_37_) );
  DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf68), .D(u2_root_416__FF_INPUT), .Q(u2_o_415_) );
  DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf67), .D(u2_root_417__FF_INPUT), .Q(u2_o_416_) );
  DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf66), .D(u2_root_418__FF_INPUT), .Q(u2_o_417_) );
  DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf65), .D(u2_root_419__FF_INPUT), .Q(u2_o_418_) );
  DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf64), .D(u2_root_420__FF_INPUT), .Q(u2_o_419_) );
  DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf63), .D(u2_root_421__FF_INPUT), .Q(u2_o_420_) );
  DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf62), .D(u2_root_422__FF_INPUT), .Q(u2_o_421_) );
  DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf61), .D(u2_root_423__FF_INPUT), .Q(u2_o_422_) );
  DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf60), .D(u2_root_424__FF_INPUT), .Q(u2_o_423_) );
  DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf59), .D(u2_root_425__FF_INPUT), .Q(u2_o_424_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf79), .D(u2_root_39__FF_INPUT), .Q(sqrto_38_) );
  DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf58), .D(u2_root_426__FF_INPUT), .Q(u2_o_425_) );
  DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf57), .D(u2_root_427__FF_INPUT), .Q(u2_o_426_) );
  DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf56), .D(u2_root_428__FF_INPUT), .Q(u2_o_427_) );
  DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf55), .D(u2_root_429__FF_INPUT), .Q(u2_o_428_) );
  DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf54), .D(u2_root_430__FF_INPUT), .Q(u2_o_429_) );
  DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf53), .D(u2_root_431__FF_INPUT), .Q(u2_o_430_) );
  DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf52), .D(u2_root_432__FF_INPUT), .Q(u2_o_431_) );
  DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf51), .D(u2_root_433__FF_INPUT), .Q(u2_o_432_) );
  DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf50), .D(u2_root_434__FF_INPUT), .Q(u2_o_433_) );
  DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf49), .D(u2_root_435__FF_INPUT), .Q(u2_o_434_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf78), .D(u2_root_40__FF_INPUT), .Q(sqrto_39_) );
  DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf48), .D(u2_root_436__FF_INPUT), .Q(u2_o_435_) );
  DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf47), .D(u2_root_437__FF_INPUT), .Q(u2_o_436_) );
  DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf46), .D(u2_root_438__FF_INPUT), .Q(u2_o_437_) );
  DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf45), .D(u2_root_439__FF_INPUT), .Q(u2_o_438_) );
  DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf44), .D(u2_root_440__FF_INPUT), .Q(u2_o_439_) );
  DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf43), .D(u2_root_441__FF_INPUT), .Q(u2_o_440_) );
  DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf42), .D(u2_root_442__FF_INPUT), .Q(u2_o_441_) );
  DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf41), .D(u2_root_443__FF_INPUT), .Q(u2_o_442_) );
  DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf40), .D(u2_root_444__FF_INPUT), .Q(u2_o_443_) );
  DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf39), .D(u2_root_445__FF_INPUT), .Q(u2_o_444_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf77), .D(u2_root_41__FF_INPUT), .Q(sqrto_40_) );
  DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf38), .D(u2_root_446__FF_INPUT), .Q(u2_o_445_) );
  DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf37), .D(u2_root_447__FF_INPUT), .Q(u2_o_446_) );
  DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf36), .D(u2_root_448__FF_INPUT), .Q(u2_o_447_) );
  DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf35), .D(u2_root_449__FF_INPUT), .Q(u2_o_448_) );
  DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf34), .D(u2_root_450__FF_INPUT), .Q(u2_o_449_) );
  DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf33), .D(u2_remLo_0__FF_INPUT), .Q(u2_remLo_0_) );
  DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf32), .D(u2_remLo_1__FF_INPUT), .Q(u2_remLo_1_) );
  DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf31), .D(u2_remLo_2__FF_INPUT), .Q(u2_remLo_2_) );
  DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf30), .D(u2_remLo_3__FF_INPUT), .Q(u2_remLo_3_) );
  DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf29), .D(u2_remLo_4__FF_INPUT), .Q(u2_remLo_4_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf76), .D(u2_root_42__FF_INPUT), .Q(sqrto_41_) );
  DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf28), .D(u2_remLo_5__FF_INPUT), .Q(u2_remLo_5_) );
  DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf27), .D(u2_remLo_6__FF_INPUT), .Q(u2_remLo_6_) );
  DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf26), .D(u2_remLo_7__FF_INPUT), .Q(u2_remLo_7_) );
  DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf25), .D(u2_remLo_8__FF_INPUT), .Q(u2_remLo_8_) );
  DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf24), .D(u2_remLo_9__FF_INPUT), .Q(u2_remLo_9_) );
  DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf23), .D(u2_remLo_10__FF_INPUT), .Q(u2_remLo_10_) );
  DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf22), .D(u2_remLo_11__FF_INPUT), .Q(u2_remLo_11_) );
  DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf21), .D(u2_remLo_12__FF_INPUT), .Q(u2_remLo_12_) );
  DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf20), .D(u2_remLo_13__FF_INPUT), .Q(u2_remLo_13_) );
  DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf19), .D(u2_remLo_14__FF_INPUT), .Q(u2_remLo_14_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf75), .D(u2_root_43__FF_INPUT), .Q(sqrto_42_) );
  DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf18), .D(u2_remLo_15__FF_INPUT), .Q(u2_remLo_15_) );
  DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf17), .D(u2_remLo_16__FF_INPUT), .Q(u2_remLo_16_) );
  DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf16), .D(u2_remLo_17__FF_INPUT), .Q(u2_remLo_17_) );
  DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf15), .D(u2_remLo_18__FF_INPUT), .Q(u2_remLo_18_) );
  DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf14), .D(u2_remLo_19__FF_INPUT), .Q(u2_remLo_19_) );
  DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf13), .D(u2_remLo_20__FF_INPUT), .Q(u2_remLo_20_) );
  DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf12), .D(u2_remLo_21__FF_INPUT), .Q(u2_remLo_21_) );
  DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf11), .D(u2_remLo_22__FF_INPUT), .Q(u2_remLo_22_) );
  DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf10), .D(u2_remLo_23__FF_INPUT), .Q(u2_remLo_23_) );
  DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf9), .D(u2_remLo_24__FF_INPUT), .Q(u2_remLo_24_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf74), .D(u2_root_44__FF_INPUT), .Q(sqrto_43_) );
  DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf8), .D(u2_remLo_25__FF_INPUT), .Q(u2_remLo_25_) );
  DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf7), .D(u2_remLo_26__FF_INPUT), .Q(u2_remLo_26_) );
  DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf6), .D(u2_remLo_27__FF_INPUT), .Q(u2_remLo_27_) );
  DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf5), .D(u2_remLo_28__FF_INPUT), .Q(u2_remLo_28_) );
  DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf4), .D(u2_remLo_29__FF_INPUT), .Q(u2_remLo_29_) );
  DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf3), .D(u2_remLo_30__FF_INPUT), .Q(u2_remLo_30_) );
  DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf2), .D(u2_remLo_31__FF_INPUT), .Q(u2_remLo_31_) );
  DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf1), .D(u2_remLo_32__FF_INPUT), .Q(u2_remLo_32_) );
  DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf0), .D(u2_remLo_33__FF_INPUT), .Q(u2_remLo_33_) );
  DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf121), .D(u2_remLo_34__FF_INPUT), .Q(u2_remLo_34_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf73), .D(u2_root_45__FF_INPUT), .Q(sqrto_44_) );
  DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf120), .D(u2_remLo_35__FF_INPUT), .Q(u2_remLo_35_) );
  DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf119), .D(u2_remLo_36__FF_INPUT), .Q(u2_remLo_36_) );
  DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf118), .D(u2_remLo_37__FF_INPUT), .Q(u2_remLo_37_) );
  DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf117), .D(u2_remLo_38__FF_INPUT), .Q(u2_remLo_38_) );
  DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf116), .D(u2_remLo_39__FF_INPUT), .Q(u2_remLo_39_) );
  DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf115), .D(u2_remLo_40__FF_INPUT), .Q(u2_remLo_40_) );
  DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf114), .D(u2_remLo_41__FF_INPUT), .Q(u2_remLo_41_) );
  DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf113), .D(u2_remLo_42__FF_INPUT), .Q(u2_remLo_42_) );
  DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf112), .D(u2_remLo_43__FF_INPUT), .Q(u2_remLo_43_) );
  DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf111), .D(u2_remLo_44__FF_INPUT), .Q(u2_remLo_44_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf117), .D(u2_root_1__FF_INPUT), .Q(sqrto_0_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf72), .D(u2_root_46__FF_INPUT), .Q(sqrto_45_) );
  DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf110), .D(u2_remLo_45__FF_INPUT), .Q(u2_remLo_45_) );
  DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf109), .D(u2_remLo_46__FF_INPUT), .Q(u2_remLo_46_) );
  DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf108), .D(u2_remLo_47__FF_INPUT), .Q(u2_remLo_47_) );
  DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf107), .D(u2_remLo_48__FF_INPUT), .Q(u2_remLo_48_) );
  DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf106), .D(u2_remLo_49__FF_INPUT), .Q(u2_remLo_49_) );
  DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf105), .D(u2_remLo_50__FF_INPUT), .Q(u2_remLo_50_) );
  DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf104), .D(u2_remLo_51__FF_INPUT), .Q(u2_remLo_51_) );
  DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf103), .D(u2_remLo_52__FF_INPUT), .Q(u2_remLo_52_) );
  DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf102), .D(u2_remLo_53__FF_INPUT), .Q(u2_remLo_53_) );
  DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf101), .D(u2_remLo_54__FF_INPUT), .Q(u2_remLo_54_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf71), .D(u2_root_47__FF_INPUT), .Q(sqrto_46_) );
  DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf100), .D(u2_remLo_55__FF_INPUT), .Q(u2_remLo_55_) );
  DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf99), .D(u2_remLo_56__FF_INPUT), .Q(u2_remLo_56_) );
  DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf98), .D(u2_remLo_57__FF_INPUT), .Q(u2_remLo_57_) );
  DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf97), .D(u2_remLo_58__FF_INPUT), .Q(u2_remLo_58_) );
  DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf96), .D(u2_remLo_59__FF_INPUT), .Q(u2_remLo_59_) );
  DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf95), .D(u2_remLo_60__FF_INPUT), .Q(u2_remLo_60_) );
  DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf94), .D(u2_remLo_61__FF_INPUT), .Q(u2_remLo_61_) );
  DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf93), .D(u2_remLo_62__FF_INPUT), .Q(u2_remLo_62_) );
  DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf92), .D(u2_remLo_63__FF_INPUT), .Q(u2_remLo_63_) );
  DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf91), .D(u2_remLo_64__FF_INPUT), .Q(u2_remLo_64_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf70), .D(u2_root_48__FF_INPUT), .Q(sqrto_47_) );
  DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf90), .D(u2_remLo_65__FF_INPUT), .Q(u2_remLo_65_) );
  DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf89), .D(u2_remLo_66__FF_INPUT), .Q(u2_remLo_66_) );
  DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf88), .D(u2_remLo_67__FF_INPUT), .Q(u2_remLo_67_) );
  DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf87), .D(u2_remLo_68__FF_INPUT), .Q(u2_remLo_68_) );
  DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf86), .D(u2_remLo_69__FF_INPUT), .Q(u2_remLo_69_) );
  DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf85), .D(u2_remLo_70__FF_INPUT), .Q(u2_remLo_70_) );
  DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf84), .D(u2_remLo_71__FF_INPUT), .Q(u2_remLo_71_) );
  DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf83), .D(u2_remLo_72__FF_INPUT), .Q(u2_remLo_72_) );
  DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf82), .D(u2_remLo_73__FF_INPUT), .Q(u2_remLo_73_) );
  DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf81), .D(u2_remLo_74__FF_INPUT), .Q(u2_remLo_74_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf69), .D(u2_root_49__FF_INPUT), .Q(sqrto_48_) );
  DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf80), .D(u2_remLo_75__FF_INPUT), .Q(u2_remLo_75_) );
  DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf79), .D(u2_remLo_76__FF_INPUT), .Q(u2_remLo_76_) );
  DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf78), .D(u2_remLo_77__FF_INPUT), .Q(u2_remLo_77_) );
  DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf77), .D(u2_remLo_78__FF_INPUT), .Q(u2_remLo_78_) );
  DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf76), .D(u2_remLo_79__FF_INPUT), .Q(u2_remLo_79_) );
  DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf75), .D(u2_remLo_80__FF_INPUT), .Q(u2_remLo_80_) );
  DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf74), .D(u2_remLo_81__FF_INPUT), .Q(u2_remLo_81_) );
  DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf73), .D(u2_remLo_82__FF_INPUT), .Q(u2_remLo_82_) );
  DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf72), .D(u2_remLo_83__FF_INPUT), .Q(u2_remLo_83_) );
  DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf71), .D(u2_remLo_84__FF_INPUT), .Q(u2_remLo_84_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf68), .D(u2_root_50__FF_INPUT), .Q(sqrto_49_) );
  DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf70), .D(u2_remLo_85__FF_INPUT), .Q(u2_remLo_85_) );
  DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf69), .D(u2_remLo_86__FF_INPUT), .Q(u2_remLo_86_) );
  DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf68), .D(u2_remLo_87__FF_INPUT), .Q(u2_remLo_87_) );
  DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf67), .D(u2_remLo_88__FF_INPUT), .Q(u2_remLo_88_) );
  DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf66), .D(u2_remLo_89__FF_INPUT), .Q(u2_remLo_89_) );
  DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf65), .D(u2_remLo_90__FF_INPUT), .Q(u2_remLo_90_) );
  DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf64), .D(u2_remLo_91__FF_INPUT), .Q(u2_remLo_91_) );
  DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf63), .D(u2_remLo_92__FF_INPUT), .Q(u2_remLo_92_) );
  DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf62), .D(u2_remLo_93__FF_INPUT), .Q(u2_remLo_93_) );
  DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf61), .D(u2_remLo_94__FF_INPUT), .Q(u2_remLo_94_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf67), .D(u2_root_51__FF_INPUT), .Q(sqrto_50_) );
  DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf60), .D(u2_remLo_95__FF_INPUT), .Q(u2_remLo_95_) );
  DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf59), .D(u2_remLo_96__FF_INPUT), .Q(u2_remLo_96_) );
  DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf58), .D(u2_remLo_97__FF_INPUT), .Q(u2_remLo_97_) );
  DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf57), .D(u2_remLo_98__FF_INPUT), .Q(u2_remLo_98_) );
  DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf56), .D(u2_remLo_99__FF_INPUT), .Q(u2_remLo_99_) );
  DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf55), .D(u2_remLo_100__FF_INPUT), .Q(u2_remLo_100_) );
  DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf54), .D(u2_remLo_101__FF_INPUT), .Q(u2_remLo_101_) );
  DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf53), .D(u2_remLo_102__FF_INPUT), .Q(u2_remLo_102_) );
  DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf52), .D(u2_remLo_103__FF_INPUT), .Q(u2_remLo_103_) );
  DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf51), .D(u2_remLo_104__FF_INPUT), .Q(u2_remLo_104_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf66), .D(u2_root_52__FF_INPUT), .Q(sqrto_51_) );
  DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf50), .D(u2_remLo_105__FF_INPUT), .Q(u2_remLo_105_) );
  DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf49), .D(u2_remLo_106__FF_INPUT), .Q(u2_remLo_106_) );
  DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf48), .D(u2_remLo_107__FF_INPUT), .Q(u2_remLo_107_) );
  DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf47), .D(u2_remLo_108__FF_INPUT), .Q(u2_remLo_108_) );
  DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf46), .D(u2_remLo_109__FF_INPUT), .Q(u2_remLo_109_) );
  DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf45), .D(u2_remLo_110__FF_INPUT), .Q(u2_remLo_110_) );
  DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf44), .D(u2_remLo_111__FF_INPUT), .Q(u2_remLo_111_) );
  DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf43), .D(u2_remLo_112__FF_INPUT), .Q(u2_remLo_112_) );
  DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf42), .D(u2_remLo_113__FF_INPUT), .Q(u2_remLo_113_) );
  DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf41), .D(u2_remLo_114__FF_INPUT), .Q(u2_remLo_114_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf65), .D(u2_root_53__FF_INPUT), .Q(sqrto_52_) );
  DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf40), .D(u2_remLo_115__FF_INPUT), .Q(u2_remLo_115_) );
  DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf39), .D(u2_remLo_116__FF_INPUT), .Q(u2_remLo_116_) );
  DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf38), .D(u2_remLo_117__FF_INPUT), .Q(u2_remLo_117_) );
  DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf37), .D(u2_remLo_118__FF_INPUT), .Q(u2_remLo_118_) );
  DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf36), .D(u2_remLo_119__FF_INPUT), .Q(u2_remLo_119_) );
  DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf35), .D(u2_remLo_120__FF_INPUT), .Q(u2_remLo_120_) );
  DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf34), .D(u2_remLo_121__FF_INPUT), .Q(u2_remLo_121_) );
  DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf33), .D(u2_remLo_122__FF_INPUT), .Q(u2_remLo_122_) );
  DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf32), .D(u2_remLo_123__FF_INPUT), .Q(u2_remLo_123_) );
  DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf31), .D(u2_remLo_124__FF_INPUT), .Q(u2_remLo_124_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf64), .D(u2_root_54__FF_INPUT), .Q(sqrto_53_) );
  DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf30), .D(u2_remLo_125__FF_INPUT), .Q(u2_remLo_125_) );
  DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf29), .D(u2_remLo_126__FF_INPUT), .Q(u2_remLo_126_) );
  DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf28), .D(u2_remLo_127__FF_INPUT), .Q(u2_remLo_127_) );
  DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf27), .D(u2_remLo_128__FF_INPUT), .Q(u2_remLo_128_) );
  DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf26), .D(u2_remLo_129__FF_INPUT), .Q(u2_remLo_129_) );
  DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf25), .D(u2_remLo_130__FF_INPUT), .Q(u2_remLo_130_) );
  DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf24), .D(u2_remLo_131__FF_INPUT), .Q(u2_remLo_131_) );
  DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf23), .D(u2_remLo_132__FF_INPUT), .Q(u2_remLo_132_) );
  DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf22), .D(u2_remLo_133__FF_INPUT), .Q(u2_remLo_133_) );
  DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf21), .D(u2_remLo_134__FF_INPUT), .Q(u2_remLo_134_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf63), .D(u2_root_55__FF_INPUT), .Q(sqrto_54_) );
  DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf20), .D(u2_remLo_135__FF_INPUT), .Q(u2_remLo_135_) );
  DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf19), .D(u2_remLo_136__FF_INPUT), .Q(u2_remLo_136_) );
  DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf18), .D(u2_remLo_137__FF_INPUT), .Q(u2_remLo_137_) );
  DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf17), .D(u2_remLo_138__FF_INPUT), .Q(u2_remLo_138_) );
  DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf16), .D(u2_remLo_139__FF_INPUT), .Q(u2_remLo_139_) );
  DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf15), .D(u2_remLo_140__FF_INPUT), .Q(u2_remLo_140_) );
  DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf14), .D(u2_remLo_141__FF_INPUT), .Q(u2_remLo_141_) );
  DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf13), .D(u2_remLo_142__FF_INPUT), .Q(u2_remLo_142_) );
  DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf12), .D(u2_remLo_143__FF_INPUT), .Q(u2_remLo_143_) );
  DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf11), .D(u2_remLo_144__FF_INPUT), .Q(u2_remLo_144_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf116), .D(u2_root_2__FF_INPUT), .Q(sqrto_1_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf62), .D(u2_root_56__FF_INPUT), .Q(sqrto_55_) );
  DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf10), .D(u2_remLo_145__FF_INPUT), .Q(u2_remLo_145_) );
  DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf9), .D(u2_remLo_146__FF_INPUT), .Q(u2_remLo_146_) );
  DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf8), .D(u2_remLo_147__FF_INPUT), .Q(u2_remLo_147_) );
  DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf7), .D(u2_remLo_148__FF_INPUT), .Q(u2_remLo_148_) );
  DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf6), .D(u2_remLo_149__FF_INPUT), .Q(u2_remLo_149_) );
  DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf5), .D(u2_remLo_150__FF_INPUT), .Q(u2_remLo_150_) );
  DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf4), .D(u2_remLo_151__FF_INPUT), .Q(u2_remLo_151_) );
  DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf3), .D(u2_remLo_152__FF_INPUT), .Q(u2_remLo_152_) );
  DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf2), .D(u2_remLo_153__FF_INPUT), .Q(u2_remLo_153_) );
  DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf1), .D(u2_remLo_154__FF_INPUT), .Q(u2_remLo_154_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf61), .D(u2_root_57__FF_INPUT), .Q(sqrto_56_) );
  DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf0), .D(u2_remLo_155__FF_INPUT), .Q(u2_remLo_155_) );
  DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf121), .D(u2_remLo_156__FF_INPUT), .Q(u2_remLo_156_) );
  DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf120), .D(u2_remLo_157__FF_INPUT), .Q(u2_remLo_157_) );
  DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf119), .D(u2_remLo_158__FF_INPUT), .Q(u2_remLo_158_) );
  DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf118), .D(u2_remLo_159__FF_INPUT), .Q(u2_remLo_159_) );
  DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf117), .D(u2_remLo_160__FF_INPUT), .Q(u2_remLo_160_) );
  DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf116), .D(u2_remLo_161__FF_INPUT), .Q(u2_remLo_161_) );
  DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf115), .D(u2_remLo_162__FF_INPUT), .Q(u2_remLo_162_) );
  DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf114), .D(u2_remLo_163__FF_INPUT), .Q(u2_remLo_163_) );
  DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf113), .D(u2_remLo_164__FF_INPUT), .Q(u2_remLo_164_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf60), .D(u2_root_58__FF_INPUT), .Q(sqrto_57_) );
  DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf112), .D(u2_remLo_165__FF_INPUT), .Q(u2_remLo_165_) );
  DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf111), .D(u2_remLo_166__FF_INPUT), .Q(u2_remLo_166_) );
  DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf110), .D(u2_remLo_167__FF_INPUT), .Q(u2_remLo_167_) );
  DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf109), .D(u2_remLo_168__FF_INPUT), .Q(u2_remLo_168_) );
  DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf108), .D(u2_remLo_169__FF_INPUT), .Q(u2_remLo_169_) );
  DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf107), .D(u2_remLo_170__FF_INPUT), .Q(u2_remLo_170_) );
  DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf106), .D(u2_remLo_171__FF_INPUT), .Q(u2_remLo_171_) );
  DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf105), .D(u2_remLo_172__FF_INPUT), .Q(u2_remLo_172_) );
  DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf104), .D(u2_remLo_173__FF_INPUT), .Q(u2_remLo_173_) );
  DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf103), .D(u2_remLo_174__FF_INPUT), .Q(u2_remLo_174_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf59), .D(u2_root_59__FF_INPUT), .Q(sqrto_58_) );
  DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf102), .D(u2_remLo_175__FF_INPUT), .Q(u2_remLo_175_) );
  DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf101), .D(u2_remLo_176__FF_INPUT), .Q(u2_remLo_176_) );
  DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf100), .D(u2_remLo_177__FF_INPUT), .Q(u2_remLo_177_) );
  DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf99), .D(u2_remLo_178__FF_INPUT), .Q(u2_remLo_178_) );
  DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf98), .D(u2_remLo_179__FF_INPUT), .Q(u2_remLo_179_) );
  DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf97), .D(u2_remLo_180__FF_INPUT), .Q(u2_remLo_180_) );
  DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf96), .D(u2_remLo_181__FF_INPUT), .Q(u2_remLo_181_) );
  DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf95), .D(u2_remLo_182__FF_INPUT), .Q(u2_remLo_182_) );
  DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf94), .D(u2_remLo_183__FF_INPUT), .Q(u2_remLo_183_) );
  DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf93), .D(u2_remLo_184__FF_INPUT), .Q(u2_remLo_184_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf58), .D(u2_root_60__FF_INPUT), .Q(sqrto_59_) );
  DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf92), .D(u2_remLo_185__FF_INPUT), .Q(u2_remLo_185_) );
  DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf91), .D(u2_remLo_186__FF_INPUT), .Q(u2_remLo_186_) );
  DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf90), .D(u2_remLo_187__FF_INPUT), .Q(u2_remLo_187_) );
  DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf89), .D(u2_remLo_188__FF_INPUT), .Q(u2_remLo_188_) );
  DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf88), .D(u2_remLo_189__FF_INPUT), .Q(u2_remLo_189_) );
  DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf87), .D(u2_remLo_190__FF_INPUT), .Q(u2_remLo_190_) );
  DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf86), .D(u2_remLo_191__FF_INPUT), .Q(u2_remLo_191_) );
  DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf85), .D(u2_remLo_192__FF_INPUT), .Q(u2_remLo_192_) );
  DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf84), .D(u2_remLo_193__FF_INPUT), .Q(u2_remLo_193_) );
  DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf83), .D(u2_remLo_194__FF_INPUT), .Q(u2_remLo_194_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf57), .D(u2_root_61__FF_INPUT), .Q(sqrto_60_) );
  DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf82), .D(u2_remLo_195__FF_INPUT), .Q(u2_remLo_195_) );
  DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf81), .D(u2_remLo_196__FF_INPUT), .Q(u2_remLo_196_) );
  DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf80), .D(u2_remLo_197__FF_INPUT), .Q(u2_remLo_197_) );
  DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf79), .D(u2_remLo_198__FF_INPUT), .Q(u2_remLo_198_) );
  DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf78), .D(u2_remLo_199__FF_INPUT), .Q(u2_remLo_199_) );
  DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf77), .D(u2_remLo_200__FF_INPUT), .Q(u2_remLo_200_) );
  DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf76), .D(u2_remLo_201__FF_INPUT), .Q(u2_remLo_201_) );
  DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf75), .D(u2_remLo_202__FF_INPUT), .Q(u2_remLo_202_) );
  DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf74), .D(u2_remLo_203__FF_INPUT), .Q(u2_remLo_203_) );
  DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf73), .D(u2_remLo_204__FF_INPUT), .Q(u2_remLo_204_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf56), .D(u2_root_62__FF_INPUT), .Q(sqrto_61_) );
  DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf72), .D(u2_remLo_205__FF_INPUT), .Q(u2_remLo_205_) );
  DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf71), .D(u2_remLo_206__FF_INPUT), .Q(u2_remLo_206_) );
  DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf70), .D(u2_remLo_207__FF_INPUT), .Q(u2_remLo_207_) );
  DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf69), .D(u2_remLo_208__FF_INPUT), .Q(u2_remLo_208_) );
  DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf68), .D(u2_remLo_209__FF_INPUT), .Q(u2_remLo_209_) );
  DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf67), .D(u2_remLo_210__FF_INPUT), .Q(u2_remLo_210_) );
  DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf66), .D(u2_remLo_211__FF_INPUT), .Q(u2_remLo_211_) );
  DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf65), .D(u2_remLo_212__FF_INPUT), .Q(u2_remLo_212_) );
  DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf64), .D(u2_remLo_213__FF_INPUT), .Q(u2_remLo_213_) );
  DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf63), .D(u2_remLo_214__FF_INPUT), .Q(u2_remLo_214_) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf55), .D(u2_root_63__FF_INPUT), .Q(sqrto_62_) );
  DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf62), .D(u2_remLo_215__FF_INPUT), .Q(u2_remLo_215_) );
  DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf61), .D(u2_remLo_216__FF_INPUT), .Q(u2_remLo_216_) );
  DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf60), .D(u2_remLo_217__FF_INPUT), .Q(u2_remLo_217_) );
  DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf59), .D(u2_remLo_218__FF_INPUT), .Q(u2_remLo_218_) );
  DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf58), .D(u2_remLo_219__FF_INPUT), .Q(u2_remLo_219_) );
  DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf57), .D(u2_remLo_220__FF_INPUT), .Q(u2_remLo_220_) );
  DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf56), .D(u2_remLo_221__FF_INPUT), .Q(u2_remLo_221_) );
  DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf55), .D(u2_remLo_222__FF_INPUT), .Q(u2_remLo_222_) );
  DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf54), .D(u2_remLo_223__FF_INPUT), .Q(u2_remLo_223_) );
  DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf53), .D(u2_remLo_224__FF_INPUT), .Q(u2_remLo_224_) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf54), .D(u2_root_64__FF_INPUT), .Q(sqrto_63_) );
  DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf52), .D(u2_remLo_225__FF_INPUT), .Q(u2_remLo_225_) );
  DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_bF_buf51), .D(u2_remLo_226__FF_INPUT), .Q(u2_remLo_226_) );
  DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_bF_buf50), .D(u2_remLo_227__FF_INPUT), .Q(u2_remLo_227_) );
  DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_bF_buf49), .D(u2_remLo_228__FF_INPUT), .Q(u2_remLo_228_) );
  DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_bF_buf48), .D(u2_remLo_229__FF_INPUT), .Q(u2_remLo_229_) );
  DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_bF_buf47), .D(u2_remLo_230__FF_INPUT), .Q(u2_remLo_230_) );
  DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_bF_buf46), .D(u2_remLo_231__FF_INPUT), .Q(u2_remLo_231_) );
  DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_bF_buf45), .D(u2_remLo_232__FF_INPUT), .Q(u2_remLo_232_) );
  DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_bF_buf44), .D(u2_remLo_233__FF_INPUT), .Q(u2_remLo_233_) );
  DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_bF_buf43), .D(u2_remLo_234__FF_INPUT), .Q(u2_remLo_234_) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf53), .D(u2_root_65__FF_INPUT), .Q(sqrto_64_) );
  DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_bF_buf42), .D(u2_remLo_235__FF_INPUT), .Q(u2_remLo_235_) );
  DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_bF_buf41), .D(u2_remLo_236__FF_INPUT), .Q(u2_remLo_236_) );
  DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_bF_buf40), .D(u2_remLo_237__FF_INPUT), .Q(u2_remLo_237_) );
  DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_bF_buf39), .D(u2_remLo_238__FF_INPUT), .Q(u2_remLo_238_) );
  DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_bF_buf38), .D(u2_remLo_239__FF_INPUT), .Q(u2_remLo_239_) );
  DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_bF_buf37), .D(u2_remLo_240__FF_INPUT), .Q(u2_remLo_240_) );
  DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_bF_buf36), .D(u2_remLo_241__FF_INPUT), .Q(u2_remLo_241_) );
  DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_bF_buf35), .D(u2_remLo_242__FF_INPUT), .Q(u2_remLo_242_) );
  DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_bF_buf34), .D(u2_remLo_243__FF_INPUT), .Q(u2_remLo_243_) );
  DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_bF_buf33), .D(u2_remLo_244__FF_INPUT), .Q(u2_remLo_244_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf115), .D(u2_root_3__FF_INPUT), .Q(sqrto_2_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf52), .D(u2_root_66__FF_INPUT), .Q(sqrto_65_) );
  DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_bF_buf32), .D(u2_remLo_245__FF_INPUT), .Q(u2_remLo_245_) );
  DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_bF_buf31), .D(u2_remLo_246__FF_INPUT), .Q(u2_remLo_246_) );
  DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_bF_buf30), .D(u2_remLo_247__FF_INPUT), .Q(u2_remLo_247_) );
  DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_bF_buf29), .D(u2_remLo_248__FF_INPUT), .Q(u2_remLo_248_) );
  DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_bF_buf28), .D(u2_remLo_249__FF_INPUT), .Q(u2_remLo_249_) );
  DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_bF_buf27), .D(u2_remLo_250__FF_INPUT), .Q(u2_remLo_250_) );
  DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_bF_buf26), .D(u2_remLo_251__FF_INPUT), .Q(u2_remLo_251_) );
  DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_bF_buf25), .D(u2_remLo_252__FF_INPUT), .Q(u2_remLo_252_) );
  DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_bF_buf24), .D(u2_remLo_253__FF_INPUT), .Q(u2_remLo_253_) );
  DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_bF_buf23), .D(u2_remLo_254__FF_INPUT), .Q(u2_remLo_254_) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf51), .D(u2_root_67__FF_INPUT), .Q(sqrto_66_) );
  DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_bF_buf22), .D(u2_remLo_255__FF_INPUT), .Q(u2_remLo_255_) );
  DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_bF_buf21), .D(u2_remLo_256__FF_INPUT), .Q(u2_remLo_256_) );
  DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_bF_buf20), .D(u2_remLo_257__FF_INPUT), .Q(u2_remLo_257_) );
  DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_bF_buf19), .D(u2_remLo_258__FF_INPUT), .Q(u2_remLo_258_) );
  DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_bF_buf18), .D(u2_remLo_259__FF_INPUT), .Q(u2_remLo_259_) );
  DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_bF_buf17), .D(u2_remLo_260__FF_INPUT), .Q(u2_remLo_260_) );
  DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_bF_buf16), .D(u2_remLo_261__FF_INPUT), .Q(u2_remLo_261_) );
  DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_bF_buf15), .D(u2_remLo_262__FF_INPUT), .Q(u2_remLo_262_) );
  DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_bF_buf14), .D(u2_remLo_263__FF_INPUT), .Q(u2_remLo_263_) );
  DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_bF_buf13), .D(u2_remLo_264__FF_INPUT), .Q(u2_remLo_264_) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf50), .D(u2_root_68__FF_INPUT), .Q(sqrto_67_) );
  DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_bF_buf12), .D(u2_remLo_265__FF_INPUT), .Q(u2_remLo_265_) );
  DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_bF_buf11), .D(u2_remLo_266__FF_INPUT), .Q(u2_remLo_266_) );
  DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_bF_buf10), .D(u2_remLo_267__FF_INPUT), .Q(u2_remLo_267_) );
  DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_bF_buf9), .D(u2_remLo_268__FF_INPUT), .Q(u2_remLo_268_) );
  DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_bF_buf8), .D(u2_remLo_269__FF_INPUT), .Q(u2_remLo_269_) );
  DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_bF_buf7), .D(u2_remLo_270__FF_INPUT), .Q(u2_remLo_270_) );
  DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_bF_buf6), .D(u2_remLo_271__FF_INPUT), .Q(u2_remLo_271_) );
  DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_bF_buf5), .D(u2_remLo_272__FF_INPUT), .Q(u2_remLo_272_) );
  DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_bF_buf4), .D(u2_remLo_273__FF_INPUT), .Q(u2_remLo_273_) );
  DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_bF_buf3), .D(u2_remLo_274__FF_INPUT), .Q(u2_remLo_274_) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf49), .D(u2_root_69__FF_INPUT), .Q(sqrto_68_) );
  DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_bF_buf2), .D(u2_remLo_275__FF_INPUT), .Q(u2_remLo_275_) );
  DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_bF_buf1), .D(u2_remLo_276__FF_INPUT), .Q(u2_remLo_276_) );
  DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_bF_buf0), .D(u2_remLo_277__FF_INPUT), .Q(u2_remLo_277_) );
  DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_bF_buf121), .D(u2_remLo_278__FF_INPUT), .Q(u2_remLo_278_) );
  DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_bF_buf120), .D(u2_remLo_279__FF_INPUT), .Q(u2_remLo_279_) );
  DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_bF_buf119), .D(u2_remLo_280__FF_INPUT), .Q(u2_remLo_280_) );
  DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_bF_buf118), .D(u2_remLo_281__FF_INPUT), .Q(u2_remLo_281_) );
  DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_bF_buf117), .D(u2_remLo_282__FF_INPUT), .Q(u2_remLo_282_) );
  DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_bF_buf116), .D(u2_remLo_283__FF_INPUT), .Q(u2_remLo_283_) );
  DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_bF_buf115), .D(u2_remLo_284__FF_INPUT), .Q(u2_remLo_284_) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf48), .D(u2_root_70__FF_INPUT), .Q(sqrto_69_) );
  DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_bF_buf114), .D(u2_remLo_285__FF_INPUT), .Q(u2_remLo_285_) );
  DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_bF_buf113), .D(u2_remLo_286__FF_INPUT), .Q(u2_remLo_286_) );
  DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_bF_buf112), .D(u2_remLo_287__FF_INPUT), .Q(u2_remLo_287_) );
  DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_bF_buf111), .D(u2_remLo_288__FF_INPUT), .Q(u2_remLo_288_) );
  DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_bF_buf110), .D(u2_remLo_289__FF_INPUT), .Q(u2_remLo_289_) );
  DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_bF_buf109), .D(u2_remLo_290__FF_INPUT), .Q(u2_remLo_290_) );
  DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_bF_buf108), .D(u2_remLo_291__FF_INPUT), .Q(u2_remLo_291_) );
  DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_bF_buf107), .D(u2_remLo_292__FF_INPUT), .Q(u2_remLo_292_) );
  DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_bF_buf106), .D(u2_remLo_293__FF_INPUT), .Q(u2_remLo_293_) );
  DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_bF_buf105), .D(u2_remLo_294__FF_INPUT), .Q(u2_remLo_294_) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf47), .D(u2_root_71__FF_INPUT), .Q(sqrto_70_) );
  DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_bF_buf104), .D(u2_remLo_295__FF_INPUT), .Q(u2_remLo_295_) );
  DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_bF_buf103), .D(u2_remLo_296__FF_INPUT), .Q(u2_remLo_296_) );
  DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_bF_buf102), .D(u2_remLo_297__FF_INPUT), .Q(u2_remLo_297_) );
  DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_bF_buf101), .D(u2_remLo_298__FF_INPUT), .Q(u2_remLo_298_) );
  DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_bF_buf100), .D(u2_remLo_299__FF_INPUT), .Q(u2_remLo_299_) );
  DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_bF_buf99), .D(u2_remLo_300__FF_INPUT), .Q(u2_remLo_300_) );
  DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_bF_buf98), .D(u2_remLo_301__FF_INPUT), .Q(u2_remLo_301_) );
  DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_bF_buf97), .D(u2_remLo_302__FF_INPUT), .Q(u2_remLo_302_) );
  DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_bF_buf96), .D(u2_remLo_303__FF_INPUT), .Q(u2_remLo_303_) );
  DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_bF_buf95), .D(u2_remLo_304__FF_INPUT), .Q(u2_remLo_304_) );
  DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf46), .D(u2_root_72__FF_INPUT), .Q(sqrto_71_) );
  DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_bF_buf94), .D(u2_remLo_305__FF_INPUT), .Q(u2_remLo_305_) );
  DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_bF_buf93), .D(u2_remLo_306__FF_INPUT), .Q(u2_remLo_306_) );
  DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_bF_buf92), .D(u2_remLo_307__FF_INPUT), .Q(u2_remLo_307_) );
  DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_bF_buf91), .D(u2_remLo_308__FF_INPUT), .Q(u2_remLo_308_) );
  DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_bF_buf90), .D(u2_remLo_309__FF_INPUT), .Q(u2_remLo_309_) );
  DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_bF_buf89), .D(u2_remLo_310__FF_INPUT), .Q(u2_remLo_310_) );
  DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_bF_buf88), .D(u2_remLo_311__FF_INPUT), .Q(u2_remLo_311_) );
  DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_bF_buf87), .D(u2_remLo_312__FF_INPUT), .Q(u2_remLo_312_) );
  DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_bF_buf86), .D(u2_remLo_313__FF_INPUT), .Q(u2_remLo_313_) );
  DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_bF_buf85), .D(u2_remLo_314__FF_INPUT), .Q(u2_remLo_314_) );
  DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf45), .D(u2_root_73__FF_INPUT), .Q(sqrto_72_) );
  DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_bF_buf84), .D(u2_remLo_315__FF_INPUT), .Q(u2_remLo_315_) );
  DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_bF_buf83), .D(u2_remLo_316__FF_INPUT), .Q(u2_remLo_316_) );
  DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_bF_buf82), .D(u2_remLo_317__FF_INPUT), .Q(u2_remLo_317_) );
  DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_bF_buf81), .D(u2_remLo_318__FF_INPUT), .Q(u2_remLo_318_) );
  DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_bF_buf80), .D(u2_remLo_319__FF_INPUT), .Q(u2_remLo_319_) );
  DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_bF_buf79), .D(u2_remLo_320__FF_INPUT), .Q(u2_remLo_320_) );
  DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_bF_buf78), .D(u2_remLo_321__FF_INPUT), .Q(u2_remLo_321_) );
  DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_bF_buf77), .D(u2_remLo_322__FF_INPUT), .Q(u2_remLo_322_) );
  DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_bF_buf76), .D(u2_remLo_323__FF_INPUT), .Q(u2_remLo_323_) );
  DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_bF_buf75), .D(u2_remLo_324__FF_INPUT), .Q(u2_remLo_324_) );
  DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf44), .D(u2_root_74__FF_INPUT), .Q(sqrto_73_) );
  DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_bF_buf74), .D(u2_remLo_325__FF_INPUT), .Q(u2_remLo_325_) );
  DFFPOSX1 DFFPOSX1_781 ( .CLK(clk_bF_buf73), .D(u2_remLo_326__FF_INPUT), .Q(u2_remLo_326_) );
  DFFPOSX1 DFFPOSX1_782 ( .CLK(clk_bF_buf72), .D(u2_remLo_327__FF_INPUT), .Q(u2_remLo_327_) );
  DFFPOSX1 DFFPOSX1_783 ( .CLK(clk_bF_buf71), .D(u2_remLo_328__FF_INPUT), .Q(u2_remLo_328_) );
  DFFPOSX1 DFFPOSX1_784 ( .CLK(clk_bF_buf70), .D(u2_remLo_329__FF_INPUT), .Q(u2_remLo_329_) );
  DFFPOSX1 DFFPOSX1_785 ( .CLK(clk_bF_buf69), .D(u2_remLo_330__FF_INPUT), .Q(u2_remLo_330_) );
  DFFPOSX1 DFFPOSX1_786 ( .CLK(clk_bF_buf68), .D(u2_remLo_331__FF_INPUT), .Q(u2_remLo_331_) );
  DFFPOSX1 DFFPOSX1_787 ( .CLK(clk_bF_buf67), .D(u2_remLo_332__FF_INPUT), .Q(u2_remLo_332_) );
  DFFPOSX1 DFFPOSX1_788 ( .CLK(clk_bF_buf66), .D(u2_remLo_333__FF_INPUT), .Q(u2_remLo_333_) );
  DFFPOSX1 DFFPOSX1_789 ( .CLK(clk_bF_buf65), .D(u2_remLo_334__FF_INPUT), .Q(u2_remLo_334_) );
  DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf43), .D(u2_root_75__FF_INPUT), .Q(sqrto_74_) );
  DFFPOSX1 DFFPOSX1_790 ( .CLK(clk_bF_buf64), .D(u2_remLo_335__FF_INPUT), .Q(u2_remLo_335_) );
  DFFPOSX1 DFFPOSX1_791 ( .CLK(clk_bF_buf63), .D(u2_remLo_336__FF_INPUT), .Q(u2_remLo_336_) );
  DFFPOSX1 DFFPOSX1_792 ( .CLK(clk_bF_buf62), .D(u2_remLo_337__FF_INPUT), .Q(u2_remLo_337_) );
  DFFPOSX1 DFFPOSX1_793 ( .CLK(clk_bF_buf61), .D(u2_remLo_338__FF_INPUT), .Q(u2_remLo_338_) );
  DFFPOSX1 DFFPOSX1_794 ( .CLK(clk_bF_buf60), .D(u2_remLo_339__FF_INPUT), .Q(u2_remLo_339_) );
  DFFPOSX1 DFFPOSX1_795 ( .CLK(clk_bF_buf59), .D(u2_remLo_340__FF_INPUT), .Q(u2_remLo_340_) );
  DFFPOSX1 DFFPOSX1_796 ( .CLK(clk_bF_buf58), .D(u2_remLo_341__FF_INPUT), .Q(u2_remLo_341_) );
  DFFPOSX1 DFFPOSX1_797 ( .CLK(clk_bF_buf57), .D(u2_remLo_342__FF_INPUT), .Q(u2_remLo_342_) );
  DFFPOSX1 DFFPOSX1_798 ( .CLK(clk_bF_buf56), .D(u2_remLo_343__FF_INPUT), .Q(u2_remLo_343_) );
  DFFPOSX1 DFFPOSX1_799 ( .CLK(clk_bF_buf55), .D(u2_remLo_344__FF_INPUT), .Q(u2_remLo_344_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf114), .D(u2_root_4__FF_INPUT), .Q(sqrto_3_) );
  DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf42), .D(u2_root_76__FF_INPUT), .Q(sqrto_75_) );
  DFFPOSX1 DFFPOSX1_800 ( .CLK(clk_bF_buf54), .D(u2_remLo_345__FF_INPUT), .Q(u2_remLo_345_) );
  DFFPOSX1 DFFPOSX1_801 ( .CLK(clk_bF_buf53), .D(u2_remLo_346__FF_INPUT), .Q(u2_remLo_346_) );
  DFFPOSX1 DFFPOSX1_802 ( .CLK(clk_bF_buf52), .D(u2_remLo_347__FF_INPUT), .Q(u2_remLo_347_) );
  DFFPOSX1 DFFPOSX1_803 ( .CLK(clk_bF_buf51), .D(u2_remLo_348__FF_INPUT), .Q(u2_remLo_348_) );
  DFFPOSX1 DFFPOSX1_804 ( .CLK(clk_bF_buf50), .D(u2_remLo_349__FF_INPUT), .Q(u2_remLo_349_) );
  DFFPOSX1 DFFPOSX1_805 ( .CLK(clk_bF_buf49), .D(u2_remLo_350__FF_INPUT), .Q(u2_remLo_350_) );
  DFFPOSX1 DFFPOSX1_806 ( .CLK(clk_bF_buf48), .D(u2_remLo_351__FF_INPUT), .Q(u2_remLo_351_) );
  DFFPOSX1 DFFPOSX1_807 ( .CLK(clk_bF_buf47), .D(u2_remLo_352__FF_INPUT), .Q(u2_remLo_352_) );
  DFFPOSX1 DFFPOSX1_808 ( .CLK(clk_bF_buf46), .D(u2_remLo_353__FF_INPUT), .Q(u2_remLo_353_) );
  DFFPOSX1 DFFPOSX1_809 ( .CLK(clk_bF_buf45), .D(u2_remLo_354__FF_INPUT), .Q(u2_remLo_354_) );
  DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf41), .D(u2_root_77__FF_INPUT), .Q(sqrto_76_) );
  DFFPOSX1 DFFPOSX1_810 ( .CLK(clk_bF_buf44), .D(u2_remLo_355__FF_INPUT), .Q(u2_remLo_355_) );
  DFFPOSX1 DFFPOSX1_811 ( .CLK(clk_bF_buf43), .D(u2_remLo_356__FF_INPUT), .Q(u2_remLo_356_) );
  DFFPOSX1 DFFPOSX1_812 ( .CLK(clk_bF_buf42), .D(u2_remLo_357__FF_INPUT), .Q(u2_remLo_357_) );
  DFFPOSX1 DFFPOSX1_813 ( .CLK(clk_bF_buf41), .D(u2_remLo_358__FF_INPUT), .Q(u2_remLo_358_) );
  DFFPOSX1 DFFPOSX1_814 ( .CLK(clk_bF_buf40), .D(u2_remLo_359__FF_INPUT), .Q(u2_remLo_359_) );
  DFFPOSX1 DFFPOSX1_815 ( .CLK(clk_bF_buf39), .D(u2_remLo_360__FF_INPUT), .Q(u2_remLo_360_) );
  DFFPOSX1 DFFPOSX1_816 ( .CLK(clk_bF_buf38), .D(u2_remLo_361__FF_INPUT), .Q(u2_remLo_361_) );
  DFFPOSX1 DFFPOSX1_817 ( .CLK(clk_bF_buf37), .D(u2_remLo_362__FF_INPUT), .Q(u2_remLo_362_) );
  DFFPOSX1 DFFPOSX1_818 ( .CLK(clk_bF_buf36), .D(u2_remLo_363__FF_INPUT), .Q(u2_remLo_363_) );
  DFFPOSX1 DFFPOSX1_819 ( .CLK(clk_bF_buf35), .D(u2_remLo_364__FF_INPUT), .Q(u2_remLo_364_) );
  DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf40), .D(u2_root_78__FF_INPUT), .Q(sqrto_77_) );
  DFFPOSX1 DFFPOSX1_820 ( .CLK(clk_bF_buf34), .D(u2_remLo_365__FF_INPUT), .Q(u2_remLo_365_) );
  DFFPOSX1 DFFPOSX1_821 ( .CLK(clk_bF_buf33), .D(u2_remLo_366__FF_INPUT), .Q(u2_remLo_366_) );
  DFFPOSX1 DFFPOSX1_822 ( .CLK(clk_bF_buf32), .D(u2_remLo_367__FF_INPUT), .Q(u2_remLo_367_) );
  DFFPOSX1 DFFPOSX1_823 ( .CLK(clk_bF_buf31), .D(u2_remLo_368__FF_INPUT), .Q(u2_remLo_368_) );
  DFFPOSX1 DFFPOSX1_824 ( .CLK(clk_bF_buf30), .D(u2_remLo_369__FF_INPUT), .Q(u2_remLo_369_) );
  DFFPOSX1 DFFPOSX1_825 ( .CLK(clk_bF_buf29), .D(u2_remLo_370__FF_INPUT), .Q(u2_remLo_370_) );
  DFFPOSX1 DFFPOSX1_826 ( .CLK(clk_bF_buf28), .D(u2_remLo_371__FF_INPUT), .Q(u2_remLo_371_) );
  DFFPOSX1 DFFPOSX1_827 ( .CLK(clk_bF_buf27), .D(u2_remLo_372__FF_INPUT), .Q(u2_remLo_372_) );
  DFFPOSX1 DFFPOSX1_828 ( .CLK(clk_bF_buf26), .D(u2_remLo_373__FF_INPUT), .Q(u2_remLo_373_) );
  DFFPOSX1 DFFPOSX1_829 ( .CLK(clk_bF_buf25), .D(u2_remLo_374__FF_INPUT), .Q(u2_remLo_374_) );
  DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf39), .D(u2_root_79__FF_INPUT), .Q(sqrto_78_) );
  DFFPOSX1 DFFPOSX1_830 ( .CLK(clk_bF_buf24), .D(u2_remLo_375__FF_INPUT), .Q(u2_remLo_375_) );
  DFFPOSX1 DFFPOSX1_831 ( .CLK(clk_bF_buf23), .D(u2_remLo_376__FF_INPUT), .Q(u2_remLo_376_) );
  DFFPOSX1 DFFPOSX1_832 ( .CLK(clk_bF_buf22), .D(u2_remLo_377__FF_INPUT), .Q(u2_remLo_377_) );
  DFFPOSX1 DFFPOSX1_833 ( .CLK(clk_bF_buf21), .D(u2_remLo_378__FF_INPUT), .Q(u2_remLo_378_) );
  DFFPOSX1 DFFPOSX1_834 ( .CLK(clk_bF_buf20), .D(u2_remLo_379__FF_INPUT), .Q(u2_remLo_379_) );
  DFFPOSX1 DFFPOSX1_835 ( .CLK(clk_bF_buf19), .D(u2_remLo_380__FF_INPUT), .Q(u2_remLo_380_) );
  DFFPOSX1 DFFPOSX1_836 ( .CLK(clk_bF_buf18), .D(u2_remLo_381__FF_INPUT), .Q(u2_remLo_381_) );
  DFFPOSX1 DFFPOSX1_837 ( .CLK(clk_bF_buf17), .D(u2_remLo_382__FF_INPUT), .Q(u2_remLo_382_) );
  DFFPOSX1 DFFPOSX1_838 ( .CLK(clk_bF_buf16), .D(u2_remLo_383__FF_INPUT), .Q(u2_remLo_383_) );
  DFFPOSX1 DFFPOSX1_839 ( .CLK(clk_bF_buf15), .D(u2_remLo_384__FF_INPUT), .Q(u2_remLo_384_) );
  DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf38), .D(u2_root_80__FF_INPUT), .Q(sqrto_79_) );
  DFFPOSX1 DFFPOSX1_840 ( .CLK(clk_bF_buf14), .D(u2_remLo_385__FF_INPUT), .Q(u2_remLo_385_) );
  DFFPOSX1 DFFPOSX1_841 ( .CLK(clk_bF_buf13), .D(u2_remLo_386__FF_INPUT), .Q(u2_remLo_386_) );
  DFFPOSX1 DFFPOSX1_842 ( .CLK(clk_bF_buf12), .D(u2_remLo_387__FF_INPUT), .Q(u2_remLo_387_) );
  DFFPOSX1 DFFPOSX1_843 ( .CLK(clk_bF_buf11), .D(u2_remLo_388__FF_INPUT), .Q(u2_remLo_388_) );
  DFFPOSX1 DFFPOSX1_844 ( .CLK(clk_bF_buf10), .D(u2_remLo_389__FF_INPUT), .Q(u2_remLo_389_) );
  DFFPOSX1 DFFPOSX1_845 ( .CLK(clk_bF_buf9), .D(u2_remLo_390__FF_INPUT), .Q(u2_remLo_390_) );
  DFFPOSX1 DFFPOSX1_846 ( .CLK(clk_bF_buf8), .D(u2_remLo_391__FF_INPUT), .Q(u2_remLo_391_) );
  DFFPOSX1 DFFPOSX1_847 ( .CLK(clk_bF_buf7), .D(u2_remLo_392__FF_INPUT), .Q(u2_remLo_392_) );
  DFFPOSX1 DFFPOSX1_848 ( .CLK(clk_bF_buf6), .D(u2_remLo_393__FF_INPUT), .Q(u2_remLo_393_) );
  DFFPOSX1 DFFPOSX1_849 ( .CLK(clk_bF_buf5), .D(u2_remLo_394__FF_INPUT), .Q(u2_remLo_394_) );
  DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf37), .D(u2_root_81__FF_INPUT), .Q(sqrto_80_) );
  DFFPOSX1 DFFPOSX1_850 ( .CLK(clk_bF_buf4), .D(u2_remLo_395__FF_INPUT), .Q(u2_remLo_395_) );
  DFFPOSX1 DFFPOSX1_851 ( .CLK(clk_bF_buf3), .D(u2_remLo_396__FF_INPUT), .Q(u2_remLo_396_) );
  DFFPOSX1 DFFPOSX1_852 ( .CLK(clk_bF_buf2), .D(u2_remLo_397__FF_INPUT), .Q(u2_remLo_397_) );
  DFFPOSX1 DFFPOSX1_853 ( .CLK(clk_bF_buf1), .D(u2_remLo_398__FF_INPUT), .Q(u2_remLo_398_) );
  DFFPOSX1 DFFPOSX1_854 ( .CLK(clk_bF_buf0), .D(u2_remLo_399__FF_INPUT), .Q(u2_remLo_399_) );
  DFFPOSX1 DFFPOSX1_855 ( .CLK(clk_bF_buf121), .D(u2_remLo_400__FF_INPUT), .Q(u2_remLo_400_) );
  DFFPOSX1 DFFPOSX1_856 ( .CLK(clk_bF_buf120), .D(u2_remLo_401__FF_INPUT), .Q(u2_remLo_401_) );
  DFFPOSX1 DFFPOSX1_857 ( .CLK(clk_bF_buf119), .D(u2_remLo_402__FF_INPUT), .Q(u2_remLo_402_) );
  DFFPOSX1 DFFPOSX1_858 ( .CLK(clk_bF_buf118), .D(u2_remLo_403__FF_INPUT), .Q(u2_remLo_403_) );
  DFFPOSX1 DFFPOSX1_859 ( .CLK(clk_bF_buf117), .D(u2_remLo_404__FF_INPUT), .Q(u2_remLo_404_) );
  DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf36), .D(u2_root_82__FF_INPUT), .Q(sqrto_81_) );
  DFFPOSX1 DFFPOSX1_860 ( .CLK(clk_bF_buf116), .D(u2_remLo_405__FF_INPUT), .Q(u2_remLo_405_) );
  DFFPOSX1 DFFPOSX1_861 ( .CLK(clk_bF_buf115), .D(u2_remLo_406__FF_INPUT), .Q(u2_remLo_406_) );
  DFFPOSX1 DFFPOSX1_862 ( .CLK(clk_bF_buf114), .D(u2_remLo_407__FF_INPUT), .Q(u2_remLo_407_) );
  DFFPOSX1 DFFPOSX1_863 ( .CLK(clk_bF_buf113), .D(u2_remLo_408__FF_INPUT), .Q(u2_remLo_408_) );
  DFFPOSX1 DFFPOSX1_864 ( .CLK(clk_bF_buf112), .D(u2_remLo_409__FF_INPUT), .Q(u2_remLo_409_) );
  DFFPOSX1 DFFPOSX1_865 ( .CLK(clk_bF_buf111), .D(u2_remLo_410__FF_INPUT), .Q(u2_remLo_410_) );
  DFFPOSX1 DFFPOSX1_866 ( .CLK(clk_bF_buf110), .D(u2_remLo_411__FF_INPUT), .Q(u2_remLo_411_) );
  DFFPOSX1 DFFPOSX1_867 ( .CLK(clk_bF_buf109), .D(u2_remLo_412__FF_INPUT), .Q(u2_remLo_412_) );
  DFFPOSX1 DFFPOSX1_868 ( .CLK(clk_bF_buf108), .D(u2_remLo_413__FF_INPUT), .Q(u2_remLo_413_) );
  DFFPOSX1 DFFPOSX1_869 ( .CLK(clk_bF_buf107), .D(u2_remLo_414__FF_INPUT), .Q(u2_remLo_414_) );
  DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf35), .D(u2_root_83__FF_INPUT), .Q(sqrto_82_) );
  DFFPOSX1 DFFPOSX1_870 ( .CLK(clk_bF_buf106), .D(u2_remLo_415__FF_INPUT), .Q(u2_remLo_415_) );
  DFFPOSX1 DFFPOSX1_871 ( .CLK(clk_bF_buf105), .D(u2_remLo_416__FF_INPUT), .Q(u2_remLo_416_) );
  DFFPOSX1 DFFPOSX1_872 ( .CLK(clk_bF_buf104), .D(u2_remLo_417__FF_INPUT), .Q(u2_remLo_417_) );
  DFFPOSX1 DFFPOSX1_873 ( .CLK(clk_bF_buf103), .D(u2_remLo_418__FF_INPUT), .Q(u2_remLo_418_) );
  DFFPOSX1 DFFPOSX1_874 ( .CLK(clk_bF_buf102), .D(u2_remLo_419__FF_INPUT), .Q(u2_remLo_419_) );
  DFFPOSX1 DFFPOSX1_875 ( .CLK(clk_bF_buf101), .D(u2_remLo_420__FF_INPUT), .Q(u2_remLo_420_) );
  DFFPOSX1 DFFPOSX1_876 ( .CLK(clk_bF_buf100), .D(u2_remLo_421__FF_INPUT), .Q(u2_remLo_421_) );
  DFFPOSX1 DFFPOSX1_877 ( .CLK(clk_bF_buf99), .D(u2_remLo_422__FF_INPUT), .Q(u2_remLo_422_) );
  DFFPOSX1 DFFPOSX1_878 ( .CLK(clk_bF_buf98), .D(u2_remLo_423__FF_INPUT), .Q(u2_remLo_423_) );
  DFFPOSX1 DFFPOSX1_879 ( .CLK(clk_bF_buf97), .D(u2_remLo_424__FF_INPUT), .Q(u2_remLo_424_) );
  DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf34), .D(u2_root_84__FF_INPUT), .Q(sqrto_83_) );
  DFFPOSX1 DFFPOSX1_880 ( .CLK(clk_bF_buf96), .D(u2_remLo_425__FF_INPUT), .Q(u2_remLo_425_) );
  DFFPOSX1 DFFPOSX1_881 ( .CLK(clk_bF_buf95), .D(u2_remLo_426__FF_INPUT), .Q(u2_remLo_426_) );
  DFFPOSX1 DFFPOSX1_882 ( .CLK(clk_bF_buf94), .D(u2_remLo_427__FF_INPUT), .Q(u2_remLo_427_) );
  DFFPOSX1 DFFPOSX1_883 ( .CLK(clk_bF_buf93), .D(u2_remLo_428__FF_INPUT), .Q(u2_remLo_428_) );
  DFFPOSX1 DFFPOSX1_884 ( .CLK(clk_bF_buf92), .D(u2_remLo_429__FF_INPUT), .Q(u2_remLo_429_) );
  DFFPOSX1 DFFPOSX1_885 ( .CLK(clk_bF_buf91), .D(u2_remLo_430__FF_INPUT), .Q(u2_remLo_430_) );
  DFFPOSX1 DFFPOSX1_886 ( .CLK(clk_bF_buf90), .D(u2_remLo_431__FF_INPUT), .Q(u2_remLo_431_) );
  DFFPOSX1 DFFPOSX1_887 ( .CLK(clk_bF_buf89), .D(u2_remLo_432__FF_INPUT), .Q(u2_remLo_432_) );
  DFFPOSX1 DFFPOSX1_888 ( .CLK(clk_bF_buf88), .D(u2_remLo_433__FF_INPUT), .Q(u2_remLo_433_) );
  DFFPOSX1 DFFPOSX1_889 ( .CLK(clk_bF_buf87), .D(u2_remLo_434__FF_INPUT), .Q(u2_remLo_434_) );
  DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf33), .D(u2_root_85__FF_INPUT), .Q(sqrto_84_) );
  DFFPOSX1 DFFPOSX1_890 ( .CLK(clk_bF_buf86), .D(u2_remLo_435__FF_INPUT), .Q(u2_remLo_435_) );
  DFFPOSX1 DFFPOSX1_891 ( .CLK(clk_bF_buf85), .D(u2_remLo_436__FF_INPUT), .Q(u2_remLo_436_) );
  DFFPOSX1 DFFPOSX1_892 ( .CLK(clk_bF_buf84), .D(u2_remLo_437__FF_INPUT), .Q(u2_remLo_437_) );
  DFFPOSX1 DFFPOSX1_893 ( .CLK(clk_bF_buf83), .D(u2_remLo_438__FF_INPUT), .Q(u2_remLo_438_) );
  DFFPOSX1 DFFPOSX1_894 ( .CLK(clk_bF_buf82), .D(u2_remLo_439__FF_INPUT), .Q(u2_remLo_439_) );
  DFFPOSX1 DFFPOSX1_895 ( .CLK(clk_bF_buf81), .D(u2_remLo_440__FF_INPUT), .Q(u2_remLo_440_) );
  DFFPOSX1 DFFPOSX1_896 ( .CLK(clk_bF_buf80), .D(u2_remLo_441__FF_INPUT), .Q(u2_remLo_441_) );
  DFFPOSX1 DFFPOSX1_897 ( .CLK(clk_bF_buf79), .D(u2_remLo_442__FF_INPUT), .Q(u2_remLo_442_) );
  DFFPOSX1 DFFPOSX1_898 ( .CLK(clk_bF_buf78), .D(u2_remLo_443__FF_INPUT), .Q(u2_remLo_443_) );
  DFFPOSX1 DFFPOSX1_899 ( .CLK(clk_bF_buf77), .D(u2_remLo_444__FF_INPUT), .Q(u2_remLo_444_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf113), .D(u2_root_5__FF_INPUT), .Q(sqrto_4_) );
  DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf32), .D(u2_root_86__FF_INPUT), .Q(sqrto_85_) );
  DFFPOSX1 DFFPOSX1_900 ( .CLK(clk_bF_buf76), .D(u2_remLo_445__FF_INPUT), .Q(u2_remLo_445_) );
  DFFPOSX1 DFFPOSX1_901 ( .CLK(clk_bF_buf75), .D(u2_remLo_446__FF_INPUT), .Q(u2_remLo_446_) );
  DFFPOSX1 DFFPOSX1_902 ( .CLK(clk_bF_buf74), .D(u2_remLo_447__FF_INPUT), .Q(u2_remLo_447_) );
  DFFPOSX1 DFFPOSX1_903 ( .CLK(clk_bF_buf73), .D(u2_remLo_448__FF_INPUT), .Q(u2_remLo_448_) );
  DFFPOSX1 DFFPOSX1_904 ( .CLK(clk_bF_buf72), .D(u2_remLo_449__FF_INPUT), .Q(u2_remLo_449_) );
  DFFPOSX1 DFFPOSX1_905 ( .CLK(clk_bF_buf71), .D(u2_remLo_450__FF_INPUT), .Q(u2_remHiShift_0_) );
  DFFPOSX1 DFFPOSX1_906 ( .CLK(clk_bF_buf70), .D(u2_remLo_451__FF_INPUT), .Q(u2_remHiShift_1_) );
  DFFPOSX1 DFFPOSX1_907 ( .CLK(clk_bF_buf69), .D(u2_remHi_0__FF_INPUT), .Q(u2_remHi_0_) );
  DFFPOSX1 DFFPOSX1_908 ( .CLK(clk_bF_buf68), .D(u2_remHi_1__FF_INPUT), .Q(u2_remHi_1_) );
  DFFPOSX1 DFFPOSX1_909 ( .CLK(clk_bF_buf67), .D(u2_remHi_2__FF_INPUT), .Q(u2_remHi_2_) );
  DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf31), .D(u2_root_87__FF_INPUT), .Q(sqrto_86_) );
  DFFPOSX1 DFFPOSX1_910 ( .CLK(clk_bF_buf66), .D(u2_remHi_3__FF_INPUT), .Q(u2_remHi_3_) );
  DFFPOSX1 DFFPOSX1_911 ( .CLK(clk_bF_buf65), .D(u2_remHi_4__FF_INPUT), .Q(u2_remHi_4_) );
  DFFPOSX1 DFFPOSX1_912 ( .CLK(clk_bF_buf64), .D(u2_remHi_5__FF_INPUT), .Q(u2_remHi_5_) );
  DFFPOSX1 DFFPOSX1_913 ( .CLK(clk_bF_buf63), .D(u2_remHi_6__FF_INPUT), .Q(u2_remHi_6_) );
  DFFPOSX1 DFFPOSX1_914 ( .CLK(clk_bF_buf62), .D(u2_remHi_7__FF_INPUT), .Q(u2_remHi_7_) );
  DFFPOSX1 DFFPOSX1_915 ( .CLK(clk_bF_buf61), .D(u2_remHi_8__FF_INPUT), .Q(u2_remHi_8_) );
  DFFPOSX1 DFFPOSX1_916 ( .CLK(clk_bF_buf60), .D(u2_remHi_9__FF_INPUT), .Q(u2_remHi_9_) );
  DFFPOSX1 DFFPOSX1_917 ( .CLK(clk_bF_buf59), .D(u2_remHi_10__FF_INPUT), .Q(u2_remHi_10_) );
  DFFPOSX1 DFFPOSX1_918 ( .CLK(clk_bF_buf58), .D(u2_remHi_11__FF_INPUT), .Q(u2_remHi_11_) );
  DFFPOSX1 DFFPOSX1_919 ( .CLK(clk_bF_buf57), .D(u2_remHi_12__FF_INPUT), .Q(u2_remHi_12_) );
  DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf30), .D(u2_root_88__FF_INPUT), .Q(sqrto_87_) );
  DFFPOSX1 DFFPOSX1_920 ( .CLK(clk_bF_buf56), .D(u2_remHi_13__FF_INPUT), .Q(u2_remHi_13_) );
  DFFPOSX1 DFFPOSX1_921 ( .CLK(clk_bF_buf55), .D(u2_remHi_14__FF_INPUT), .Q(u2_remHi_14_) );
  DFFPOSX1 DFFPOSX1_922 ( .CLK(clk_bF_buf54), .D(u2_remHi_15__FF_INPUT), .Q(u2_remHi_15_) );
  DFFPOSX1 DFFPOSX1_923 ( .CLK(clk_bF_buf53), .D(u2_remHi_16__FF_INPUT), .Q(u2_remHi_16_) );
  DFFPOSX1 DFFPOSX1_924 ( .CLK(clk_bF_buf52), .D(u2_remHi_17__FF_INPUT), .Q(u2_remHi_17_) );
  DFFPOSX1 DFFPOSX1_925 ( .CLK(clk_bF_buf51), .D(u2_remHi_18__FF_INPUT), .Q(u2_remHi_18_) );
  DFFPOSX1 DFFPOSX1_926 ( .CLK(clk_bF_buf50), .D(u2_remHi_19__FF_INPUT), .Q(u2_remHi_19_) );
  DFFPOSX1 DFFPOSX1_927 ( .CLK(clk_bF_buf49), .D(u2_remHi_20__FF_INPUT), .Q(u2_remHi_20_) );
  DFFPOSX1 DFFPOSX1_928 ( .CLK(clk_bF_buf48), .D(u2_remHi_21__FF_INPUT), .Q(u2_remHi_21_) );
  DFFPOSX1 DFFPOSX1_929 ( .CLK(clk_bF_buf47), .D(u2_remHi_22__FF_INPUT), .Q(u2_remHi_22_) );
  DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf29), .D(u2_root_89__FF_INPUT), .Q(sqrto_88_) );
  DFFPOSX1 DFFPOSX1_930 ( .CLK(clk_bF_buf46), .D(u2_remHi_23__FF_INPUT), .Q(u2_remHi_23_) );
  DFFPOSX1 DFFPOSX1_931 ( .CLK(clk_bF_buf45), .D(u2_remHi_24__FF_INPUT), .Q(u2_remHi_24_) );
  DFFPOSX1 DFFPOSX1_932 ( .CLK(clk_bF_buf44), .D(u2_remHi_25__FF_INPUT), .Q(u2_remHi_25_) );
  DFFPOSX1 DFFPOSX1_933 ( .CLK(clk_bF_buf43), .D(u2_remHi_26__FF_INPUT), .Q(u2_remHi_26_) );
  DFFPOSX1 DFFPOSX1_934 ( .CLK(clk_bF_buf42), .D(u2_remHi_27__FF_INPUT), .Q(u2_remHi_27_) );
  DFFPOSX1 DFFPOSX1_935 ( .CLK(clk_bF_buf41), .D(u2_remHi_28__FF_INPUT), .Q(u2_remHi_28_) );
  DFFPOSX1 DFFPOSX1_936 ( .CLK(clk_bF_buf40), .D(u2_remHi_29__FF_INPUT), .Q(u2_remHi_29_) );
  DFFPOSX1 DFFPOSX1_937 ( .CLK(clk_bF_buf39), .D(u2_remHi_30__FF_INPUT), .Q(u2_remHi_30_) );
  DFFPOSX1 DFFPOSX1_938 ( .CLK(clk_bF_buf38), .D(u2_remHi_31__FF_INPUT), .Q(u2_remHi_31_) );
  DFFPOSX1 DFFPOSX1_939 ( .CLK(clk_bF_buf37), .D(u2_remHi_32__FF_INPUT), .Q(u2_remHi_32_) );
  DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf28), .D(u2_root_90__FF_INPUT), .Q(sqrto_89_) );
  DFFPOSX1 DFFPOSX1_940 ( .CLK(clk_bF_buf36), .D(u2_remHi_33__FF_INPUT), .Q(u2_remHi_33_) );
  DFFPOSX1 DFFPOSX1_941 ( .CLK(clk_bF_buf35), .D(u2_remHi_34__FF_INPUT), .Q(u2_remHi_34_) );
  DFFPOSX1 DFFPOSX1_942 ( .CLK(clk_bF_buf34), .D(u2_remHi_35__FF_INPUT), .Q(u2_remHi_35_) );
  DFFPOSX1 DFFPOSX1_943 ( .CLK(clk_bF_buf33), .D(u2_remHi_36__FF_INPUT), .Q(u2_remHi_36_) );
  DFFPOSX1 DFFPOSX1_944 ( .CLK(clk_bF_buf32), .D(u2_remHi_37__FF_INPUT), .Q(u2_remHi_37_) );
  DFFPOSX1 DFFPOSX1_945 ( .CLK(clk_bF_buf31), .D(u2_remHi_38__FF_INPUT), .Q(u2_remHi_38_) );
  DFFPOSX1 DFFPOSX1_946 ( .CLK(clk_bF_buf30), .D(u2_remHi_39__FF_INPUT), .Q(u2_remHi_39_) );
  DFFPOSX1 DFFPOSX1_947 ( .CLK(clk_bF_buf29), .D(u2_remHi_40__FF_INPUT), .Q(u2_remHi_40_) );
  DFFPOSX1 DFFPOSX1_948 ( .CLK(clk_bF_buf28), .D(u2_remHi_41__FF_INPUT), .Q(u2_remHi_41_) );
  DFFPOSX1 DFFPOSX1_949 ( .CLK(clk_bF_buf27), .D(u2_remHi_42__FF_INPUT), .Q(u2_remHi_42_) );
  DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf27), .D(u2_root_91__FF_INPUT), .Q(sqrto_90_) );
  DFFPOSX1 DFFPOSX1_950 ( .CLK(clk_bF_buf26), .D(u2_remHi_43__FF_INPUT), .Q(u2_remHi_43_) );
  DFFPOSX1 DFFPOSX1_951 ( .CLK(clk_bF_buf25), .D(u2_remHi_44__FF_INPUT), .Q(u2_remHi_44_) );
  DFFPOSX1 DFFPOSX1_952 ( .CLK(clk_bF_buf24), .D(u2_remHi_45__FF_INPUT), .Q(u2_remHi_45_) );
  DFFPOSX1 DFFPOSX1_953 ( .CLK(clk_bF_buf23), .D(u2_remHi_46__FF_INPUT), .Q(u2_remHi_46_) );
  DFFPOSX1 DFFPOSX1_954 ( .CLK(clk_bF_buf22), .D(u2_remHi_47__FF_INPUT), .Q(u2_remHi_47_) );
  DFFPOSX1 DFFPOSX1_955 ( .CLK(clk_bF_buf21), .D(u2_remHi_48__FF_INPUT), .Q(u2_remHi_48_) );
  DFFPOSX1 DFFPOSX1_956 ( .CLK(clk_bF_buf20), .D(u2_remHi_49__FF_INPUT), .Q(u2_remHi_49_) );
  DFFPOSX1 DFFPOSX1_957 ( .CLK(clk_bF_buf19), .D(u2_remHi_50__FF_INPUT), .Q(u2_remHi_50_) );
  DFFPOSX1 DFFPOSX1_958 ( .CLK(clk_bF_buf18), .D(u2_remHi_51__FF_INPUT), .Q(u2_remHi_51_) );
  DFFPOSX1 DFFPOSX1_959 ( .CLK(clk_bF_buf17), .D(u2_remHi_52__FF_INPUT), .Q(u2_remHi_52_) );
  DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf26), .D(u2_root_92__FF_INPUT), .Q(sqrto_91_) );
  DFFPOSX1 DFFPOSX1_960 ( .CLK(clk_bF_buf16), .D(u2_remHi_53__FF_INPUT), .Q(u2_remHi_53_) );
  DFFPOSX1 DFFPOSX1_961 ( .CLK(clk_bF_buf15), .D(u2_remHi_54__FF_INPUT), .Q(u2_remHi_54_) );
  DFFPOSX1 DFFPOSX1_962 ( .CLK(clk_bF_buf14), .D(u2_remHi_55__FF_INPUT), .Q(u2_remHi_55_) );
  DFFPOSX1 DFFPOSX1_963 ( .CLK(clk_bF_buf13), .D(u2_remHi_56__FF_INPUT), .Q(u2_remHi_56_) );
  DFFPOSX1 DFFPOSX1_964 ( .CLK(clk_bF_buf12), .D(u2_remHi_57__FF_INPUT), .Q(u2_remHi_57_) );
  DFFPOSX1 DFFPOSX1_965 ( .CLK(clk_bF_buf11), .D(u2_remHi_58__FF_INPUT), .Q(u2_remHi_58_) );
  DFFPOSX1 DFFPOSX1_966 ( .CLK(clk_bF_buf10), .D(u2_remHi_59__FF_INPUT), .Q(u2_remHi_59_) );
  DFFPOSX1 DFFPOSX1_967 ( .CLK(clk_bF_buf9), .D(u2_remHi_60__FF_INPUT), .Q(u2_remHi_60_) );
  DFFPOSX1 DFFPOSX1_968 ( .CLK(clk_bF_buf8), .D(u2_remHi_61__FF_INPUT), .Q(u2_remHi_61_) );
  DFFPOSX1 DFFPOSX1_969 ( .CLK(clk_bF_buf7), .D(u2_remHi_62__FF_INPUT), .Q(u2_remHi_62_) );
  DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf25), .D(u2_root_93__FF_INPUT), .Q(sqrto_92_) );
  DFFPOSX1 DFFPOSX1_970 ( .CLK(clk_bF_buf6), .D(u2_remHi_63__FF_INPUT), .Q(u2_remHi_63_) );
  DFFPOSX1 DFFPOSX1_971 ( .CLK(clk_bF_buf5), .D(u2_remHi_64__FF_INPUT), .Q(u2_remHi_64_) );
  DFFPOSX1 DFFPOSX1_972 ( .CLK(clk_bF_buf4), .D(u2_remHi_65__FF_INPUT), .Q(u2_remHi_65_) );
  DFFPOSX1 DFFPOSX1_973 ( .CLK(clk_bF_buf3), .D(u2_remHi_66__FF_INPUT), .Q(u2_remHi_66_) );
  DFFPOSX1 DFFPOSX1_974 ( .CLK(clk_bF_buf2), .D(u2_remHi_67__FF_INPUT), .Q(u2_remHi_67_) );
  DFFPOSX1 DFFPOSX1_975 ( .CLK(clk_bF_buf1), .D(u2_remHi_68__FF_INPUT), .Q(u2_remHi_68_) );
  DFFPOSX1 DFFPOSX1_976 ( .CLK(clk_bF_buf0), .D(u2_remHi_69__FF_INPUT), .Q(u2_remHi_69_) );
  DFFPOSX1 DFFPOSX1_977 ( .CLK(clk_bF_buf121), .D(u2_remHi_70__FF_INPUT), .Q(u2_remHi_70_) );
  DFFPOSX1 DFFPOSX1_978 ( .CLK(clk_bF_buf120), .D(u2_remHi_71__FF_INPUT), .Q(u2_remHi_71_) );
  DFFPOSX1 DFFPOSX1_979 ( .CLK(clk_bF_buf119), .D(u2_remHi_72__FF_INPUT), .Q(u2_remHi_72_) );
  DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf24), .D(u2_root_94__FF_INPUT), .Q(sqrto_93_) );
  DFFPOSX1 DFFPOSX1_980 ( .CLK(clk_bF_buf118), .D(u2_remHi_73__FF_INPUT), .Q(u2_remHi_73_) );
  DFFPOSX1 DFFPOSX1_981 ( .CLK(clk_bF_buf117), .D(u2_remHi_74__FF_INPUT), .Q(u2_remHi_74_) );
  DFFPOSX1 DFFPOSX1_982 ( .CLK(clk_bF_buf116), .D(u2_remHi_75__FF_INPUT), .Q(u2_remHi_75_) );
  DFFPOSX1 DFFPOSX1_983 ( .CLK(clk_bF_buf115), .D(u2_remHi_76__FF_INPUT), .Q(u2_remHi_76_) );
  DFFPOSX1 DFFPOSX1_984 ( .CLK(clk_bF_buf114), .D(u2_remHi_77__FF_INPUT), .Q(u2_remHi_77_) );
  DFFPOSX1 DFFPOSX1_985 ( .CLK(clk_bF_buf113), .D(u2_remHi_78__FF_INPUT), .Q(u2_remHi_78_) );
  DFFPOSX1 DFFPOSX1_986 ( .CLK(clk_bF_buf112), .D(u2_remHi_79__FF_INPUT), .Q(u2_remHi_79_) );
  DFFPOSX1 DFFPOSX1_987 ( .CLK(clk_bF_buf111), .D(u2_remHi_80__FF_INPUT), .Q(u2_remHi_80_) );
  DFFPOSX1 DFFPOSX1_988 ( .CLK(clk_bF_buf110), .D(u2_remHi_81__FF_INPUT), .Q(u2_remHi_81_) );
  DFFPOSX1 DFFPOSX1_989 ( .CLK(clk_bF_buf109), .D(u2_remHi_82__FF_INPUT), .Q(u2_remHi_82_) );
  DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf23), .D(u2_root_95__FF_INPUT), .Q(sqrto_94_) );
  DFFPOSX1 DFFPOSX1_990 ( .CLK(clk_bF_buf108), .D(u2_remHi_83__FF_INPUT), .Q(u2_remHi_83_) );
  DFFPOSX1 DFFPOSX1_991 ( .CLK(clk_bF_buf107), .D(u2_remHi_84__FF_INPUT), .Q(u2_remHi_84_) );
  DFFPOSX1 DFFPOSX1_992 ( .CLK(clk_bF_buf106), .D(u2_remHi_85__FF_INPUT), .Q(u2_remHi_85_) );
  DFFPOSX1 DFFPOSX1_993 ( .CLK(clk_bF_buf105), .D(u2_remHi_86__FF_INPUT), .Q(u2_remHi_86_) );
  DFFPOSX1 DFFPOSX1_994 ( .CLK(clk_bF_buf104), .D(u2_remHi_87__FF_INPUT), .Q(u2_remHi_87_) );
  DFFPOSX1 DFFPOSX1_995 ( .CLK(clk_bF_buf103), .D(u2_remHi_88__FF_INPUT), .Q(u2_remHi_88_) );
  DFFPOSX1 DFFPOSX1_996 ( .CLK(clk_bF_buf102), .D(u2_remHi_89__FF_INPUT), .Q(u2_remHi_89_) );
  DFFPOSX1 DFFPOSX1_997 ( .CLK(clk_bF_buf101), .D(u2_remHi_90__FF_INPUT), .Q(u2_remHi_90_) );
  DFFPOSX1 DFFPOSX1_998 ( .CLK(clk_bF_buf100), .D(u2_remHi_91__FF_INPUT), .Q(u2_remHi_91_) );
  DFFPOSX1 DFFPOSX1_999 ( .CLK(clk_bF_buf99), .D(u2_remHi_92__FF_INPUT), .Q(u2_remHi_92_) );
  INVX1 INVX1_1 ( .A(\a[113] ), .Y(_abc_64468_n1508) );
  INVX1 INVX1_10 ( .A(_abc_64468_n1531), .Y(_abc_64468_n1545) );
  INVX1 INVX1_100 ( .A(\a[14] ), .Y(u1__abc_43968_n261) );
  INVX1 INVX1_1000 ( .A(u2_remHi_159_), .Y(u2__abc_44228_n5010) );
  INVX1 INVX1_1001 ( .A(u2__abc_44228_n5011), .Y(u2__abc_44228_n5012) );
  INVX1 INVX1_1002 ( .A(sqrto_157_), .Y(u2__abc_44228_n5019) );
  INVX1 INVX1_1003 ( .A(u2__abc_44228_n5020), .Y(u2__abc_44228_n5021) );
  INVX1 INVX1_1004 ( .A(u2_remHi_157_), .Y(u2__abc_44228_n5022) );
  INVX1 INVX1_1005 ( .A(u2__abc_44228_n5023_1), .Y(u2__abc_44228_n5024) );
  INVX1 INVX1_1006 ( .A(sqrto_156_), .Y(u2__abc_44228_n5026) );
  INVX1 INVX1_1007 ( .A(u2_remHi_156_), .Y(u2__abc_44228_n5028) );
  INVX1 INVX1_1008 ( .A(u2__abc_44228_n5030), .Y(u2__abc_44228_n5031) );
  INVX1 INVX1_1009 ( .A(sqrto_155_), .Y(u2__abc_44228_n5033) );
  INVX1 INVX1_101 ( .A(\a[15] ), .Y(u1__abc_43968_n262) );
  INVX1 INVX1_1010 ( .A(u2__abc_44228_n5034), .Y(u2__abc_44228_n5035) );
  INVX1 INVX1_1011 ( .A(u2_remHi_155_), .Y(u2__abc_44228_n5036) );
  INVX1 INVX1_1012 ( .A(u2__abc_44228_n5037), .Y(u2__abc_44228_n5038) );
  INVX1 INVX1_1013 ( .A(sqrto_154_), .Y(u2__abc_44228_n5040) );
  INVX1 INVX1_1014 ( .A(u2_remHi_154_), .Y(u2__abc_44228_n5042_1) );
  INVX1 INVX1_1015 ( .A(u2__abc_44228_n5044), .Y(u2__abc_44228_n5045) );
  INVX1 INVX1_1016 ( .A(sqrto_153_), .Y(u2__abc_44228_n5048) );
  INVX1 INVX1_1017 ( .A(u2__abc_44228_n5049), .Y(u2__abc_44228_n5050) );
  INVX1 INVX1_1018 ( .A(u2_remHi_153_), .Y(u2__abc_44228_n5051_1) );
  INVX1 INVX1_1019 ( .A(u2__abc_44228_n5052), .Y(u2__abc_44228_n5053) );
  INVX1 INVX1_102 ( .A(\a[12] ), .Y(u1__abc_43968_n264) );
  INVX1 INVX1_1020 ( .A(sqrto_152_), .Y(u2__abc_44228_n5055) );
  INVX1 INVX1_1021 ( .A(u2_remHi_152_), .Y(u2__abc_44228_n5057) );
  INVX1 INVX1_1022 ( .A(u2__abc_44228_n5059), .Y(u2__abc_44228_n5060) );
  INVX1 INVX1_1023 ( .A(sqrto_150_), .Y(u2__abc_44228_n5062) );
  INVX1 INVX1_1024 ( .A(u2_remHi_150_), .Y(u2__abc_44228_n5064) );
  INVX1 INVX1_1025 ( .A(u2__abc_44228_n5066), .Y(u2__abc_44228_n5067) );
  INVX1 INVX1_1026 ( .A(sqrto_151_), .Y(u2__abc_44228_n5068) );
  INVX1 INVX1_1027 ( .A(u2__abc_44228_n5069), .Y(u2__abc_44228_n5070) );
  INVX1 INVX1_1028 ( .A(u2_remHi_151_), .Y(u2__abc_44228_n5071_1) );
  INVX1 INVX1_1029 ( .A(u2__abc_44228_n5072), .Y(u2__abc_44228_n5073) );
  INVX1 INVX1_103 ( .A(\a[13] ), .Y(u1__abc_43968_n265) );
  INVX1 INVX1_1030 ( .A(sqrto_149_), .Y(u2__abc_44228_n5078) );
  INVX1 INVX1_1031 ( .A(u2__abc_44228_n5079), .Y(u2__abc_44228_n5080_1) );
  INVX1 INVX1_1032 ( .A(u2_remHi_149_), .Y(u2__abc_44228_n5081) );
  INVX1 INVX1_1033 ( .A(u2__abc_44228_n5082), .Y(u2__abc_44228_n5083) );
  INVX1 INVX1_1034 ( .A(sqrto_148_), .Y(u2__abc_44228_n5085) );
  INVX1 INVX1_1035 ( .A(u2_remHi_148_), .Y(u2__abc_44228_n5087) );
  INVX1 INVX1_1036 ( .A(u2__abc_44228_n5089_1), .Y(u2__abc_44228_n5090) );
  INVX1 INVX1_1037 ( .A(sqrto_146_), .Y(u2__abc_44228_n5092) );
  INVX1 INVX1_1038 ( .A(u2_remHi_146_), .Y(u2__abc_44228_n5094) );
  INVX1 INVX1_1039 ( .A(u2__abc_44228_n5096), .Y(u2__abc_44228_n5097) );
  INVX1 INVX1_104 ( .A(\a[10] ), .Y(u1__abc_43968_n268_1) );
  INVX1 INVX1_1040 ( .A(sqrto_147_), .Y(u2__abc_44228_n5098) );
  INVX1 INVX1_1041 ( .A(u2__abc_44228_n5099_1), .Y(u2__abc_44228_n5100) );
  INVX1 INVX1_1042 ( .A(u2_remHi_147_), .Y(u2__abc_44228_n5101) );
  INVX1 INVX1_1043 ( .A(u2__abc_44228_n5102), .Y(u2__abc_44228_n5103) );
  INVX1 INVX1_1044 ( .A(sqrto_145_), .Y(u2__abc_44228_n5107) );
  INVX1 INVX1_1045 ( .A(u2__abc_44228_n5108), .Y(u2__abc_44228_n5109_1) );
  INVX1 INVX1_1046 ( .A(u2_remHi_145_), .Y(u2__abc_44228_n5110) );
  INVX1 INVX1_1047 ( .A(u2__abc_44228_n5111), .Y(u2__abc_44228_n5112) );
  INVX1 INVX1_1048 ( .A(sqrto_144_), .Y(u2__abc_44228_n5114) );
  INVX1 INVX1_1049 ( .A(u2_remHi_144_), .Y(u2__abc_44228_n5116) );
  INVX1 INVX1_105 ( .A(\a[11] ), .Y(u1__abc_43968_n269_1) );
  INVX1 INVX1_1050 ( .A(u2__abc_44228_n5118_1), .Y(u2__abc_44228_n5119) );
  INVX1 INVX1_1051 ( .A(sqrto_143_), .Y(u2__abc_44228_n5121) );
  INVX1 INVX1_1052 ( .A(u2__abc_44228_n5122), .Y(u2__abc_44228_n5123) );
  INVX1 INVX1_1053 ( .A(u2_remHi_143_), .Y(u2__abc_44228_n5124) );
  INVX1 INVX1_1054 ( .A(u2__abc_44228_n5125), .Y(u2__abc_44228_n5126) );
  INVX1 INVX1_1055 ( .A(sqrto_142_), .Y(u2__abc_44228_n5128) );
  INVX1 INVX1_1056 ( .A(u2_remHi_142_), .Y(u2__abc_44228_n5130) );
  INVX1 INVX1_1057 ( .A(u2__abc_44228_n5132), .Y(u2__abc_44228_n5133) );
  INVX1 INVX1_1058 ( .A(sqrto_141_), .Y(u2__abc_44228_n5138) );
  INVX1 INVX1_1059 ( .A(u2__abc_44228_n5139), .Y(u2__abc_44228_n5140) );
  INVX1 INVX1_106 ( .A(\a[8] ), .Y(u1__abc_43968_n271) );
  INVX1 INVX1_1060 ( .A(u2_remHi_141_), .Y(u2__abc_44228_n5141) );
  INVX1 INVX1_1061 ( .A(u2__abc_44228_n5142), .Y(u2__abc_44228_n5143) );
  INVX1 INVX1_1062 ( .A(sqrto_140_), .Y(u2__abc_44228_n5145) );
  INVX1 INVX1_1063 ( .A(u2_remHi_140_), .Y(u2__abc_44228_n5147) );
  INVX1 INVX1_1064 ( .A(u2__abc_44228_n5149), .Y(u2__abc_44228_n5150) );
  INVX1 INVX1_1065 ( .A(sqrto_139_), .Y(u2__abc_44228_n5152) );
  INVX1 INVX1_1066 ( .A(u2__abc_44228_n5153), .Y(u2__abc_44228_n5154) );
  INVX1 INVX1_1067 ( .A(u2_remHi_139_), .Y(u2__abc_44228_n5155_1) );
  INVX1 INVX1_1068 ( .A(u2__abc_44228_n5156), .Y(u2__abc_44228_n5157) );
  INVX1 INVX1_1069 ( .A(sqrto_138_), .Y(u2__abc_44228_n5159) );
  INVX1 INVX1_107 ( .A(\a[9] ), .Y(u1__abc_43968_n272_1) );
  INVX1 INVX1_1070 ( .A(u2_remHi_138_), .Y(u2__abc_44228_n5161) );
  INVX1 INVX1_1071 ( .A(u2__abc_44228_n5163), .Y(u2__abc_44228_n5164_1) );
  INVX1 INVX1_1072 ( .A(sqrto_135_), .Y(u2__abc_44228_n5167) );
  INVX1 INVX1_1073 ( .A(u2__abc_44228_n5168), .Y(u2__abc_44228_n5169) );
  INVX1 INVX1_1074 ( .A(u2_remHi_135_), .Y(u2__abc_44228_n5170) );
  INVX1 INVX1_1075 ( .A(u2__abc_44228_n5171), .Y(u2__abc_44228_n5172) );
  INVX1 INVX1_1076 ( .A(sqrto_134_), .Y(u2__abc_44228_n5174) );
  INVX1 INVX1_1077 ( .A(u2_remHi_134_), .Y(u2__abc_44228_n5176) );
  INVX1 INVX1_1078 ( .A(u2__abc_44228_n5178), .Y(u2__abc_44228_n5179) );
  INVX1 INVX1_1079 ( .A(sqrto_137_), .Y(u2__abc_44228_n5181) );
  INVX1 INVX1_108 ( .A(\a[6] ), .Y(u1__abc_43968_n276) );
  INVX1 INVX1_1080 ( .A(u2__abc_44228_n5182_1), .Y(u2__abc_44228_n5183) );
  INVX1 INVX1_1081 ( .A(u2_remHi_137_), .Y(u2__abc_44228_n5184) );
  INVX1 INVX1_1082 ( .A(u2__abc_44228_n5185), .Y(u2__abc_44228_n5186) );
  INVX1 INVX1_1083 ( .A(sqrto_136_), .Y(u2__abc_44228_n5188) );
  INVX1 INVX1_1084 ( .A(u2_remHi_136_), .Y(u2__abc_44228_n5190) );
  INVX1 INVX1_1085 ( .A(u2__abc_44228_n5192_1), .Y(u2__abc_44228_n5193) );
  INVX1 INVX1_1086 ( .A(sqrto_133_), .Y(u2__abc_44228_n5197) );
  INVX1 INVX1_1087 ( .A(u2__abc_44228_n5198), .Y(u2__abc_44228_n5199) );
  INVX1 INVX1_1088 ( .A(u2_remHi_133_), .Y(u2__abc_44228_n5200) );
  INVX1 INVX1_1089 ( .A(u2__abc_44228_n5201_1), .Y(u2__abc_44228_n5202) );
  INVX1 INVX1_109 ( .A(\a[7] ), .Y(u1__abc_43968_n277) );
  INVX1 INVX1_1090 ( .A(sqrto_132_), .Y(u2__abc_44228_n5204) );
  INVX1 INVX1_1091 ( .A(u2_remHi_132_), .Y(u2__abc_44228_n5206) );
  INVX1 INVX1_1092 ( .A(u2__abc_44228_n5208), .Y(u2__abc_44228_n5209) );
  INVX1 INVX1_1093 ( .A(sqrto_131_), .Y(u2__abc_44228_n5211_1) );
  INVX1 INVX1_1094 ( .A(u2__abc_44228_n5212), .Y(u2__abc_44228_n5213) );
  INVX1 INVX1_1095 ( .A(u2_remHi_131_), .Y(u2__abc_44228_n5214) );
  INVX1 INVX1_1096 ( .A(u2__abc_44228_n5215), .Y(u2__abc_44228_n5216) );
  INVX1 INVX1_1097 ( .A(sqrto_130_), .Y(u2__abc_44228_n5218) );
  INVX1 INVX1_1098 ( .A(u2_remHi_130_), .Y(u2__abc_44228_n5220) );
  INVX1 INVX1_1099 ( .A(u2__abc_44228_n5222), .Y(u2__abc_44228_n5223) );
  INVX1 INVX1_11 ( .A(_abc_64468_n1543), .Y(_abc_64468_n1546) );
  INVX1 INVX1_110 ( .A(\a[4] ), .Y(u1__abc_43968_n279) );
  INVX1 INVX1_1100 ( .A(u2_remHi_129_), .Y(u2__abc_44228_n5226) );
  INVX1 INVX1_1101 ( .A(sqrto_129_), .Y(u2__abc_44228_n5228) );
  INVX1 INVX1_1102 ( .A(u2_remHi_128_), .Y(u2__abc_44228_n5231) );
  INVX1 INVX1_1103 ( .A(sqrto_128_), .Y(u2__abc_44228_n5233) );
  INVX1 INVX1_1104 ( .A(sqrto_127_), .Y(u2__abc_44228_n5237) );
  INVX1 INVX1_1105 ( .A(u2__abc_44228_n5238), .Y(u2__abc_44228_n5239_1) );
  INVX1 INVX1_1106 ( .A(u2_remHi_127_), .Y(u2__abc_44228_n5240) );
  INVX1 INVX1_1107 ( .A(u2__abc_44228_n5241), .Y(u2__abc_44228_n5242) );
  INVX1 INVX1_1108 ( .A(sqrto_126_), .Y(u2__abc_44228_n5244) );
  INVX1 INVX1_1109 ( .A(u2_remHi_126_), .Y(u2__abc_44228_n5246) );
  INVX1 INVX1_111 ( .A(\a[5] ), .Y(u1__abc_43968_n280) );
  INVX1 INVX1_1110 ( .A(u2__abc_44228_n5248), .Y(u2__abc_44228_n5249) );
  INVX1 INVX1_1111 ( .A(u2__abc_44228_n5227), .Y(u2__abc_44228_n5261) );
  INVX1 INVX1_1112 ( .A(u2__abc_44228_n5232), .Y(u2__abc_44228_n5262) );
  INVX1 INVX1_1113 ( .A(u2__abc_44228_n5160), .Y(u2__abc_44228_n5282) );
  INVX1 INVX1_1114 ( .A(u2__abc_44228_n5283), .Y(u2__abc_44228_n5284) );
  INVX1 INVX1_1115 ( .A(u2__abc_44228_n5115), .Y(u2__abc_44228_n5296) );
  INVX1 INVX1_1116 ( .A(u2__abc_44228_n5297_1), .Y(u2__abc_44228_n5298) );
  INVX1 INVX1_1117 ( .A(u2__abc_44228_n5093), .Y(u2__abc_44228_n5302) );
  INVX1 INVX1_1118 ( .A(u2__abc_44228_n5303), .Y(u2__abc_44228_n5304) );
  INVX1 INVX1_1119 ( .A(u2__abc_44228_n5063), .Y(u2__abc_44228_n5314) );
  INVX1 INVX1_112 ( .A(\a[2] ), .Y(u1__abc_43968_n283) );
  INVX1 INVX1_1120 ( .A(u2__abc_44228_n5315_1), .Y(u2__abc_44228_n5316) );
  INVX1 INVX1_1121 ( .A(u2__abc_44228_n5041), .Y(u2__abc_44228_n5323) );
  INVX1 INVX1_1122 ( .A(u2__abc_44228_n5325), .Y(u2__abc_44228_n5326) );
  INVX1 INVX1_1123 ( .A(u2__abc_44228_n4973), .Y(u2__abc_44228_n5340) );
  INVX1 INVX1_1124 ( .A(u2__abc_44228_n5341), .Y(u2__abc_44228_n5342) );
  INVX1 INVX1_1125 ( .A(u2__abc_44228_n4943), .Y(u2__abc_44228_n5352_1) );
  INVX1 INVX1_1126 ( .A(u2__abc_44228_n5353), .Y(u2__abc_44228_n5354) );
  INVX1 INVX1_1127 ( .A(u2__abc_44228_n4914), .Y(u2__abc_44228_n5359) );
  INVX1 INVX1_1128 ( .A(u2__abc_44228_n5360), .Y(u2__abc_44228_n5361) );
  INVX1 INVX1_1129 ( .A(u2__abc_44228_n4890), .Y(u2__abc_44228_n5370) );
  INVX1 INVX1_113 ( .A(\a[3] ), .Y(u1__abc_43968_n284) );
  INVX1 INVX1_1130 ( .A(u2__abc_44228_n5372_1), .Y(u2__abc_44228_n5373) );
  INVX1 INVX1_1131 ( .A(u2__abc_44228_n4861), .Y(u2__abc_44228_n5379) );
  INVX1 INVX1_1132 ( .A(u2__abc_44228_n5381_1), .Y(u2__abc_44228_n5382) );
  INVX1 INVX1_1133 ( .A(u2__abc_44228_n4802), .Y(u2__abc_44228_n5389) );
  INVX1 INVX1_1134 ( .A(u2__abc_44228_n5391), .Y(u2__abc_44228_n5392) );
  INVX1 INVX1_1135 ( .A(u2__abc_44228_n4817), .Y(u2__abc_44228_n5397) );
  INVX1 INVX1_1136 ( .A(u2__abc_44228_n5399), .Y(u2__abc_44228_n5400_1) );
  INVX1 INVX1_1137 ( .A(u2__abc_44228_n4831), .Y(u2__abc_44228_n5402) );
  INVX1 INVX1_1138 ( .A(u2__abc_44228_n5403), .Y(u2__abc_44228_n5404) );
  INVX1 INVX1_1139 ( .A(u2__abc_44228_n4740), .Y(u2__abc_44228_n5420) );
  INVX1 INVX1_114 ( .A(\a[0] ), .Y(u1__abc_43968_n286) );
  INVX1 INVX1_1140 ( .A(u2__abc_44228_n5422), .Y(u2__abc_44228_n5423) );
  INVX1 INVX1_1141 ( .A(u2__abc_44228_n4703), .Y(u2__abc_44228_n5430) );
  INVX1 INVX1_1142 ( .A(u2__abc_44228_n5431), .Y(u2__abc_44228_n5432) );
  INVX1 INVX1_1143 ( .A(u2__abc_44228_n4681), .Y(u2__abc_44228_n5439) );
  INVX1 INVX1_1144 ( .A(u2__abc_44228_n5441), .Y(u2__abc_44228_n5442) );
  INVX1 INVX1_1145 ( .A(u2__abc_44228_n4650), .Y(u2__abc_44228_n5450) );
  INVX1 INVX1_1146 ( .A(u2__abc_44228_n5452), .Y(u2__abc_44228_n5453) );
  INVX1 INVX1_1147 ( .A(u2__abc_44228_n4614), .Y(u2__abc_44228_n5459) );
  INVX1 INVX1_1148 ( .A(u2__abc_44228_n5460), .Y(u2__abc_44228_n5461) );
  INVX1 INVX1_1149 ( .A(u2__abc_44228_n4584), .Y(u2__abc_44228_n5469) );
  INVX1 INVX1_115 ( .A(\a[1] ), .Y(u1__abc_43968_n287) );
  INVX1 INVX1_1150 ( .A(u2__abc_44228_n5470), .Y(u2__abc_44228_n5471) );
  INVX1 INVX1_1151 ( .A(u2__abc_44228_n4555), .Y(u2__abc_44228_n5480) );
  INVX1 INVX1_1152 ( .A(u2__abc_44228_n5481), .Y(u2__abc_44228_n5482) );
  INVX1 INVX1_1153 ( .A(u2__abc_44228_n4523), .Y(u2__abc_44228_n5490) );
  INVX1 INVX1_1154 ( .A(u2__abc_44228_n5492), .Y(u2__abc_44228_n5493_1) );
  INVX1 INVX1_1155 ( .A(u2__abc_44228_n4494), .Y(u2__abc_44228_n5499) );
  INVX1 INVX1_1156 ( .A(u2__abc_44228_n5500), .Y(u2__abc_44228_n5501) );
  INVX1 INVX1_1157 ( .A(u2__abc_44228_n4457), .Y(u2__abc_44228_n5509) );
  INVX1 INVX1_1158 ( .A(u2__abc_44228_n5511), .Y(u2__abc_44228_n5512_1) );
  INVX1 INVX1_1159 ( .A(u2__abc_44228_n4471_1), .Y(u2__abc_44228_n5514) );
  INVX1 INVX1_116 ( .A(\a[30] ), .Y(u1__abc_43968_n292) );
  INVX1 INVX1_1160 ( .A(u2__abc_44228_n5515), .Y(u2__abc_44228_n5516) );
  INVX1 INVX1_1161 ( .A(u2__abc_44228_n4435), .Y(u2__abc_44228_n5520) );
  INVX1 INVX1_1162 ( .A(u2__abc_44228_n5521), .Y(u2__abc_44228_n5522_1) );
  INVX1 INVX1_1163 ( .A(u2__abc_44228_n4345), .Y(u2__abc_44228_n5531_1) );
  INVX1 INVX1_1164 ( .A(u2__abc_44228_n5532), .Y(u2__abc_44228_n5533) );
  INVX1 INVX1_1165 ( .A(u2__abc_44228_n4316), .Y(u2__abc_44228_n5542) );
  INVX1 INVX1_1166 ( .A(u2__abc_44228_n5543), .Y(u2__abc_44228_n5544) );
  INVX1 INVX1_1167 ( .A(u2__abc_44228_n4404), .Y(u2__abc_44228_n5549_1) );
  INVX1 INVX1_1168 ( .A(u2__abc_44228_n5550), .Y(u2__abc_44228_n5551) );
  INVX1 INVX1_1169 ( .A(u2__abc_44228_n4375), .Y(u2__abc_44228_n5558_1) );
  INVX1 INVX1_117 ( .A(\a[31] ), .Y(u1__abc_43968_n293) );
  INVX1 INVX1_1170 ( .A(u2__abc_44228_n5559), .Y(u2__abc_44228_n5560) );
  INVX1 INVX1_1171 ( .A(u2_o_381_), .Y(u2__abc_44228_n5573) );
  INVX1 INVX1_1172 ( .A(u2__abc_44228_n5574), .Y(u2__abc_44228_n5575) );
  INVX1 INVX1_1173 ( .A(u2_remHi_381_), .Y(u2__abc_44228_n5576) );
  INVX1 INVX1_1174 ( .A(u2__abc_44228_n5577_1), .Y(u2__abc_44228_n5578) );
  INVX1 INVX1_1175 ( .A(u2_o_380_), .Y(u2__abc_44228_n5580) );
  INVX1 INVX1_1176 ( .A(u2_remHi_380_), .Y(u2__abc_44228_n5582) );
  INVX1 INVX1_1177 ( .A(u2__abc_44228_n5584), .Y(u2__abc_44228_n5585) );
  INVX1 INVX1_1178 ( .A(u2_o_379_), .Y(u2__abc_44228_n5587_1) );
  INVX1 INVX1_1179 ( .A(u2__abc_44228_n5588), .Y(u2__abc_44228_n5589) );
  INVX1 INVX1_118 ( .A(\a[28] ), .Y(u1__abc_43968_n295) );
  INVX1 INVX1_1180 ( .A(u2_remHi_379_), .Y(u2__abc_44228_n5590) );
  INVX1 INVX1_1181 ( .A(u2__abc_44228_n5591), .Y(u2__abc_44228_n5592) );
  INVX1 INVX1_1182 ( .A(u2_o_378_), .Y(u2__abc_44228_n5594) );
  INVX1 INVX1_1183 ( .A(u2_remHi_378_), .Y(u2__abc_44228_n5596) );
  INVX1 INVX1_1184 ( .A(u2__abc_44228_n5598), .Y(u2__abc_44228_n5599) );
  INVX1 INVX1_1185 ( .A(u2_o_375_), .Y(u2__abc_44228_n5602) );
  INVX1 INVX1_1186 ( .A(u2__abc_44228_n5603), .Y(u2__abc_44228_n5604) );
  INVX1 INVX1_1187 ( .A(u2_remHi_375_), .Y(u2__abc_44228_n5605) );
  INVX1 INVX1_1188 ( .A(u2__abc_44228_n5606_1), .Y(u2__abc_44228_n5607) );
  INVX1 INVX1_1189 ( .A(u2_o_374_), .Y(u2__abc_44228_n5609) );
  INVX1 INVX1_119 ( .A(\a[29] ), .Y(u1__abc_43968_n296) );
  INVX1 INVX1_1190 ( .A(u2_remHi_374_), .Y(u2__abc_44228_n5611) );
  INVX1 INVX1_1191 ( .A(u2__abc_44228_n5613), .Y(u2__abc_44228_n5614) );
  INVX1 INVX1_1192 ( .A(u2_o_377_), .Y(u2__abc_44228_n5616) );
  INVX1 INVX1_1193 ( .A(u2__abc_44228_n5617), .Y(u2__abc_44228_n5618) );
  INVX1 INVX1_1194 ( .A(u2_remHi_377_), .Y(u2__abc_44228_n5619) );
  INVX1 INVX1_1195 ( .A(u2__abc_44228_n5620), .Y(u2__abc_44228_n5621) );
  INVX1 INVX1_1196 ( .A(u2_o_376_), .Y(u2__abc_44228_n5623) );
  INVX1 INVX1_1197 ( .A(u2_remHi_376_), .Y(u2__abc_44228_n5625) );
  INVX1 INVX1_1198 ( .A(u2__abc_44228_n5627), .Y(u2__abc_44228_n5628) );
  INVX1 INVX1_1199 ( .A(u2_o_373_), .Y(u2__abc_44228_n5632) );
  INVX1 INVX1_12 ( .A(_abc_64468_n1544), .Y(_abc_64468_n1552) );
  INVX1 INVX1_120 ( .A(\a[26] ), .Y(u1__abc_43968_n299) );
  INVX1 INVX1_1200 ( .A(u2__abc_44228_n5633_1), .Y(u2__abc_44228_n5634) );
  INVX1 INVX1_1201 ( .A(u2_remHi_373_), .Y(u2__abc_44228_n5635) );
  INVX1 INVX1_1202 ( .A(u2__abc_44228_n5636), .Y(u2__abc_44228_n5637) );
  INVX1 INVX1_1203 ( .A(u2_o_372_), .Y(u2__abc_44228_n5639) );
  INVX1 INVX1_1204 ( .A(u2_remHi_372_), .Y(u2__abc_44228_n5641) );
  INVX1 INVX1_1205 ( .A(u2__abc_44228_n5643_1), .Y(u2__abc_44228_n5644) );
  INVX1 INVX1_1206 ( .A(u2_o_370_), .Y(u2__abc_44228_n5646) );
  INVX1 INVX1_1207 ( .A(u2_remHi_370_), .Y(u2__abc_44228_n5648) );
  INVX1 INVX1_1208 ( .A(u2__abc_44228_n5650), .Y(u2__abc_44228_n5651) );
  INVX1 INVX1_1209 ( .A(u2_o_371_), .Y(u2__abc_44228_n5652_1) );
  INVX1 INVX1_121 ( .A(\a[27] ), .Y(u1__abc_43968_n300) );
  INVX1 INVX1_1210 ( .A(u2__abc_44228_n5653), .Y(u2__abc_44228_n5654) );
  INVX1 INVX1_1211 ( .A(u2_remHi_371_), .Y(u2__abc_44228_n5655) );
  INVX1 INVX1_1212 ( .A(u2__abc_44228_n5656), .Y(u2__abc_44228_n5657) );
  INVX1 INVX1_1213 ( .A(u2_o_367_), .Y(u2__abc_44228_n5661) );
  INVX1 INVX1_1214 ( .A(u2__abc_44228_n5662_1), .Y(u2__abc_44228_n5663) );
  INVX1 INVX1_1215 ( .A(u2_remHi_367_), .Y(u2__abc_44228_n5664) );
  INVX1 INVX1_1216 ( .A(u2__abc_44228_n5665), .Y(u2__abc_44228_n5666) );
  INVX1 INVX1_1217 ( .A(u2_o_366_), .Y(u2__abc_44228_n5668) );
  INVX1 INVX1_1218 ( .A(u2_remHi_366_), .Y(u2__abc_44228_n5670) );
  INVX1 INVX1_1219 ( .A(u2__abc_44228_n5672_1), .Y(u2__abc_44228_n5673) );
  INVX1 INVX1_122 ( .A(\a[24] ), .Y(u1__abc_43968_n302) );
  INVX1 INVX1_1220 ( .A(u2_o_369_), .Y(u2__abc_44228_n5675) );
  INVX1 INVX1_1221 ( .A(u2__abc_44228_n5676), .Y(u2__abc_44228_n5677) );
  INVX1 INVX1_1222 ( .A(u2_remHi_369_), .Y(u2__abc_44228_n5678) );
  INVX1 INVX1_1223 ( .A(u2__abc_44228_n5679), .Y(u2__abc_44228_n5680) );
  INVX1 INVX1_1224 ( .A(u2_o_368_), .Y(u2__abc_44228_n5682) );
  INVX1 INVX1_1225 ( .A(u2_remHi_368_), .Y(u2__abc_44228_n5684) );
  INVX1 INVX1_1226 ( .A(u2__abc_44228_n5686), .Y(u2__abc_44228_n5687) );
  INVX1 INVX1_1227 ( .A(u2_o_365_), .Y(u2__abc_44228_n5692) );
  INVX1 INVX1_1228 ( .A(u2__abc_44228_n5693), .Y(u2__abc_44228_n5694) );
  INVX1 INVX1_1229 ( .A(u2_remHi_365_), .Y(u2__abc_44228_n5695) );
  INVX1 INVX1_123 ( .A(\a[25] ), .Y(u1__abc_43968_n303) );
  INVX1 INVX1_1230 ( .A(u2__abc_44228_n5696), .Y(u2__abc_44228_n5697) );
  INVX1 INVX1_1231 ( .A(u2_o_364_), .Y(u2__abc_44228_n5699) );
  INVX1 INVX1_1232 ( .A(u2_remHi_364_), .Y(u2__abc_44228_n5701) );
  INVX1 INVX1_1233 ( .A(u2__abc_44228_n5703), .Y(u2__abc_44228_n5704) );
  INVX1 INVX1_1234 ( .A(u2_o_363_), .Y(u2__abc_44228_n5706) );
  INVX1 INVX1_1235 ( .A(u2__abc_44228_n5707), .Y(u2__abc_44228_n5708) );
  INVX1 INVX1_1236 ( .A(u2_remHi_363_), .Y(u2__abc_44228_n5709) );
  INVX1 INVX1_1237 ( .A(u2__abc_44228_n5710_1), .Y(u2__abc_44228_n5711) );
  INVX1 INVX1_1238 ( .A(u2_o_362_), .Y(u2__abc_44228_n5713) );
  INVX1 INVX1_1239 ( .A(u2_remHi_362_), .Y(u2__abc_44228_n5715) );
  INVX1 INVX1_124 ( .A(\a[22] ), .Y(u1__abc_43968_n307) );
  INVX1 INVX1_1240 ( .A(u2__abc_44228_n5717), .Y(u2__abc_44228_n5718) );
  INVX1 INVX1_1241 ( .A(u2_o_359_), .Y(u2__abc_44228_n5721) );
  INVX1 INVX1_1242 ( .A(u2__abc_44228_n5722), .Y(u2__abc_44228_n5723) );
  INVX1 INVX1_1243 ( .A(u2_remHi_359_), .Y(u2__abc_44228_n5724) );
  INVX1 INVX1_1244 ( .A(u2__abc_44228_n5725), .Y(u2__abc_44228_n5726) );
  INVX1 INVX1_1245 ( .A(u2_o_358_), .Y(u2__abc_44228_n5728_1) );
  INVX1 INVX1_1246 ( .A(u2_remHi_358_), .Y(u2__abc_44228_n5730) );
  INVX1 INVX1_1247 ( .A(u2__abc_44228_n5732), .Y(u2__abc_44228_n5733) );
  INVX1 INVX1_1248 ( .A(u2_o_361_), .Y(u2__abc_44228_n5735) );
  INVX1 INVX1_1249 ( .A(u2__abc_44228_n5736), .Y(u2__abc_44228_n5737_1) );
  INVX1 INVX1_125 ( .A(\a[23] ), .Y(u1__abc_43968_n308) );
  INVX1 INVX1_1250 ( .A(u2_remHi_361_), .Y(u2__abc_44228_n5738) );
  INVX1 INVX1_1251 ( .A(u2__abc_44228_n5739), .Y(u2__abc_44228_n5740) );
  INVX1 INVX1_1252 ( .A(u2_o_360_), .Y(u2__abc_44228_n5742) );
  INVX1 INVX1_1253 ( .A(u2_remHi_360_), .Y(u2__abc_44228_n5744) );
  INVX1 INVX1_1254 ( .A(u2__abc_44228_n5746), .Y(u2__abc_44228_n5747_1) );
  INVX1 INVX1_1255 ( .A(u2_o_357_), .Y(u2__abc_44228_n5751) );
  INVX1 INVX1_1256 ( .A(u2__abc_44228_n5752), .Y(u2__abc_44228_n5753) );
  INVX1 INVX1_1257 ( .A(u2_remHi_357_), .Y(u2__abc_44228_n5754) );
  INVX1 INVX1_1258 ( .A(u2__abc_44228_n5755), .Y(u2__abc_44228_n5756_1) );
  INVX1 INVX1_1259 ( .A(u2_o_356_), .Y(u2__abc_44228_n5758) );
  INVX1 INVX1_126 ( .A(\a[20] ), .Y(u1__abc_43968_n310) );
  INVX1 INVX1_1260 ( .A(u2_remHi_356_), .Y(u2__abc_44228_n5760) );
  INVX1 INVX1_1261 ( .A(u2__abc_44228_n5762), .Y(u2__abc_44228_n5763) );
  INVX1 INVX1_1262 ( .A(u2_o_354_), .Y(u2__abc_44228_n5765_1) );
  INVX1 INVX1_1263 ( .A(u2_remHi_354_), .Y(u2__abc_44228_n5767) );
  INVX1 INVX1_1264 ( .A(u2__abc_44228_n5769), .Y(u2__abc_44228_n5770) );
  INVX1 INVX1_1265 ( .A(u2_o_355_), .Y(u2__abc_44228_n5771) );
  INVX1 INVX1_1266 ( .A(u2__abc_44228_n5772), .Y(u2__abc_44228_n5773) );
  INVX1 INVX1_1267 ( .A(u2_remHi_355_), .Y(u2__abc_44228_n5774_1) );
  INVX1 INVX1_1268 ( .A(u2__abc_44228_n5775), .Y(u2__abc_44228_n5776) );
  INVX1 INVX1_1269 ( .A(u2_o_353_), .Y(u2__abc_44228_n5780) );
  INVX1 INVX1_127 ( .A(\a[21] ), .Y(u1__abc_43968_n311) );
  INVX1 INVX1_1270 ( .A(u2__abc_44228_n5781), .Y(u2__abc_44228_n5782) );
  INVX1 INVX1_1271 ( .A(u2_remHi_353_), .Y(u2__abc_44228_n5783_1) );
  INVX1 INVX1_1272 ( .A(u2__abc_44228_n5784), .Y(u2__abc_44228_n5785) );
  INVX1 INVX1_1273 ( .A(u2_o_352_), .Y(u2__abc_44228_n5787) );
  INVX1 INVX1_1274 ( .A(u2_remHi_352_), .Y(u2__abc_44228_n5789) );
  INVX1 INVX1_1275 ( .A(u2__abc_44228_n5791), .Y(u2__abc_44228_n5792) );
  INVX1 INVX1_1276 ( .A(u2_o_351_), .Y(u2__abc_44228_n5794) );
  INVX1 INVX1_1277 ( .A(u2__abc_44228_n5795), .Y(u2__abc_44228_n5796) );
  INVX1 INVX1_1278 ( .A(u2_remHi_351_), .Y(u2__abc_44228_n5797) );
  INVX1 INVX1_1279 ( .A(u2__abc_44228_n5798), .Y(u2__abc_44228_n5799) );
  INVX1 INVX1_128 ( .A(\a[18] ), .Y(u1__abc_43968_n314) );
  INVX1 INVX1_1280 ( .A(u2_o_350_), .Y(u2__abc_44228_n5801) );
  INVX1 INVX1_1281 ( .A(u2_remHi_350_), .Y(u2__abc_44228_n5803) );
  INVX1 INVX1_1282 ( .A(u2__abc_44228_n5805), .Y(u2__abc_44228_n5806) );
  INVX1 INVX1_1283 ( .A(u2_o_349_), .Y(u2__abc_44228_n5812_1) );
  INVX1 INVX1_1284 ( .A(u2__abc_44228_n5813), .Y(u2__abc_44228_n5814) );
  INVX1 INVX1_1285 ( .A(u2_remHi_349_), .Y(u2__abc_44228_n5815) );
  INVX1 INVX1_1286 ( .A(u2__abc_44228_n5816), .Y(u2__abc_44228_n5817) );
  INVX1 INVX1_1287 ( .A(u2_o_348_), .Y(u2__abc_44228_n5819) );
  INVX1 INVX1_1288 ( .A(u2_remHi_348_), .Y(u2__abc_44228_n5821) );
  INVX1 INVX1_1289 ( .A(u2__abc_44228_n5823), .Y(u2__abc_44228_n5824) );
  INVX1 INVX1_129 ( .A(\a[19] ), .Y(u1__abc_43968_n315) );
  INVX1 INVX1_1290 ( .A(u2_o_346_), .Y(u2__abc_44228_n5826) );
  INVX1 INVX1_1291 ( .A(u2_remHi_346_), .Y(u2__abc_44228_n5828) );
  INVX1 INVX1_1292 ( .A(u2__abc_44228_n5830_1), .Y(u2__abc_44228_n5831) );
  INVX1 INVX1_1293 ( .A(u2_o_347_), .Y(u2__abc_44228_n5832) );
  INVX1 INVX1_1294 ( .A(u2__abc_44228_n5833), .Y(u2__abc_44228_n5834) );
  INVX1 INVX1_1295 ( .A(u2_remHi_347_), .Y(u2__abc_44228_n5835) );
  INVX1 INVX1_1296 ( .A(u2__abc_44228_n5836), .Y(u2__abc_44228_n5837) );
  INVX1 INVX1_1297 ( .A(u2_o_343_), .Y(u2__abc_44228_n5841) );
  INVX1 INVX1_1298 ( .A(u2__abc_44228_n5842), .Y(u2__abc_44228_n5843) );
  INVX1 INVX1_1299 ( .A(u2_remHi_343_), .Y(u2__abc_44228_n5844) );
  INVX1 INVX1_13 ( .A(\a[117] ), .Y(_abc_64468_n1555) );
  INVX1 INVX1_130 ( .A(\a[16] ), .Y(u1__abc_43968_n317) );
  INVX1 INVX1_1300 ( .A(u2__abc_44228_n5845_1), .Y(u2__abc_44228_n5846) );
  INVX1 INVX1_1301 ( .A(u2_o_342_), .Y(u2__abc_44228_n5848) );
  INVX1 INVX1_1302 ( .A(u2_remHi_342_), .Y(u2__abc_44228_n5850) );
  INVX1 INVX1_1303 ( .A(u2__abc_44228_n5852), .Y(u2__abc_44228_n5853) );
  INVX1 INVX1_1304 ( .A(u2_o_345_), .Y(u2__abc_44228_n5855) );
  INVX1 INVX1_1305 ( .A(u2__abc_44228_n5856), .Y(u2__abc_44228_n5857) );
  INVX1 INVX1_1306 ( .A(u2_remHi_345_), .Y(u2__abc_44228_n5858) );
  INVX1 INVX1_1307 ( .A(u2__abc_44228_n5859), .Y(u2__abc_44228_n5860) );
  INVX1 INVX1_1308 ( .A(u2_o_344_), .Y(u2__abc_44228_n5862) );
  INVX1 INVX1_1309 ( .A(u2_remHi_344_), .Y(u2__abc_44228_n5864) );
  INVX1 INVX1_131 ( .A(\a[17] ), .Y(u1__abc_43968_n318) );
  INVX1 INVX1_1310 ( .A(u2__abc_44228_n5866), .Y(u2__abc_44228_n5867) );
  INVX1 INVX1_1311 ( .A(u2_o_341_), .Y(u2__abc_44228_n5871) );
  INVX1 INVX1_1312 ( .A(u2__abc_44228_n5872), .Y(u2__abc_44228_n5873_1) );
  INVX1 INVX1_1313 ( .A(u2_remHi_341_), .Y(u2__abc_44228_n5874) );
  INVX1 INVX1_1314 ( .A(u2__abc_44228_n5875), .Y(u2__abc_44228_n5876) );
  INVX1 INVX1_1315 ( .A(u2_o_340_), .Y(u2__abc_44228_n5878) );
  INVX1 INVX1_1316 ( .A(u2_remHi_340_), .Y(u2__abc_44228_n5880) );
  INVX1 INVX1_1317 ( .A(u2__abc_44228_n5882), .Y(u2__abc_44228_n5883_1) );
  INVX1 INVX1_1318 ( .A(u2_o_338_), .Y(u2__abc_44228_n5885) );
  INVX1 INVX1_1319 ( .A(u2_remHi_338_), .Y(u2__abc_44228_n5887) );
  INVX1 INVX1_132 ( .A(\a[94] ), .Y(u1__abc_43968_n324) );
  INVX1 INVX1_1320 ( .A(u2__abc_44228_n5889), .Y(u2__abc_44228_n5890) );
  INVX1 INVX1_1321 ( .A(u2_o_339_), .Y(u2__abc_44228_n5891) );
  INVX1 INVX1_1322 ( .A(u2__abc_44228_n5892_1), .Y(u2__abc_44228_n5893) );
  INVX1 INVX1_1323 ( .A(u2_remHi_339_), .Y(u2__abc_44228_n5894) );
  INVX1 INVX1_1324 ( .A(u2__abc_44228_n5895), .Y(u2__abc_44228_n5896) );
  INVX1 INVX1_1325 ( .A(u2_o_337_), .Y(u2__abc_44228_n5900) );
  INVX1 INVX1_1326 ( .A(u2__abc_44228_n5901_1), .Y(u2__abc_44228_n5902) );
  INVX1 INVX1_1327 ( .A(u2_remHi_337_), .Y(u2__abc_44228_n5903) );
  INVX1 INVX1_1328 ( .A(u2__abc_44228_n5904), .Y(u2__abc_44228_n5905) );
  INVX1 INVX1_1329 ( .A(u2_o_336_), .Y(u2__abc_44228_n5907) );
  INVX1 INVX1_133 ( .A(\a[95] ), .Y(u1__abc_43968_n325) );
  INVX1 INVX1_1330 ( .A(u2_remHi_336_), .Y(u2__abc_44228_n5909) );
  INVX1 INVX1_1331 ( .A(u2__abc_44228_n5911_1), .Y(u2__abc_44228_n5912) );
  INVX1 INVX1_1332 ( .A(u2_o_335_), .Y(u2__abc_44228_n5914) );
  INVX1 INVX1_1333 ( .A(u2__abc_44228_n5915), .Y(u2__abc_44228_n5916) );
  INVX1 INVX1_1334 ( .A(u2_remHi_335_), .Y(u2__abc_44228_n5917) );
  INVX1 INVX1_1335 ( .A(u2__abc_44228_n5918), .Y(u2__abc_44228_n5919) );
  INVX1 INVX1_1336 ( .A(u2_o_334_), .Y(u2__abc_44228_n5921) );
  INVX1 INVX1_1337 ( .A(u2_remHi_334_), .Y(u2__abc_44228_n5923) );
  INVX1 INVX1_1338 ( .A(u2__abc_44228_n5925), .Y(u2__abc_44228_n5926) );
  INVX1 INVX1_1339 ( .A(u2_o_333_), .Y(u2__abc_44228_n5931) );
  INVX1 INVX1_134 ( .A(\a[92] ), .Y(u1__abc_43968_n327) );
  INVX1 INVX1_1340 ( .A(u2__abc_44228_n5932), .Y(u2__abc_44228_n5933) );
  INVX1 INVX1_1341 ( .A(u2_remHi_333_), .Y(u2__abc_44228_n5934) );
  INVX1 INVX1_1342 ( .A(u2__abc_44228_n5935), .Y(u2__abc_44228_n5936) );
  INVX1 INVX1_1343 ( .A(u2_o_332_), .Y(u2__abc_44228_n5938_1) );
  INVX1 INVX1_1344 ( .A(u2_remHi_332_), .Y(u2__abc_44228_n5940) );
  INVX1 INVX1_1345 ( .A(u2__abc_44228_n5942), .Y(u2__abc_44228_n5943) );
  INVX1 INVX1_1346 ( .A(u2_o_331_), .Y(u2__abc_44228_n5945) );
  INVX1 INVX1_1347 ( .A(u2__abc_44228_n5946), .Y(u2__abc_44228_n5947) );
  INVX1 INVX1_1348 ( .A(u2_remHi_331_), .Y(u2__abc_44228_n5948_1) );
  INVX1 INVX1_1349 ( .A(u2__abc_44228_n5949), .Y(u2__abc_44228_n5950) );
  INVX1 INVX1_135 ( .A(\a[93] ), .Y(u1__abc_43968_n328) );
  INVX1 INVX1_1350 ( .A(u2_o_330_), .Y(u2__abc_44228_n5952) );
  INVX1 INVX1_1351 ( .A(u2_remHi_330_), .Y(u2__abc_44228_n5954) );
  INVX1 INVX1_1352 ( .A(u2__abc_44228_n5956), .Y(u2__abc_44228_n5957_1) );
  INVX1 INVX1_1353 ( .A(u2_o_329_), .Y(u2__abc_44228_n5960) );
  INVX1 INVX1_1354 ( .A(u2__abc_44228_n5961), .Y(u2__abc_44228_n5962) );
  INVX1 INVX1_1355 ( .A(u2_remHi_329_), .Y(u2__abc_44228_n5963) );
  INVX1 INVX1_1356 ( .A(u2__abc_44228_n5964), .Y(u2__abc_44228_n5965) );
  INVX1 INVX1_1357 ( .A(u2_o_328_), .Y(u2__abc_44228_n5967) );
  INVX1 INVX1_1358 ( .A(u2_remHi_328_), .Y(u2__abc_44228_n5969) );
  INVX1 INVX1_1359 ( .A(u2__abc_44228_n5971), .Y(u2__abc_44228_n5972) );
  INVX1 INVX1_136 ( .A(\a[90] ), .Y(u1__abc_43968_n331) );
  INVX1 INVX1_1360 ( .A(u2_o_327_), .Y(u2__abc_44228_n5974) );
  INVX1 INVX1_1361 ( .A(u2__abc_44228_n5975_1), .Y(u2__abc_44228_n5976) );
  INVX1 INVX1_1362 ( .A(u2_remHi_327_), .Y(u2__abc_44228_n5977) );
  INVX1 INVX1_1363 ( .A(u2__abc_44228_n5978), .Y(u2__abc_44228_n5979) );
  INVX1 INVX1_1364 ( .A(u2_o_326_), .Y(u2__abc_44228_n5981) );
  INVX1 INVX1_1365 ( .A(u2_remHi_326_), .Y(u2__abc_44228_n5983) );
  INVX1 INVX1_1366 ( .A(u2__abc_44228_n5985_1), .Y(u2__abc_44228_n5986) );
  INVX1 INVX1_1367 ( .A(u2_o_325_), .Y(u2__abc_44228_n5990) );
  INVX1 INVX1_1368 ( .A(u2__abc_44228_n5991), .Y(u2__abc_44228_n5992) );
  INVX1 INVX1_1369 ( .A(u2_remHi_325_), .Y(u2__abc_44228_n5993) );
  INVX1 INVX1_137 ( .A(\a[91] ), .Y(u1__abc_43968_n332) );
  INVX1 INVX1_1370 ( .A(u2__abc_44228_n5994_1), .Y(u2__abc_44228_n5995) );
  INVX1 INVX1_1371 ( .A(u2_o_324_), .Y(u2__abc_44228_n5997) );
  INVX1 INVX1_1372 ( .A(u2_remHi_324_), .Y(u2__abc_44228_n5999) );
  INVX1 INVX1_1373 ( .A(u2__abc_44228_n6001), .Y(u2__abc_44228_n6002) );
  INVX1 INVX1_1374 ( .A(u2_o_322_), .Y(u2__abc_44228_n6004) );
  INVX1 INVX1_1375 ( .A(u2_remHi_322_), .Y(u2__abc_44228_n6006) );
  INVX1 INVX1_1376 ( .A(u2__abc_44228_n6008), .Y(u2__abc_44228_n6009) );
  INVX1 INVX1_1377 ( .A(u2_o_323_), .Y(u2__abc_44228_n6010) );
  INVX1 INVX1_1378 ( .A(u2__abc_44228_n6011), .Y(u2__abc_44228_n6012_1) );
  INVX1 INVX1_1379 ( .A(u2_remHi_323_), .Y(u2__abc_44228_n6013) );
  INVX1 INVX1_138 ( .A(\a[88] ), .Y(u1__abc_43968_n334) );
  INVX1 INVX1_1380 ( .A(u2__abc_44228_n6014), .Y(u2__abc_44228_n6015) );
  INVX1 INVX1_1381 ( .A(u2_o_321_), .Y(u2__abc_44228_n6019) );
  INVX1 INVX1_1382 ( .A(u2__abc_44228_n6020), .Y(u2__abc_44228_n6021) );
  INVX1 INVX1_1383 ( .A(u2_remHi_321_), .Y(u2__abc_44228_n6022_1) );
  INVX1 INVX1_1384 ( .A(u2__abc_44228_n6023), .Y(u2__abc_44228_n6024) );
  INVX1 INVX1_1385 ( .A(u2_o_320_), .Y(u2__abc_44228_n6026) );
  INVX1 INVX1_1386 ( .A(u2_remHi_320_), .Y(u2__abc_44228_n6028) );
  INVX1 INVX1_1387 ( .A(u2__abc_44228_n6030), .Y(u2__abc_44228_n6031_1) );
  INVX1 INVX1_1388 ( .A(u2_o_318_), .Y(u2__abc_44228_n6033) );
  INVX1 INVX1_1389 ( .A(u2_remHi_318_), .Y(u2__abc_44228_n6035) );
  INVX1 INVX1_139 ( .A(\a[89] ), .Y(u1__abc_43968_n335) );
  INVX1 INVX1_1390 ( .A(u2__abc_44228_n6037), .Y(u2__abc_44228_n6038) );
  INVX1 INVX1_1391 ( .A(u2_o_319_), .Y(u2__abc_44228_n6039) );
  INVX1 INVX1_1392 ( .A(u2__abc_44228_n6040_1), .Y(u2__abc_44228_n6041) );
  INVX1 INVX1_1393 ( .A(u2_remHi_319_), .Y(u2__abc_44228_n6042) );
  INVX1 INVX1_1394 ( .A(u2__abc_44228_n6043), .Y(u2__abc_44228_n6044) );
  INVX1 INVX1_1395 ( .A(u2_o_317_), .Y(u2__abc_44228_n6052) );
  INVX1 INVX1_1396 ( .A(u2__abc_44228_n6053), .Y(u2__abc_44228_n6054) );
  INVX1 INVX1_1397 ( .A(u2_remHi_317_), .Y(u2__abc_44228_n6055) );
  INVX1 INVX1_1398 ( .A(u2__abc_44228_n6056), .Y(u2__abc_44228_n6057) );
  INVX1 INVX1_1399 ( .A(u2_o_316_), .Y(u2__abc_44228_n6059_1) );
  INVX1 INVX1_14 ( .A(_abc_64468_n1553), .Y(_abc_64468_n1556) );
  INVX1 INVX1_140 ( .A(\a[86] ), .Y(u1__abc_43968_n339) );
  INVX1 INVX1_1400 ( .A(u2_remHi_316_), .Y(u2__abc_44228_n6061) );
  INVX1 INVX1_1401 ( .A(u2__abc_44228_n6063), .Y(u2__abc_44228_n6064) );
  INVX1 INVX1_1402 ( .A(u2_o_315_), .Y(u2__abc_44228_n6066) );
  INVX1 INVX1_1403 ( .A(u2__abc_44228_n6067), .Y(u2__abc_44228_n6068_1) );
  INVX1 INVX1_1404 ( .A(u2_remHi_315_), .Y(u2__abc_44228_n6069) );
  INVX1 INVX1_1405 ( .A(u2__abc_44228_n6070), .Y(u2__abc_44228_n6071) );
  INVX1 INVX1_1406 ( .A(u2_o_314_), .Y(u2__abc_44228_n6073) );
  INVX1 INVX1_1407 ( .A(u2_remHi_314_), .Y(u2__abc_44228_n6075) );
  INVX1 INVX1_1408 ( .A(u2__abc_44228_n6077), .Y(u2__abc_44228_n6078_1) );
  INVX1 INVX1_1409 ( .A(u2_o_313_), .Y(u2__abc_44228_n6081) );
  INVX1 INVX1_141 ( .A(\a[87] ), .Y(u1__abc_43968_n340) );
  INVX1 INVX1_1410 ( .A(u2__abc_44228_n6082), .Y(u2__abc_44228_n6083) );
  INVX1 INVX1_1411 ( .A(u2_remHi_313_), .Y(u2__abc_44228_n6084) );
  INVX1 INVX1_1412 ( .A(u2__abc_44228_n6085), .Y(u2__abc_44228_n6086_1) );
  INVX1 INVX1_1413 ( .A(u2_o_312_), .Y(u2__abc_44228_n6088) );
  INVX1 INVX1_1414 ( .A(u2_remHi_312_), .Y(u2__abc_44228_n6090) );
  INVX1 INVX1_1415 ( .A(u2__abc_44228_n6092), .Y(u2__abc_44228_n6093) );
  INVX1 INVX1_1416 ( .A(u2_o_311_), .Y(u2__abc_44228_n6095) );
  INVX1 INVX1_1417 ( .A(u2__abc_44228_n6096_1), .Y(u2__abc_44228_n6097) );
  INVX1 INVX1_1418 ( .A(u2_remHi_311_), .Y(u2__abc_44228_n6098) );
  INVX1 INVX1_1419 ( .A(u2__abc_44228_n6099), .Y(u2__abc_44228_n6100) );
  INVX1 INVX1_142 ( .A(\a[84] ), .Y(u1__abc_43968_n342) );
  INVX1 INVX1_1420 ( .A(u2_o_310_), .Y(u2__abc_44228_n6102) );
  INVX1 INVX1_1421 ( .A(u2_remHi_310_), .Y(u2__abc_44228_n6104_1) );
  INVX1 INVX1_1422 ( .A(u2__abc_44228_n6106), .Y(u2__abc_44228_n6107) );
  INVX1 INVX1_1423 ( .A(u2_o_309_), .Y(u2__abc_44228_n6111) );
  INVX1 INVX1_1424 ( .A(u2__abc_44228_n6112), .Y(u2__abc_44228_n6113_1) );
  INVX1 INVX1_1425 ( .A(u2_remHi_309_), .Y(u2__abc_44228_n6114) );
  INVX1 INVX1_1426 ( .A(u2__abc_44228_n6115), .Y(u2__abc_44228_n6116) );
  INVX1 INVX1_1427 ( .A(u2_o_308_), .Y(u2__abc_44228_n6118) );
  INVX1 INVX1_1428 ( .A(u2_remHi_308_), .Y(u2__abc_44228_n6120) );
  INVX1 INVX1_1429 ( .A(u2__abc_44228_n6122_1), .Y(u2__abc_44228_n6123) );
  INVX1 INVX1_143 ( .A(\a[85] ), .Y(u1__abc_43968_n343) );
  INVX1 INVX1_1430 ( .A(u2_o_306_), .Y(u2__abc_44228_n6125) );
  INVX1 INVX1_1431 ( .A(u2_remHi_306_), .Y(u2__abc_44228_n6127) );
  INVX1 INVX1_1432 ( .A(u2__abc_44228_n6129), .Y(u2__abc_44228_n6130) );
  INVX1 INVX1_1433 ( .A(u2_o_307_), .Y(u2__abc_44228_n6131) );
  INVX1 INVX1_1434 ( .A(u2__abc_44228_n6132_1), .Y(u2__abc_44228_n6133) );
  INVX1 INVX1_1435 ( .A(u2_remHi_307_), .Y(u2__abc_44228_n6134) );
  INVX1 INVX1_1436 ( .A(u2__abc_44228_n6135), .Y(u2__abc_44228_n6136) );
  INVX1 INVX1_1437 ( .A(u2_o_305_), .Y(u2__abc_44228_n6140) );
  INVX1 INVX1_1438 ( .A(u2__abc_44228_n6141_1), .Y(u2__abc_44228_n6142) );
  INVX1 INVX1_1439 ( .A(u2_remHi_305_), .Y(u2__abc_44228_n6143) );
  INVX1 INVX1_144 ( .A(\a[82] ), .Y(u1__abc_43968_n346) );
  INVX1 INVX1_1440 ( .A(u2__abc_44228_n6144), .Y(u2__abc_44228_n6145) );
  INVX1 INVX1_1441 ( .A(u2_o_304_), .Y(u2__abc_44228_n6147) );
  INVX1 INVX1_1442 ( .A(u2_remHi_304_), .Y(u2__abc_44228_n6149) );
  INVX1 INVX1_1443 ( .A(u2__abc_44228_n6151_1), .Y(u2__abc_44228_n6152) );
  INVX1 INVX1_1444 ( .A(u2_o_302_), .Y(u2__abc_44228_n6154) );
  INVX1 INVX1_1445 ( .A(u2_remHi_302_), .Y(u2__abc_44228_n6156) );
  INVX1 INVX1_1446 ( .A(u2__abc_44228_n6158), .Y(u2__abc_44228_n6159_1) );
  INVX1 INVX1_1447 ( .A(u2_o_303_), .Y(u2__abc_44228_n6160) );
  INVX1 INVX1_1448 ( .A(u2__abc_44228_n6161), .Y(u2__abc_44228_n6162) );
  INVX1 INVX1_1449 ( .A(u2_remHi_303_), .Y(u2__abc_44228_n6163) );
  INVX1 INVX1_145 ( .A(\a[83] ), .Y(u1__abc_43968_n347) );
  INVX1 INVX1_1450 ( .A(u2__abc_44228_n6164), .Y(u2__abc_44228_n6165) );
  INVX1 INVX1_1451 ( .A(u2_o_301_), .Y(u2__abc_44228_n6171) );
  INVX1 INVX1_1452 ( .A(u2__abc_44228_n6172), .Y(u2__abc_44228_n6173) );
  INVX1 INVX1_1453 ( .A(u2_remHi_301_), .Y(u2__abc_44228_n6174) );
  INVX1 INVX1_1454 ( .A(u2__abc_44228_n6175), .Y(u2__abc_44228_n6176) );
  INVX1 INVX1_1455 ( .A(u2_o_300_), .Y(u2__abc_44228_n6178_1) );
  INVX1 INVX1_1456 ( .A(u2_remHi_300_), .Y(u2__abc_44228_n6180) );
  INVX1 INVX1_1457 ( .A(u2__abc_44228_n6182), .Y(u2__abc_44228_n6183) );
  INVX1 INVX1_1458 ( .A(u2_o_299_), .Y(u2__abc_44228_n6185) );
  INVX1 INVX1_1459 ( .A(u2__abc_44228_n6186), .Y(u2__abc_44228_n6187_1) );
  INVX1 INVX1_146 ( .A(\a[80] ), .Y(u1__abc_43968_n349) );
  INVX1 INVX1_1460 ( .A(u2_remHi_299_), .Y(u2__abc_44228_n6188) );
  INVX1 INVX1_1461 ( .A(u2__abc_44228_n6189), .Y(u2__abc_44228_n6190) );
  INVX1 INVX1_1462 ( .A(u2_o_298_), .Y(u2__abc_44228_n6192) );
  INVX1 INVX1_1463 ( .A(u2_remHi_298_), .Y(u2__abc_44228_n6194) );
  INVX1 INVX1_1464 ( .A(u2__abc_44228_n6196_1), .Y(u2__abc_44228_n6197) );
  INVX1 INVX1_1465 ( .A(u2_o_295_), .Y(u2__abc_44228_n6200) );
  INVX1 INVX1_1466 ( .A(u2__abc_44228_n6201), .Y(u2__abc_44228_n6202) );
  INVX1 INVX1_1467 ( .A(u2_remHi_295_), .Y(u2__abc_44228_n6203) );
  INVX1 INVX1_1468 ( .A(u2__abc_44228_n6204), .Y(u2__abc_44228_n6205) );
  INVX1 INVX1_1469 ( .A(u2_o_294_), .Y(u2__abc_44228_n6207) );
  INVX1 INVX1_147 ( .A(\a[81] ), .Y(u1__abc_43968_n350) );
  INVX1 INVX1_1470 ( .A(u2_remHi_294_), .Y(u2__abc_44228_n6209) );
  INVX1 INVX1_1471 ( .A(u2__abc_44228_n6211), .Y(u2__abc_44228_n6212) );
  INVX1 INVX1_1472 ( .A(u2_o_297_), .Y(u2__abc_44228_n6214_1) );
  INVX1 INVX1_1473 ( .A(u2__abc_44228_n6215), .Y(u2__abc_44228_n6216) );
  INVX1 INVX1_1474 ( .A(u2_remHi_297_), .Y(u2__abc_44228_n6217) );
  INVX1 INVX1_1475 ( .A(u2__abc_44228_n6218), .Y(u2__abc_44228_n6219) );
  INVX1 INVX1_1476 ( .A(u2_o_296_), .Y(u2__abc_44228_n6221) );
  INVX1 INVX1_1477 ( .A(u2_remHi_296_), .Y(u2__abc_44228_n6223) );
  INVX1 INVX1_1478 ( .A(u2__abc_44228_n6225), .Y(u2__abc_44228_n6226) );
  INVX1 INVX1_1479 ( .A(u2_o_293_), .Y(u2__abc_44228_n6230) );
  INVX1 INVX1_148 ( .A(\a[46] ), .Y(u1__abc_43968_n355) );
  INVX1 INVX1_1480 ( .A(u2__abc_44228_n6231), .Y(u2__abc_44228_n6232_1) );
  INVX1 INVX1_1481 ( .A(u2_remHi_293_), .Y(u2__abc_44228_n6233) );
  INVX1 INVX1_1482 ( .A(u2__abc_44228_n6234), .Y(u2__abc_44228_n6235) );
  INVX1 INVX1_1483 ( .A(u2_o_292_), .Y(u2__abc_44228_n6237) );
  INVX1 INVX1_1484 ( .A(u2_remHi_292_), .Y(u2__abc_44228_n6239) );
  INVX1 INVX1_1485 ( .A(u2__abc_44228_n6241), .Y(u2__abc_44228_n6242_1) );
  INVX1 INVX1_1486 ( .A(u2_o_291_), .Y(u2__abc_44228_n6244) );
  INVX1 INVX1_1487 ( .A(u2__abc_44228_n6245), .Y(u2__abc_44228_n6246) );
  INVX1 INVX1_1488 ( .A(u2_remHi_291_), .Y(u2__abc_44228_n6247) );
  INVX1 INVX1_1489 ( .A(u2__abc_44228_n6248), .Y(u2__abc_44228_n6249) );
  INVX1 INVX1_149 ( .A(\a[47] ), .Y(u1__abc_43968_n356) );
  INVX1 INVX1_1490 ( .A(u2_o_290_), .Y(u2__abc_44228_n6251_1) );
  INVX1 INVX1_1491 ( .A(u2_remHi_290_), .Y(u2__abc_44228_n6253) );
  INVX1 INVX1_1492 ( .A(u2__abc_44228_n6255), .Y(u2__abc_44228_n6256) );
  INVX1 INVX1_1493 ( .A(u2_o_289_), .Y(u2__abc_44228_n6259) );
  INVX1 INVX1_1494 ( .A(u2__abc_44228_n6260_1), .Y(u2__abc_44228_n6261) );
  INVX1 INVX1_1495 ( .A(u2_remHi_289_), .Y(u2__abc_44228_n6262) );
  INVX1 INVX1_1496 ( .A(u2__abc_44228_n6263), .Y(u2__abc_44228_n6264) );
  INVX1 INVX1_1497 ( .A(u2_o_288_), .Y(u2__abc_44228_n6266) );
  INVX1 INVX1_1498 ( .A(u2_remHi_288_), .Y(u2__abc_44228_n6268) );
  INVX1 INVX1_1499 ( .A(u2__abc_44228_n6270), .Y(u2__abc_44228_n6271) );
  INVX1 INVX1_15 ( .A(_abc_64468_n1558), .Y(_abc_64468_n1559) );
  INVX1 INVX1_150 ( .A(\a[44] ), .Y(u1__abc_43968_n358) );
  INVX1 INVX1_1500 ( .A(u2_o_287_), .Y(u2__abc_44228_n6273) );
  INVX1 INVX1_1501 ( .A(u2__abc_44228_n6274), .Y(u2__abc_44228_n6275) );
  INVX1 INVX1_1502 ( .A(u2_remHi_287_), .Y(u2__abc_44228_n6276) );
  INVX1 INVX1_1503 ( .A(u2__abc_44228_n6277), .Y(u2__abc_44228_n6278) );
  INVX1 INVX1_1504 ( .A(u2_o_286_), .Y(u2__abc_44228_n6280) );
  INVX1 INVX1_1505 ( .A(u2_remHi_286_), .Y(u2__abc_44228_n6282) );
  INVX1 INVX1_1506 ( .A(u2__abc_44228_n6284), .Y(u2__abc_44228_n6285) );
  INVX1 INVX1_1507 ( .A(u2_o_285_), .Y(u2__abc_44228_n6291) );
  INVX1 INVX1_1508 ( .A(u2__abc_44228_n6292), .Y(u2__abc_44228_n6293) );
  INVX1 INVX1_1509 ( .A(u2_remHi_285_), .Y(u2__abc_44228_n6294) );
  INVX1 INVX1_151 ( .A(\a[45] ), .Y(u1__abc_43968_n359) );
  INVX1 INVX1_1510 ( .A(u2__abc_44228_n6295), .Y(u2__abc_44228_n6296_1) );
  INVX1 INVX1_1511 ( .A(u2_o_284_), .Y(u2__abc_44228_n6298) );
  INVX1 INVX1_1512 ( .A(u2_remHi_284_), .Y(u2__abc_44228_n6300) );
  INVX1 INVX1_1513 ( .A(u2__abc_44228_n6302), .Y(u2__abc_44228_n6303) );
  INVX1 INVX1_1514 ( .A(u2_o_283_), .Y(u2__abc_44228_n6305_1) );
  INVX1 INVX1_1515 ( .A(u2__abc_44228_n6306), .Y(u2__abc_44228_n6307) );
  INVX1 INVX1_1516 ( .A(u2_remHi_283_), .Y(u2__abc_44228_n6308) );
  INVX1 INVX1_1517 ( .A(u2__abc_44228_n6309), .Y(u2__abc_44228_n6310) );
  INVX1 INVX1_1518 ( .A(u2_o_282_), .Y(u2__abc_44228_n6312) );
  INVX1 INVX1_1519 ( .A(u2_remHi_282_), .Y(u2__abc_44228_n6314) );
  INVX1 INVX1_152 ( .A(\a[42] ), .Y(u1__abc_43968_n362) );
  INVX1 INVX1_1520 ( .A(u2__abc_44228_n6316), .Y(u2__abc_44228_n6317) );
  INVX1 INVX1_1521 ( .A(u2_o_279_), .Y(u2__abc_44228_n6320) );
  INVX1 INVX1_1522 ( .A(u2__abc_44228_n6321), .Y(u2__abc_44228_n6322) );
  INVX1 INVX1_1523 ( .A(u2_remHi_279_), .Y(u2__abc_44228_n6323) );
  INVX1 INVX1_1524 ( .A(u2__abc_44228_n6324_1), .Y(u2__abc_44228_n6325) );
  INVX1 INVX1_1525 ( .A(u2_o_278_), .Y(u2__abc_44228_n6327) );
  INVX1 INVX1_1526 ( .A(u2_remHi_278_), .Y(u2__abc_44228_n6329) );
  INVX1 INVX1_1527 ( .A(u2__abc_44228_n6331), .Y(u2__abc_44228_n6332) );
  INVX1 INVX1_1528 ( .A(u2_o_281_), .Y(u2__abc_44228_n6334) );
  INVX1 INVX1_1529 ( .A(u2__abc_44228_n6335), .Y(u2__abc_44228_n6336) );
  INVX1 INVX1_153 ( .A(\a[43] ), .Y(u1__abc_43968_n363) );
  INVX1 INVX1_1530 ( .A(u2_remHi_281_), .Y(u2__abc_44228_n6337) );
  INVX1 INVX1_1531 ( .A(u2__abc_44228_n6338), .Y(u2__abc_44228_n6339) );
  INVX1 INVX1_1532 ( .A(u2_o_280_), .Y(u2__abc_44228_n6341) );
  INVX1 INVX1_1533 ( .A(u2_remHi_280_), .Y(u2__abc_44228_n6343) );
  INVX1 INVX1_1534 ( .A(u2__abc_44228_n6345), .Y(u2__abc_44228_n6346) );
  INVX1 INVX1_1535 ( .A(u2_o_277_), .Y(u2__abc_44228_n6350) );
  INVX1 INVX1_1536 ( .A(u2__abc_44228_n6351), .Y(u2__abc_44228_n6352_1) );
  INVX1 INVX1_1537 ( .A(u2_remHi_277_), .Y(u2__abc_44228_n6353) );
  INVX1 INVX1_1538 ( .A(u2__abc_44228_n6354), .Y(u2__abc_44228_n6355) );
  INVX1 INVX1_1539 ( .A(u2_o_276_), .Y(u2__abc_44228_n6357) );
  INVX1 INVX1_154 ( .A(\a[40] ), .Y(u1__abc_43968_n365) );
  INVX1 INVX1_1540 ( .A(u2_remHi_276_), .Y(u2__abc_44228_n6359) );
  INVX1 INVX1_1541 ( .A(u2__abc_44228_n6361_1), .Y(u2__abc_44228_n6362) );
  INVX1 INVX1_1542 ( .A(u2_o_275_), .Y(u2__abc_44228_n6364) );
  INVX1 INVX1_1543 ( .A(u2__abc_44228_n6365), .Y(u2__abc_44228_n6366) );
  INVX1 INVX1_1544 ( .A(u2_remHi_275_), .Y(u2__abc_44228_n6367) );
  INVX1 INVX1_1545 ( .A(u2__abc_44228_n6368), .Y(u2__abc_44228_n6369) );
  INVX1 INVX1_1546 ( .A(u2_o_274_), .Y(u2__abc_44228_n6371_1) );
  INVX1 INVX1_1547 ( .A(u2_remHi_274_), .Y(u2__abc_44228_n6373) );
  INVX1 INVX1_1548 ( .A(u2__abc_44228_n6375), .Y(u2__abc_44228_n6376) );
  INVX1 INVX1_1549 ( .A(u2_o_273_), .Y(u2__abc_44228_n6379_1) );
  INVX1 INVX1_155 ( .A(\a[41] ), .Y(u1__abc_43968_n366) );
  INVX1 INVX1_1550 ( .A(u2__abc_44228_n6380), .Y(u2__abc_44228_n6381) );
  INVX1 INVX1_1551 ( .A(u2_remHi_273_), .Y(u2__abc_44228_n6382) );
  INVX1 INVX1_1552 ( .A(u2__abc_44228_n6383), .Y(u2__abc_44228_n6384) );
  INVX1 INVX1_1553 ( .A(u2_o_272_), .Y(u2__abc_44228_n6386) );
  INVX1 INVX1_1554 ( .A(u2_remHi_272_), .Y(u2__abc_44228_n6388) );
  INVX1 INVX1_1555 ( .A(u2__abc_44228_n6390), .Y(u2__abc_44228_n6391) );
  INVX1 INVX1_1556 ( .A(u2_o_270_), .Y(u2__abc_44228_n6393) );
  INVX1 INVX1_1557 ( .A(u2_remHi_270_), .Y(u2__abc_44228_n6395) );
  INVX1 INVX1_1558 ( .A(u2__abc_44228_n6397_1), .Y(u2__abc_44228_n6398) );
  INVX1 INVX1_1559 ( .A(u2_o_271_), .Y(u2__abc_44228_n6399) );
  INVX1 INVX1_156 ( .A(\a[38] ), .Y(u1__abc_43968_n370) );
  INVX1 INVX1_1560 ( .A(u2__abc_44228_n6400), .Y(u2__abc_44228_n6401) );
  INVX1 INVX1_1561 ( .A(u2_remHi_271_), .Y(u2__abc_44228_n6402) );
  INVX1 INVX1_1562 ( .A(u2__abc_44228_n6403), .Y(u2__abc_44228_n6404) );
  INVX1 INVX1_1563 ( .A(u2_o_269_), .Y(u2__abc_44228_n6410) );
  INVX1 INVX1_1564 ( .A(u2__abc_44228_n6411), .Y(u2__abc_44228_n6412) );
  INVX1 INVX1_1565 ( .A(u2_remHi_269_), .Y(u2__abc_44228_n6413) );
  INVX1 INVX1_1566 ( .A(u2__abc_44228_n6414), .Y(u2__abc_44228_n6415_1) );
  INVX1 INVX1_1567 ( .A(u2_o_268_), .Y(u2__abc_44228_n6417) );
  INVX1 INVX1_1568 ( .A(u2_remHi_268_), .Y(u2__abc_44228_n6419) );
  INVX1 INVX1_1569 ( .A(u2__abc_44228_n6421), .Y(u2__abc_44228_n6422) );
  INVX1 INVX1_157 ( .A(\a[39] ), .Y(u1__abc_43968_n371) );
  INVX1 INVX1_1570 ( .A(u2_o_267_), .Y(u2__abc_44228_n6424) );
  INVX1 INVX1_1571 ( .A(u2__abc_44228_n6425_1), .Y(u2__abc_44228_n6426) );
  INVX1 INVX1_1572 ( .A(u2_remHi_267_), .Y(u2__abc_44228_n6427) );
  INVX1 INVX1_1573 ( .A(u2__abc_44228_n6428), .Y(u2__abc_44228_n6429) );
  INVX1 INVX1_1574 ( .A(u2_o_266_), .Y(u2__abc_44228_n6431) );
  INVX1 INVX1_1575 ( .A(u2_remHi_266_), .Y(u2__abc_44228_n6433) );
  INVX1 INVX1_1576 ( .A(u2__abc_44228_n6435_1), .Y(u2__abc_44228_n6436) );
  INVX1 INVX1_1577 ( .A(u2_o_265_), .Y(u2__abc_44228_n6439) );
  INVX1 INVX1_1578 ( .A(u2__abc_44228_n6440), .Y(u2__abc_44228_n6441) );
  INVX1 INVX1_1579 ( .A(u2_remHi_265_), .Y(u2__abc_44228_n6442) );
  INVX1 INVX1_158 ( .A(\a[36] ), .Y(u1__abc_43968_n373) );
  INVX1 INVX1_1580 ( .A(u2__abc_44228_n6443), .Y(u2__abc_44228_n6444) );
  INVX1 INVX1_1581 ( .A(u2_o_264_), .Y(u2__abc_44228_n6446) );
  INVX1 INVX1_1582 ( .A(u2_remHi_264_), .Y(u2__abc_44228_n6448) );
  INVX1 INVX1_1583 ( .A(u2__abc_44228_n6450), .Y(u2__abc_44228_n6451) );
  INVX1 INVX1_1584 ( .A(u2_o_263_), .Y(u2__abc_44228_n6453_1) );
  INVX1 INVX1_1585 ( .A(u2__abc_44228_n6454), .Y(u2__abc_44228_n6455) );
  INVX1 INVX1_1586 ( .A(u2_remHi_263_), .Y(u2__abc_44228_n6456) );
  INVX1 INVX1_1587 ( .A(u2__abc_44228_n6457), .Y(u2__abc_44228_n6458) );
  INVX1 INVX1_1588 ( .A(u2_o_262_), .Y(u2__abc_44228_n6460) );
  INVX1 INVX1_1589 ( .A(u2_remHi_262_), .Y(u2__abc_44228_n6462) );
  INVX1 INVX1_159 ( .A(\a[37] ), .Y(u1__abc_43968_n374) );
  INVX1 INVX1_1590 ( .A(u2__abc_44228_n6464), .Y(u2__abc_44228_n6465) );
  INVX1 INVX1_1591 ( .A(u2_o_261_), .Y(u2__abc_44228_n6469) );
  INVX1 INVX1_1592 ( .A(u2__abc_44228_n6470), .Y(u2__abc_44228_n6471_1) );
  INVX1 INVX1_1593 ( .A(u2_remHi_261_), .Y(u2__abc_44228_n6472) );
  INVX1 INVX1_1594 ( .A(u2__abc_44228_n6473), .Y(u2__abc_44228_n6474) );
  INVX1 INVX1_1595 ( .A(u2_o_260_), .Y(u2__abc_44228_n6476) );
  INVX1 INVX1_1596 ( .A(u2_remHi_260_), .Y(u2__abc_44228_n6478) );
  INVX1 INVX1_1597 ( .A(u2__abc_44228_n6480_1), .Y(u2__abc_44228_n6481) );
  INVX1 INVX1_1598 ( .A(u2_o_259_), .Y(u2__abc_44228_n6483) );
  INVX1 INVX1_1599 ( .A(u2__abc_44228_n6484), .Y(u2__abc_44228_n6485) );
  INVX1 INVX1_16 ( .A(_abc_64468_n1561), .Y(_abc_64468_n1567) );
  INVX1 INVX1_160 ( .A(\a[34] ), .Y(u1__abc_43968_n377) );
  INVX1 INVX1_1600 ( .A(u2_remHi_259_), .Y(u2__abc_44228_n6486) );
  INVX1 INVX1_1601 ( .A(u2__abc_44228_n6487), .Y(u2__abc_44228_n6488) );
  INVX1 INVX1_1602 ( .A(u2_o_258_), .Y(u2__abc_44228_n6490) );
  INVX1 INVX1_1603 ( .A(u2_remHi_258_), .Y(u2__abc_44228_n6492) );
  INVX1 INVX1_1604 ( .A(u2__abc_44228_n6494), .Y(u2__abc_44228_n6495) );
  INVX1 INVX1_1605 ( .A(u2_o_257_), .Y(u2__abc_44228_n6498) );
  INVX1 INVX1_1606 ( .A(u2__abc_44228_n6499_1), .Y(u2__abc_44228_n6500) );
  INVX1 INVX1_1607 ( .A(u2_remHi_257_), .Y(u2__abc_44228_n6501) );
  INVX1 INVX1_1608 ( .A(u2__abc_44228_n6502), .Y(u2__abc_44228_n6503) );
  INVX1 INVX1_1609 ( .A(u2_o_256_), .Y(u2__abc_44228_n6505) );
  INVX1 INVX1_161 ( .A(\a[35] ), .Y(u1__abc_43968_n378) );
  INVX1 INVX1_1610 ( .A(u2_remHi_256_), .Y(u2__abc_44228_n6507_1) );
  INVX1 INVX1_1611 ( .A(u2__abc_44228_n6509), .Y(u2__abc_44228_n6510) );
  INVX1 INVX1_1612 ( .A(u2_o_255_), .Y(u2__abc_44228_n6512) );
  INVX1 INVX1_1613 ( .A(u2__abc_44228_n6513), .Y(u2__abc_44228_n6514) );
  INVX1 INVX1_1614 ( .A(u2_remHi_255_), .Y(u2__abc_44228_n6515) );
  INVX1 INVX1_1615 ( .A(u2__abc_44228_n6516), .Y(u2__abc_44228_n6517_1) );
  INVX1 INVX1_1616 ( .A(u2_o_254_), .Y(u2__abc_44228_n6519) );
  INVX1 INVX1_1617 ( .A(u2_remHi_254_), .Y(u2__abc_44228_n6521) );
  INVX1 INVX1_1618 ( .A(u2__abc_44228_n6523), .Y(u2__abc_44228_n6524) );
  INVX1 INVX1_1619 ( .A(u2__abc_44228_n6520), .Y(u2__abc_44228_n6533) );
  INVX1 INVX1_162 ( .A(\a[32] ), .Y(u1__abc_43968_n380) );
  INVX1 INVX1_1620 ( .A(u2__abc_44228_n6535_1), .Y(u2__abc_44228_n6536) );
  INVX1 INVX1_1621 ( .A(u2__abc_44228_n6491), .Y(u2__abc_44228_n6542) );
  INVX1 INVX1_1622 ( .A(u2__abc_44228_n6544), .Y(u2__abc_44228_n6545) );
  INVX1 INVX1_1623 ( .A(u2__abc_44228_n6461), .Y(u2__abc_44228_n6554) );
  INVX1 INVX1_1624 ( .A(u2__abc_44228_n6555), .Y(u2__abc_44228_n6556) );
  INVX1 INVX1_1625 ( .A(u2__abc_44228_n6432), .Y(u2__abc_44228_n6561_1) );
  INVX1 INVX1_1626 ( .A(u2__abc_44228_n6563), .Y(u2__abc_44228_n6564) );
  INVX1 INVX1_1627 ( .A(u2__abc_44228_n6394), .Y(u2__abc_44228_n6572) );
  INVX1 INVX1_1628 ( .A(u2__abc_44228_n6573), .Y(u2__abc_44228_n6574) );
  INVX1 INVX1_1629 ( .A(u2__abc_44228_n6372), .Y(u2__abc_44228_n6581) );
  INVX1 INVX1_163 ( .A(\a[33] ), .Y(u1__abc_43968_n381) );
  INVX1 INVX1_1630 ( .A(u2__abc_44228_n6583), .Y(u2__abc_44228_n6584) );
  INVX1 INVX1_1631 ( .A(u2__abc_44228_n6328), .Y(u2__abc_44228_n6591) );
  INVX1 INVX1_1632 ( .A(u2__abc_44228_n6593), .Y(u2__abc_44228_n6594) );
  INVX1 INVX1_1633 ( .A(u2__abc_44228_n6342_1), .Y(u2__abc_44228_n6596) );
  INVX1 INVX1_1634 ( .A(u2__abc_44228_n6597_1), .Y(u2__abc_44228_n6598) );
  INVX1 INVX1_1635 ( .A(u2__abc_44228_n6313), .Y(u2__abc_44228_n6604) );
  INVX1 INVX1_1636 ( .A(u2__abc_44228_n6605), .Y(u2__abc_44228_n6606) );
  INVX1 INVX1_1637 ( .A(u2__abc_44228_n6281), .Y(u2__abc_44228_n6614) );
  INVX1 INVX1_1638 ( .A(u2__abc_44228_n6616_1), .Y(u2__abc_44228_n6617) );
  INVX1 INVX1_1639 ( .A(u2__abc_44228_n6252), .Y(u2__abc_44228_n6623) );
  INVX1 INVX1_164 ( .A(u1_mz), .Y(u1__abc_43968_n392) );
  INVX1 INVX1_1640 ( .A(u2__abc_44228_n6625_1), .Y(u2__abc_44228_n6626) );
  INVX1 INVX1_1641 ( .A(u2__abc_44228_n6208), .Y(u2__abc_44228_n6633) );
  INVX1 INVX1_1642 ( .A(u2__abc_44228_n6635), .Y(u2__abc_44228_n6636) );
  INVX1 INVX1_1643 ( .A(u2__abc_44228_n6222), .Y(u2__abc_44228_n6638) );
  INVX1 INVX1_1644 ( .A(u2__abc_44228_n6639), .Y(u2__abc_44228_n6640) );
  INVX1 INVX1_1645 ( .A(u2__abc_44228_n6193), .Y(u2__abc_44228_n6644_1) );
  INVX1 INVX1_1646 ( .A(u2__abc_44228_n6645), .Y(u2__abc_44228_n6646) );
  INVX1 INVX1_1647 ( .A(u2__abc_44228_n6155), .Y(u2__abc_44228_n6655) );
  INVX1 INVX1_1648 ( .A(u2__abc_44228_n6657), .Y(u2__abc_44228_n6658) );
  INVX1 INVX1_1649 ( .A(u2__abc_44228_n6126), .Y(u2__abc_44228_n6664) );
  INVX1 INVX1_165 ( .A(ld), .Y(u2__abc_44228_n2962) );
  INVX1 INVX1_1650 ( .A(u2__abc_44228_n6666), .Y(u2__abc_44228_n6667) );
  INVX1 INVX1_1651 ( .A(u2__abc_44228_n6103), .Y(u2__abc_44228_n6674) );
  INVX1 INVX1_1652 ( .A(u2__abc_44228_n6676), .Y(u2__abc_44228_n6677) );
  INVX1 INVX1_1653 ( .A(u2__abc_44228_n6089), .Y(u2__abc_44228_n6679) );
  INVX1 INVX1_1654 ( .A(u2__abc_44228_n6680), .Y(u2__abc_44228_n6681_1) );
  INVX1 INVX1_1655 ( .A(u2__abc_44228_n6074), .Y(u2__abc_44228_n6687) );
  INVX1 INVX1_1656 ( .A(u2__abc_44228_n6689_1), .Y(u2__abc_44228_n6690) );
  INVX1 INVX1_1657 ( .A(u2__abc_44228_n6034), .Y(u2__abc_44228_n6698_1) );
  INVX1 INVX1_1658 ( .A(u2__abc_44228_n6699), .Y(u2__abc_44228_n6700) );
  INVX1 INVX1_1659 ( .A(u2__abc_44228_n6005), .Y(u2__abc_44228_n6707_1) );
  INVX1 INVX1_166 ( .A(ce), .Y(u2__abc_44228_n2967) );
  INVX1 INVX1_1660 ( .A(u2__abc_44228_n6708), .Y(u2__abc_44228_n6709) );
  INVX1 INVX1_1661 ( .A(u2__abc_44228_n5982), .Y(u2__abc_44228_n6719) );
  INVX1 INVX1_1662 ( .A(u2__abc_44228_n6720), .Y(u2__abc_44228_n6721) );
  INVX1 INVX1_1663 ( .A(u2__abc_44228_n5953), .Y(u2__abc_44228_n6726) );
  INVX1 INVX1_1664 ( .A(u2__abc_44228_n6727), .Y(u2__abc_44228_n6728) );
  INVX1 INVX1_1665 ( .A(u2__abc_44228_n5922), .Y(u2__abc_44228_n6737) );
  INVX1 INVX1_1666 ( .A(u2__abc_44228_n6739), .Y(u2__abc_44228_n6740) );
  INVX1 INVX1_1667 ( .A(u2__abc_44228_n5886), .Y(u2__abc_44228_n6746) );
  INVX1 INVX1_1668 ( .A(u2__abc_44228_n6747), .Y(u2__abc_44228_n6748) );
  INVX1 INVX1_1669 ( .A(u2__abc_44228_n5849), .Y(u2__abc_44228_n6756) );
  INVX1 INVX1_167 ( .A(u2_cnt_0_), .Y(u2__abc_44228_n2974) );
  INVX1 INVX1_1670 ( .A(u2__abc_44228_n6758), .Y(u2__abc_44228_n6759) );
  INVX1 INVX1_1671 ( .A(u2__abc_44228_n5863_1), .Y(u2__abc_44228_n6761_1) );
  INVX1 INVX1_1672 ( .A(u2__abc_44228_n6762), .Y(u2__abc_44228_n6763) );
  INVX1 INVX1_1673 ( .A(u2__abc_44228_n5827), .Y(u2__abc_44228_n6769) );
  INVX1 INVX1_1674 ( .A(u2__abc_44228_n6770_1), .Y(u2__abc_44228_n6771) );
  INVX1 INVX1_1675 ( .A(u2__abc_44228_n5802_1), .Y(u2__abc_44228_n6779_1) );
  INVX1 INVX1_1676 ( .A(u2__abc_44228_n6781), .Y(u2__abc_44228_n6782) );
  INVX1 INVX1_1677 ( .A(u2__abc_44228_n5766), .Y(u2__abc_44228_n6788) );
  INVX1 INVX1_1678 ( .A(u2__abc_44228_n6789_1), .Y(u2__abc_44228_n6790) );
  INVX1 INVX1_1679 ( .A(u2__abc_44228_n5729), .Y(u2__abc_44228_n6798) );
  INVX1 INVX1_168 ( .A(u2__abc_44228_n2976), .Y(u2__abc_44228_n2977) );
  INVX1 INVX1_1680 ( .A(u2__abc_44228_n6800), .Y(u2__abc_44228_n6801) );
  INVX1 INVX1_1681 ( .A(u2__abc_44228_n5743), .Y(u2__abc_44228_n6803) );
  INVX1 INVX1_1682 ( .A(u2__abc_44228_n6804), .Y(u2__abc_44228_n6805) );
  INVX1 INVX1_1683 ( .A(u2__abc_44228_n5714), .Y(u2__abc_44228_n6811) );
  INVX1 INVX1_1684 ( .A(u2__abc_44228_n6813), .Y(u2__abc_44228_n6814) );
  INVX1 INVX1_1685 ( .A(u2__abc_44228_n5669), .Y(u2__abc_44228_n6820) );
  INVX1 INVX1_1686 ( .A(u2__abc_44228_n6822), .Y(u2__abc_44228_n6823) );
  INVX1 INVX1_1687 ( .A(u2__abc_44228_n5683), .Y(u2__abc_44228_n6825_1) );
  INVX1 INVX1_1688 ( .A(u2__abc_44228_n6826), .Y(u2__abc_44228_n6827) );
  INVX1 INVX1_1689 ( .A(u2__abc_44228_n5647), .Y(u2__abc_44228_n6831) );
  INVX1 INVX1_169 ( .A(u2_cnt_4_), .Y(u2__abc_44228_n2979) );
  INVX1 INVX1_1690 ( .A(u2__abc_44228_n6832), .Y(u2__abc_44228_n6833_1) );
  INVX1 INVX1_1691 ( .A(u2__abc_44228_n5610), .Y(u2__abc_44228_n6841) );
  INVX1 INVX1_1692 ( .A(u2__abc_44228_n6843), .Y(u2__abc_44228_n6844) );
  INVX1 INVX1_1693 ( .A(u2__abc_44228_n5624_1), .Y(u2__abc_44228_n6846) );
  INVX1 INVX1_1694 ( .A(u2__abc_44228_n6847), .Y(u2__abc_44228_n6848) );
  INVX1 INVX1_1695 ( .A(u2__abc_44228_n5595), .Y(u2__abc_44228_n6854) );
  INVX1 INVX1_1696 ( .A(u2__abc_44228_n6855), .Y(u2__abc_44228_n6856) );
  INVX1 INVX1_1697 ( .A(u2_o_445_), .Y(u2__abc_44228_n6866) );
  INVX1 INVX1_1698 ( .A(u2__abc_44228_n6867), .Y(u2__abc_44228_n6868) );
  INVX1 INVX1_1699 ( .A(u2_remHi_445_), .Y(u2__abc_44228_n6869_1) );
  INVX1 INVX1_17 ( .A(\a[118] ), .Y(_abc_64468_n1568) );
  INVX1 INVX1_170 ( .A(u2__abc_44228_n2988_bF_buf12), .Y(u2__abc_44228_n2995) );
  INVX1 INVX1_1700 ( .A(u2__abc_44228_n6870), .Y(u2__abc_44228_n6871) );
  INVX1 INVX1_1701 ( .A(u2_o_444_), .Y(u2__abc_44228_n6873) );
  INVX1 INVX1_1702 ( .A(u2_remHi_444_), .Y(u2__abc_44228_n6875) );
  INVX1 INVX1_1703 ( .A(u2__abc_44228_n6877), .Y(u2__abc_44228_n6878_1) );
  INVX1 INVX1_1704 ( .A(u2_o_443_), .Y(u2__abc_44228_n6880) );
  INVX1 INVX1_1705 ( .A(u2__abc_44228_n6881), .Y(u2__abc_44228_n6882) );
  INVX1 INVX1_1706 ( .A(u2_remHi_443_), .Y(u2__abc_44228_n6883) );
  INVX1 INVX1_1707 ( .A(u2__abc_44228_n6884), .Y(u2__abc_44228_n6885) );
  INVX1 INVX1_1708 ( .A(u2_o_442_), .Y(u2__abc_44228_n6887_1) );
  INVX1 INVX1_1709 ( .A(u2_remHi_442_), .Y(u2__abc_44228_n6889) );
  INVX1 INVX1_171 ( .A(u2__abc_44228_n3003), .Y(u2__abc_44228_n3004) );
  INVX1 INVX1_1710 ( .A(u2__abc_44228_n6891), .Y(u2__abc_44228_n6892) );
  INVX1 INVX1_1711 ( .A(u2_o_441_), .Y(u2__abc_44228_n6895) );
  INVX1 INVX1_1712 ( .A(u2__abc_44228_n6896), .Y(u2__abc_44228_n6897_1) );
  INVX1 INVX1_1713 ( .A(u2_remHi_441_), .Y(u2__abc_44228_n6898) );
  INVX1 INVX1_1714 ( .A(u2__abc_44228_n6899), .Y(u2__abc_44228_n6900) );
  INVX1 INVX1_1715 ( .A(u2_o_440_), .Y(u2__abc_44228_n6902) );
  INVX1 INVX1_1716 ( .A(u2_remHi_440_), .Y(u2__abc_44228_n6904) );
  INVX1 INVX1_1717 ( .A(u2__abc_44228_n6906_1), .Y(u2__abc_44228_n6907) );
  INVX1 INVX1_1718 ( .A(u2_o_439_), .Y(u2__abc_44228_n6909) );
  INVX1 INVX1_1719 ( .A(u2__abc_44228_n6910), .Y(u2__abc_44228_n6911) );
  INVX1 INVX1_172 ( .A(u2__abc_44228_n2968), .Y(u2__abc_44228_n3008) );
  INVX1 INVX1_1720 ( .A(u2_remHi_439_), .Y(u2__abc_44228_n6912) );
  INVX1 INVX1_1721 ( .A(u2__abc_44228_n6913), .Y(u2__abc_44228_n6914) );
  INVX1 INVX1_1722 ( .A(u2_o_438_), .Y(u2__abc_44228_n6916) );
  INVX1 INVX1_1723 ( .A(u2_remHi_438_), .Y(u2__abc_44228_n6918) );
  INVX1 INVX1_1724 ( .A(u2__abc_44228_n6920), .Y(u2__abc_44228_n6921) );
  INVX1 INVX1_1725 ( .A(u2_o_437_), .Y(u2__abc_44228_n6925) );
  INVX1 INVX1_1726 ( .A(u2__abc_44228_n6926), .Y(u2__abc_44228_n6927) );
  INVX1 INVX1_1727 ( .A(u2_remHi_437_), .Y(u2__abc_44228_n6928) );
  INVX1 INVX1_1728 ( .A(u2__abc_44228_n6929), .Y(u2__abc_44228_n6930) );
  INVX1 INVX1_1729 ( .A(u2_o_436_), .Y(u2__abc_44228_n6932) );
  INVX1 INVX1_173 ( .A(u2__abc_44228_n2987_bF_buf12), .Y(u2__abc_44228_n3010) );
  INVX1 INVX1_1730 ( .A(u2_remHi_436_), .Y(u2__abc_44228_n6934_1) );
  INVX1 INVX1_1731 ( .A(u2__abc_44228_n6936), .Y(u2__abc_44228_n6937) );
  INVX1 INVX1_1732 ( .A(u2_o_434_), .Y(u2__abc_44228_n6939) );
  INVX1 INVX1_1733 ( .A(u2_remHi_434_), .Y(u2__abc_44228_n6941) );
  INVX1 INVX1_1734 ( .A(u2__abc_44228_n6943_1), .Y(u2__abc_44228_n6944) );
  INVX1 INVX1_1735 ( .A(u2_o_435_), .Y(u2__abc_44228_n6945) );
  INVX1 INVX1_1736 ( .A(u2__abc_44228_n6946), .Y(u2__abc_44228_n6947) );
  INVX1 INVX1_1737 ( .A(u2_remHi_435_), .Y(u2__abc_44228_n6948) );
  INVX1 INVX1_1738 ( .A(u2__abc_44228_n6949), .Y(u2__abc_44228_n6950) );
  INVX1 INVX1_1739 ( .A(u2_o_431_), .Y(u2__abc_44228_n6954) );
  INVX1 INVX1_174 ( .A(u2__abc_44228_n3011), .Y(u2__abc_44228_n3012) );
  INVX1 INVX1_1740 ( .A(u2__abc_44228_n6955), .Y(u2__abc_44228_n6956) );
  INVX1 INVX1_1741 ( .A(u2_remHi_431_), .Y(u2__abc_44228_n6957) );
  INVX1 INVX1_1742 ( .A(u2__abc_44228_n6958), .Y(u2__abc_44228_n6959) );
  INVX1 INVX1_1743 ( .A(u2_o_430_), .Y(u2__abc_44228_n6961_1) );
  INVX1 INVX1_1744 ( .A(u2_remHi_430_), .Y(u2__abc_44228_n6963) );
  INVX1 INVX1_1745 ( .A(u2__abc_44228_n6965), .Y(u2__abc_44228_n6966) );
  INVX1 INVX1_1746 ( .A(u2_o_433_), .Y(u2__abc_44228_n6968) );
  INVX1 INVX1_1747 ( .A(u2__abc_44228_n6969), .Y(u2__abc_44228_n6970) );
  INVX1 INVX1_1748 ( .A(u2_remHi_433_), .Y(u2__abc_44228_n6971_1) );
  INVX1 INVX1_1749 ( .A(u2__abc_44228_n6972), .Y(u2__abc_44228_n6973) );
  INVX1 INVX1_175 ( .A(u2__abc_44228_n3020), .Y(u2__abc_44228_n3021) );
  INVX1 INVX1_1750 ( .A(u2_o_432_), .Y(u2__abc_44228_n6975) );
  INVX1 INVX1_1751 ( .A(u2_remHi_432_), .Y(u2__abc_44228_n6977) );
  INVX1 INVX1_1752 ( .A(u2__abc_44228_n6979_1), .Y(u2__abc_44228_n6980) );
  INVX1 INVX1_1753 ( .A(u2_o_429_), .Y(u2__abc_44228_n6985) );
  INVX1 INVX1_1754 ( .A(u2__abc_44228_n6986), .Y(u2__abc_44228_n6987) );
  INVX1 INVX1_1755 ( .A(u2_remHi_429_), .Y(u2__abc_44228_n6988_1) );
  INVX1 INVX1_1756 ( .A(u2__abc_44228_n6989), .Y(u2__abc_44228_n6990) );
  INVX1 INVX1_1757 ( .A(u2_o_428_), .Y(u2__abc_44228_n6992) );
  INVX1 INVX1_1758 ( .A(u2_remHi_428_), .Y(u2__abc_44228_n6994) );
  INVX1 INVX1_1759 ( .A(u2__abc_44228_n6996), .Y(u2__abc_44228_n6997_1) );
  INVX1 INVX1_176 ( .A(u2__abc_44228_n3026), .Y(u2__abc_44228_n3027) );
  INVX1 INVX1_1760 ( .A(u2_o_427_), .Y(u2__abc_44228_n6999) );
  INVX1 INVX1_1761 ( .A(u2__abc_44228_n7000), .Y(u2__abc_44228_n7001) );
  INVX1 INVX1_1762 ( .A(u2_remHi_427_), .Y(u2__abc_44228_n7002) );
  INVX1 INVX1_1763 ( .A(u2__abc_44228_n7003), .Y(u2__abc_44228_n7004) );
  INVX1 INVX1_1764 ( .A(u2_o_426_), .Y(u2__abc_44228_n7006) );
  INVX1 INVX1_1765 ( .A(u2_remHi_426_), .Y(u2__abc_44228_n7008) );
  INVX1 INVX1_1766 ( .A(u2__abc_44228_n7010), .Y(u2__abc_44228_n7011) );
  INVX1 INVX1_1767 ( .A(u2_o_425_), .Y(u2__abc_44228_n7014_1) );
  INVX1 INVX1_1768 ( .A(u2__abc_44228_n7015), .Y(u2__abc_44228_n7016) );
  INVX1 INVX1_1769 ( .A(u2_remHi_425_), .Y(u2__abc_44228_n7017) );
  INVX1 INVX1_177 ( .A(u2__abc_44228_n3034), .Y(u2__abc_44228_n3035) );
  INVX1 INVX1_1770 ( .A(u2__abc_44228_n7018), .Y(u2__abc_44228_n7019) );
  INVX1 INVX1_1771 ( .A(u2_o_424_), .Y(u2__abc_44228_n7021) );
  INVX1 INVX1_1772 ( .A(u2_remHi_424_), .Y(u2__abc_44228_n7023) );
  INVX1 INVX1_1773 ( .A(u2__abc_44228_n7025), .Y(u2__abc_44228_n7026) );
  INVX1 INVX1_1774 ( .A(u2_o_423_), .Y(u2__abc_44228_n7028) );
  INVX1 INVX1_1775 ( .A(u2__abc_44228_n7029), .Y(u2__abc_44228_n7030) );
  INVX1 INVX1_1776 ( .A(u2_remHi_423_), .Y(u2__abc_44228_n7031) );
  INVX1 INVX1_1777 ( .A(u2__abc_44228_n7032_1), .Y(u2__abc_44228_n7033) );
  INVX1 INVX1_1778 ( .A(u2_o_422_), .Y(u2__abc_44228_n7035) );
  INVX1 INVX1_1779 ( .A(u2_remHi_422_), .Y(u2__abc_44228_n7037) );
  INVX1 INVX1_178 ( .A(u2__abc_44228_n3042), .Y(u2__abc_44228_n3043) );
  INVX1 INVX1_1780 ( .A(u2__abc_44228_n7039), .Y(u2__abc_44228_n7040) );
  INVX1 INVX1_1781 ( .A(u2_o_421_), .Y(u2__abc_44228_n7044) );
  INVX1 INVX1_1782 ( .A(u2__abc_44228_n7045), .Y(u2__abc_44228_n7046) );
  INVX1 INVX1_1783 ( .A(u2_remHi_421_), .Y(u2__abc_44228_n7047) );
  INVX1 INVX1_1784 ( .A(u2__abc_44228_n7048), .Y(u2__abc_44228_n7049) );
  INVX1 INVX1_1785 ( .A(u2_o_420_), .Y(u2__abc_44228_n7051) );
  INVX1 INVX1_1786 ( .A(u2_remHi_420_), .Y(u2__abc_44228_n7053) );
  INVX1 INVX1_1787 ( .A(u2__abc_44228_n7055), .Y(u2__abc_44228_n7056) );
  INVX1 INVX1_1788 ( .A(u2_o_419_), .Y(u2__abc_44228_n7058) );
  INVX1 INVX1_1789 ( .A(u2__abc_44228_n7059_1), .Y(u2__abc_44228_n7060) );
  INVX1 INVX1_179 ( .A(u2__abc_44228_n2989_bF_buf2), .Y(u2__abc_44228_n3047) );
  INVX1 INVX1_1790 ( .A(u2_remHi_419_), .Y(u2__abc_44228_n7061) );
  INVX1 INVX1_1791 ( .A(u2__abc_44228_n7062), .Y(u2__abc_44228_n7063) );
  INVX1 INVX1_1792 ( .A(u2_o_418_), .Y(u2__abc_44228_n7065) );
  INVX1 INVX1_1793 ( .A(u2_remHi_418_), .Y(u2__abc_44228_n7067) );
  INVX1 INVX1_1794 ( .A(u2__abc_44228_n7069), .Y(u2__abc_44228_n7070) );
  INVX1 INVX1_1795 ( .A(u2_o_417_), .Y(u2__abc_44228_n7073) );
  INVX1 INVX1_1796 ( .A(u2__abc_44228_n7074), .Y(u2__abc_44228_n7075) );
  INVX1 INVX1_1797 ( .A(u2_remHi_417_), .Y(u2__abc_44228_n7076) );
  INVX1 INVX1_1798 ( .A(u2__abc_44228_n7077), .Y(u2__abc_44228_n7078_1) );
  INVX1 INVX1_1799 ( .A(u2_o_416_), .Y(u2__abc_44228_n7080) );
  INVX1 INVX1_18 ( .A(_abc_64468_n1570), .Y(_abc_64468_n1571) );
  INVX1 INVX1_180 ( .A(u2__abc_44228_n3050), .Y(u2__abc_44228_n3051) );
  INVX1 INVX1_1800 ( .A(u2_remHi_416_), .Y(u2__abc_44228_n7082) );
  INVX1 INVX1_1801 ( .A(u2__abc_44228_n7084), .Y(u2__abc_44228_n7085) );
  INVX1 INVX1_1802 ( .A(u2_o_414_), .Y(u2__abc_44228_n7087) );
  INVX1 INVX1_1803 ( .A(u2_remHi_414_), .Y(u2__abc_44228_n7089) );
  INVX1 INVX1_1804 ( .A(u2__abc_44228_n7091), .Y(u2__abc_44228_n7092) );
  INVX1 INVX1_1805 ( .A(u2_o_415_), .Y(u2__abc_44228_n7093) );
  INVX1 INVX1_1806 ( .A(u2__abc_44228_n7094), .Y(u2__abc_44228_n7095) );
  INVX1 INVX1_1807 ( .A(u2_remHi_415_), .Y(u2__abc_44228_n7096) );
  INVX1 INVX1_1808 ( .A(u2__abc_44228_n7097), .Y(u2__abc_44228_n7098_1) );
  INVX1 INVX1_1809 ( .A(u2_o_413_), .Y(u2__abc_44228_n7105) );
  INVX1 INVX1_181 ( .A(u2_cnt_7_), .Y(u2__abc_44228_n3053) );
  INVX1 INVX1_1810 ( .A(u2__abc_44228_n7106_1), .Y(u2__abc_44228_n7107) );
  INVX1 INVX1_1811 ( .A(u2_remHi_413_), .Y(u2__abc_44228_n7108) );
  INVX1 INVX1_1812 ( .A(u2__abc_44228_n7109), .Y(u2__abc_44228_n7110) );
  INVX1 INVX1_1813 ( .A(u2_o_412_), .Y(u2__abc_44228_n7112) );
  INVX1 INVX1_1814 ( .A(u2_remHi_412_), .Y(u2__abc_44228_n7114) );
  INVX1 INVX1_1815 ( .A(u2__abc_44228_n7116_1), .Y(u2__abc_44228_n7117) );
  INVX1 INVX1_1816 ( .A(u2_o_411_), .Y(u2__abc_44228_n7119) );
  INVX1 INVX1_1817 ( .A(u2__abc_44228_n7120), .Y(u2__abc_44228_n7121) );
  INVX1 INVX1_1818 ( .A(u2_remHi_411_), .Y(u2__abc_44228_n7122) );
  INVX1 INVX1_1819 ( .A(u2__abc_44228_n7123), .Y(u2__abc_44228_n7124) );
  INVX1 INVX1_182 ( .A(u2__abc_44228_n2972_bF_buf106), .Y(u2__abc_44228_n3058) );
  INVX1 INVX1_1820 ( .A(u2_o_410_), .Y(u2__abc_44228_n7126) );
  INVX1 INVX1_1821 ( .A(u2_remHi_410_), .Y(u2__abc_44228_n7128) );
  INVX1 INVX1_1822 ( .A(u2__abc_44228_n7130), .Y(u2__abc_44228_n7131) );
  INVX1 INVX1_1823 ( .A(u2_o_409_), .Y(u2__abc_44228_n7134_1) );
  INVX1 INVX1_1824 ( .A(u2__abc_44228_n7135), .Y(u2__abc_44228_n7136) );
  INVX1 INVX1_1825 ( .A(u2_remHi_409_), .Y(u2__abc_44228_n7137) );
  INVX1 INVX1_1826 ( .A(u2__abc_44228_n7138), .Y(u2__abc_44228_n7139) );
  INVX1 INVX1_1827 ( .A(u2_o_408_), .Y(u2__abc_44228_n7141) );
  INVX1 INVX1_1828 ( .A(u2_remHi_408_), .Y(u2__abc_44228_n7143_1) );
  INVX1 INVX1_1829 ( .A(u2__abc_44228_n7145), .Y(u2__abc_44228_n7146) );
  INVX1 INVX1_183 ( .A(u2__abc_44228_n3059), .Y(u2__abc_44228_n3060) );
  INVX1 INVX1_1830 ( .A(u2_o_407_), .Y(u2__abc_44228_n7148) );
  INVX1 INVX1_1831 ( .A(u2__abc_44228_n7149), .Y(u2__abc_44228_n7150) );
  INVX1 INVX1_1832 ( .A(u2_remHi_407_), .Y(u2__abc_44228_n7151) );
  INVX1 INVX1_1833 ( .A(u2__abc_44228_n7152), .Y(u2__abc_44228_n7153_1) );
  INVX1 INVX1_1834 ( .A(u2_o_406_), .Y(u2__abc_44228_n7155) );
  INVX1 INVX1_1835 ( .A(u2_remHi_406_), .Y(u2__abc_44228_n7157) );
  INVX1 INVX1_1836 ( .A(u2__abc_44228_n7159), .Y(u2__abc_44228_n7160) );
  INVX1 INVX1_1837 ( .A(u2_o_405_), .Y(u2__abc_44228_n7164) );
  INVX1 INVX1_1838 ( .A(u2__abc_44228_n7165), .Y(u2__abc_44228_n7166) );
  INVX1 INVX1_1839 ( .A(u2_remHi_405_), .Y(u2__abc_44228_n7167) );
  INVX1 INVX1_184 ( .A(u2_remHiShift_1_), .Y(u2__abc_44228_n3064) );
  INVX1 INVX1_1840 ( .A(u2__abc_44228_n7168), .Y(u2__abc_44228_n7169) );
  INVX1 INVX1_1841 ( .A(u2_o_404_), .Y(u2__abc_44228_n7171) );
  INVX1 INVX1_1842 ( .A(u2_remHi_404_), .Y(u2__abc_44228_n7173) );
  INVX1 INVX1_1843 ( .A(u2__abc_44228_n7175), .Y(u2__abc_44228_n7176) );
  INVX1 INVX1_1844 ( .A(u2_o_403_), .Y(u2__abc_44228_n7178) );
  INVX1 INVX1_1845 ( .A(u2__abc_44228_n7179_1), .Y(u2__abc_44228_n7180) );
  INVX1 INVX1_1846 ( .A(u2_remHi_403_), .Y(u2__abc_44228_n7181) );
  INVX1 INVX1_1847 ( .A(u2__abc_44228_n7182), .Y(u2__abc_44228_n7183) );
  INVX1 INVX1_1848 ( .A(u2_o_402_), .Y(u2__abc_44228_n7185) );
  INVX1 INVX1_1849 ( .A(u2_remHi_402_), .Y(u2__abc_44228_n7187) );
  INVX1 INVX1_185 ( .A(u2__abc_44228_n3065), .Y(u2__abc_44228_n3066) );
  INVX1 INVX1_1850 ( .A(u2__abc_44228_n7189_1), .Y(u2__abc_44228_n7190) );
  INVX1 INVX1_1851 ( .A(u2_o_401_), .Y(u2__abc_44228_n7193) );
  INVX1 INVX1_1852 ( .A(u2__abc_44228_n7194), .Y(u2__abc_44228_n7195) );
  INVX1 INVX1_1853 ( .A(u2_remHi_401_), .Y(u2__abc_44228_n7196) );
  INVX1 INVX1_1854 ( .A(u2__abc_44228_n7197_1), .Y(u2__abc_44228_n7198) );
  INVX1 INVX1_1855 ( .A(u2_o_400_), .Y(u2__abc_44228_n7200) );
  INVX1 INVX1_1856 ( .A(u2_remHi_400_), .Y(u2__abc_44228_n7202) );
  INVX1 INVX1_1857 ( .A(u2__abc_44228_n7204), .Y(u2__abc_44228_n7205) );
  INVX1 INVX1_1858 ( .A(u2_o_398_), .Y(u2__abc_44228_n7207) );
  INVX1 INVX1_1859 ( .A(u2_remHi_398_), .Y(u2__abc_44228_n7209) );
  INVX1 INVX1_186 ( .A(u2_root_0_), .Y(u2__abc_44228_n3067) );
  INVX1 INVX1_1860 ( .A(u2__abc_44228_n7211), .Y(u2__abc_44228_n7212) );
  INVX1 INVX1_1861 ( .A(u2_o_399_), .Y(u2__abc_44228_n7213) );
  INVX1 INVX1_1862 ( .A(u2__abc_44228_n7214), .Y(u2__abc_44228_n7215_1) );
  INVX1 INVX1_1863 ( .A(u2_remHi_399_), .Y(u2__abc_44228_n7216) );
  INVX1 INVX1_1864 ( .A(u2__abc_44228_n7217), .Y(u2__abc_44228_n7218) );
  INVX1 INVX1_1865 ( .A(u2_o_397_), .Y(u2__abc_44228_n7224) );
  INVX1 INVX1_1866 ( .A(u2__abc_44228_n7225_1), .Y(u2__abc_44228_n7226) );
  INVX1 INVX1_1867 ( .A(u2_remHi_397_), .Y(u2__abc_44228_n7227) );
  INVX1 INVX1_1868 ( .A(u2__abc_44228_n7228), .Y(u2__abc_44228_n7229) );
  INVX1 INVX1_1869 ( .A(u2_o_396_), .Y(u2__abc_44228_n7231) );
  INVX1 INVX1_187 ( .A(u2_remHi_1_), .Y(u2__abc_44228_n3072) );
  INVX1 INVX1_1870 ( .A(u2_remHi_396_), .Y(u2__abc_44228_n7233) );
  INVX1 INVX1_1871 ( .A(u2__abc_44228_n7235), .Y(u2__abc_44228_n7236) );
  INVX1 INVX1_1872 ( .A(u2_o_394_), .Y(u2__abc_44228_n7238) );
  INVX1 INVX1_1873 ( .A(u2_remHi_394_), .Y(u2__abc_44228_n7240) );
  INVX1 INVX1_1874 ( .A(u2__abc_44228_n7242), .Y(u2__abc_44228_n7243) );
  INVX1 INVX1_1875 ( .A(u2_o_395_), .Y(u2__abc_44228_n7244_1) );
  INVX1 INVX1_1876 ( .A(u2__abc_44228_n7245), .Y(u2__abc_44228_n7246) );
  INVX1 INVX1_1877 ( .A(u2_remHi_395_), .Y(u2__abc_44228_n7247) );
  INVX1 INVX1_1878 ( .A(u2__abc_44228_n7248), .Y(u2__abc_44228_n7249) );
  INVX1 INVX1_1879 ( .A(u2_o_393_), .Y(u2__abc_44228_n7253) );
  INVX1 INVX1_188 ( .A(sqrto_1_), .Y(u2__abc_44228_n3074) );
  INVX1 INVX1_1880 ( .A(u2__abc_44228_n7254), .Y(u2__abc_44228_n7255) );
  INVX1 INVX1_1881 ( .A(u2_remHi_393_), .Y(u2__abc_44228_n7256) );
  INVX1 INVX1_1882 ( .A(u2__abc_44228_n7257), .Y(u2__abc_44228_n7258) );
  INVX1 INVX1_1883 ( .A(u2_o_392_), .Y(u2__abc_44228_n7260) );
  INVX1 INVX1_1884 ( .A(u2_remHi_392_), .Y(u2__abc_44228_n7262_1) );
  INVX1 INVX1_1885 ( .A(u2__abc_44228_n7264), .Y(u2__abc_44228_n7265) );
  INVX1 INVX1_1886 ( .A(u2_o_390_), .Y(u2__abc_44228_n7267) );
  INVX1 INVX1_1887 ( .A(u2_remHi_390_), .Y(u2__abc_44228_n7269) );
  INVX1 INVX1_1888 ( .A(u2__abc_44228_n7271_1), .Y(u2__abc_44228_n7272) );
  INVX1 INVX1_1889 ( .A(u2_o_391_), .Y(u2__abc_44228_n7273) );
  INVX1 INVX1_189 ( .A(sqrto_0_), .Y(u2__abc_44228_n3077) );
  INVX1 INVX1_1890 ( .A(u2__abc_44228_n7274), .Y(u2__abc_44228_n7275) );
  INVX1 INVX1_1891 ( .A(u2_remHi_391_), .Y(u2__abc_44228_n7276) );
  INVX1 INVX1_1892 ( .A(u2__abc_44228_n7277), .Y(u2__abc_44228_n7278) );
  INVX1 INVX1_1893 ( .A(u2_o_389_), .Y(u2__abc_44228_n7283) );
  INVX1 INVX1_1894 ( .A(u2__abc_44228_n7284), .Y(u2__abc_44228_n7285) );
  INVX1 INVX1_1895 ( .A(u2_remHi_389_), .Y(u2__abc_44228_n7286) );
  INVX1 INVX1_1896 ( .A(u2__abc_44228_n7287), .Y(u2__abc_44228_n7288) );
  INVX1 INVX1_1897 ( .A(u2_o_388_), .Y(u2__abc_44228_n7290) );
  INVX1 INVX1_1898 ( .A(u2_remHi_388_), .Y(u2__abc_44228_n7292) );
  INVX1 INVX1_1899 ( .A(u2__abc_44228_n7294), .Y(u2__abc_44228_n7295) );
  INVX1 INVX1_19 ( .A(_abc_64468_n1572), .Y(_abc_64468_n1573) );
  INVX1 INVX1_190 ( .A(u2__abc_44228_n3078), .Y(u2__abc_44228_n3079) );
  INVX1 INVX1_1900 ( .A(u2_o_386_), .Y(u2__abc_44228_n7297) );
  INVX1 INVX1_1901 ( .A(u2_remHi_386_), .Y(u2__abc_44228_n7299_1) );
  INVX1 INVX1_1902 ( .A(u2__abc_44228_n7301), .Y(u2__abc_44228_n7302) );
  INVX1 INVX1_1903 ( .A(u2_o_387_), .Y(u2__abc_44228_n7303) );
  INVX1 INVX1_1904 ( .A(u2__abc_44228_n7304), .Y(u2__abc_44228_n7305) );
  INVX1 INVX1_1905 ( .A(u2_remHi_387_), .Y(u2__abc_44228_n7306) );
  INVX1 INVX1_1906 ( .A(u2__abc_44228_n7307), .Y(u2__abc_44228_n7308) );
  INVX1 INVX1_1907 ( .A(u2_o_385_), .Y(u2__abc_44228_n7312) );
  INVX1 INVX1_1908 ( .A(u2__abc_44228_n7313), .Y(u2__abc_44228_n7314) );
  INVX1 INVX1_1909 ( .A(u2_remHi_385_), .Y(u2__abc_44228_n7315) );
  INVX1 INVX1_191 ( .A(u2__abc_44228_n3073), .Y(u2__abc_44228_n3084) );
  INVX1 INVX1_1910 ( .A(u2__abc_44228_n7316), .Y(u2__abc_44228_n7317) );
  INVX1 INVX1_1911 ( .A(u2_o_384_), .Y(u2__abc_44228_n7319_1) );
  INVX1 INVX1_1912 ( .A(u2_remHi_384_), .Y(u2__abc_44228_n7321) );
  INVX1 INVX1_1913 ( .A(u2__abc_44228_n7323), .Y(u2__abc_44228_n7324) );
  INVX1 INVX1_1914 ( .A(u2_o_383_), .Y(u2__abc_44228_n7326) );
  INVX1 INVX1_1915 ( .A(u2__abc_44228_n7327_1), .Y(u2__abc_44228_n7328) );
  INVX1 INVX1_1916 ( .A(u2_remHi_383_), .Y(u2__abc_44228_n7329) );
  INVX1 INVX1_1917 ( .A(u2__abc_44228_n7330), .Y(u2__abc_44228_n7331) );
  INVX1 INVX1_1918 ( .A(u2_o_382_), .Y(u2__abc_44228_n7333) );
  INVX1 INVX1_1919 ( .A(u2_remHi_382_), .Y(u2__abc_44228_n7335) );
  INVX1 INVX1_192 ( .A(u2_remHi_5_), .Y(u2__abc_44228_n3088) );
  INVX1 INVX1_1920 ( .A(u2__abc_44228_n7337_1), .Y(u2__abc_44228_n7338) );
  INVX1 INVX1_1921 ( .A(u2__abc_44228_n7334), .Y(u2__abc_44228_n7346_1) );
  INVX1 INVX1_1922 ( .A(u2__abc_44228_n7348), .Y(u2__abc_44228_n7349) );
  INVX1 INVX1_1923 ( .A(u2__abc_44228_n7298), .Y(u2__abc_44228_n7355_1) );
  INVX1 INVX1_1924 ( .A(u2__abc_44228_n7356), .Y(u2__abc_44228_n7357) );
  INVX1 INVX1_1925 ( .A(u2__abc_44228_n7268), .Y(u2__abc_44228_n7365) );
  INVX1 INVX1_1926 ( .A(u2__abc_44228_n7366), .Y(u2__abc_44228_n7367) );
  INVX1 INVX1_1927 ( .A(u2__abc_44228_n7239), .Y(u2__abc_44228_n7376) );
  INVX1 INVX1_1928 ( .A(u2__abc_44228_n7377), .Y(u2__abc_44228_n7378) );
  INVX1 INVX1_1929 ( .A(u2__abc_44228_n7208), .Y(u2__abc_44228_n7385) );
  INVX1 INVX1_193 ( .A(sqrto_5_), .Y(u2__abc_44228_n3090) );
  INVX1 INVX1_1930 ( .A(u2__abc_44228_n7386), .Y(u2__abc_44228_n7387) );
  INVX1 INVX1_1931 ( .A(u2__abc_44228_n7186), .Y(u2__abc_44228_n7394) );
  INVX1 INVX1_1932 ( .A(u2__abc_44228_n7396), .Y(u2__abc_44228_n7397) );
  INVX1 INVX1_1933 ( .A(u2__abc_44228_n7156), .Y(u2__abc_44228_n7406) );
  INVX1 INVX1_1934 ( .A(u2__abc_44228_n7407), .Y(u2__abc_44228_n7408) );
  INVX1 INVX1_1935 ( .A(u2__abc_44228_n7127), .Y(u2__abc_44228_n7413) );
  INVX1 INVX1_1936 ( .A(u2__abc_44228_n7414), .Y(u2__abc_44228_n7415) );
  INVX1 INVX1_1937 ( .A(u2__abc_44228_n7088_1), .Y(u2__abc_44228_n7425) );
  INVX1 INVX1_1938 ( .A(u2__abc_44228_n7426), .Y(u2__abc_44228_n7427) );
  INVX1 INVX1_1939 ( .A(u2__abc_44228_n7066), .Y(u2__abc_44228_n7434) );
  INVX1 INVX1_194 ( .A(u2_remHi_4_), .Y(u2__abc_44228_n3093) );
  INVX1 INVX1_1940 ( .A(u2__abc_44228_n7436), .Y(u2__abc_44228_n7437_1) );
  INVX1 INVX1_1941 ( .A(u2__abc_44228_n7036), .Y(u2__abc_44228_n7444) );
  INVX1 INVX1_1942 ( .A(u2__abc_44228_n7446), .Y(u2__abc_44228_n7447_1) );
  INVX1 INVX1_1943 ( .A(u2__abc_44228_n7022_1), .Y(u2__abc_44228_n7449) );
  INVX1 INVX1_1944 ( .A(u2__abc_44228_n7450), .Y(u2__abc_44228_n7451) );
  INVX1 INVX1_1945 ( .A(u2__abc_44228_n7007_1), .Y(u2__abc_44228_n7457) );
  INVX1 INVX1_1946 ( .A(u2__abc_44228_n7458), .Y(u2__abc_44228_n7459) );
  INVX1 INVX1_1947 ( .A(u2__abc_44228_n6962), .Y(u2__abc_44228_n7466) );
  INVX1 INVX1_1948 ( .A(u2__abc_44228_n7468), .Y(u2__abc_44228_n7469) );
  INVX1 INVX1_1949 ( .A(u2__abc_44228_n6976), .Y(u2__abc_44228_n7471) );
  INVX1 INVX1_195 ( .A(sqrto_4_), .Y(u2__abc_44228_n3095) );
  INVX1 INVX1_1950 ( .A(u2__abc_44228_n7472), .Y(u2__abc_44228_n7473_1) );
  INVX1 INVX1_1951 ( .A(u2__abc_44228_n6940), .Y(u2__abc_44228_n7477) );
  INVX1 INVX1_1952 ( .A(u2__abc_44228_n7478), .Y(u2__abc_44228_n7479) );
  INVX1 INVX1_1953 ( .A(u2__abc_44228_n6917), .Y(u2__abc_44228_n7489) );
  INVX1 INVX1_1954 ( .A(u2__abc_44228_n7490), .Y(u2__abc_44228_n7491) );
  INVX1 INVX1_1955 ( .A(u2__abc_44228_n6888), .Y(u2__abc_44228_n7496) );
  INVX1 INVX1_1956 ( .A(u2__abc_44228_n7498), .Y(u2__abc_44228_n7499) );
  INVX1 INVX1_1957 ( .A(u2_o_449_), .Y(u2__abc_44228_n7509) );
  INVX1 INVX1_1958 ( .A(u2__abc_44228_n7510), .Y(u2__abc_44228_n7511_1) );
  INVX1 INVX1_1959 ( .A(u2_remHi_449_), .Y(u2__abc_44228_n7512) );
  INVX1 INVX1_196 ( .A(sqrto_3_), .Y(u2__abc_44228_n3099) );
  INVX1 INVX1_1960 ( .A(u2__abc_44228_n7513), .Y(u2__abc_44228_n7514) );
  INVX1 INVX1_1961 ( .A(u2_o_448_), .Y(u2__abc_44228_n7516) );
  INVX1 INVX1_1962 ( .A(u2_remHi_448_), .Y(u2__abc_44228_n7518) );
  INVX1 INVX1_1963 ( .A(u2__abc_44228_n7520), .Y(u2__abc_44228_n7521_1) );
  INVX1 INVX1_1964 ( .A(u2_o_446_), .Y(u2__abc_44228_n7523) );
  INVX1 INVX1_1965 ( .A(u2_remHi_446_), .Y(u2__abc_44228_n7525) );
  INVX1 INVX1_1966 ( .A(u2__abc_44228_n7527), .Y(u2__abc_44228_n7528) );
  INVX1 INVX1_1967 ( .A(u2_o_447_), .Y(u2__abc_44228_n7529) );
  INVX1 INVX1_1968 ( .A(u2__abc_44228_n7530_1), .Y(u2__abc_44228_n7531) );
  INVX1 INVX1_1969 ( .A(u2_remHi_447_), .Y(u2__abc_44228_n7532) );
  INVX1 INVX1_197 ( .A(u2__abc_44228_n3100), .Y(u2__abc_44228_n3101) );
  INVX1 INVX1_1970 ( .A(u2__abc_44228_n7533), .Y(u2__abc_44228_n7534) );
  INVX1 INVX1_1971 ( .A(u2__abc_44228_n7524), .Y(u2__abc_44228_n7539) );
  INVX1 INVX1_1972 ( .A(u2__abc_44228_n7541), .Y(u2__abc_44228_n7542) );
  INVX1 INVX1_1973 ( .A(u2_remHiShift_0_), .Y(u2__abc_44228_n7550) );
  INVX1 INVX1_1974 ( .A(u2_remHi_0_), .Y(u2__abc_44228_n7554) );
  INVX1 INVX1_1975 ( .A(u2__abc_44228_n7555), .Y(u2__abc_44228_n7556) );
  INVX1 INVX1_1976 ( .A(u2__abc_44228_n3070), .Y(u2__abc_44228_n7562) );
  INVX1 INVX1_1977 ( .A(u2__abc_44228_n7569), .Y(u2__abc_44228_n7570) );
  INVX1 INVX1_1978 ( .A(u2__abc_44228_n7576_1), .Y(u2__abc_44228_n7577) );
  INVX1 INVX1_1979 ( .A(u2_remHi_2_), .Y(u2__abc_44228_n7584) );
  INVX1 INVX1_198 ( .A(sqrto_2_), .Y(u2__abc_44228_n3104) );
  INVX1 INVX1_1980 ( .A(u2__abc_44228_n7585), .Y(u2__abc_44228_n7586_1) );
  INVX1 INVX1_1981 ( .A(u2__abc_44228_n7592), .Y(u2__abc_44228_n7593) );
  INVX1 INVX1_1982 ( .A(u2__abc_44228_n3076), .Y(u2__abc_44228_n7595) );
  INVX1 INVX1_1983 ( .A(u2_remHi_3_), .Y(u2__abc_44228_n7602) );
  INVX1 INVX1_1984 ( .A(u2__abc_44228_n7603), .Y(u2__abc_44228_n7604) );
  INVX1 INVX1_1985 ( .A(u2__abc_44228_n7611), .Y(u2__abc_44228_n7612) );
  INVX1 INVX1_1986 ( .A(u2__abc_44228_n7618), .Y(u2__abc_44228_n7619) );
  INVX1 INVX1_1987 ( .A(u2__abc_44228_n3103), .Y(u2__abc_44228_n7625) );
  INVX1 INVX1_1988 ( .A(u2__abc_44228_n7626), .Y(u2__abc_44228_n7628) );
  INVX1 INVX1_1989 ( .A(u2__abc_44228_n7635), .Y(u2__abc_44228_n7636_1) );
  INVX1 INVX1_199 ( .A(u2__abc_44228_n3105), .Y(u2__abc_44228_n3106) );
  INVX1 INVX1_1990 ( .A(u2__abc_44228_n7644_1), .Y(u2__abc_44228_n7645) );
  INVX1 INVX1_1991 ( .A(u2__abc_44228_n7652), .Y(u2__abc_44228_n7653) );
  INVX1 INVX1_1992 ( .A(u2__abc_44228_n7659), .Y(u2__abc_44228_n7660) );
  INVX1 INVX1_1993 ( .A(u2__abc_44228_n3092), .Y(u2__abc_44228_n7662) );
  INVX1 INVX1_1994 ( .A(u2__abc_44228_n7669), .Y(u2__abc_44228_n7670) );
  INVX1 INVX1_1995 ( .A(u2__abc_44228_n7676), .Y(u2__abc_44228_n7677) );
  INVX1 INVX1_1996 ( .A(u2__abc_44228_n7684), .Y(u2__abc_44228_n7685_1) );
  INVX1 INVX1_1997 ( .A(u2__abc_44228_n3173), .Y(u2__abc_44228_n7691) );
  INVX1 INVX1_1998 ( .A(u2__abc_44228_n7692_1), .Y(u2__abc_44228_n7694) );
  INVX1 INVX1_1999 ( .A(u2__abc_44228_n7701), .Y(u2__abc_44228_n7702) );
  INVX1 INVX1_2 ( .A(_abc_64468_n1514), .Y(_abc_64468_n1515) );
  INVX1 INVX1_20 ( .A(_abc_64468_n1575), .Y(_abc_64468_n1579) );
  INVX1 INVX1_200 ( .A(u2__abc_44228_n3089), .Y(u2__abc_44228_n3115) );
  INVX1 INVX1_2000 ( .A(u2__abc_44228_n7711), .Y(u2__abc_44228_n7712) );
  INVX1 INVX1_2001 ( .A(u2__abc_44228_n7718), .Y(u2__abc_44228_n7719) );
  INVX1 INVX1_2002 ( .A(u2__abc_44228_n7725), .Y(u2__abc_44228_n7726) );
  INVX1 INVX1_2003 ( .A(u2__abc_44228_n3154), .Y(u2__abc_44228_n7728_1) );
  INVX1 INVX1_2004 ( .A(u2__abc_44228_n7735_1), .Y(u2__abc_44228_n7736) );
  INVX1 INVX1_2005 ( .A(u2__abc_44228_n7744), .Y(u2__abc_44228_n7745) );
  INVX1 INVX1_2006 ( .A(u2__abc_44228_n7752), .Y(u2__abc_44228_n7753) );
  INVX1 INVX1_2007 ( .A(u2__abc_44228_n3141), .Y(u2__abc_44228_n7761) );
  INVX1 INVX1_2008 ( .A(u2__abc_44228_n7759), .Y(u2__abc_44228_n7762_1) );
  INVX1 INVX1_2009 ( .A(u2__abc_44228_n7769_1), .Y(u2__abc_44228_n7770_1) );
  INVX1 INVX1_201 ( .A(u2__abc_44228_n3094), .Y(u2__abc_44228_n3116) );
  INVX1 INVX1_2010 ( .A(u2__abc_44228_n7779), .Y(u2__abc_44228_n7780) );
  INVX1 INVX1_2011 ( .A(u2__abc_44228_n7786), .Y(u2__abc_44228_n7787) );
  INVX1 INVX1_2012 ( .A(u2__abc_44228_n3127), .Y(u2__abc_44228_n7793) );
  INVX1 INVX1_2013 ( .A(u2__abc_44228_n7794), .Y(u2__abc_44228_n7795) );
  INVX1 INVX1_2014 ( .A(u2__abc_44228_n7803), .Y(u2__abc_44228_n7804_1) );
  INVX1 INVX1_2015 ( .A(u2__abc_44228_n7811_1), .Y(u2__abc_44228_n7812_1) );
  INVX1 INVX1_2016 ( .A(u2__abc_44228_n7818_1), .Y(u2__abc_44228_n7819_1) );
  INVX1 INVX1_2017 ( .A(u2__abc_44228_n3300), .Y(u2__abc_44228_n7827) );
  INVX1 INVX1_2018 ( .A(u2__abc_44228_n7825_1), .Y(u2__abc_44228_n7828) );
  INVX1 INVX1_2019 ( .A(u2__abc_44228_n7835), .Y(u2__abc_44228_n7836) );
  INVX1 INVX1_202 ( .A(sqrto_13_), .Y(u2__abc_44228_n3121) );
  INVX1 INVX1_2020 ( .A(u2__abc_44228_n7845_1), .Y(u2__abc_44228_n7846) );
  INVX1 INVX1_2021 ( .A(u2__abc_44228_n7852), .Y(u2__abc_44228_n7853) );
  INVX1 INVX1_2022 ( .A(u2__abc_44228_n7859), .Y(u2__abc_44228_n7860) );
  INVX1 INVX1_2023 ( .A(u2__abc_44228_n3287), .Y(u2__abc_44228_n7862_1) );
  INVX1 INVX1_2024 ( .A(u2__abc_44228_n7869), .Y(u2__abc_44228_n7870) );
  INVX1 INVX1_2025 ( .A(u2__abc_44228_n7878_1), .Y(u2__abc_44228_n7879) );
  INVX1 INVX1_2026 ( .A(u2__abc_44228_n7886), .Y(u2__abc_44228_n7887) );
  INVX1 INVX1_2027 ( .A(u2__abc_44228_n3280), .Y(u2__abc_44228_n7893) );
  INVX1 INVX1_2028 ( .A(u2__abc_44228_n7894_1), .Y(u2__abc_44228_n7896) );
  INVX1 INVX1_2029 ( .A(u2__abc_44228_n7903), .Y(u2__abc_44228_n7904) );
  INVX1 INVX1_203 ( .A(u2__abc_44228_n3122), .Y(u2__abc_44228_n3123) );
  INVX1 INVX1_2030 ( .A(u2__abc_44228_n7913), .Y(u2__abc_44228_n7914) );
  INVX1 INVX1_2031 ( .A(u2__abc_44228_n7920), .Y(u2__abc_44228_n7921) );
  INVX1 INVX1_2032 ( .A(u2__abc_44228_n3260), .Y(u2__abc_44228_n7927_1) );
  INVX1 INVX1_2033 ( .A(u2__abc_44228_n7928_1), .Y(u2__abc_44228_n7930) );
  INVX1 INVX1_2034 ( .A(u2__abc_44228_n7937), .Y(u2__abc_44228_n7938_1) );
  INVX1 INVX1_2035 ( .A(u2__abc_44228_n7947), .Y(u2__abc_44228_n7948) );
  INVX1 INVX1_2036 ( .A(u2__abc_44228_n7954), .Y(u2__abc_44228_n7955_1) );
  INVX1 INVX1_2037 ( .A(u2__abc_44228_n3230), .Y(u2__abc_44228_n7961_1) );
  INVX1 INVX1_2038 ( .A(u2__abc_44228_n7962), .Y(u2__abc_44228_n7963) );
  INVX1 INVX1_2039 ( .A(u2__abc_44228_n7971_1), .Y(u2__abc_44228_n7972_1) );
  INVX1 INVX1_204 ( .A(u2_remHi_13_), .Y(u2__abc_44228_n3124) );
  INVX1 INVX1_2040 ( .A(u2__abc_44228_n7981), .Y(u2__abc_44228_n7982_1) );
  INVX1 INVX1_2041 ( .A(u2__abc_44228_n7988_1), .Y(u2__abc_44228_n7989) );
  INVX1 INVX1_2042 ( .A(u2__abc_44228_n7995), .Y(u2__abc_44228_n7996) );
  INVX1 INVX1_2043 ( .A(u2__abc_44228_n3244), .Y(u2__abc_44228_n7998) );
  INVX1 INVX1_2044 ( .A(u2__abc_44228_n8005_1), .Y(u2__abc_44228_n8006) );
  INVX1 INVX1_2045 ( .A(u2__abc_44228_n8014), .Y(u2__abc_44228_n8015_1) );
  INVX1 INVX1_2046 ( .A(u2__abc_44228_n8016_1), .Y(u2__abc_44228_n8017) );
  INVX1 INVX1_2047 ( .A(u2__abc_44228_n8023), .Y(u2__abc_44228_n8024) );
  INVX1 INVX1_2048 ( .A(u2__abc_44228_n3221), .Y(u2__abc_44228_n8031) );
  INVX1 INVX1_2049 ( .A(u2__abc_44228_n8032_1), .Y(u2__abc_44228_n8033) );
  INVX1 INVX1_205 ( .A(u2__abc_44228_n3125), .Y(u2__abc_44228_n3126) );
  INVX1 INVX1_2050 ( .A(u2__abc_44228_n8040), .Y(u2__abc_44228_n8041) );
  INVX1 INVX1_2051 ( .A(u2__abc_44228_n8048_1), .Y(u2__abc_44228_n8049_1) );
  INVX1 INVX1_2052 ( .A(u2__abc_44228_n8051), .Y(u2__abc_44228_n8052) );
  INVX1 INVX1_2053 ( .A(u2__abc_44228_n8058), .Y(u2__abc_44228_n8059_1) );
  INVX1 INVX1_2054 ( .A(u2__abc_44228_n3201), .Y(u2__abc_44228_n8065_1) );
  INVX1 INVX1_2055 ( .A(u2__abc_44228_n8066), .Y(u2__abc_44228_n8067) );
  INVX1 INVX1_2056 ( .A(u2__abc_44228_n8075), .Y(u2__abc_44228_n8076_1) );
  INVX1 INVX1_2057 ( .A(u2__abc_44228_n8082_1), .Y(u2__abc_44228_n8083) );
  INVX1 INVX1_2058 ( .A(u2__abc_44228_n8090), .Y(u2__abc_44228_n8091) );
  INVX1 INVX1_2059 ( .A(u2__abc_44228_n3579), .Y(u2__abc_44228_n8099) );
  INVX1 INVX1_206 ( .A(sqrto_12_), .Y(u2__abc_44228_n3128) );
  INVX1 INVX1_2060 ( .A(u2__abc_44228_n8097), .Y(u2__abc_44228_n8100) );
  INVX1 INVX1_2061 ( .A(u2__abc_44228_n8107), .Y(u2__abc_44228_n8108) );
  INVX1 INVX1_2062 ( .A(u2__abc_44228_n8117), .Y(u2__abc_44228_n8118) );
  INVX1 INVX1_2063 ( .A(u2__abc_44228_n8124), .Y(u2__abc_44228_n8125_1) );
  INVX1 INVX1_2064 ( .A(u2__abc_44228_n3560), .Y(u2__abc_44228_n8132) );
  INVX1 INVX1_2065 ( .A(u2__abc_44228_n8133), .Y(u2__abc_44228_n8135) );
  INVX1 INVX1_2066 ( .A(u2__abc_44228_n8141), .Y(u2__abc_44228_n8142_1) );
  INVX1 INVX1_2067 ( .A(u2__abc_44228_n8150), .Y(u2__abc_44228_n8151) );
  INVX1 INVX1_2068 ( .A(u2__abc_44228_n8158_1), .Y(u2__abc_44228_n8159_1) );
  INVX1 INVX1_2069 ( .A(u2__abc_44228_n3553), .Y(u2__abc_44228_n8165) );
  INVX1 INVX1_207 ( .A(u2_remHi_12_), .Y(u2__abc_44228_n3130) );
  INVX1 INVX1_2070 ( .A(u2__abc_44228_n8166), .Y(u2__abc_44228_n8168) );
  INVX1 INVX1_2071 ( .A(u2__abc_44228_n8175_1), .Y(u2__abc_44228_n8176) );
  INVX1 INVX1_2072 ( .A(u2__abc_44228_n8184), .Y(u2__abc_44228_n8185) );
  INVX1 INVX1_2073 ( .A(u2__abc_44228_n8187), .Y(u2__abc_44228_n8188) );
  INVX1 INVX1_2074 ( .A(u2__abc_44228_n8193), .Y(u2__abc_44228_n8194) );
  INVX1 INVX1_2075 ( .A(u2__abc_44228_n3533), .Y(u2__abc_44228_n8200) );
  INVX1 INVX1_2076 ( .A(u2__abc_44228_n8201), .Y(u2__abc_44228_n8203_1) );
  INVX1 INVX1_2077 ( .A(u2__abc_44228_n8213_1), .Y(u2__abc_44228_n8214_1) );
  INVX1 INVX1_2078 ( .A(u2__abc_44228_n8223), .Y(u2__abc_44228_n8224_1) );
  INVX1 INVX1_2079 ( .A(u2__abc_44228_n8230_1), .Y(u2__abc_44228_n8231) );
  INVX1 INVX1_208 ( .A(u2__abc_44228_n3132), .Y(u2__abc_44228_n3133) );
  INVX1 INVX1_2080 ( .A(u2__abc_44228_n3503), .Y(u2__abc_44228_n8237) );
  INVX1 INVX1_2081 ( .A(u2__abc_44228_n8238), .Y(u2__abc_44228_n8239) );
  INVX1 INVX1_2082 ( .A(u2__abc_44228_n8247_1), .Y(u2__abc_44228_n8248) );
  INVX1 INVX1_2083 ( .A(u2__abc_44228_n8257_1), .Y(u2__abc_44228_n8258_1) );
  INVX1 INVX1_2084 ( .A(u2__abc_44228_n8264), .Y(u2__abc_44228_n8265) );
  INVX1 INVX1_2085 ( .A(u2__abc_44228_n3517), .Y(u2__abc_44228_n8271) );
  INVX1 INVX1_2086 ( .A(u2__abc_44228_n8272), .Y(u2__abc_44228_n8273) );
  INVX1 INVX1_2087 ( .A(u2__abc_44228_n8281), .Y(u2__abc_44228_n8282) );
  INVX1 INVX1_2088 ( .A(u2__abc_44228_n8289), .Y(u2__abc_44228_n8290_1) );
  INVX1 INVX1_2089 ( .A(u2__abc_44228_n8291_1), .Y(u2__abc_44228_n8292) );
  INVX1 INVX1_209 ( .A(sqrto_11_), .Y(u2__abc_44228_n3135) );
  INVX1 INVX1_2090 ( .A(u2__abc_44228_n8299), .Y(u2__abc_44228_n8300) );
  INVX1 INVX1_2091 ( .A(u2__abc_44228_n3494), .Y(u2__abc_44228_n8306) );
  INVX1 INVX1_2092 ( .A(u2__abc_44228_n8307_1), .Y(u2__abc_44228_n8309) );
  INVX1 INVX1_2093 ( .A(u2__abc_44228_n8316), .Y(u2__abc_44228_n8317) );
  INVX1 INVX1_2094 ( .A(u2__abc_44228_n8324_1), .Y(u2__abc_44228_n8325) );
  INVX1 INVX1_2095 ( .A(u2__abc_44228_n8327), .Y(u2__abc_44228_n8328) );
  INVX1 INVX1_2096 ( .A(u2__abc_44228_n8334_1), .Y(u2__abc_44228_n8335_1) );
  INVX1 INVX1_2097 ( .A(u2__abc_44228_n3474), .Y(u2__abc_44228_n8341) );
  INVX1 INVX1_2098 ( .A(u2__abc_44228_n8342), .Y(u2__abc_44228_n8343) );
  INVX1 INVX1_2099 ( .A(u2__abc_44228_n8351_1), .Y(u2__abc_44228_n8352) );
  INVX1 INVX1_21 ( .A(\a[119] ), .Y(_abc_64468_n1580) );
  INVX1 INVX1_210 ( .A(u2__abc_44228_n3136), .Y(u2__abc_44228_n3137) );
  INVX1 INVX1_2100 ( .A(u2__abc_44228_n8360), .Y(u2__abc_44228_n8361) );
  INVX1 INVX1_2101 ( .A(u2__abc_44228_n8368_1), .Y(u2__abc_44228_n8369) );
  INVX1 INVX1_2102 ( .A(u2__abc_44228_n3457_1), .Y(u2__abc_44228_n8375) );
  INVX1 INVX1_2103 ( .A(u2__abc_44228_n8376), .Y(u2__abc_44228_n8377) );
  INVX1 INVX1_2104 ( .A(u2__abc_44228_n8385), .Y(u2__abc_44228_n8386) );
  INVX1 INVX1_2105 ( .A(u2__abc_44228_n8395_1), .Y(u2__abc_44228_n8396) );
  INVX1 INVX1_2106 ( .A(u2__abc_44228_n8402), .Y(u2__abc_44228_n8403) );
  INVX1 INVX1_2107 ( .A(u2__abc_44228_n3443), .Y(u2__abc_44228_n8409) );
  INVX1 INVX1_2108 ( .A(u2__abc_44228_n8410), .Y(u2__abc_44228_n8412_1) );
  INVX1 INVX1_2109 ( .A(u2__abc_44228_n8419), .Y(u2__abc_44228_n8420) );
  INVX1 INVX1_211 ( .A(u2_remHi_11_), .Y(u2__abc_44228_n3138) );
  INVX1 INVX1_2110 ( .A(u2__abc_44228_n8428_1), .Y(u2__abc_44228_n8429) );
  INVX1 INVX1_2111 ( .A(u2__abc_44228_n8436), .Y(u2__abc_44228_n8437) );
  INVX1 INVX1_2112 ( .A(u2__abc_44228_n3434), .Y(u2__abc_44228_n8445_1) );
  INVX1 INVX1_2113 ( .A(u2__abc_44228_n8443), .Y(u2__abc_44228_n8446) );
  INVX1 INVX1_2114 ( .A(u2__abc_44228_n8453), .Y(u2__abc_44228_n8454) );
  INVX1 INVX1_2115 ( .A(u2__abc_44228_n8461_1), .Y(u2__abc_44228_n8462) );
  INVX1 INVX1_2116 ( .A(u2__abc_44228_n8464), .Y(u2__abc_44228_n8465) );
  INVX1 INVX1_2117 ( .A(u2__abc_44228_n8471), .Y(u2__abc_44228_n8472_1) );
  INVX1 INVX1_2118 ( .A(u2__abc_44228_n3414), .Y(u2__abc_44228_n8478_1) );
  INVX1 INVX1_2119 ( .A(u2__abc_44228_n8479), .Y(u2__abc_44228_n8480) );
  INVX1 INVX1_212 ( .A(u2__abc_44228_n3139), .Y(u2__abc_44228_n3140) );
  INVX1 INVX1_2120 ( .A(u2__abc_44228_n8488_1), .Y(u2__abc_44228_n8489_1) );
  INVX1 INVX1_2121 ( .A(u2__abc_44228_n8498), .Y(u2__abc_44228_n8499_1) );
  INVX1 INVX1_2122 ( .A(u2__abc_44228_n8505_1), .Y(u2__abc_44228_n8506) );
  INVX1 INVX1_2123 ( .A(u2__abc_44228_n3398), .Y(u2__abc_44228_n8513) );
  INVX1 INVX1_2124 ( .A(u2__abc_44228_n8514), .Y(u2__abc_44228_n8516_1) );
  INVX1 INVX1_2125 ( .A(u2__abc_44228_n8522_1), .Y(u2__abc_44228_n8523) );
  INVX1 INVX1_2126 ( .A(u2__abc_44228_n8532_1), .Y(u2__abc_44228_n8533_1) );
  INVX1 INVX1_2127 ( .A(u2__abc_44228_n8539), .Y(u2__abc_44228_n8540) );
  INVX1 INVX1_2128 ( .A(u2__abc_44228_n8546), .Y(u2__abc_44228_n8547) );
  INVX1 INVX1_2129 ( .A(u2__abc_44228_n3384), .Y(u2__abc_44228_n8549_1) );
  INVX1 INVX1_213 ( .A(sqrto_10_), .Y(u2__abc_44228_n3142) );
  INVX1 INVX1_2130 ( .A(u2__abc_44228_n8556), .Y(u2__abc_44228_n8557) );
  INVX1 INVX1_2131 ( .A(u2__abc_44228_n8564), .Y(u2__abc_44228_n8565_1) );
  INVX1 INVX1_2132 ( .A(u2__abc_44228_n8566_1), .Y(u2__abc_44228_n8567) );
  INVX1 INVX1_2133 ( .A(u2__abc_44228_n8574), .Y(u2__abc_44228_n8575) );
  INVX1 INVX1_2134 ( .A(u2__abc_44228_n8581), .Y(u2__abc_44228_n8582_1) );
  INVX1 INVX1_2135 ( .A(u2__abc_44228_n3375), .Y(u2__abc_44228_n8584) );
  INVX1 INVX1_2136 ( .A(u2__abc_44228_n8591), .Y(u2__abc_44228_n8592) );
  INVX1 INVX1_2137 ( .A(u2__abc_44228_n8599_1), .Y(u2__abc_44228_n8600) );
  INVX1 INVX1_2138 ( .A(u2__abc_44228_n8602), .Y(u2__abc_44228_n8603) );
  INVX1 INVX1_2139 ( .A(u2__abc_44228_n8609_1), .Y(u2__abc_44228_n8610_1) );
  INVX1 INVX1_214 ( .A(u2_remHi_10_), .Y(u2__abc_44228_n3144) );
  INVX1 INVX1_2140 ( .A(u2__abc_44228_n3355), .Y(u2__abc_44228_n8616) );
  INVX1 INVX1_2141 ( .A(u2__abc_44228_n8617), .Y(u2__abc_44228_n8618) );
  INVX1 INVX1_2142 ( .A(u2__abc_44228_n8626_1), .Y(u2__abc_44228_n8627) );
  INVX1 INVX1_2143 ( .A(u2__abc_44228_n8634), .Y(u2__abc_44228_n8635) );
  INVX1 INVX1_2144 ( .A(u2__abc_44228_n8641), .Y(u2__abc_44228_n8642_1) );
  INVX1 INVX1_2145 ( .A(u2__abc_44228_n4128_1), .Y(u2__abc_44228_n8648_1) );
  INVX1 INVX1_2146 ( .A(u2__abc_44228_n8649), .Y(u2__abc_44228_n8650) );
  INVX1 INVX1_2147 ( .A(u2__abc_44228_n8658), .Y(u2__abc_44228_n8659_1) );
  INVX1 INVX1_2148 ( .A(u2__abc_44228_n8668), .Y(u2__abc_44228_n8669) );
  INVX1 INVX1_2149 ( .A(u2__abc_44228_n8675_1), .Y(u2__abc_44228_n8676_1) );
  INVX1 INVX1_215 ( .A(u2__abc_44228_n3146), .Y(u2__abc_44228_n3147) );
  INVX1 INVX1_2150 ( .A(u2__abc_44228_n4115), .Y(u2__abc_44228_n8682) );
  INVX1 INVX1_2151 ( .A(u2__abc_44228_n8683), .Y(u2__abc_44228_n8684) );
  INVX1 INVX1_2152 ( .A(u2__abc_44228_n8692_1), .Y(u2__abc_44228_n8693) );
  INVX1 INVX1_2153 ( .A(u2__abc_44228_n8701), .Y(u2__abc_44228_n8702) );
  INVX1 INVX1_2154 ( .A(u2__abc_44228_n8709_1), .Y(u2__abc_44228_n8710) );
  INVX1 INVX1_2155 ( .A(u2__abc_44228_n4102), .Y(u2__abc_44228_n8716) );
  INVX1 INVX1_2156 ( .A(u2__abc_44228_n8717), .Y(u2__abc_44228_n8719_1) );
  INVX1 INVX1_2157 ( .A(u2__abc_44228_n8726), .Y(u2__abc_44228_n8727) );
  INVX1 INVX1_2158 ( .A(u2__abc_44228_n8737), .Y(u2__abc_44228_n8738) );
  INVX1 INVX1_2159 ( .A(u2__abc_44228_n8743), .Y(u2__abc_44228_n8744) );
  INVX1 INVX1_216 ( .A(u2_remHi_9_), .Y(u2__abc_44228_n3150) );
  INVX1 INVX1_2160 ( .A(u2__abc_44228_n4088), .Y(u2__abc_44228_n8751) );
  INVX1 INVX1_2161 ( .A(u2__abc_44228_n8752_1), .Y(u2__abc_44228_n8754) );
  INVX1 INVX1_2162 ( .A(u2__abc_44228_n8760), .Y(u2__abc_44228_n8761) );
  INVX1 INVX1_2163 ( .A(u2__abc_44228_n8770), .Y(u2__abc_44228_n8771) );
  INVX1 INVX1_2164 ( .A(u2__abc_44228_n8777), .Y(u2__abc_44228_n8778) );
  INVX1 INVX1_2165 ( .A(u2__abc_44228_n4058), .Y(u2__abc_44228_n8784) );
  INVX1 INVX1_2166 ( .A(u2__abc_44228_n8785_1), .Y(u2__abc_44228_n8787) );
  INVX1 INVX1_2167 ( .A(u2__abc_44228_n8794), .Y(u2__abc_44228_n8795) );
  INVX1 INVX1_2168 ( .A(u2__abc_44228_n8805), .Y(u2__abc_44228_n8806) );
  INVX1 INVX1_2169 ( .A(u2__abc_44228_n8811), .Y(u2__abc_44228_n8812) );
  INVX1 INVX1_217 ( .A(sqrto_9_), .Y(u2__abc_44228_n3152) );
  INVX1 INVX1_2170 ( .A(u2__abc_44228_n4072), .Y(u2__abc_44228_n8819_1) );
  INVX1 INVX1_2171 ( .A(u2__abc_44228_n8820), .Y(u2__abc_44228_n8821) );
  INVX1 INVX1_2172 ( .A(u2__abc_44228_n8828), .Y(u2__abc_44228_n8829_1) );
  INVX1 INVX1_2173 ( .A(u2__abc_44228_n8836), .Y(u2__abc_44228_n8837) );
  INVX1 INVX1_2174 ( .A(u2__abc_44228_n8838), .Y(u2__abc_44228_n8839) );
  INVX1 INVX1_2175 ( .A(u2__abc_44228_n8846_1), .Y(u2__abc_44228_n8847) );
  INVX1 INVX1_2176 ( .A(u2__abc_44228_n8853), .Y(u2__abc_44228_n8854) );
  INVX1 INVX1_2177 ( .A(u2__abc_44228_n4049), .Y(u2__abc_44228_n8856) );
  INVX1 INVX1_2178 ( .A(u2__abc_44228_n8863_1), .Y(u2__abc_44228_n8864) );
  INVX1 INVX1_2179 ( .A(u2__abc_44228_n8871), .Y(u2__abc_44228_n8872) );
  INVX1 INVX1_218 ( .A(u2_remHi_8_), .Y(u2__abc_44228_n3155) );
  INVX1 INVX1_2180 ( .A(u2__abc_44228_n8874_1), .Y(u2__abc_44228_n8875) );
  INVX1 INVX1_2181 ( .A(u2__abc_44228_n8881), .Y(u2__abc_44228_n8882) );
  INVX1 INVX1_2182 ( .A(u2__abc_44228_n4029), .Y(u2__abc_44228_n8888) );
  INVX1 INVX1_2183 ( .A(u2__abc_44228_n4031), .Y(u2__abc_44228_n8889) );
  INVX1 INVX1_2184 ( .A(u2__abc_44228_n8890_1), .Y(u2__abc_44228_n8892) );
  INVX1 INVX1_2185 ( .A(u2__abc_44228_n8899), .Y(u2__abc_44228_n8900) );
  INVX1 INVX1_2186 ( .A(u2__abc_44228_n8908), .Y(u2__abc_44228_n8909) );
  INVX1 INVX1_2187 ( .A(u2__abc_44228_n8916), .Y(u2__abc_44228_n8917_1) );
  INVX1 INVX1_2188 ( .A(u2__abc_44228_n4018), .Y(u2__abc_44228_n8923_1) );
  INVX1 INVX1_2189 ( .A(u2__abc_44228_n8924), .Y(u2__abc_44228_n8925) );
  INVX1 INVX1_219 ( .A(sqrto_8_), .Y(u2__abc_44228_n3157) );
  INVX1 INVX1_2190 ( .A(u2__abc_44228_n8933), .Y(u2__abc_44228_n8934_1) );
  INVX1 INVX1_2191 ( .A(u2__abc_44228_n8941), .Y(u2__abc_44228_n8942) );
  INVX1 INVX1_2192 ( .A(u2__abc_44228_n8944), .Y(u2__abc_44228_n8945_1) );
  INVX1 INVX1_2193 ( .A(u2__abc_44228_n8951_1), .Y(u2__abc_44228_n8952) );
  INVX1 INVX1_2194 ( .A(u2__abc_44228_n3998), .Y(u2__abc_44228_n8960) );
  INVX1 INVX1_2195 ( .A(u2__abc_44228_n8958), .Y(u2__abc_44228_n8961_1) );
  INVX1 INVX1_2196 ( .A(u2__abc_44228_n8968), .Y(u2__abc_44228_n8969) );
  INVX1 INVX1_2197 ( .A(u2__abc_44228_n8978_1), .Y(u2__abc_44228_n8979) );
  INVX1 INVX1_2198 ( .A(u2__abc_44228_n8985), .Y(u2__abc_44228_n8986) );
  INVX1 INVX1_2199 ( .A(u2__abc_44228_n3989), .Y(u2__abc_44228_n8992) );
  INVX1 INVX1_22 ( .A(_abc_64468_n1583), .Y(_abc_64468_n1584) );
  INVX1 INVX1_220 ( .A(sqrto_6_), .Y(u2__abc_44228_n3161) );
  INVX1 INVX1_2200 ( .A(u2__abc_44228_n8993), .Y(u2__abc_44228_n8995_1) );
  INVX1 INVX1_2201 ( .A(u2__abc_44228_n9002), .Y(u2__abc_44228_n9003) );
  INVX1 INVX1_2202 ( .A(u2__abc_44228_n9012), .Y(u2__abc_44228_n9013) );
  INVX1 INVX1_2203 ( .A(u2__abc_44228_n9019), .Y(u2__abc_44228_n9020) );
  INVX1 INVX1_2204 ( .A(u2__abc_44228_n3969), .Y(u2__abc_44228_n9028_1) );
  INVX1 INVX1_2205 ( .A(u2__abc_44228_n9026), .Y(u2__abc_44228_n9029) );
  INVX1 INVX1_2206 ( .A(u2__abc_44228_n9036), .Y(u2__abc_44228_n9037) );
  INVX1 INVX1_2207 ( .A(u2__abc_44228_n9047), .Y(u2__abc_44228_n9048) );
  INVX1 INVX1_2208 ( .A(u2__abc_44228_n9053), .Y(u2__abc_44228_n9054) );
  INVX1 INVX1_2209 ( .A(u2__abc_44228_n3959), .Y(u2__abc_44228_n9061_1) );
  INVX1 INVX1_221 ( .A(u2_remHi_6_), .Y(u2__abc_44228_n3163) );
  INVX1 INVX1_2210 ( .A(u2__abc_44228_n9062), .Y(u2__abc_44228_n9063) );
  INVX1 INVX1_2211 ( .A(u2__abc_44228_n9070), .Y(u2__abc_44228_n9071_1) );
  INVX1 INVX1_2212 ( .A(u2__abc_44228_n9078), .Y(u2__abc_44228_n9079) );
  INVX1 INVX1_2213 ( .A(u2__abc_44228_n9081), .Y(u2__abc_44228_n9082_1) );
  INVX1 INVX1_2214 ( .A(u2__abc_44228_n9088_1), .Y(u2__abc_44228_n9089) );
  INVX1 INVX1_2215 ( .A(u2__abc_44228_n3939), .Y(u2__abc_44228_n9095) );
  INVX1 INVX1_2216 ( .A(u2__abc_44228_n9096), .Y(u2__abc_44228_n9097) );
  INVX1 INVX1_2217 ( .A(u2__abc_44228_n9105_1), .Y(u2__abc_44228_n9106) );
  INVX1 INVX1_2218 ( .A(u2__abc_44228_n9114), .Y(u2__abc_44228_n9115_1) );
  INVX1 INVX1_2219 ( .A(u2__abc_44228_n9122), .Y(u2__abc_44228_n9123) );
  INVX1 INVX1_222 ( .A(u2__abc_44228_n3165), .Y(u2__abc_44228_n3166) );
  INVX1 INVX1_2220 ( .A(u2__abc_44228_n3930_1), .Y(u2__abc_44228_n9131) );
  INVX1 INVX1_2221 ( .A(u2__abc_44228_n9129), .Y(u2__abc_44228_n9132_1) );
  INVX1 INVX1_2222 ( .A(u2__abc_44228_n9139), .Y(u2__abc_44228_n9140) );
  INVX1 INVX1_2223 ( .A(u2__abc_44228_n9147), .Y(u2__abc_44228_n9148_1) );
  INVX1 INVX1_2224 ( .A(u2__abc_44228_n9150), .Y(u2__abc_44228_n9151) );
  INVX1 INVX1_2225 ( .A(u2__abc_44228_n9157), .Y(u2__abc_44228_n9158) );
  INVX1 INVX1_2226 ( .A(u2__abc_44228_n3910), .Y(u2__abc_44228_n9164) );
  INVX1 INVX1_2227 ( .A(u2__abc_44228_n9165_1), .Y(u2__abc_44228_n9166) );
  INVX1 INVX1_2228 ( .A(u2__abc_44228_n9174), .Y(u2__abc_44228_n9175) );
  INVX1 INVX1_2229 ( .A(u2__abc_44228_n9183), .Y(u2__abc_44228_n9184) );
  INVX1 INVX1_223 ( .A(sqrto_7_), .Y(u2__abc_44228_n3167) );
  INVX1 INVX1_2230 ( .A(u2__abc_44228_n9191), .Y(u2__abc_44228_n9192_1) );
  INVX1 INVX1_2231 ( .A(u2__abc_44228_n3898), .Y(u2__abc_44228_n9200) );
  INVX1 INVX1_2232 ( .A(u2__abc_44228_n9198_1), .Y(u2__abc_44228_n9201) );
  INVX1 INVX1_2233 ( .A(u2__abc_44228_n9208), .Y(u2__abc_44228_n9209_1) );
  INVX1 INVX1_2234 ( .A(u2__abc_44228_n9216), .Y(u2__abc_44228_n9217) );
  INVX1 INVX1_2235 ( .A(u2__abc_44228_n9219), .Y(u2__abc_44228_n9220_1) );
  INVX1 INVX1_2236 ( .A(u2__abc_44228_n9226_1), .Y(u2__abc_44228_n9227) );
  INVX1 INVX1_2237 ( .A(u2__abc_44228_n3878), .Y(u2__abc_44228_n9235) );
  INVX1 INVX1_2238 ( .A(u2__abc_44228_n9233), .Y(u2__abc_44228_n9236_1) );
  INVX1 INVX1_2239 ( .A(u2__abc_44228_n9243), .Y(u2__abc_44228_n9244) );
  INVX1 INVX1_224 ( .A(u2__abc_44228_n3168), .Y(u2__abc_44228_n3169) );
  INVX1 INVX1_2240 ( .A(u2__abc_44228_n9253_1), .Y(u2__abc_44228_n9254) );
  INVX1 INVX1_2241 ( .A(u2__abc_44228_n9260), .Y(u2__abc_44228_n9261) );
  INVX1 INVX1_2242 ( .A(u2__abc_44228_n3869), .Y(u2__abc_44228_n9267) );
  INVX1 INVX1_2243 ( .A(u2__abc_44228_n9268), .Y(u2__abc_44228_n9270_1) );
  INVX1 INVX1_2244 ( .A(u2__abc_44228_n9277), .Y(u2__abc_44228_n9278) );
  INVX1 INVX1_2245 ( .A(u2__abc_44228_n9287), .Y(u2__abc_44228_n9288) );
  INVX1 INVX1_2246 ( .A(u2__abc_44228_n9294), .Y(u2__abc_44228_n9295) );
  INVX1 INVX1_2247 ( .A(u2__abc_44228_n3849), .Y(u2__abc_44228_n9303_1) );
  INVX1 INVX1_2248 ( .A(u2__abc_44228_n9301), .Y(u2__abc_44228_n9304) );
  INVX1 INVX1_2249 ( .A(u2__abc_44228_n9311), .Y(u2__abc_44228_n9312) );
  INVX1 INVX1_225 ( .A(u2_remHi_7_), .Y(u2__abc_44228_n3170) );
  INVX1 INVX1_2250 ( .A(u2__abc_44228_n9322), .Y(u2__abc_44228_n9323) );
  INVX1 INVX1_2251 ( .A(u2__abc_44228_n9328), .Y(u2__abc_44228_n9329) );
  INVX1 INVX1_2252 ( .A(u2__abc_44228_n3819), .Y(u2__abc_44228_n9336_1) );
  INVX1 INVX1_2253 ( .A(u2__abc_44228_n9337), .Y(u2__abc_44228_n9338) );
  INVX1 INVX1_2254 ( .A(u2__abc_44228_n9345), .Y(u2__abc_44228_n9346_1) );
  INVX1 INVX1_2255 ( .A(u2__abc_44228_n9355), .Y(u2__abc_44228_n9356) );
  INVX1 INVX1_2256 ( .A(u2__abc_44228_n9362), .Y(u2__abc_44228_n9363_1) );
  INVX1 INVX1_2257 ( .A(u2__abc_44228_n3833), .Y(u2__abc_44228_n9369_1) );
  INVX1 INVX1_2258 ( .A(u2__abc_44228_n9370), .Y(u2__abc_44228_n9372) );
  INVX1 INVX1_2259 ( .A(u2__abc_44228_n9379_1), .Y(u2__abc_44228_n9380_1) );
  INVX1 INVX1_226 ( .A(u2__abc_44228_n3171), .Y(u2__abc_44228_n3172) );
  INVX1 INVX1_2260 ( .A(u2__abc_44228_n9387), .Y(u2__abc_44228_n9388) );
  INVX1 INVX1_2261 ( .A(u2__abc_44228_n9389), .Y(u2__abc_44228_n9390_1) );
  INVX1 INVX1_2262 ( .A(u2__abc_44228_n9397), .Y(u2__abc_44228_n9398) );
  INVX1 INVX1_2263 ( .A(u2__abc_44228_n3810), .Y(u2__abc_44228_n9406) );
  INVX1 INVX1_2264 ( .A(u2__abc_44228_n9404), .Y(u2__abc_44228_n9407_1) );
  INVX1 INVX1_2265 ( .A(u2__abc_44228_n9414), .Y(u2__abc_44228_n9415) );
  INVX1 INVX1_2266 ( .A(u2__abc_44228_n9422), .Y(u2__abc_44228_n9423_1) );
  INVX1 INVX1_2267 ( .A(u2__abc_44228_n9425), .Y(u2__abc_44228_n9426) );
  INVX1 INVX1_2268 ( .A(u2__abc_44228_n9432), .Y(u2__abc_44228_n9433) );
  INVX1 INVX1_2269 ( .A(u2__abc_44228_n3790), .Y(u2__abc_44228_n9439) );
  INVX1 INVX1_227 ( .A(u2__abc_44228_n3151), .Y(u2__abc_44228_n3181) );
  INVX1 INVX1_2270 ( .A(u2__abc_44228_n9440_1), .Y(u2__abc_44228_n9441) );
  INVX1 INVX1_2271 ( .A(u2__abc_44228_n9449), .Y(u2__abc_44228_n9450) );
  INVX1 INVX1_2272 ( .A(u2__abc_44228_n9459), .Y(u2__abc_44228_n9460) );
  INVX1 INVX1_2273 ( .A(u2__abc_44228_n9466), .Y(u2__abc_44228_n9467_1) );
  INVX1 INVX1_2274 ( .A(u2__abc_44228_n3779_1), .Y(u2__abc_44228_n9474) );
  INVX1 INVX1_2275 ( .A(u2__abc_44228_n9475), .Y(u2__abc_44228_n9476) );
  INVX1 INVX1_2276 ( .A(u2__abc_44228_n9483), .Y(u2__abc_44228_n9484_1) );
  INVX1 INVX1_2277 ( .A(u2__abc_44228_n9491), .Y(u2__abc_44228_n9492) );
  INVX1 INVX1_2278 ( .A(u2__abc_44228_n9494), .Y(u2__abc_44228_n9495_1) );
  INVX1 INVX1_2279 ( .A(u2__abc_44228_n9501_1), .Y(u2__abc_44228_n9502) );
  INVX1 INVX1_228 ( .A(u2__abc_44228_n3156), .Y(u2__abc_44228_n3182) );
  INVX1 INVX1_2280 ( .A(u2__abc_44228_n3759_1), .Y(u2__abc_44228_n9508) );
  INVX1 INVX1_2281 ( .A(u2__abc_44228_n9509), .Y(u2__abc_44228_n9510) );
  INVX1 INVX1_2282 ( .A(u2__abc_44228_n9518), .Y(u2__abc_44228_n9519) );
  INVX1 INVX1_2283 ( .A(u2__abc_44228_n9527), .Y(u2__abc_44228_n9528_1) );
  INVX1 INVX1_2284 ( .A(u2__abc_44228_n9535), .Y(u2__abc_44228_n9536) );
  INVX1 INVX1_2285 ( .A(u2__abc_44228_n9542), .Y(u2__abc_44228_n9543) );
  INVX1 INVX1_2286 ( .A(u2__abc_44228_n3744), .Y(u2__abc_44228_n9545_1) );
  INVX1 INVX1_2287 ( .A(u2__abc_44228_n9552), .Y(u2__abc_44228_n9553) );
  INVX1 INVX1_2288 ( .A(u2__abc_44228_n9562), .Y(u2__abc_44228_n9563) );
  INVX1 INVX1_2289 ( .A(u2__abc_44228_n9569), .Y(u2__abc_44228_n9570) );
  INVX1 INVX1_229 ( .A(sqrto_29_), .Y(u2__abc_44228_n3195) );
  INVX1 INVX1_2290 ( .A(u2__abc_44228_n3730), .Y(u2__abc_44228_n9576) );
  INVX1 INVX1_2291 ( .A(u2__abc_44228_n9577_1), .Y(u2__abc_44228_n9578_1) );
  INVX1 INVX1_2292 ( .A(u2__abc_44228_n9586), .Y(u2__abc_44228_n9587) );
  INVX1 INVX1_2293 ( .A(u2__abc_44228_n9596), .Y(u2__abc_44228_n9597) );
  INVX1 INVX1_2294 ( .A(u2__abc_44228_n9603), .Y(u2__abc_44228_n9604) );
  INVX1 INVX1_2295 ( .A(u2__abc_44228_n3700), .Y(u2__abc_44228_n9610_1) );
  INVX1 INVX1_2296 ( .A(u2__abc_44228_n9611_1), .Y(u2__abc_44228_n9613) );
  INVX1 INVX1_2297 ( .A(u2__abc_44228_n9620), .Y(u2__abc_44228_n9621_1) );
  INVX1 INVX1_2298 ( .A(u2__abc_44228_n9630), .Y(u2__abc_44228_n9631) );
  INVX1 INVX1_2299 ( .A(u2__abc_44228_n9637), .Y(u2__abc_44228_n9638_1) );
  INVX1 INVX1_23 ( .A(_abc_64468_n1585), .Y(_abc_64468_n1586) );
  INVX1 INVX1_230 ( .A(u2__abc_44228_n3196), .Y(u2__abc_44228_n3197) );
  INVX1 INVX1_2300 ( .A(u2__abc_44228_n3714_1), .Y(u2__abc_44228_n9644_1) );
  INVX1 INVX1_2301 ( .A(u2__abc_44228_n9645), .Y(u2__abc_44228_n9646) );
  INVX1 INVX1_2302 ( .A(u2__abc_44228_n9654_1), .Y(u2__abc_44228_n9655_1) );
  INVX1 INVX1_2303 ( .A(u2__abc_44228_n9663), .Y(u2__abc_44228_n9664) );
  INVX1 INVX1_2304 ( .A(u2__abc_44228_n9671_1), .Y(u2__abc_44228_n9672) );
  INVX1 INVX1_2305 ( .A(u2__abc_44228_n3691), .Y(u2__abc_44228_n9680) );
  INVX1 INVX1_2306 ( .A(u2__abc_44228_n9678), .Y(u2__abc_44228_n9681) );
  INVX1 INVX1_2307 ( .A(u2__abc_44228_n9688_1), .Y(u2__abc_44228_n9689) );
  INVX1 INVX1_2308 ( .A(u2__abc_44228_n9696), .Y(u2__abc_44228_n9697) );
  INVX1 INVX1_2309 ( .A(u2__abc_44228_n9699_1), .Y(u2__abc_44228_n9700) );
  INVX1 INVX1_231 ( .A(u2_remHi_29_), .Y(u2__abc_44228_n3198) );
  INVX1 INVX1_2310 ( .A(u2__abc_44228_n9706), .Y(u2__abc_44228_n9707) );
  INVX1 INVX1_2311 ( .A(u2__abc_44228_n3671), .Y(u2__abc_44228_n9713) );
  INVX1 INVX1_2312 ( .A(u2__abc_44228_n9714), .Y(u2__abc_44228_n9715_1) );
  INVX1 INVX1_2313 ( .A(u2__abc_44228_n9723), .Y(u2__abc_44228_n9724) );
  INVX1 INVX1_2314 ( .A(u2__abc_44228_n9730), .Y(u2__abc_44228_n9731_1) );
  INVX1 INVX1_2315 ( .A(u2__abc_44228_n9738), .Y(u2__abc_44228_n9739) );
  INVX1 INVX1_2316 ( .A(u2__abc_44228_n5243), .Y(u2__abc_44228_n9745) );
  INVX1 INVX1_2317 ( .A(u2__abc_44228_n9746), .Y(u2__abc_44228_n9748_1) );
  INVX1 INVX1_2318 ( .A(u2__abc_44228_n9755), .Y(u2__abc_44228_n9756) );
  INVX1 INVX1_2319 ( .A(u2__abc_44228_n9766), .Y(u2__abc_44228_n9767) );
  INVX1 INVX1_232 ( .A(u2__abc_44228_n3199), .Y(u2__abc_44228_n3200) );
  INVX1 INVX1_2320 ( .A(u2__abc_44228_n9772), .Y(u2__abc_44228_n9773) );
  INVX1 INVX1_2321 ( .A(u2__abc_44228_n5230_1), .Y(u2__abc_44228_n9780) );
  INVX1 INVX1_2322 ( .A(u2__abc_44228_n9781_1), .Y(u2__abc_44228_n9782) );
  INVX1 INVX1_2323 ( .A(u2__abc_44228_n9789), .Y(u2__abc_44228_n9790) );
  INVX1 INVX1_2324 ( .A(u2__abc_44228_n9799), .Y(u2__abc_44228_n9800) );
  INVX1 INVX1_2325 ( .A(u2__abc_44228_n9806), .Y(u2__abc_44228_n9807) );
  INVX1 INVX1_2326 ( .A(u2__abc_44228_n5217), .Y(u2__abc_44228_n9814_1) );
  INVX1 INVX1_2327 ( .A(u2__abc_44228_n9815), .Y(u2__abc_44228_n9817) );
  INVX1 INVX1_2328 ( .A(u2__abc_44228_n9823), .Y(u2__abc_44228_n9824) );
  INVX1 INVX1_2329 ( .A(u2__abc_44228_n9833), .Y(u2__abc_44228_n9834) );
  INVX1 INVX1_233 ( .A(sqrto_28_), .Y(u2__abc_44228_n3202) );
  INVX1 INVX1_2330 ( .A(u2__abc_44228_n9840), .Y(u2__abc_44228_n9841_1) );
  INVX1 INVX1_2331 ( .A(u2__abc_44228_n5203), .Y(u2__abc_44228_n9849) );
  INVX1 INVX1_2332 ( .A(u2__abc_44228_n9847_1), .Y(u2__abc_44228_n9850) );
  INVX1 INVX1_2333 ( .A(u2__abc_44228_n9857), .Y(u2__abc_44228_n9858_1) );
  INVX1 INVX1_2334 ( .A(u2__abc_44228_n9868), .Y(u2__abc_44228_n9869_1) );
  INVX1 INVX1_2335 ( .A(u2__abc_44228_n9874_1), .Y(u2__abc_44228_n9875_1) );
  INVX1 INVX1_2336 ( .A(u2__abc_44228_n5173_1), .Y(u2__abc_44228_n9882) );
  INVX1 INVX1_2337 ( .A(u2__abc_44228_n9883), .Y(u2__abc_44228_n9885_1) );
  INVX1 INVX1_2338 ( .A(u2__abc_44228_n9891_1), .Y(u2__abc_44228_n9892) );
  INVX1 INVX1_2339 ( .A(u2__abc_44228_n9901), .Y(u2__abc_44228_n9902_1) );
  INVX1 INVX1_234 ( .A(u2_remHi_28_), .Y(u2__abc_44228_n3204) );
  INVX1 INVX1_2340 ( .A(u2__abc_44228_n9908_1), .Y(u2__abc_44228_n9909) );
  INVX1 INVX1_2341 ( .A(u2__abc_44228_n5187), .Y(u2__abc_44228_n9915) );
  INVX1 INVX1_2342 ( .A(u2__abc_44228_n9916), .Y(u2__abc_44228_n9917) );
  INVX1 INVX1_2343 ( .A(u2__abc_44228_n9925), .Y(u2__abc_44228_n9926) );
  INVX1 INVX1_2344 ( .A(u2__abc_44228_n9934), .Y(u2__abc_44228_n9935_1) );
  INVX1 INVX1_2345 ( .A(u2__abc_44228_n9942), .Y(u2__abc_44228_n9943) );
  INVX1 INVX1_2346 ( .A(u2__abc_44228_n5158), .Y(u2__abc_44228_n9951_1) );
  INVX1 INVX1_2347 ( .A(u2__abc_44228_n9949), .Y(u2__abc_44228_n9952_1) );
  INVX1 INVX1_2348 ( .A(u2__abc_44228_n9959), .Y(u2__abc_44228_n9960) );
  INVX1 INVX1_2349 ( .A(u2__abc_44228_n9967), .Y(u2__abc_44228_n9968_1) );
  INVX1 INVX1_235 ( .A(u2__abc_44228_n3206), .Y(u2__abc_44228_n3207) );
  INVX1 INVX1_2350 ( .A(u2__abc_44228_n9970), .Y(u2__abc_44228_n9971) );
  INVX1 INVX1_2351 ( .A(u2__abc_44228_n9977), .Y(u2__abc_44228_n9978) );
  INVX1 INVX1_2352 ( .A(u2__abc_44228_n5144), .Y(u2__abc_44228_n9984_1) );
  INVX1 INVX1_2353 ( .A(u2__abc_44228_n9985_1), .Y(u2__abc_44228_n9986) );
  INVX1 INVX1_2354 ( .A(u2__abc_44228_n9994), .Y(u2__abc_44228_n9995_1) );
  INVX1 INVX1_2355 ( .A(u2__abc_44228_n10004), .Y(u2__abc_44228_n10005) );
  INVX1 INVX1_2356 ( .A(u2__abc_44228_n10011), .Y(u2__abc_44228_n10012_1) );
  INVX1 INVX1_2357 ( .A(u2__abc_44228_n5127_1), .Y(u2__abc_44228_n10018_1) );
  INVX1 INVX1_2358 ( .A(u2__abc_44228_n10019), .Y(u2__abc_44228_n10020) );
  INVX1 INVX1_2359 ( .A(u2__abc_44228_n10028_1), .Y(u2__abc_44228_n10029_1) );
  INVX1 INVX1_236 ( .A(sqrto_26_), .Y(u2__abc_44228_n3209) );
  INVX1 INVX1_2360 ( .A(u2__abc_44228_n10038), .Y(u2__abc_44228_n10039_1) );
  INVX1 INVX1_2361 ( .A(u2__abc_44228_n10045_1), .Y(u2__abc_44228_n10046) );
  INVX1 INVX1_2362 ( .A(u2__abc_44228_n5113), .Y(u2__abc_44228_n10054) );
  INVX1 INVX1_2363 ( .A(u2__abc_44228_n10052), .Y(u2__abc_44228_n10055) );
  INVX1 INVX1_2364 ( .A(u2__abc_44228_n10062_1), .Y(u2__abc_44228_n10063) );
  INVX1 INVX1_2365 ( .A(u2__abc_44228_n10070), .Y(u2__abc_44228_n10071) );
  INVX1 INVX1_2366 ( .A(u2__abc_44228_n10072_1), .Y(u2__abc_44228_n10073_1) );
  INVX1 INVX1_2367 ( .A(u2__abc_44228_n10080), .Y(u2__abc_44228_n10081) );
  INVX1 INVX1_2368 ( .A(u2__abc_44228_n10087), .Y(u2__abc_44228_n10088) );
  INVX1 INVX1_2369 ( .A(u2__abc_44228_n5104), .Y(u2__abc_44228_n10090) );
  INVX1 INVX1_237 ( .A(u2_remHi_26_), .Y(u2__abc_44228_n3211) );
  INVX1 INVX1_2370 ( .A(u2__abc_44228_n10097), .Y(u2__abc_44228_n10098) );
  INVX1 INVX1_2371 ( .A(u2__abc_44228_n10105_1), .Y(u2__abc_44228_n10106_1) );
  INVX1 INVX1_2372 ( .A(u2__abc_44228_n10108), .Y(u2__abc_44228_n10109) );
  INVX1 INVX1_2373 ( .A(u2__abc_44228_n10115), .Y(u2__abc_44228_n10116_1) );
  INVX1 INVX1_2374 ( .A(u2__abc_44228_n5084), .Y(u2__abc_44228_n10122_1) );
  INVX1 INVX1_2375 ( .A(u2__abc_44228_n10123), .Y(u2__abc_44228_n10124) );
  INVX1 INVX1_2376 ( .A(u2__abc_44228_n10132), .Y(u2__abc_44228_n10133_1) );
  INVX1 INVX1_2377 ( .A(u2__abc_44228_n10142), .Y(u2__abc_44228_n10143) );
  INVX1 INVX1_2378 ( .A(u2__abc_44228_n10149_1), .Y(u2__abc_44228_n10150_1) );
  INVX1 INVX1_2379 ( .A(u2__abc_44228_n5074), .Y(u2__abc_44228_n10158) );
  INVX1 INVX1_238 ( .A(u2__abc_44228_n3213), .Y(u2__abc_44228_n3214) );
  INVX1 INVX1_2380 ( .A(u2__abc_44228_n10156), .Y(u2__abc_44228_n10159) );
  INVX1 INVX1_2381 ( .A(u2__abc_44228_n10166_1), .Y(u2__abc_44228_n10167) );
  INVX1 INVX1_2382 ( .A(u2__abc_44228_n10174), .Y(u2__abc_44228_n10175) );
  INVX1 INVX1_2383 ( .A(u2__abc_44228_n10177_1), .Y(u2__abc_44228_n10178) );
  INVX1 INVX1_2384 ( .A(u2__abc_44228_n10184), .Y(u2__abc_44228_n10185) );
  INVX1 INVX1_2385 ( .A(u2__abc_44228_n5054), .Y(u2__abc_44228_n10191) );
  INVX1 INVX1_2386 ( .A(u2__abc_44228_n10192), .Y(u2__abc_44228_n10193_1) );
  INVX1 INVX1_2387 ( .A(u2__abc_44228_n10201), .Y(u2__abc_44228_n10202) );
  INVX1 INVX1_2388 ( .A(u2__abc_44228_n10210_1), .Y(u2__abc_44228_n10211) );
  INVX1 INVX1_2389 ( .A(u2__abc_44228_n10218), .Y(u2__abc_44228_n10219) );
  INVX1 INVX1_239 ( .A(sqrto_27_), .Y(u2__abc_44228_n3215) );
  INVX1 INVX1_2390 ( .A(u2__abc_44228_n5039), .Y(u2__abc_44228_n10225) );
  INVX1 INVX1_2391 ( .A(u2__abc_44228_n10226_1), .Y(u2__abc_44228_n10228) );
  INVX1 INVX1_2392 ( .A(u2__abc_44228_n10235), .Y(u2__abc_44228_n10236) );
  INVX1 INVX1_2393 ( .A(u2__abc_44228_n10245), .Y(u2__abc_44228_n10246) );
  INVX1 INVX1_2394 ( .A(u2__abc_44228_n10252), .Y(u2__abc_44228_n10253) );
  INVX1 INVX1_2395 ( .A(u2__abc_44228_n5025), .Y(u2__abc_44228_n10259_1) );
  INVX1 INVX1_2396 ( .A(u2__abc_44228_n10260_1), .Y(u2__abc_44228_n10261) );
  INVX1 INVX1_2397 ( .A(u2__abc_44228_n10269), .Y(u2__abc_44228_n10270_1) );
  INVX1 INVX1_2398 ( .A(u2__abc_44228_n10280), .Y(u2__abc_44228_n10281_1) );
  INVX1 INVX1_2399 ( .A(u2__abc_44228_n10286), .Y(u2__abc_44228_n10287_1) );
  INVX1 INVX1_24 ( .A(_abc_64468_n1588), .Y(_abc_64468_n1594) );
  INVX1 INVX1_240 ( .A(u2__abc_44228_n3216), .Y(u2__abc_44228_n3217) );
  INVX1 INVX1_2400 ( .A(u2__abc_44228_n5013), .Y(u2__abc_44228_n10293_1) );
  INVX1 INVX1_2401 ( .A(u2__abc_44228_n10294), .Y(u2__abc_44228_n10295) );
  INVX1 INVX1_2402 ( .A(u2__abc_44228_n10303_1), .Y(u2__abc_44228_n10304_1) );
  INVX1 INVX1_2403 ( .A(u2__abc_44228_n10313), .Y(u2__abc_44228_n10314_1) );
  INVX1 INVX1_2404 ( .A(u2__abc_44228_n10320_1), .Y(u2__abc_44228_n10321) );
  INVX1 INVX1_2405 ( .A(u2__abc_44228_n4993), .Y(u2__abc_44228_n10329) );
  INVX1 INVX1_2406 ( .A(u2__abc_44228_n10327), .Y(u2__abc_44228_n10330) );
  INVX1 INVX1_2407 ( .A(u2__abc_44228_n10337), .Y(u2__abc_44228_n10338) );
  INVX1 INVX1_2408 ( .A(u2__abc_44228_n10346_1), .Y(u2__abc_44228_n10347_1) );
  INVX1 INVX1_2409 ( .A(u2__abc_44228_n10354_1), .Y(u2__abc_44228_n10355) );
  INVX1 INVX1_241 ( .A(u2_remHi_27_), .Y(u2__abc_44228_n3218) );
  INVX1 INVX1_2410 ( .A(u2__abc_44228_n4984), .Y(u2__abc_44228_n10363) );
  INVX1 INVX1_2411 ( .A(u2__abc_44228_n10361_1), .Y(u2__abc_44228_n10364) );
  INVX1 INVX1_2412 ( .A(u2__abc_44228_n10371), .Y(u2__abc_44228_n10372) );
  INVX1 INVX1_2413 ( .A(u2__abc_44228_n10379), .Y(u2__abc_44228_n10380) );
  INVX1 INVX1_2414 ( .A(u2__abc_44228_n10382_1), .Y(u2__abc_44228_n10383) );
  INVX1 INVX1_2415 ( .A(u2__abc_44228_n10389_1), .Y(u2__abc_44228_n10390) );
  INVX1 INVX1_2416 ( .A(u2__abc_44228_n4964), .Y(u2__abc_44228_n10396_1) );
  INVX1 INVX1_2417 ( .A(u2__abc_44228_n10397), .Y(u2__abc_44228_n10398) );
  INVX1 INVX1_2418 ( .A(u2__abc_44228_n10406), .Y(u2__abc_44228_n10407) );
  INVX1 INVX1_2419 ( .A(u2__abc_44228_n10416_1), .Y(u2__abc_44228_n10417_1) );
  INVX1 INVX1_242 ( .A(u2__abc_44228_n3219), .Y(u2__abc_44228_n3220) );
  INVX1 INVX1_2420 ( .A(u2__abc_44228_n10423_1), .Y(u2__abc_44228_n10424_1) );
  INVX1 INVX1_2421 ( .A(u2__abc_44228_n4954), .Y(u2__abc_44228_n10432) );
  INVX1 INVX1_2422 ( .A(u2__abc_44228_n10430_1), .Y(u2__abc_44228_n10433) );
  INVX1 INVX1_2423 ( .A(u2__abc_44228_n10440), .Y(u2__abc_44228_n10441) );
  INVX1 INVX1_2424 ( .A(u2__abc_44228_n10448), .Y(u2__abc_44228_n10449) );
  INVX1 INVX1_2425 ( .A(u2__abc_44228_n10451_1), .Y(u2__abc_44228_n10452_1) );
  INVX1 INVX1_2426 ( .A(u2__abc_44228_n10458_1), .Y(u2__abc_44228_n10459_1) );
  INVX1 INVX1_2427 ( .A(u2__abc_44228_n4934), .Y(u2__abc_44228_n10465_1) );
  INVX1 INVX1_2428 ( .A(u2__abc_44228_n10466_1), .Y(u2__abc_44228_n10467) );
  INVX1 INVX1_2429 ( .A(u2__abc_44228_n10475), .Y(u2__abc_44228_n10476) );
  INVX1 INVX1_243 ( .A(sqrto_23_), .Y(u2__abc_44228_n3224) );
  INVX1 INVX1_2430 ( .A(u2__abc_44228_n10484), .Y(u2__abc_44228_n10485) );
  INVX1 INVX1_2431 ( .A(u2__abc_44228_n10492), .Y(u2__abc_44228_n10493_1) );
  INVX1 INVX1_2432 ( .A(u2__abc_44228_n10499), .Y(u2__abc_44228_n10500_1) );
  INVX1 INVX1_2433 ( .A(u2__abc_44228_n4925), .Y(u2__abc_44228_n10502) );
  INVX1 INVX1_2434 ( .A(u2__abc_44228_n10509), .Y(u2__abc_44228_n10510) );
  INVX1 INVX1_2435 ( .A(u2__abc_44228_n10517), .Y(u2__abc_44228_n10518) );
  INVX1 INVX1_2436 ( .A(u2__abc_44228_n10520), .Y(u2__abc_44228_n10521_1) );
  INVX1 INVX1_2437 ( .A(u2__abc_44228_n10527), .Y(u2__abc_44228_n10528_1) );
  INVX1 INVX1_2438 ( .A(u2__abc_44228_n4905), .Y(u2__abc_44228_n10534) );
  INVX1 INVX1_2439 ( .A(u2__abc_44228_n10535_1), .Y(u2__abc_44228_n10536_1) );
  INVX1 INVX1_244 ( .A(u2__abc_44228_n3225), .Y(u2__abc_44228_n3226) );
  INVX1 INVX1_2440 ( .A(u2__abc_44228_n10544), .Y(u2__abc_44228_n10545) );
  INVX1 INVX1_2441 ( .A(u2__abc_44228_n10553), .Y(u2__abc_44228_n10554) );
  INVX1 INVX1_2442 ( .A(u2__abc_44228_n10561), .Y(u2__abc_44228_n10562) );
  INVX1 INVX1_2443 ( .A(u2__abc_44228_n10568), .Y(u2__abc_44228_n10569) );
  INVX1 INVX1_2444 ( .A(u2__abc_44228_n4888), .Y(u2__abc_44228_n10571_1) );
  INVX1 INVX1_2445 ( .A(u2__abc_44228_n10578_1), .Y(u2__abc_44228_n10579) );
  INVX1 INVX1_2446 ( .A(u2__abc_44228_n10588), .Y(u2__abc_44228_n10589) );
  INVX1 INVX1_2447 ( .A(u2__abc_44228_n10595), .Y(u2__abc_44228_n10596) );
  INVX1 INVX1_2448 ( .A(u2__abc_44228_n4874), .Y(u2__abc_44228_n10602) );
  INVX1 INVX1_2449 ( .A(u2__abc_44228_n10603), .Y(u2__abc_44228_n10604) );
  INVX1 INVX1_245 ( .A(u2_remHi_23_), .Y(u2__abc_44228_n3227) );
  INVX1 INVX1_2450 ( .A(u2__abc_44228_n10612_1), .Y(u2__abc_44228_n10613_1) );
  INVX1 INVX1_2451 ( .A(u2__abc_44228_n10621), .Y(u2__abc_44228_n10622) );
  INVX1 INVX1_2452 ( .A(u2__abc_44228_n10629), .Y(u2__abc_44228_n10630) );
  INVX1 INVX1_2453 ( .A(u2__abc_44228_n4859), .Y(u2__abc_44228_n10636) );
  INVX1 INVX1_2454 ( .A(u2__abc_44228_n10637), .Y(u2__abc_44228_n10639) );
  INVX1 INVX1_2455 ( .A(u2__abc_44228_n10646), .Y(u2__abc_44228_n10647_1) );
  INVX1 INVX1_2456 ( .A(u2__abc_44228_n10656), .Y(u2__abc_44228_n10657) );
  INVX1 INVX1_2457 ( .A(u2__abc_44228_n10663), .Y(u2__abc_44228_n10664) );
  INVX1 INVX1_2458 ( .A(u2__abc_44228_n4845), .Y(u2__abc_44228_n10670) );
  INVX1 INVX1_2459 ( .A(u2__abc_44228_n10671), .Y(u2__abc_44228_n10672) );
  INVX1 INVX1_246 ( .A(u2__abc_44228_n3228), .Y(u2__abc_44228_n3229) );
  INVX1 INVX1_2460 ( .A(u2__abc_44228_n10680), .Y(u2__abc_44228_n10681) );
  INVX1 INVX1_2461 ( .A(u2__abc_44228_n10690_1), .Y(u2__abc_44228_n10691) );
  INVX1 INVX1_2462 ( .A(u2__abc_44228_n10697_1), .Y(u2__abc_44228_n10698) );
  INVX1 INVX1_2463 ( .A(u2__abc_44228_n4815), .Y(u2__abc_44228_n10704_1) );
  INVX1 INVX1_2464 ( .A(u2__abc_44228_n10705), .Y(u2__abc_44228_n10707) );
  INVX1 INVX1_2465 ( .A(u2__abc_44228_n10714), .Y(u2__abc_44228_n10715) );
  INVX1 INVX1_2466 ( .A(u2__abc_44228_n10724_1), .Y(u2__abc_44228_n10725_1) );
  INVX1 INVX1_2467 ( .A(u2__abc_44228_n10731_1), .Y(u2__abc_44228_n10732_1) );
  INVX1 INVX1_2468 ( .A(u2__abc_44228_n4829), .Y(u2__abc_44228_n10738_1) );
  INVX1 INVX1_2469 ( .A(u2__abc_44228_n10739_1), .Y(u2__abc_44228_n10741) );
  INVX1 INVX1_247 ( .A(sqrto_22_), .Y(u2__abc_44228_n3231) );
  INVX1 INVX1_2470 ( .A(u2__abc_44228_n10748), .Y(u2__abc_44228_n10749) );
  INVX1 INVX1_2471 ( .A(u2__abc_44228_n10756), .Y(u2__abc_44228_n10757) );
  INVX1 INVX1_2472 ( .A(u2__abc_44228_n10758), .Y(u2__abc_44228_n10759_1) );
  INVX1 INVX1_2473 ( .A(u2__abc_44228_n10766_1), .Y(u2__abc_44228_n10767_1) );
  INVX1 INVX1_2474 ( .A(u2__abc_44228_n4800), .Y(u2__abc_44228_n10773_1) );
  INVX1 INVX1_2475 ( .A(u2__abc_44228_n10774_1), .Y(u2__abc_44228_n10776) );
  INVX1 INVX1_2476 ( .A(u2__abc_44228_n10783), .Y(u2__abc_44228_n10784) );
  INVX1 INVX1_2477 ( .A(u2__abc_44228_n10793), .Y(u2__abc_44228_n10794_1) );
  INVX1 INVX1_2478 ( .A(u2__abc_44228_n10800), .Y(u2__abc_44228_n10801_1) );
  INVX1 INVX1_2479 ( .A(u2__abc_44228_n4786), .Y(u2__abc_44228_n10807) );
  INVX1 INVX1_248 ( .A(u2_remHi_22_), .Y(u2__abc_44228_n3233) );
  INVX1 INVX1_2480 ( .A(u2__abc_44228_n10808_1), .Y(u2__abc_44228_n10809_1) );
  INVX1 INVX1_2481 ( .A(u2__abc_44228_n10817), .Y(u2__abc_44228_n10818) );
  INVX1 INVX1_2482 ( .A(u2__abc_44228_n10827), .Y(u2__abc_44228_n10828) );
  INVX1 INVX1_2483 ( .A(u2__abc_44228_n10834), .Y(u2__abc_44228_n10835) );
  INVX1 INVX1_2484 ( .A(u2__abc_44228_n4773), .Y(u2__abc_44228_n10841) );
  INVX1 INVX1_2485 ( .A(u2__abc_44228_n10842), .Y(u2__abc_44228_n10843_1) );
  INVX1 INVX1_2486 ( .A(u2__abc_44228_n10851_1), .Y(u2__abc_44228_n10852) );
  INVX1 INVX1_2487 ( .A(u2__abc_44228_n10861), .Y(u2__abc_44228_n10862) );
  INVX1 INVX1_2488 ( .A(u2__abc_44228_n10868), .Y(u2__abc_44228_n10869) );
  INVX1 INVX1_2489 ( .A(u2__abc_44228_n10875), .Y(u2__abc_44228_n10876) );
  INVX1 INVX1_249 ( .A(u2__abc_44228_n3235), .Y(u2__abc_44228_n3236) );
  INVX1 INVX1_2490 ( .A(u2__abc_44228_n4753), .Y(u2__abc_44228_n10878_1) );
  INVX1 INVX1_2491 ( .A(u2__abc_44228_n10885_1), .Y(u2__abc_44228_n10886_1) );
  INVX1 INVX1_2492 ( .A(u2__abc_44228_n10894), .Y(u2__abc_44228_n10895) );
  INVX1 INVX1_2493 ( .A(u2__abc_44228_n10902), .Y(u2__abc_44228_n10903) );
  INVX1 INVX1_2494 ( .A(u2__abc_44228_n4738), .Y(u2__abc_44228_n10909) );
  INVX1 INVX1_2495 ( .A(u2__abc_44228_n10910), .Y(u2__abc_44228_n10912) );
  INVX1 INVX1_2496 ( .A(u2__abc_44228_n10919), .Y(u2__abc_44228_n10920_1) );
  INVX1 INVX1_2497 ( .A(u2__abc_44228_n10929), .Y(u2__abc_44228_n10930) );
  INVX1 INVX1_2498 ( .A(u2__abc_44228_n10936), .Y(u2__abc_44228_n10937) );
  INVX1 INVX1_2499 ( .A(u2__abc_44228_n4724), .Y(u2__abc_44228_n10943) );
  INVX1 INVX1_25 ( .A(\a[120] ), .Y(_abc_64468_n1595) );
  INVX1 INVX1_250 ( .A(sqrto_25_), .Y(u2__abc_44228_n3238) );
  INVX1 INVX1_2500 ( .A(u2__abc_44228_n10944), .Y(u2__abc_44228_n10945) );
  INVX1 INVX1_2501 ( .A(u2__abc_44228_n10953), .Y(u2__abc_44228_n10954) );
  INVX1 INVX1_2502 ( .A(u2__abc_44228_n10963_1), .Y(u2__abc_44228_n10964) );
  INVX1 INVX1_2503 ( .A(u2__abc_44228_n10970_1), .Y(u2__abc_44228_n10971) );
  INVX1 INVX1_2504 ( .A(u2__abc_44228_n10977_1), .Y(u2__abc_44228_n10978) );
  INVX1 INVX1_2505 ( .A(u2__abc_44228_n4714), .Y(u2__abc_44228_n10980) );
  INVX1 INVX1_2506 ( .A(u2__abc_44228_n10987), .Y(u2__abc_44228_n10988) );
  INVX1 INVX1_2507 ( .A(u2__abc_44228_n10995), .Y(u2__abc_44228_n10996) );
  INVX1 INVX1_2508 ( .A(u2__abc_44228_n10998_1), .Y(u2__abc_44228_n10999) );
  INVX1 INVX1_2509 ( .A(u2__abc_44228_n11005_1), .Y(u2__abc_44228_n11006) );
  INVX1 INVX1_251 ( .A(u2__abc_44228_n3239), .Y(u2__abc_44228_n3240) );
  INVX1 INVX1_2510 ( .A(u2__abc_44228_n4694), .Y(u2__abc_44228_n11012_1) );
  INVX1 INVX1_2511 ( .A(u2__abc_44228_n11013), .Y(u2__abc_44228_n11014) );
  INVX1 INVX1_2512 ( .A(u2__abc_44228_n11022), .Y(u2__abc_44228_n11023) );
  INVX1 INVX1_2513 ( .A(u2__abc_44228_n11031), .Y(u2__abc_44228_n11032_1) );
  INVX1 INVX1_2514 ( .A(u2__abc_44228_n11039_1), .Y(u2__abc_44228_n11040_1) );
  INVX1 INVX1_2515 ( .A(u2__abc_44228_n4679), .Y(u2__abc_44228_n11046_1) );
  INVX1 INVX1_2516 ( .A(u2__abc_44228_n11047_1), .Y(u2__abc_44228_n11049) );
  INVX1 INVX1_2517 ( .A(u2__abc_44228_n11056), .Y(u2__abc_44228_n11057) );
  INVX1 INVX1_2518 ( .A(u2__abc_44228_n11066), .Y(u2__abc_44228_n11067_1) );
  INVX1 INVX1_2519 ( .A(u2__abc_44228_n11073), .Y(u2__abc_44228_n11074_1) );
  INVX1 INVX1_252 ( .A(u2_remHi_25_), .Y(u2__abc_44228_n3241) );
  INVX1 INVX1_2520 ( .A(u2__abc_44228_n4665_1), .Y(u2__abc_44228_n11080) );
  INVX1 INVX1_2521 ( .A(u2__abc_44228_n11081_1), .Y(u2__abc_44228_n11082_1) );
  INVX1 INVX1_2522 ( .A(u2__abc_44228_n11090), .Y(u2__abc_44228_n11091) );
  INVX1 INVX1_2523 ( .A(u2__abc_44228_n11099), .Y(u2__abc_44228_n11100) );
  INVX1 INVX1_2524 ( .A(u2__abc_44228_n11107), .Y(u2__abc_44228_n11108) );
  INVX1 INVX1_2525 ( .A(u2__abc_44228_n11114), .Y(u2__abc_44228_n11115) );
  INVX1 INVX1_2526 ( .A(u2__abc_44228_n4648), .Y(u2__abc_44228_n11117_1) );
  INVX1 INVX1_2527 ( .A(u2__abc_44228_n11124_1), .Y(u2__abc_44228_n11125) );
  INVX1 INVX1_2528 ( .A(u2__abc_44228_n11134), .Y(u2__abc_44228_n11135) );
  INVX1 INVX1_2529 ( .A(u2__abc_44228_n11141), .Y(u2__abc_44228_n11142) );
  INVX1 INVX1_253 ( .A(u2__abc_44228_n3242), .Y(u2__abc_44228_n3243) );
  INVX1 INVX1_2530 ( .A(u2__abc_44228_n4634), .Y(u2__abc_44228_n11148) );
  INVX1 INVX1_2531 ( .A(u2__abc_44228_n11149), .Y(u2__abc_44228_n11150) );
  INVX1 INVX1_2532 ( .A(u2__abc_44228_n11158_1), .Y(u2__abc_44228_n11159_1) );
  INVX1 INVX1_2533 ( .A(u2__abc_44228_n11167), .Y(u2__abc_44228_n11168) );
  INVX1 INVX1_2534 ( .A(u2__abc_44228_n11175), .Y(u2__abc_44228_n11176) );
  INVX1 INVX1_2535 ( .A(u2__abc_44228_n4625), .Y(u2__abc_44228_n11184) );
  INVX1 INVX1_2536 ( .A(u2__abc_44228_n11182), .Y(u2__abc_44228_n11185) );
  INVX1 INVX1_2537 ( .A(u2__abc_44228_n11192), .Y(u2__abc_44228_n11193_1) );
  INVX1 INVX1_2538 ( .A(u2__abc_44228_n11200_1), .Y(u2__abc_44228_n11201_1) );
  INVX1 INVX1_2539 ( .A(u2__abc_44228_n11203), .Y(u2__abc_44228_n11204) );
  INVX1 INVX1_254 ( .A(sqrto_24_), .Y(u2__abc_44228_n3245) );
  INVX1 INVX1_2540 ( .A(u2__abc_44228_n11210), .Y(u2__abc_44228_n11211) );
  INVX1 INVX1_2541 ( .A(u2__abc_44228_n4605), .Y(u2__abc_44228_n11217) );
  INVX1 INVX1_2542 ( .A(u2__abc_44228_n11218), .Y(u2__abc_44228_n11219) );
  INVX1 INVX1_2543 ( .A(u2__abc_44228_n11227), .Y(u2__abc_44228_n11228_1) );
  INVX1 INVX1_2544 ( .A(u2__abc_44228_n11237), .Y(u2__abc_44228_n11238) );
  INVX1 INVX1_2545 ( .A(u2__abc_44228_n11244), .Y(u2__abc_44228_n11245) );
  INVX1 INVX1_2546 ( .A(u2__abc_44228_n4595), .Y(u2__abc_44228_n11253) );
  INVX1 INVX1_2547 ( .A(u2__abc_44228_n11251), .Y(u2__abc_44228_n11254) );
  INVX1 INVX1_2548 ( .A(u2__abc_44228_n11261), .Y(u2__abc_44228_n11262) );
  INVX1 INVX1_2549 ( .A(u2__abc_44228_n11269), .Y(u2__abc_44228_n11270_1) );
  INVX1 INVX1_255 ( .A(u2_remHi_24_), .Y(u2__abc_44228_n3247) );
  INVX1 INVX1_2550 ( .A(u2__abc_44228_n11272), .Y(u2__abc_44228_n11273) );
  INVX1 INVX1_2551 ( .A(u2__abc_44228_n11279), .Y(u2__abc_44228_n11280) );
  INVX1 INVX1_2552 ( .A(u2__abc_44228_n4575), .Y(u2__abc_44228_n11286) );
  INVX1 INVX1_2553 ( .A(u2__abc_44228_n11287), .Y(u2__abc_44228_n11288) );
  INVX1 INVX1_2554 ( .A(u2__abc_44228_n11296), .Y(u2__abc_44228_n11297) );
  INVX1 INVX1_2555 ( .A(u2__abc_44228_n11305_1), .Y(u2__abc_44228_n11306_1) );
  INVX1 INVX1_2556 ( .A(u2__abc_44228_n11313_1), .Y(u2__abc_44228_n11314) );
  INVX1 INVX1_2557 ( .A(u2__abc_44228_n11320_1), .Y(u2__abc_44228_n11321) );
  INVX1 INVX1_2558 ( .A(u2__abc_44228_n4566), .Y(u2__abc_44228_n11323) );
  INVX1 INVX1_2559 ( .A(u2__abc_44228_n11330), .Y(u2__abc_44228_n11331) );
  INVX1 INVX1_256 ( .A(u2__abc_44228_n3249), .Y(u2__abc_44228_n3250) );
  INVX1 INVX1_2560 ( .A(u2__abc_44228_n11338), .Y(u2__abc_44228_n11339) );
  INVX1 INVX1_2561 ( .A(u2__abc_44228_n11341_1), .Y(u2__abc_44228_n11342) );
  INVX1 INVX1_2562 ( .A(u2__abc_44228_n11348_1), .Y(u2__abc_44228_n11349) );
  INVX1 INVX1_2563 ( .A(u2__abc_44228_n4546), .Y(u2__abc_44228_n11355_1) );
  INVX1 INVX1_2564 ( .A(u2__abc_44228_n11356), .Y(u2__abc_44228_n11357) );
  INVX1 INVX1_2565 ( .A(u2__abc_44228_n11365), .Y(u2__abc_44228_n11366) );
  INVX1 INVX1_2566 ( .A(u2__abc_44228_n11375_1), .Y(u2__abc_44228_n11376_1) );
  INVX1 INVX1_2567 ( .A(u2__abc_44228_n11382_1), .Y(u2__abc_44228_n11383_1) );
  INVX1 INVX1_2568 ( .A(u2__abc_44228_n4534), .Y(u2__abc_44228_n11389_1) );
  INVX1 INVX1_2569 ( .A(u2__abc_44228_n11390_1), .Y(u2__abc_44228_n11392) );
  INVX1 INVX1_257 ( .A(sqrto_21_), .Y(u2__abc_44228_n3254) );
  INVX1 INVX1_2570 ( .A(u2__abc_44228_n11399), .Y(u2__abc_44228_n11400) );
  INVX1 INVX1_2571 ( .A(u2__abc_44228_n11409), .Y(u2__abc_44228_n11410_1) );
  INVX1 INVX1_2572 ( .A(u2__abc_44228_n11416), .Y(u2__abc_44228_n11417_1) );
  INVX1 INVX1_2573 ( .A(u2__abc_44228_n4514), .Y(u2__abc_44228_n11423) );
  INVX1 INVX1_2574 ( .A(u2__abc_44228_n11424_1), .Y(u2__abc_44228_n11425_1) );
  INVX1 INVX1_2575 ( .A(u2__abc_44228_n11433), .Y(u2__abc_44228_n11434) );
  INVX1 INVX1_2576 ( .A(u2__abc_44228_n11442), .Y(u2__abc_44228_n11443) );
  INVX1 INVX1_2577 ( .A(u2__abc_44228_n11450), .Y(u2__abc_44228_n11451) );
  INVX1 INVX1_2578 ( .A(u2__abc_44228_n11457), .Y(u2__abc_44228_n11458) );
  INVX1 INVX1_2579 ( .A(u2__abc_44228_n4505), .Y(u2__abc_44228_n11460_1) );
  INVX1 INVX1_258 ( .A(u2__abc_44228_n3255), .Y(u2__abc_44228_n3256) );
  INVX1 INVX1_2580 ( .A(u2__abc_44228_n11467_1), .Y(u2__abc_44228_n11468) );
  INVX1 INVX1_2581 ( .A(u2__abc_44228_n11475), .Y(u2__abc_44228_n11476) );
  INVX1 INVX1_2582 ( .A(u2__abc_44228_n11478), .Y(u2__abc_44228_n11479) );
  INVX1 INVX1_2583 ( .A(u2__abc_44228_n11485), .Y(u2__abc_44228_n11486) );
  INVX1 INVX1_2584 ( .A(u2__abc_44228_n4485), .Y(u2__abc_44228_n11492) );
  INVX1 INVX1_2585 ( .A(u2__abc_44228_n11493), .Y(u2__abc_44228_n11494_1) );
  INVX1 INVX1_2586 ( .A(u2__abc_44228_n11502_1), .Y(u2__abc_44228_n11503) );
  INVX1 INVX1_2587 ( .A(u2__abc_44228_n11512), .Y(u2__abc_44228_n11513) );
  INVX1 INVX1_2588 ( .A(u2__abc_44228_n11519), .Y(u2__abc_44228_n11520) );
  INVX1 INVX1_2589 ( .A(u2__abc_44228_n4455), .Y(u2__abc_44228_n11526) );
  INVX1 INVX1_259 ( .A(u2_remHi_21_), .Y(u2__abc_44228_n3257) );
  INVX1 INVX1_2590 ( .A(u2__abc_44228_n11527), .Y(u2__abc_44228_n11529_1) );
  INVX1 INVX1_2591 ( .A(u2__abc_44228_n11536_1), .Y(u2__abc_44228_n11537_1) );
  INVX1 INVX1_2592 ( .A(u2__abc_44228_n11546), .Y(u2__abc_44228_n11547) );
  INVX1 INVX1_2593 ( .A(u2__abc_44228_n11553), .Y(u2__abc_44228_n11554) );
  INVX1 INVX1_2594 ( .A(u2__abc_44228_n4469), .Y(u2__abc_44228_n11560) );
  INVX1 INVX1_2595 ( .A(u2__abc_44228_n11561), .Y(u2__abc_44228_n11563) );
  INVX1 INVX1_2596 ( .A(u2__abc_44228_n11570), .Y(u2__abc_44228_n11571_1) );
  INVX1 INVX1_2597 ( .A(u2__abc_44228_n11578_1), .Y(u2__abc_44228_n11579_1) );
  INVX1 INVX1_2598 ( .A(u2__abc_44228_n11580), .Y(u2__abc_44228_n11581) );
  INVX1 INVX1_2599 ( .A(u2__abc_44228_n11588), .Y(u2__abc_44228_n11589) );
  INVX1 INVX1_26 ( .A(_abc_64468_n1598), .Y(_abc_64468_n1599) );
  INVX1 INVX1_260 ( .A(u2__abc_44228_n3258), .Y(u2__abc_44228_n3259) );
  INVX1 INVX1_2600 ( .A(u2__abc_44228_n11595), .Y(u2__abc_44228_n11596) );
  INVX1 INVX1_2601 ( .A(u2__abc_44228_n4446), .Y(u2__abc_44228_n11598) );
  INVX1 INVX1_2602 ( .A(u2__abc_44228_n11605), .Y(u2__abc_44228_n11606_1) );
  INVX1 INVX1_2603 ( .A(u2__abc_44228_n11613_1), .Y(u2__abc_44228_n11614_1) );
  INVX1 INVX1_2604 ( .A(u2__abc_44228_n11615), .Y(u2__abc_44228_n11616) );
  INVX1 INVX1_2605 ( .A(u2__abc_44228_n11623), .Y(u2__abc_44228_n11624) );
  INVX1 INVX1_2606 ( .A(u2__abc_44228_n4426), .Y(u2__abc_44228_n11630) );
  INVX1 INVX1_2607 ( .A(u2__abc_44228_n11631), .Y(u2__abc_44228_n11632) );
  INVX1 INVX1_2608 ( .A(u2__abc_44228_n11640), .Y(u2__abc_44228_n11641_1) );
  INVX1 INVX1_2609 ( .A(u2__abc_44228_n11649_1), .Y(u2__abc_44228_n11650) );
  INVX1 INVX1_261 ( .A(sqrto_20_), .Y(u2__abc_44228_n3261) );
  INVX1 INVX1_2610 ( .A(u2__abc_44228_n11657), .Y(u2__abc_44228_n11658) );
  INVX1 INVX1_2611 ( .A(u2__abc_44228_n4415), .Y(u2__abc_44228_n11664) );
  INVX1 INVX1_2612 ( .A(u2__abc_44228_n11665), .Y(u2__abc_44228_n11667) );
  INVX1 INVX1_2613 ( .A(u2__abc_44228_n11674_1), .Y(u2__abc_44228_n11675) );
  INVX1 INVX1_2614 ( .A(u2__abc_44228_n11682), .Y(u2__abc_44228_n11683) );
  INVX1 INVX1_2615 ( .A(u2__abc_44228_n11685), .Y(u2__abc_44228_n11686) );
  INVX1 INVX1_2616 ( .A(u2__abc_44228_n11692), .Y(u2__abc_44228_n11693) );
  INVX1 INVX1_2617 ( .A(u2__abc_44228_n4395), .Y(u2__abc_44228_n11699) );
  INVX1 INVX1_2618 ( .A(u2__abc_44228_n11700), .Y(u2__abc_44228_n11701) );
  INVX1 INVX1_2619 ( .A(u2__abc_44228_n11709), .Y(u2__abc_44228_n11710) );
  INVX1 INVX1_262 ( .A(u2_remHi_20_), .Y(u2__abc_44228_n3263) );
  INVX1 INVX1_2620 ( .A(u2__abc_44228_n11718), .Y(u2__abc_44228_n11719_1) );
  INVX1 INVX1_2621 ( .A(u2__abc_44228_n11726_1), .Y(u2__abc_44228_n11727) );
  INVX1 INVX1_2622 ( .A(u2__abc_44228_n11733), .Y(u2__abc_44228_n11734_1) );
  INVX1 INVX1_2623 ( .A(u2__abc_44228_n4386_1), .Y(u2__abc_44228_n11736) );
  INVX1 INVX1_2624 ( .A(u2__abc_44228_n11743), .Y(u2__abc_44228_n11744) );
  INVX1 INVX1_2625 ( .A(u2__abc_44228_n11751), .Y(u2__abc_44228_n11752) );
  INVX1 INVX1_2626 ( .A(u2__abc_44228_n11754), .Y(u2__abc_44228_n11755) );
  INVX1 INVX1_2627 ( .A(u2__abc_44228_n11761), .Y(u2__abc_44228_n11762) );
  INVX1 INVX1_2628 ( .A(u2__abc_44228_n4366), .Y(u2__abc_44228_n11768) );
  INVX1 INVX1_2629 ( .A(u2__abc_44228_n11769), .Y(u2__abc_44228_n11770) );
  INVX1 INVX1_263 ( .A(u2__abc_44228_n3265), .Y(u2__abc_44228_n3266) );
  INVX1 INVX1_2630 ( .A(u2__abc_44228_n11778), .Y(u2__abc_44228_n11779) );
  INVX1 INVX1_2631 ( .A(u2__abc_44228_n11788_1), .Y(u2__abc_44228_n11789) );
  INVX1 INVX1_2632 ( .A(u2__abc_44228_n11795), .Y(u2__abc_44228_n11796_1) );
  INVX1 INVX1_2633 ( .A(u2__abc_44228_n4356), .Y(u2__abc_44228_n11804) );
  INVX1 INVX1_2634 ( .A(u2__abc_44228_n11802), .Y(u2__abc_44228_n11805) );
  INVX1 INVX1_2635 ( .A(u2__abc_44228_n11812), .Y(u2__abc_44228_n11813_1) );
  INVX1 INVX1_2636 ( .A(u2__abc_44228_n11820_1), .Y(u2__abc_44228_n11821) );
  INVX1 INVX1_2637 ( .A(u2__abc_44228_n11823), .Y(u2__abc_44228_n11824) );
  INVX1 INVX1_2638 ( .A(u2__abc_44228_n11830), .Y(u2__abc_44228_n11831) );
  INVX1 INVX1_2639 ( .A(u2__abc_44228_n4336), .Y(u2__abc_44228_n11837) );
  INVX1 INVX1_264 ( .A(sqrto_18_), .Y(u2__abc_44228_n3268) );
  INVX1 INVX1_2640 ( .A(u2__abc_44228_n11838), .Y(u2__abc_44228_n11839) );
  INVX1 INVX1_2641 ( .A(u2__abc_44228_n11847), .Y(u2__abc_44228_n11848) );
  INVX1 INVX1_2642 ( .A(u2__abc_44228_n11856), .Y(u2__abc_44228_n11857) );
  INVX1 INVX1_2643 ( .A(u2__abc_44228_n11864), .Y(u2__abc_44228_n11865) );
  INVX1 INVX1_2644 ( .A(u2__abc_44228_n4327), .Y(u2__abc_44228_n11873) );
  INVX1 INVX1_2645 ( .A(u2__abc_44228_n11871), .Y(u2__abc_44228_n11874) );
  INVX1 INVX1_2646 ( .A(u2__abc_44228_n11881), .Y(u2__abc_44228_n11882) );
  INVX1 INVX1_2647 ( .A(u2__abc_44228_n11889), .Y(u2__abc_44228_n11890) );
  INVX1 INVX1_2648 ( .A(u2__abc_44228_n11892), .Y(u2__abc_44228_n11893) );
  INVX1 INVX1_2649 ( .A(u2__abc_44228_n11899), .Y(u2__abc_44228_n11900) );
  INVX1 INVX1_265 ( .A(u2_remHi_18_), .Y(u2__abc_44228_n3270) );
  INVX1 INVX1_2650 ( .A(u2__abc_44228_n4307), .Y(u2__abc_44228_n11906) );
  INVX1 INVX1_2651 ( .A(u2__abc_44228_n11907_1), .Y(u2__abc_44228_n11908) );
  INVX1 INVX1_2652 ( .A(u2__abc_44228_n11916), .Y(u2__abc_44228_n11917) );
  INVX1 INVX1_2653 ( .A(u2__abc_44228_n11925), .Y(u2__abc_44228_n11926) );
  INVX1 INVX1_2654 ( .A(u2__abc_44228_n11931), .Y(u2__abc_44228_n11932) );
  INVX1 INVX1_2655 ( .A(u2__abc_44228_n6518), .Y(u2__abc_44228_n11939) );
  INVX1 INVX1_2656 ( .A(u2__abc_44228_n11940_1), .Y(u2__abc_44228_n11941) );
  INVX1 INVX1_2657 ( .A(u2__abc_44228_n11948), .Y(u2__abc_44228_n11949) );
  INVX1 INVX1_2658 ( .A(u2__abc_44228_n11957), .Y(u2__abc_44228_n11958) );
  INVX1 INVX1_2659 ( .A(u2__abc_44228_n11965), .Y(u2__abc_44228_n11966) );
  INVX1 INVX1_266 ( .A(u2__abc_44228_n3272), .Y(u2__abc_44228_n3273) );
  INVX1 INVX1_2660 ( .A(u2__abc_44228_n6504), .Y(u2__abc_44228_n11974) );
  INVX1 INVX1_2661 ( .A(u2__abc_44228_n11972), .Y(u2__abc_44228_n11975) );
  INVX1 INVX1_2662 ( .A(u2__abc_44228_n11982), .Y(u2__abc_44228_n11983) );
  INVX1 INVX1_2663 ( .A(u2__abc_44228_n11992), .Y(u2__abc_44228_n11993_1) );
  INVX1 INVX1_2664 ( .A(u2__abc_44228_n11999), .Y(u2__abc_44228_n12000) );
  INVX1 INVX1_2665 ( .A(u2__abc_44228_n6489_1), .Y(u2__abc_44228_n12006) );
  INVX1 INVX1_2666 ( .A(u2__abc_44228_n12007), .Y(u2__abc_44228_n12009) );
  INVX1 INVX1_2667 ( .A(u2__abc_44228_n12016), .Y(u2__abc_44228_n12017) );
  INVX1 INVX1_2668 ( .A(u2__abc_44228_n12025_1), .Y(u2__abc_44228_n12026) );
  INVX1 INVX1_2669 ( .A(u2__abc_44228_n12033), .Y(u2__abc_44228_n12034_1) );
  INVX1 INVX1_267 ( .A(sqrto_19_), .Y(u2__abc_44228_n3274) );
  INVX1 INVX1_2670 ( .A(u2__abc_44228_n6475), .Y(u2__abc_44228_n12040) );
  INVX1 INVX1_2671 ( .A(u2__abc_44228_n12041_1), .Y(u2__abc_44228_n12042) );
  INVX1 INVX1_2672 ( .A(u2__abc_44228_n12050), .Y(u2__abc_44228_n12051) );
  INVX1 INVX1_2673 ( .A(u2__abc_44228_n12059), .Y(u2__abc_44228_n12060) );
  INVX1 INVX1_2674 ( .A(u2__abc_44228_n12067_1), .Y(u2__abc_44228_n12068) );
  INVX1 INVX1_2675 ( .A(u2__abc_44228_n6459), .Y(u2__abc_44228_n12074_1) );
  INVX1 INVX1_2676 ( .A(u2__abc_44228_n12075), .Y(u2__abc_44228_n12077) );
  INVX1 INVX1_2677 ( .A(u2__abc_44228_n12084), .Y(u2__abc_44228_n12085) );
  INVX1 INVX1_2678 ( .A(u2__abc_44228_n12092), .Y(u2__abc_44228_n12093) );
  INVX1 INVX1_2679 ( .A(u2__abc_44228_n12094), .Y(u2__abc_44228_n12095) );
  INVX1 INVX1_268 ( .A(u2__abc_44228_n3275), .Y(u2__abc_44228_n3276) );
  INVX1 INVX1_2680 ( .A(u2__abc_44228_n12102), .Y(u2__abc_44228_n12103) );
  INVX1 INVX1_2681 ( .A(u2__abc_44228_n6445_1), .Y(u2__abc_44228_n12109) );
  INVX1 INVX1_2682 ( .A(u2__abc_44228_n12110), .Y(u2__abc_44228_n12111) );
  INVX1 INVX1_2683 ( .A(u2__abc_44228_n12119), .Y(u2__abc_44228_n12120_1) );
  INVX1 INVX1_2684 ( .A(u2__abc_44228_n12129), .Y(u2__abc_44228_n12130_1) );
  INVX1 INVX1_2685 ( .A(u2__abc_44228_n12136), .Y(u2__abc_44228_n12137_1) );
  INVX1 INVX1_2686 ( .A(u2__abc_44228_n6430), .Y(u2__abc_44228_n12143) );
  INVX1 INVX1_2687 ( .A(u2__abc_44228_n12144), .Y(u2__abc_44228_n12146) );
  INVX1 INVX1_2688 ( .A(u2__abc_44228_n12153), .Y(u2__abc_44228_n12154) );
  INVX1 INVX1_2689 ( .A(u2__abc_44228_n12162), .Y(u2__abc_44228_n12163) );
  INVX1 INVX1_269 ( .A(u2_remHi_19_), .Y(u2__abc_44228_n3277) );
  INVX1 INVX1_2690 ( .A(u2__abc_44228_n12170), .Y(u2__abc_44228_n12171) );
  INVX1 INVX1_2691 ( .A(u2__abc_44228_n6416), .Y(u2__abc_44228_n12177) );
  INVX1 INVX1_2692 ( .A(u2__abc_44228_n12178), .Y(u2__abc_44228_n12179) );
  INVX1 INVX1_2693 ( .A(u2__abc_44228_n12187), .Y(u2__abc_44228_n12188) );
  INVX1 INVX1_2694 ( .A(u2__abc_44228_n12197), .Y(u2__abc_44228_n12198) );
  INVX1 INVX1_2695 ( .A(u2__abc_44228_n12204), .Y(u2__abc_44228_n12205) );
  INVX1 INVX1_2696 ( .A(u2__abc_44228_n6405), .Y(u2__abc_44228_n12211) );
  INVX1 INVX1_2697 ( .A(u2__abc_44228_n12212), .Y(u2__abc_44228_n12214) );
  INVX1 INVX1_2698 ( .A(u2__abc_44228_n12221), .Y(u2__abc_44228_n12222) );
  INVX1 INVX1_2699 ( .A(u2__abc_44228_n12229), .Y(u2__abc_44228_n12230) );
  INVX1 INVX1_27 ( .A(_abc_64468_n1600), .Y(_abc_64468_n1601) );
  INVX1 INVX1_270 ( .A(u2__abc_44228_n3278), .Y(u2__abc_44228_n3279) );
  INVX1 INVX1_2700 ( .A(u2__abc_44228_n12231), .Y(u2__abc_44228_n12232) );
  INVX1 INVX1_2701 ( .A(u2__abc_44228_n12239), .Y(u2__abc_44228_n12240) );
  INVX1 INVX1_2702 ( .A(u2__abc_44228_n6385), .Y(u2__abc_44228_n12246) );
  INVX1 INVX1_2703 ( .A(u2__abc_44228_n12247), .Y(u2__abc_44228_n12248_1) );
  INVX1 INVX1_2704 ( .A(u2__abc_44228_n12256), .Y(u2__abc_44228_n12257) );
  INVX1 INVX1_2705 ( .A(u2__abc_44228_n12266), .Y(u2__abc_44228_n12267) );
  INVX1 INVX1_2706 ( .A(u2__abc_44228_n12273_1), .Y(u2__abc_44228_n12274) );
  INVX1 INVX1_2707 ( .A(u2__abc_44228_n6370), .Y(u2__abc_44228_n12280_1) );
  INVX1 INVX1_2708 ( .A(u2__abc_44228_n12281), .Y(u2__abc_44228_n12283) );
  INVX1 INVX1_2709 ( .A(u2__abc_44228_n12290), .Y(u2__abc_44228_n12291) );
  INVX1 INVX1_271 ( .A(u2_remHi_17_), .Y(u2__abc_44228_n3283) );
  INVX1 INVX1_2710 ( .A(u2__abc_44228_n12299), .Y(u2__abc_44228_n12300) );
  INVX1 INVX1_2711 ( .A(u2__abc_44228_n12307), .Y(u2__abc_44228_n12308) );
  INVX1 INVX1_2712 ( .A(u2__abc_44228_n6356), .Y(u2__abc_44228_n12314) );
  INVX1 INVX1_2713 ( .A(u2__abc_44228_n12315), .Y(u2__abc_44228_n12316) );
  INVX1 INVX1_2714 ( .A(u2__abc_44228_n12324), .Y(u2__abc_44228_n12325) );
  INVX1 INVX1_2715 ( .A(u2__abc_44228_n12333), .Y(u2__abc_44228_n12334) );
  INVX1 INVX1_2716 ( .A(u2__abc_44228_n12341), .Y(u2__abc_44228_n12342) );
  INVX1 INVX1_2717 ( .A(u2__abc_44228_n6326), .Y(u2__abc_44228_n12348) );
  INVX1 INVX1_2718 ( .A(u2__abc_44228_n12349), .Y(u2__abc_44228_n12351) );
  INVX1 INVX1_2719 ( .A(u2__abc_44228_n12358), .Y(u2__abc_44228_n12359) );
  INVX1 INVX1_272 ( .A(sqrto_17_), .Y(u2__abc_44228_n3285) );
  INVX1 INVX1_2720 ( .A(u2__abc_44228_n12367), .Y(u2__abc_44228_n12368_1) );
  INVX1 INVX1_2721 ( .A(u2__abc_44228_n12375_1), .Y(u2__abc_44228_n12376) );
  INVX1 INVX1_2722 ( .A(u2__abc_44228_n6340), .Y(u2__abc_44228_n12382) );
  INVX1 INVX1_2723 ( .A(u2__abc_44228_n12383), .Y(u2__abc_44228_n12385_1) );
  INVX1 INVX1_2724 ( .A(u2__abc_44228_n12392_1), .Y(u2__abc_44228_n12393) );
  INVX1 INVX1_2725 ( .A(u2__abc_44228_n12400_1), .Y(u2__abc_44228_n12401) );
  INVX1 INVX1_2726 ( .A(u2__abc_44228_n12403), .Y(u2__abc_44228_n12404) );
  INVX1 INVX1_2727 ( .A(u2__abc_44228_n12410), .Y(u2__abc_44228_n12411) );
  INVX1 INVX1_2728 ( .A(u2__abc_44228_n6311), .Y(u2__abc_44228_n12419) );
  INVX1 INVX1_2729 ( .A(u2__abc_44228_n12417), .Y(u2__abc_44228_n12420) );
  INVX1 INVX1_273 ( .A(u2_remHi_16_), .Y(u2__abc_44228_n3288) );
  INVX1 INVX1_2730 ( .A(u2__abc_44228_n12427), .Y(u2__abc_44228_n12428) );
  INVX1 INVX1_2731 ( .A(u2__abc_44228_n12435), .Y(u2__abc_44228_n12436) );
  INVX1 INVX1_2732 ( .A(u2__abc_44228_n12437), .Y(u2__abc_44228_n12438_1) );
  INVX1 INVX1_2733 ( .A(u2__abc_44228_n12445), .Y(u2__abc_44228_n12446) );
  INVX1 INVX1_2734 ( .A(u2__abc_44228_n6297), .Y(u2__abc_44228_n12452) );
  INVX1 INVX1_2735 ( .A(u2__abc_44228_n12453), .Y(u2__abc_44228_n12454) );
  INVX1 INVX1_2736 ( .A(u2__abc_44228_n12462), .Y(u2__abc_44228_n12463) );
  INVX1 INVX1_2737 ( .A(u2__abc_44228_n12471), .Y(u2__abc_44228_n12472_1) );
  INVX1 INVX1_2738 ( .A(u2__abc_44228_n12479), .Y(u2__abc_44228_n12480) );
  INVX1 INVX1_2739 ( .A(u2__abc_44228_n6279_1), .Y(u2__abc_44228_n12486) );
  INVX1 INVX1_274 ( .A(sqrto_16_), .Y(u2__abc_44228_n3290) );
  INVX1 INVX1_2740 ( .A(u2__abc_44228_n12487), .Y(u2__abc_44228_n12489) );
  INVX1 INVX1_2741 ( .A(u2__abc_44228_n12496_1), .Y(u2__abc_44228_n12497) );
  INVX1 INVX1_2742 ( .A(u2__abc_44228_n12505), .Y(u2__abc_44228_n12506) );
  INVX1 INVX1_2743 ( .A(u2__abc_44228_n12513_1), .Y(u2__abc_44228_n12514) );
  INVX1 INVX1_2744 ( .A(u2__abc_44228_n6265), .Y(u2__abc_44228_n12520_1) );
  INVX1 INVX1_2745 ( .A(u2__abc_44228_n12521), .Y(u2__abc_44228_n12522) );
  INVX1 INVX1_2746 ( .A(u2__abc_44228_n12530), .Y(u2__abc_44228_n12531) );
  INVX1 INVX1_2747 ( .A(u2__abc_44228_n12540), .Y(u2__abc_44228_n12541) );
  INVX1 INVX1_2748 ( .A(u2__abc_44228_n12547), .Y(u2__abc_44228_n12548) );
  INVX1 INVX1_2749 ( .A(u2__abc_44228_n6250), .Y(u2__abc_44228_n12554) );
  INVX1 INVX1_275 ( .A(sqrto_15_), .Y(u2__abc_44228_n3294) );
  INVX1 INVX1_2750 ( .A(u2__abc_44228_n12555), .Y(u2__abc_44228_n12557) );
  INVX1 INVX1_2751 ( .A(u2__abc_44228_n12564), .Y(u2__abc_44228_n12565) );
  INVX1 INVX1_2752 ( .A(u2__abc_44228_n12573), .Y(u2__abc_44228_n12574) );
  INVX1 INVX1_2753 ( .A(u2__abc_44228_n12581), .Y(u2__abc_44228_n12582) );
  INVX1 INVX1_2754 ( .A(u2__abc_44228_n6236), .Y(u2__abc_44228_n12588) );
  INVX1 INVX1_2755 ( .A(u2__abc_44228_n12589), .Y(u2__abc_44228_n12590) );
  INVX1 INVX1_2756 ( .A(u2__abc_44228_n12598), .Y(u2__abc_44228_n12599_1) );
  INVX1 INVX1_2757 ( .A(u2__abc_44228_n12607), .Y(u2__abc_44228_n12608_1) );
  INVX1 INVX1_2758 ( .A(u2__abc_44228_n12615_1), .Y(u2__abc_44228_n12616) );
  INVX1 INVX1_2759 ( .A(u2__abc_44228_n6206_1), .Y(u2__abc_44228_n12622) );
  INVX1 INVX1_276 ( .A(u2__abc_44228_n3295), .Y(u2__abc_44228_n3296) );
  INVX1 INVX1_2760 ( .A(u2__abc_44228_n12623_1), .Y(u2__abc_44228_n12625) );
  INVX1 INVX1_2761 ( .A(u2__abc_44228_n12632), .Y(u2__abc_44228_n12633) );
  INVX1 INVX1_2762 ( .A(u2__abc_44228_n12641), .Y(u2__abc_44228_n12642) );
  INVX1 INVX1_2763 ( .A(u2__abc_44228_n12649), .Y(u2__abc_44228_n12650) );
  INVX1 INVX1_2764 ( .A(u2__abc_44228_n6220), .Y(u2__abc_44228_n12656) );
  INVX1 INVX1_2765 ( .A(u2__abc_44228_n12657), .Y(u2__abc_44228_n12659) );
  INVX1 INVX1_2766 ( .A(u2__abc_44228_n12666), .Y(u2__abc_44228_n12667) );
  INVX1 INVX1_2767 ( .A(u2__abc_44228_n12674), .Y(u2__abc_44228_n12675) );
  INVX1 INVX1_2768 ( .A(u2__abc_44228_n12677), .Y(u2__abc_44228_n12678_1) );
  INVX1 INVX1_2769 ( .A(u2__abc_44228_n12684), .Y(u2__abc_44228_n12685) );
  INVX1 INVX1_277 ( .A(u2_remHi_15_), .Y(u2__abc_44228_n3297) );
  INVX1 INVX1_2770 ( .A(u2__abc_44228_n12691), .Y(u2__abc_44228_n12692) );
  INVX1 INVX1_2771 ( .A(u2__abc_44228_n6191), .Y(u2__abc_44228_n12694) );
  INVX1 INVX1_2772 ( .A(u2__abc_44228_n12701), .Y(u2__abc_44228_n12702) );
  INVX1 INVX1_2773 ( .A(u2__abc_44228_n12709), .Y(u2__abc_44228_n12710) );
  INVX1 INVX1_2774 ( .A(u2__abc_44228_n12711), .Y(u2__abc_44228_n12712) );
  INVX1 INVX1_2775 ( .A(u2__abc_44228_n12719), .Y(u2__abc_44228_n12720) );
  INVX1 INVX1_2776 ( .A(u2__abc_44228_n6177), .Y(u2__abc_44228_n12726) );
  INVX1 INVX1_2777 ( .A(u2__abc_44228_n12727), .Y(u2__abc_44228_n12728_1) );
  INVX1 INVX1_2778 ( .A(u2__abc_44228_n12736), .Y(u2__abc_44228_n12737_1) );
  INVX1 INVX1_2779 ( .A(u2__abc_44228_n12746), .Y(u2__abc_44228_n12747) );
  INVX1 INVX1_278 ( .A(u2__abc_44228_n3298), .Y(u2__abc_44228_n3299) );
  INVX1 INVX1_2780 ( .A(u2__abc_44228_n12753), .Y(u2__abc_44228_n12754) );
  INVX1 INVX1_2781 ( .A(u2__abc_44228_n6166), .Y(u2__abc_44228_n12762) );
  INVX1 INVX1_2782 ( .A(u2__abc_44228_n12763), .Y(u2__abc_44228_n12765) );
  INVX1 INVX1_2783 ( .A(u2__abc_44228_n12770), .Y(u2__abc_44228_n12771) );
  INVX1 INVX1_2784 ( .A(u2__abc_44228_n12779), .Y(u2__abc_44228_n12780) );
  INVX1 INVX1_2785 ( .A(u2__abc_44228_n12787), .Y(u2__abc_44228_n12788) );
  INVX1 INVX1_2786 ( .A(u2__abc_44228_n6146), .Y(u2__abc_44228_n12794) );
  INVX1 INVX1_2787 ( .A(u2__abc_44228_n12795), .Y(u2__abc_44228_n12796) );
  INVX1 INVX1_2788 ( .A(u2__abc_44228_n12804), .Y(u2__abc_44228_n12805) );
  INVX1 INVX1_2789 ( .A(u2__abc_44228_n12814), .Y(u2__abc_44228_n12815_1) );
  INVX1 INVX1_279 ( .A(sqrto_14_), .Y(u2__abc_44228_n3301) );
  INVX1 INVX1_2790 ( .A(u2__abc_44228_n12821), .Y(u2__abc_44228_n12822_1) );
  INVX1 INVX1_2791 ( .A(u2__abc_44228_n6137), .Y(u2__abc_44228_n12830) );
  INVX1 INVX1_2792 ( .A(u2__abc_44228_n12831), .Y(u2__abc_44228_n12833_1) );
  INVX1 INVX1_2793 ( .A(u2__abc_44228_n12838), .Y(u2__abc_44228_n12839) );
  INVX1 INVX1_2794 ( .A(u2__abc_44228_n12847), .Y(u2__abc_44228_n12848_1) );
  INVX1 INVX1_2795 ( .A(u2__abc_44228_n12855_1), .Y(u2__abc_44228_n12856) );
  INVX1 INVX1_2796 ( .A(u2__abc_44228_n6117), .Y(u2__abc_44228_n12862) );
  INVX1 INVX1_2797 ( .A(u2__abc_44228_n12863), .Y(u2__abc_44228_n12864_1) );
  INVX1 INVX1_2798 ( .A(u2__abc_44228_n12872), .Y(u2__abc_44228_n12873) );
  INVX1 INVX1_2799 ( .A(u2__abc_44228_n12881), .Y(u2__abc_44228_n12882) );
  INVX1 INVX1_28 ( .A(_abc_64468_n1603), .Y(_abc_64468_n1607) );
  INVX1 INVX1_280 ( .A(u2_remHi_14_), .Y(u2__abc_44228_n3303) );
  INVX1 INVX1_2800 ( .A(u2__abc_44228_n12889), .Y(u2__abc_44228_n12890) );
  INVX1 INVX1_2801 ( .A(u2__abc_44228_n6101), .Y(u2__abc_44228_n12898) );
  INVX1 INVX1_2802 ( .A(u2__abc_44228_n12899), .Y(u2__abc_44228_n12901) );
  INVX1 INVX1_2803 ( .A(u2__abc_44228_n12906), .Y(u2__abc_44228_n12907) );
  INVX1 INVX1_2804 ( .A(u2__abc_44228_n12915), .Y(u2__abc_44228_n12916) );
  INVX1 INVX1_2805 ( .A(u2__abc_44228_n12923), .Y(u2__abc_44228_n12924) );
  INVX1 INVX1_2806 ( .A(u2__abc_44228_n6087), .Y(u2__abc_44228_n12930) );
  INVX1 INVX1_2807 ( .A(u2__abc_44228_n12931), .Y(u2__abc_44228_n12933) );
  INVX1 INVX1_2808 ( .A(u2__abc_44228_n12940), .Y(u2__abc_44228_n12941) );
  INVX1 INVX1_2809 ( .A(u2__abc_44228_n12948), .Y(u2__abc_44228_n12949_1) );
  INVX1 INVX1_281 ( .A(u2__abc_44228_n3305), .Y(u2__abc_44228_n3306) );
  INVX1 INVX1_2810 ( .A(u2__abc_44228_n12950), .Y(u2__abc_44228_n12951) );
  INVX1 INVX1_2811 ( .A(u2__abc_44228_n12958), .Y(u2__abc_44228_n12959) );
  INVX1 INVX1_2812 ( .A(u2__abc_44228_n6072), .Y(u2__abc_44228_n12965) );
  INVX1 INVX1_2813 ( .A(u2__abc_44228_n12966), .Y(u2__abc_44228_n12968_1) );
  INVX1 INVX1_2814 ( .A(u2__abc_44228_n12975), .Y(u2__abc_44228_n12976_1) );
  INVX1 INVX1_2815 ( .A(u2__abc_44228_n12984), .Y(u2__abc_44228_n12985) );
  INVX1 INVX1_2816 ( .A(u2__abc_44228_n12992_1), .Y(u2__abc_44228_n12993) );
  INVX1 INVX1_2817 ( .A(u2__abc_44228_n6058), .Y(u2__abc_44228_n12999_1) );
  INVX1 INVX1_2818 ( .A(u2__abc_44228_n13000), .Y(u2__abc_44228_n13001) );
  INVX1 INVX1_2819 ( .A(u2__abc_44228_n13009), .Y(u2__abc_44228_n13010) );
  INVX1 INVX1_282 ( .A(u2__abc_44228_n3284), .Y(u2__abc_44228_n3315) );
  INVX1 INVX1_2820 ( .A(u2__abc_44228_n13018), .Y(u2__abc_44228_n13019) );
  INVX1 INVX1_2821 ( .A(u2__abc_44228_n13026), .Y(u2__abc_44228_n13027) );
  INVX1 INVX1_2822 ( .A(u2__abc_44228_n6045), .Y(u2__abc_44228_n13035) );
  INVX1 INVX1_2823 ( .A(u2__abc_44228_n13033), .Y(u2__abc_44228_n13036) );
  INVX1 INVX1_2824 ( .A(u2__abc_44228_n13043), .Y(u2__abc_44228_n13044) );
  INVX1 INVX1_2825 ( .A(u2__abc_44228_n13051), .Y(u2__abc_44228_n13052) );
  INVX1 INVX1_2826 ( .A(u2__abc_44228_n13053), .Y(u2__abc_44228_n13054) );
  INVX1 INVX1_2827 ( .A(u2__abc_44228_n13061), .Y(u2__abc_44228_n13062_1) );
  INVX1 INVX1_2828 ( .A(u2__abc_44228_n6025), .Y(u2__abc_44228_n13068) );
  INVX1 INVX1_2829 ( .A(u2__abc_44228_n13069), .Y(u2__abc_44228_n13070_1) );
  INVX1 INVX1_283 ( .A(u2__abc_44228_n3289), .Y(u2__abc_44228_n3316) );
  INVX1 INVX1_2830 ( .A(u2__abc_44228_n13078), .Y(u2__abc_44228_n13079) );
  INVX1 INVX1_2831 ( .A(u2__abc_44228_n13088_1), .Y(u2__abc_44228_n13089) );
  INVX1 INVX1_2832 ( .A(u2__abc_44228_n13095_1), .Y(u2__abc_44228_n13096) );
  INVX1 INVX1_2833 ( .A(u2__abc_44228_n13102), .Y(u2__abc_44228_n13103_1) );
  INVX1 INVX1_2834 ( .A(u2__abc_44228_n6016), .Y(u2__abc_44228_n13105) );
  INVX1 INVX1_2835 ( .A(u2__abc_44228_n13112), .Y(u2__abc_44228_n13113) );
  INVX1 INVX1_2836 ( .A(u2__abc_44228_n13120), .Y(u2__abc_44228_n13121) );
  INVX1 INVX1_2837 ( .A(u2__abc_44228_n13122), .Y(u2__abc_44228_n13123) );
  INVX1 INVX1_2838 ( .A(u2__abc_44228_n13130), .Y(u2__abc_44228_n13131) );
  INVX1 INVX1_2839 ( .A(u2__abc_44228_n5996), .Y(u2__abc_44228_n13137) );
  INVX1 INVX1_284 ( .A(u2__abc_44228_n3246), .Y(u2__abc_44228_n3332) );
  INVX1 INVX1_2840 ( .A(u2__abc_44228_n13138), .Y(u2__abc_44228_n13139) );
  INVX1 INVX1_2841 ( .A(u2__abc_44228_n13147), .Y(u2__abc_44228_n13148) );
  INVX1 INVX1_2842 ( .A(u2__abc_44228_n13156), .Y(u2__abc_44228_n13157) );
  INVX1 INVX1_2843 ( .A(u2__abc_44228_n13164), .Y(u2__abc_44228_n13165) );
  INVX1 INVX1_2844 ( .A(u2__abc_44228_n5980), .Y(u2__abc_44228_n13173_1) );
  INVX1 INVX1_2845 ( .A(u2__abc_44228_n13171), .Y(u2__abc_44228_n13174) );
  INVX1 INVX1_2846 ( .A(u2__abc_44228_n13181), .Y(u2__abc_44228_n13182_1) );
  INVX1 INVX1_2847 ( .A(u2__abc_44228_n13189_1), .Y(u2__abc_44228_n13190) );
  INVX1 INVX1_2848 ( .A(u2__abc_44228_n13191), .Y(u2__abc_44228_n13192) );
  INVX1 INVX1_2849 ( .A(u2__abc_44228_n13199), .Y(u2__abc_44228_n13200) );
  INVX1 INVX1_285 ( .A(u2__abc_44228_n3333), .Y(u2__abc_44228_n3334) );
  INVX1 INVX1_2850 ( .A(u2__abc_44228_n5966_1), .Y(u2__abc_44228_n13206) );
  INVX1 INVX1_2851 ( .A(u2__abc_44228_n13207), .Y(u2__abc_44228_n13208) );
  INVX1 INVX1_2852 ( .A(u2__abc_44228_n13216), .Y(u2__abc_44228_n13217_1) );
  INVX1 INVX1_2853 ( .A(u2__abc_44228_n13226), .Y(u2__abc_44228_n13227) );
  INVX1 INVX1_2854 ( .A(u2__abc_44228_n13233), .Y(u2__abc_44228_n13234) );
  INVX1 INVX1_2855 ( .A(u2__abc_44228_n5951), .Y(u2__abc_44228_n13242) );
  INVX1 INVX1_2856 ( .A(u2__abc_44228_n13240), .Y(u2__abc_44228_n13243) );
  INVX1 INVX1_2857 ( .A(u2__abc_44228_n13250), .Y(u2__abc_44228_n13251) );
  INVX1 INVX1_2858 ( .A(u2__abc_44228_n13258), .Y(u2__abc_44228_n13259) );
  INVX1 INVX1_2859 ( .A(u2__abc_44228_n13260), .Y(u2__abc_44228_n13261) );
  INVX1 INVX1_286 ( .A(u2__abc_44228_n3210), .Y(u2__abc_44228_n3338) );
  INVX1 INVX1_2860 ( .A(u2__abc_44228_n13268), .Y(u2__abc_44228_n13269) );
  INVX1 INVX1_2861 ( .A(u2__abc_44228_n5937), .Y(u2__abc_44228_n13275) );
  INVX1 INVX1_2862 ( .A(u2__abc_44228_n13276), .Y(u2__abc_44228_n13277) );
  INVX1 INVX1_2863 ( .A(u2__abc_44228_n13285), .Y(u2__abc_44228_n13286) );
  INVX1 INVX1_2864 ( .A(u2__abc_44228_n13295_1), .Y(u2__abc_44228_n13296) );
  INVX1 INVX1_2865 ( .A(u2__abc_44228_n13302_1), .Y(u2__abc_44228_n13303) );
  INVX1 INVX1_2866 ( .A(u2__abc_44228_n5920_1), .Y(u2__abc_44228_n13309) );
  INVX1 INVX1_2867 ( .A(u2__abc_44228_n13310), .Y(u2__abc_44228_n13312) );
  INVX1 INVX1_2868 ( .A(u2__abc_44228_n13319), .Y(u2__abc_44228_n13320) );
  INVX1 INVX1_2869 ( .A(u2__abc_44228_n13328), .Y(u2__abc_44228_n13329) );
  INVX1 INVX1_287 ( .A(u2__abc_44228_n3339), .Y(u2__abc_44228_n3340) );
  INVX1 INVX1_2870 ( .A(u2__abc_44228_n13336), .Y(u2__abc_44228_n13337) );
  INVX1 INVX1_2871 ( .A(u2__abc_44228_n5906), .Y(u2__abc_44228_n13343) );
  INVX1 INVX1_2872 ( .A(u2__abc_44228_n13344_1), .Y(u2__abc_44228_n13345) );
  INVX1 INVX1_2873 ( .A(u2__abc_44228_n13353), .Y(u2__abc_44228_n13354) );
  INVX1 INVX1_2874 ( .A(u2__abc_44228_n13363), .Y(u2__abc_44228_n13364) );
  INVX1 INVX1_2875 ( .A(u2__abc_44228_n13370), .Y(u2__abc_44228_n13371) );
  INVX1 INVX1_2876 ( .A(u2__abc_44228_n5897), .Y(u2__abc_44228_n13379) );
  INVX1 INVX1_2877 ( .A(u2__abc_44228_n13377), .Y(u2__abc_44228_n13380) );
  INVX1 INVX1_2878 ( .A(u2__abc_44228_n13387), .Y(u2__abc_44228_n13388) );
  INVX1 INVX1_2879 ( .A(u2__abc_44228_n13395), .Y(u2__abc_44228_n13396) );
  INVX1 INVX1_288 ( .A(sqrto_61_), .Y(u2__abc_44228_n3349) );
  INVX1 INVX1_2880 ( .A(u2__abc_44228_n13397_1), .Y(u2__abc_44228_n13398) );
  INVX1 INVX1_2881 ( .A(u2__abc_44228_n13405), .Y(u2__abc_44228_n13406) );
  INVX1 INVX1_2882 ( .A(u2__abc_44228_n5877), .Y(u2__abc_44228_n13412) );
  INVX1 INVX1_2883 ( .A(u2__abc_44228_n13413), .Y(u2__abc_44228_n13414_1) );
  INVX1 INVX1_2884 ( .A(u2__abc_44228_n13422_1), .Y(u2__abc_44228_n13423) );
  INVX1 INVX1_2885 ( .A(u2__abc_44228_n13431), .Y(u2__abc_44228_n13432) );
  INVX1 INVX1_2886 ( .A(u2__abc_44228_n13439), .Y(u2__abc_44228_n13440) );
  INVX1 INVX1_2887 ( .A(u2__abc_44228_n5847), .Y(u2__abc_44228_n13446) );
  INVX1 INVX1_2888 ( .A(u2__abc_44228_n13447), .Y(u2__abc_44228_n13449) );
  INVX1 INVX1_2889 ( .A(u2__abc_44228_n13456), .Y(u2__abc_44228_n13457) );
  INVX1 INVX1_289 ( .A(u2__abc_44228_n3350), .Y(u2__abc_44228_n3351) );
  INVX1 INVX1_2890 ( .A(u2__abc_44228_n13465), .Y(u2__abc_44228_n13466) );
  INVX1 INVX1_2891 ( .A(u2__abc_44228_n13473), .Y(u2__abc_44228_n13474) );
  INVX1 INVX1_2892 ( .A(u2__abc_44228_n5861), .Y(u2__abc_44228_n13480) );
  INVX1 INVX1_2893 ( .A(u2__abc_44228_n13481), .Y(u2__abc_44228_n13483) );
  INVX1 INVX1_2894 ( .A(u2__abc_44228_n13490), .Y(u2__abc_44228_n13491) );
  INVX1 INVX1_2895 ( .A(u2__abc_44228_n13498), .Y(u2__abc_44228_n13499) );
  INVX1 INVX1_2896 ( .A(u2__abc_44228_n13501), .Y(u2__abc_44228_n13502) );
  INVX1 INVX1_2897 ( .A(u2__abc_44228_n13508), .Y(u2__abc_44228_n13509) );
  INVX1 INVX1_2898 ( .A(u2__abc_44228_n13515), .Y(u2__abc_44228_n13516) );
  INVX1 INVX1_2899 ( .A(u2__abc_44228_n5838_1), .Y(u2__abc_44228_n13518_1) );
  INVX1 INVX1_29 ( .A(\a[121] ), .Y(_abc_64468_n1608) );
  INVX1 INVX1_290 ( .A(u2_remHi_61_), .Y(u2__abc_44228_n3352) );
  INVX1 INVX1_2900 ( .A(u2__abc_44228_n13525_1), .Y(u2__abc_44228_n13526) );
  INVX1 INVX1_2901 ( .A(u2__abc_44228_n13533), .Y(u2__abc_44228_n13534) );
  INVX1 INVX1_2902 ( .A(u2__abc_44228_n13535_1), .Y(u2__abc_44228_n13536) );
  INVX1 INVX1_2903 ( .A(u2__abc_44228_n13543), .Y(u2__abc_44228_n13544) );
  INVX1 INVX1_2904 ( .A(u2__abc_44228_n5818), .Y(u2__abc_44228_n13550_1) );
  INVX1 INVX1_2905 ( .A(u2__abc_44228_n13551), .Y(u2__abc_44228_n13552) );
  INVX1 INVX1_2906 ( .A(u2__abc_44228_n13560), .Y(u2__abc_44228_n13561) );
  INVX1 INVX1_2907 ( .A(u2__abc_44228_n13569), .Y(u2__abc_44228_n13570) );
  INVX1 INVX1_2908 ( .A(u2__abc_44228_n13577), .Y(u2__abc_44228_n13578) );
  INVX1 INVX1_2909 ( .A(u2__abc_44228_n5800), .Y(u2__abc_44228_n13584) );
  INVX1 INVX1_291 ( .A(u2__abc_44228_n3353), .Y(u2__abc_44228_n3354) );
  INVX1 INVX1_2910 ( .A(u2__abc_44228_n13585), .Y(u2__abc_44228_n13587) );
  INVX1 INVX1_2911 ( .A(u2__abc_44228_n13594), .Y(u2__abc_44228_n13595) );
  INVX1 INVX1_2912 ( .A(u2__abc_44228_n13603), .Y(u2__abc_44228_n13604) );
  INVX1 INVX1_2913 ( .A(u2__abc_44228_n13611), .Y(u2__abc_44228_n13612) );
  INVX1 INVX1_2914 ( .A(u2__abc_44228_n5786), .Y(u2__abc_44228_n13618) );
  INVX1 INVX1_2915 ( .A(u2__abc_44228_n13619), .Y(u2__abc_44228_n13620) );
  INVX1 INVX1_2916 ( .A(u2__abc_44228_n13628), .Y(u2__abc_44228_n13629) );
  INVX1 INVX1_2917 ( .A(u2__abc_44228_n13638), .Y(u2__abc_44228_n13639) );
  INVX1 INVX1_2918 ( .A(u2__abc_44228_n13645_1), .Y(u2__abc_44228_n13646) );
  INVX1 INVX1_2919 ( .A(u2__abc_44228_n5777), .Y(u2__abc_44228_n13654) );
  INVX1 INVX1_292 ( .A(sqrto_60_), .Y(u2__abc_44228_n3356) );
  INVX1 INVX1_2920 ( .A(u2__abc_44228_n13652_1), .Y(u2__abc_44228_n13655) );
  INVX1 INVX1_2921 ( .A(u2__abc_44228_n13662_1), .Y(u2__abc_44228_n13663) );
  INVX1 INVX1_2922 ( .A(u2__abc_44228_n13670), .Y(u2__abc_44228_n13671) );
  INVX1 INVX1_2923 ( .A(u2__abc_44228_n13672), .Y(u2__abc_44228_n13673) );
  INVX1 INVX1_2924 ( .A(u2__abc_44228_n13680), .Y(u2__abc_44228_n13681) );
  INVX1 INVX1_2925 ( .A(u2__abc_44228_n5757), .Y(u2__abc_44228_n13687) );
  INVX1 INVX1_2926 ( .A(u2__abc_44228_n13688), .Y(u2__abc_44228_n13689) );
  INVX1 INVX1_2927 ( .A(u2__abc_44228_n13697), .Y(u2__abc_44228_n13698) );
  INVX1 INVX1_2928 ( .A(u2__abc_44228_n13706), .Y(u2__abc_44228_n13707) );
  INVX1 INVX1_2929 ( .A(u2__abc_44228_n13714), .Y(u2__abc_44228_n13715) );
  INVX1 INVX1_293 ( .A(u2_remHi_60_), .Y(u2__abc_44228_n3358) );
  INVX1 INVX1_2930 ( .A(u2__abc_44228_n5727), .Y(u2__abc_44228_n13721) );
  INVX1 INVX1_2931 ( .A(u2__abc_44228_n13722), .Y(u2__abc_44228_n13724) );
  INVX1 INVX1_2932 ( .A(u2__abc_44228_n13731), .Y(u2__abc_44228_n13732_1) );
  INVX1 INVX1_2933 ( .A(u2__abc_44228_n13740_1), .Y(u2__abc_44228_n13741) );
  INVX1 INVX1_2934 ( .A(u2__abc_44228_n13748), .Y(u2__abc_44228_n13749_1) );
  INVX1 INVX1_2935 ( .A(u2__abc_44228_n5741), .Y(u2__abc_44228_n13755) );
  INVX1 INVX1_2936 ( .A(u2__abc_44228_n13756), .Y(u2__abc_44228_n13758) );
  INVX1 INVX1_2937 ( .A(u2__abc_44228_n13765), .Y(u2__abc_44228_n13766) );
  INVX1 INVX1_2938 ( .A(u2__abc_44228_n13773), .Y(u2__abc_44228_n13774) );
  INVX1 INVX1_2939 ( .A(u2__abc_44228_n13776), .Y(u2__abc_44228_n13777) );
  INVX1 INVX1_294 ( .A(u2__abc_44228_n3360), .Y(u2__abc_44228_n3361) );
  INVX1 INVX1_2940 ( .A(u2__abc_44228_n13783), .Y(u2__abc_44228_n13784_1) );
  INVX1 INVX1_2941 ( .A(u2__abc_44228_n5712), .Y(u2__abc_44228_n13790) );
  INVX1 INVX1_2942 ( .A(u2__abc_44228_n13791), .Y(u2__abc_44228_n13793) );
  INVX1 INVX1_2943 ( .A(u2__abc_44228_n13800), .Y(u2__abc_44228_n13801) );
  INVX1 INVX1_2944 ( .A(u2__abc_44228_n13809), .Y(u2__abc_44228_n13810) );
  INVX1 INVX1_2945 ( .A(u2__abc_44228_n13817), .Y(u2__abc_44228_n13818) );
  INVX1 INVX1_2946 ( .A(u2__abc_44228_n5698), .Y(u2__abc_44228_n13824) );
  INVX1 INVX1_2947 ( .A(u2__abc_44228_n13825), .Y(u2__abc_44228_n13826) );
  INVX1 INVX1_2948 ( .A(u2__abc_44228_n13834), .Y(u2__abc_44228_n13835) );
  INVX1 INVX1_2949 ( .A(u2__abc_44228_n13844), .Y(u2__abc_44228_n13845) );
  INVX1 INVX1_295 ( .A(sqrto_58_), .Y(u2__abc_44228_n3363) );
  INVX1 INVX1_2950 ( .A(u2__abc_44228_n13851), .Y(u2__abc_44228_n13852) );
  INVX1 INVX1_2951 ( .A(u2__abc_44228_n5667), .Y(u2__abc_44228_n13860) );
  INVX1 INVX1_2952 ( .A(u2__abc_44228_n13861), .Y(u2__abc_44228_n13863_1) );
  INVX1 INVX1_2953 ( .A(u2__abc_44228_n13868), .Y(u2__abc_44228_n13869) );
  INVX1 INVX1_2954 ( .A(u2__abc_44228_n13877), .Y(u2__abc_44228_n13878) );
  INVX1 INVX1_2955 ( .A(u2__abc_44228_n13885), .Y(u2__abc_44228_n13886) );
  INVX1 INVX1_2956 ( .A(u2__abc_44228_n5681_1), .Y(u2__abc_44228_n13892_1) );
  INVX1 INVX1_2957 ( .A(u2__abc_44228_n13893), .Y(u2__abc_44228_n13895) );
  INVX1 INVX1_2958 ( .A(u2__abc_44228_n13902), .Y(u2__abc_44228_n13903) );
  INVX1 INVX1_2959 ( .A(u2__abc_44228_n13910_1), .Y(u2__abc_44228_n13911) );
  INVX1 INVX1_296 ( .A(u2_remHi_58_), .Y(u2__abc_44228_n3365) );
  INVX1 INVX1_2960 ( .A(u2__abc_44228_n13912), .Y(u2__abc_44228_n13913) );
  INVX1 INVX1_2961 ( .A(u2__abc_44228_n13920), .Y(u2__abc_44228_n13921) );
  INVX1 INVX1_2962 ( .A(u2__abc_44228_n5658), .Y(u2__abc_44228_n13929) );
  INVX1 INVX1_2963 ( .A(u2__abc_44228_n13927_1), .Y(u2__abc_44228_n13930) );
  INVX1 INVX1_2964 ( .A(u2__abc_44228_n13937), .Y(u2__abc_44228_n13938) );
  INVX1 INVX1_2965 ( .A(u2__abc_44228_n13945), .Y(u2__abc_44228_n13946_1) );
  INVX1 INVX1_2966 ( .A(u2__abc_44228_n13947), .Y(u2__abc_44228_n13948) );
  INVX1 INVX1_2967 ( .A(u2__abc_44228_n13955), .Y(u2__abc_44228_n13956) );
  INVX1 INVX1_2968 ( .A(u2__abc_44228_n5638), .Y(u2__abc_44228_n13962) );
  INVX1 INVX1_2969 ( .A(u2__abc_44228_n13963_1), .Y(u2__abc_44228_n13964) );
  INVX1 INVX1_297 ( .A(u2__abc_44228_n3367), .Y(u2__abc_44228_n3368) );
  INVX1 INVX1_2970 ( .A(u2__abc_44228_n13972), .Y(u2__abc_44228_n13973) );
  INVX1 INVX1_2971 ( .A(u2__abc_44228_n13981_1), .Y(u2__abc_44228_n13982) );
  INVX1 INVX1_2972 ( .A(u2__abc_44228_n13989_1), .Y(u2__abc_44228_n13990) );
  INVX1 INVX1_2973 ( .A(u2__abc_44228_n5608), .Y(u2__abc_44228_n13996) );
  INVX1 INVX1_2974 ( .A(u2__abc_44228_n13997), .Y(u2__abc_44228_n13999) );
  INVX1 INVX1_2975 ( .A(u2__abc_44228_n14006_1), .Y(u2__abc_44228_n14007) );
  INVX1 INVX1_2976 ( .A(u2__abc_44228_n14015), .Y(u2__abc_44228_n14016) );
  INVX1 INVX1_2977 ( .A(u2__abc_44228_n14023), .Y(u2__abc_44228_n14024) );
  INVX1 INVX1_2978 ( .A(u2__abc_44228_n5622), .Y(u2__abc_44228_n14030) );
  INVX1 INVX1_2979 ( .A(u2__abc_44228_n14031), .Y(u2__abc_44228_n14033) );
  INVX1 INVX1_298 ( .A(sqrto_59_), .Y(u2__abc_44228_n3369) );
  INVX1 INVX1_2980 ( .A(u2__abc_44228_n14040), .Y(u2__abc_44228_n14041) );
  INVX1 INVX1_2981 ( .A(u2__abc_44228_n14048), .Y(u2__abc_44228_n14049) );
  INVX1 INVX1_2982 ( .A(u2__abc_44228_n14050), .Y(u2__abc_44228_n14051) );
  INVX1 INVX1_2983 ( .A(u2__abc_44228_n14058), .Y(u2__abc_44228_n14059) );
  INVX1 INVX1_2984 ( .A(u2__abc_44228_n5593), .Y(u2__abc_44228_n14067) );
  INVX1 INVX1_2985 ( .A(u2__abc_44228_n14065), .Y(u2__abc_44228_n14068) );
  INVX1 INVX1_2986 ( .A(u2__abc_44228_n14075), .Y(u2__abc_44228_n14076) );
  INVX1 INVX1_2987 ( .A(u2__abc_44228_n14083), .Y(u2__abc_44228_n14084) );
  INVX1 INVX1_2988 ( .A(u2__abc_44228_n14085), .Y(u2__abc_44228_n14086) );
  INVX1 INVX1_2989 ( .A(u2__abc_44228_n14093), .Y(u2__abc_44228_n14094) );
  INVX1 INVX1_299 ( .A(u2__abc_44228_n3370), .Y(u2__abc_44228_n3371) );
  INVX1 INVX1_2990 ( .A(u2__abc_44228_n5579), .Y(u2__abc_44228_n14100) );
  INVX1 INVX1_2991 ( .A(u2__abc_44228_n14101), .Y(u2__abc_44228_n14102) );
  INVX1 INVX1_2992 ( .A(u2__abc_44228_n14110), .Y(u2__abc_44228_n14111) );
  INVX1 INVX1_2993 ( .A(u2__abc_44228_n14117), .Y(u2__abc_44228_n14118) );
  INVX1 INVX1_2994 ( .A(u2__abc_44228_n14125_1), .Y(u2__abc_44228_n14126) );
  INVX1 INVX1_2995 ( .A(u2__abc_44228_n7332), .Y(u2__abc_44228_n14132) );
  INVX1 INVX1_2996 ( .A(u2__abc_44228_n14133_1), .Y(u2__abc_44228_n14135) );
  INVX1 INVX1_2997 ( .A(u2__abc_44228_n14142_1), .Y(u2__abc_44228_n14143) );
  INVX1 INVX1_2998 ( .A(u2__abc_44228_n14151), .Y(u2__abc_44228_n14152) );
  INVX1 INVX1_2999 ( .A(u2__abc_44228_n14159), .Y(u2__abc_44228_n14160) );
  INVX1 INVX1_3 ( .A(_abc_64468_n1516), .Y(_abc_64468_n1517) );
  INVX1 INVX1_30 ( .A(_abc_64468_n1611), .Y(_abc_64468_n1612) );
  INVX1 INVX1_300 ( .A(u2_remHi_59_), .Y(u2__abc_44228_n3372) );
  INVX1 INVX1_3000 ( .A(u2__abc_44228_n7318), .Y(u2__abc_44228_n14166) );
  INVX1 INVX1_3001 ( .A(u2__abc_44228_n14167), .Y(u2__abc_44228_n14168) );
  INVX1 INVX1_3002 ( .A(u2__abc_44228_n14176), .Y(u2__abc_44228_n14177) );
  INVX1 INVX1_3003 ( .A(u2__abc_44228_n14186), .Y(u2__abc_44228_n14187_1) );
  INVX1 INVX1_3004 ( .A(u2__abc_44228_n14193), .Y(u2__abc_44228_n14194) );
  INVX1 INVX1_3005 ( .A(u2__abc_44228_n14200), .Y(u2__abc_44228_n14201) );
  INVX1 INVX1_3006 ( .A(u2__abc_44228_n7309_1), .Y(u2__abc_44228_n14203) );
  INVX1 INVX1_3007 ( .A(u2__abc_44228_n14210), .Y(u2__abc_44228_n14211) );
  INVX1 INVX1_3008 ( .A(u2__abc_44228_n14218), .Y(u2__abc_44228_n14219) );
  INVX1 INVX1_3009 ( .A(u2__abc_44228_n14220), .Y(u2__abc_44228_n14221) );
  INVX1 INVX1_301 ( .A(u2__abc_44228_n3373), .Y(u2__abc_44228_n3374) );
  INVX1 INVX1_3010 ( .A(u2__abc_44228_n14228), .Y(u2__abc_44228_n14229) );
  INVX1 INVX1_3011 ( .A(u2__abc_44228_n7289_1), .Y(u2__abc_44228_n14235) );
  INVX1 INVX1_3012 ( .A(u2__abc_44228_n14236), .Y(u2__abc_44228_n14237) );
  INVX1 INVX1_3013 ( .A(u2__abc_44228_n14245), .Y(u2__abc_44228_n14246) );
  INVX1 INVX1_3014 ( .A(u2__abc_44228_n14254), .Y(u2__abc_44228_n14255) );
  INVX1 INVX1_3015 ( .A(u2__abc_44228_n14262), .Y(u2__abc_44228_n14263) );
  INVX1 INVX1_3016 ( .A(u2__abc_44228_n7279), .Y(u2__abc_44228_n14269) );
  INVX1 INVX1_3017 ( .A(u2__abc_44228_n14270), .Y(u2__abc_44228_n14272) );
  INVX1 INVX1_3018 ( .A(u2__abc_44228_n14279), .Y(u2__abc_44228_n14280) );
  INVX1 INVX1_3019 ( .A(u2__abc_44228_n14287), .Y(u2__abc_44228_n14288) );
  INVX1 INVX1_302 ( .A(sqrto_57_), .Y(u2__abc_44228_n3378) );
  INVX1 INVX1_3020 ( .A(u2__abc_44228_n14289), .Y(u2__abc_44228_n14290) );
  INVX1 INVX1_3021 ( .A(u2__abc_44228_n14297), .Y(u2__abc_44228_n14298) );
  INVX1 INVX1_3022 ( .A(u2__abc_44228_n7259), .Y(u2__abc_44228_n14304) );
  INVX1 INVX1_3023 ( .A(u2__abc_44228_n14305), .Y(u2__abc_44228_n14306) );
  INVX1 INVX1_3024 ( .A(u2__abc_44228_n14314), .Y(u2__abc_44228_n14315_1) );
  INVX1 INVX1_3025 ( .A(u2__abc_44228_n14324_1), .Y(u2__abc_44228_n14325) );
  INVX1 INVX1_3026 ( .A(u2__abc_44228_n14331), .Y(u2__abc_44228_n14332_1) );
  INVX1 INVX1_3027 ( .A(u2__abc_44228_n7250), .Y(u2__abc_44228_n14340) );
  INVX1 INVX1_3028 ( .A(u2__abc_44228_n14338), .Y(u2__abc_44228_n14341) );
  INVX1 INVX1_3029 ( .A(u2__abc_44228_n14348), .Y(u2__abc_44228_n14349) );
  INVX1 INVX1_303 ( .A(u2__abc_44228_n3379), .Y(u2__abc_44228_n3380) );
  INVX1 INVX1_3030 ( .A(u2__abc_44228_n14356), .Y(u2__abc_44228_n14357) );
  INVX1 INVX1_3031 ( .A(u2__abc_44228_n14358), .Y(u2__abc_44228_n14359_1) );
  INVX1 INVX1_3032 ( .A(u2__abc_44228_n14366), .Y(u2__abc_44228_n14367_1) );
  INVX1 INVX1_3033 ( .A(u2__abc_44228_n7230), .Y(u2__abc_44228_n14373) );
  INVX1 INVX1_3034 ( .A(u2__abc_44228_n14374), .Y(u2__abc_44228_n14375) );
  INVX1 INVX1_3035 ( .A(u2__abc_44228_n14383), .Y(u2__abc_44228_n14384) );
  INVX1 INVX1_3036 ( .A(u2__abc_44228_n14393), .Y(u2__abc_44228_n14394) );
  INVX1 INVX1_3037 ( .A(u2__abc_44228_n14400), .Y(u2__abc_44228_n14401) );
  INVX1 INVX1_3038 ( .A(u2__abc_44228_n7219), .Y(u2__abc_44228_n14409) );
  INVX1 INVX1_3039 ( .A(u2__abc_44228_n14407), .Y(u2__abc_44228_n14410) );
  INVX1 INVX1_304 ( .A(u2_remHi_57_), .Y(u2__abc_44228_n3381) );
  INVX1 INVX1_3040 ( .A(u2__abc_44228_n14417), .Y(u2__abc_44228_n14418) );
  INVX1 INVX1_3041 ( .A(u2__abc_44228_n14425), .Y(u2__abc_44228_n14426) );
  INVX1 INVX1_3042 ( .A(u2__abc_44228_n14427), .Y(u2__abc_44228_n14428) );
  INVX1 INVX1_3043 ( .A(u2__abc_44228_n14435), .Y(u2__abc_44228_n14436) );
  INVX1 INVX1_3044 ( .A(u2__abc_44228_n7199), .Y(u2__abc_44228_n14442) );
  INVX1 INVX1_3045 ( .A(u2__abc_44228_n14443), .Y(u2__abc_44228_n14444) );
  INVX1 INVX1_3046 ( .A(u2__abc_44228_n14452), .Y(u2__abc_44228_n14453) );
  INVX1 INVX1_3047 ( .A(u2__abc_44228_n14462), .Y(u2__abc_44228_n14463) );
  INVX1 INVX1_3048 ( .A(u2__abc_44228_n14469), .Y(u2__abc_44228_n14470) );
  INVX1 INVX1_3049 ( .A(u2__abc_44228_n7184), .Y(u2__abc_44228_n14476) );
  INVX1 INVX1_305 ( .A(u2__abc_44228_n3382), .Y(u2__abc_44228_n3383) );
  INVX1 INVX1_3050 ( .A(u2__abc_44228_n14477), .Y(u2__abc_44228_n14479) );
  INVX1 INVX1_3051 ( .A(u2__abc_44228_n14486), .Y(u2__abc_44228_n14487) );
  INVX1 INVX1_3052 ( .A(u2__abc_44228_n14495), .Y(u2__abc_44228_n14496) );
  INVX1 INVX1_3053 ( .A(u2__abc_44228_n14503), .Y(u2__abc_44228_n14504) );
  INVX1 INVX1_3054 ( .A(u2__abc_44228_n7170_1), .Y(u2__abc_44228_n14510_1) );
  INVX1 INVX1_3055 ( .A(u2__abc_44228_n14511), .Y(u2__abc_44228_n14512) );
  INVX1 INVX1_3056 ( .A(u2__abc_44228_n14520), .Y(u2__abc_44228_n14521_1) );
  INVX1 INVX1_3057 ( .A(u2__abc_44228_n14529_1), .Y(u2__abc_44228_n14530) );
  INVX1 INVX1_3058 ( .A(u2__abc_44228_n14537), .Y(u2__abc_44228_n14538_1) );
  INVX1 INVX1_3059 ( .A(u2__abc_44228_n7154), .Y(u2__abc_44228_n14544) );
  INVX1 INVX1_306 ( .A(sqrto_56_), .Y(u2__abc_44228_n3385) );
  INVX1 INVX1_3060 ( .A(u2__abc_44228_n14545), .Y(u2__abc_44228_n14547) );
  INVX1 INVX1_3061 ( .A(u2__abc_44228_n14554), .Y(u2__abc_44228_n14555) );
  INVX1 INVX1_3062 ( .A(u2__abc_44228_n14562), .Y(u2__abc_44228_n14563) );
  INVX1 INVX1_3063 ( .A(u2__abc_44228_n14564_1), .Y(u2__abc_44228_n14565) );
  INVX1 INVX1_3064 ( .A(u2__abc_44228_n14572), .Y(u2__abc_44228_n14573_1) );
  INVX1 INVX1_3065 ( .A(u2__abc_44228_n7140), .Y(u2__abc_44228_n14579) );
  INVX1 INVX1_3066 ( .A(u2__abc_44228_n14580), .Y(u2__abc_44228_n14581_1) );
  INVX1 INVX1_3067 ( .A(u2__abc_44228_n14589), .Y(u2__abc_44228_n14590) );
  INVX1 INVX1_3068 ( .A(u2__abc_44228_n14599), .Y(u2__abc_44228_n14600) );
  INVX1 INVX1_3069 ( .A(u2__abc_44228_n14606), .Y(u2__abc_44228_n14607) );
  INVX1 INVX1_307 ( .A(u2_remHi_56_), .Y(u2__abc_44228_n3387) );
  INVX1 INVX1_3070 ( .A(u2__abc_44228_n14613), .Y(u2__abc_44228_n14614) );
  INVX1 INVX1_3071 ( .A(u2__abc_44228_n7125_1), .Y(u2__abc_44228_n14616) );
  INVX1 INVX1_3072 ( .A(u2__abc_44228_n14623), .Y(u2__abc_44228_n14624) );
  INVX1 INVX1_3073 ( .A(u2__abc_44228_n14631), .Y(u2__abc_44228_n14632) );
  INVX1 INVX1_3074 ( .A(u2__abc_44228_n14633), .Y(u2__abc_44228_n14634) );
  INVX1 INVX1_3075 ( .A(u2__abc_44228_n14641), .Y(u2__abc_44228_n14642) );
  INVX1 INVX1_3076 ( .A(u2__abc_44228_n7111), .Y(u2__abc_44228_n14648) );
  INVX1 INVX1_3077 ( .A(u2__abc_44228_n14649), .Y(u2__abc_44228_n14650) );
  INVX1 INVX1_3078 ( .A(u2__abc_44228_n14658), .Y(u2__abc_44228_n14659) );
  INVX1 INVX1_3079 ( .A(u2__abc_44228_n14667), .Y(u2__abc_44228_n14668) );
  INVX1 INVX1_308 ( .A(u2__abc_44228_n3389), .Y(u2__abc_44228_n3390) );
  INVX1 INVX1_3080 ( .A(u2__abc_44228_n14675), .Y(u2__abc_44228_n14676) );
  INVX1 INVX1_3081 ( .A(u2__abc_44228_n7099), .Y(u2__abc_44228_n14684) );
  INVX1 INVX1_3082 ( .A(u2__abc_44228_n14682_1), .Y(u2__abc_44228_n14685) );
  INVX1 INVX1_3083 ( .A(u2__abc_44228_n14692), .Y(u2__abc_44228_n14693) );
  INVX1 INVX1_3084 ( .A(u2__abc_44228_n14700_1), .Y(u2__abc_44228_n14701) );
  INVX1 INVX1_3085 ( .A(u2__abc_44228_n14702), .Y(u2__abc_44228_n14703) );
  INVX1 INVX1_3086 ( .A(u2__abc_44228_n14710), .Y(u2__abc_44228_n14711) );
  INVX1 INVX1_3087 ( .A(u2__abc_44228_n7079), .Y(u2__abc_44228_n14717_1) );
  INVX1 INVX1_3088 ( .A(u2__abc_44228_n14718), .Y(u2__abc_44228_n14719) );
  INVX1 INVX1_3089 ( .A(u2__abc_44228_n14727), .Y(u2__abc_44228_n14728) );
  INVX1 INVX1_309 ( .A(sqrto_55_), .Y(u2__abc_44228_n3392) );
  INVX1 INVX1_3090 ( .A(u2__abc_44228_n14737_1), .Y(u2__abc_44228_n14738) );
  INVX1 INVX1_3091 ( .A(u2__abc_44228_n14744), .Y(u2__abc_44228_n14745_1) );
  INVX1 INVX1_3092 ( .A(u2__abc_44228_n7064), .Y(u2__abc_44228_n14751) );
  INVX1 INVX1_3093 ( .A(u2__abc_44228_n14752), .Y(u2__abc_44228_n14754_1) );
  INVX1 INVX1_3094 ( .A(u2__abc_44228_n14761), .Y(u2__abc_44228_n14762_1) );
  INVX1 INVX1_3095 ( .A(u2__abc_44228_n14770), .Y(u2__abc_44228_n14771) );
  INVX1 INVX1_3096 ( .A(u2__abc_44228_n14778), .Y(u2__abc_44228_n14779) );
  INVX1 INVX1_3097 ( .A(u2__abc_44228_n7050_1), .Y(u2__abc_44228_n14785) );
  INVX1 INVX1_3098 ( .A(u2__abc_44228_n14786), .Y(u2__abc_44228_n14787) );
  INVX1 INVX1_3099 ( .A(u2__abc_44228_n14795), .Y(u2__abc_44228_n14796) );
  INVX1 INVX1_31 ( .A(_abc_64468_n1613), .Y(_abc_64468_n1614) );
  INVX1 INVX1_310 ( .A(u2__abc_44228_n3393), .Y(u2__abc_44228_n3394) );
  INVX1 INVX1_3100 ( .A(u2__abc_44228_n14804), .Y(u2__abc_44228_n14805) );
  INVX1 INVX1_3101 ( .A(u2__abc_44228_n14812), .Y(u2__abc_44228_n14813) );
  INVX1 INVX1_3102 ( .A(u2__abc_44228_n7034), .Y(u2__abc_44228_n14821) );
  INVX1 INVX1_3103 ( .A(u2__abc_44228_n14822), .Y(u2__abc_44228_n14824) );
  INVX1 INVX1_3104 ( .A(u2__abc_44228_n14829), .Y(u2__abc_44228_n14830) );
  INVX1 INVX1_3105 ( .A(u2__abc_44228_n14838), .Y(u2__abc_44228_n14839) );
  INVX1 INVX1_3106 ( .A(u2__abc_44228_n14846), .Y(u2__abc_44228_n14847) );
  INVX1 INVX1_3107 ( .A(u2__abc_44228_n7020), .Y(u2__abc_44228_n14853) );
  INVX1 INVX1_3108 ( .A(u2__abc_44228_n14854), .Y(u2__abc_44228_n14856) );
  INVX1 INVX1_3109 ( .A(u2__abc_44228_n14863), .Y(u2__abc_44228_n14864) );
  INVX1 INVX1_311 ( .A(u2_remHi_55_), .Y(u2__abc_44228_n3395) );
  INVX1 INVX1_3110 ( .A(u2__abc_44228_n14871), .Y(u2__abc_44228_n14872) );
  INVX1 INVX1_3111 ( .A(u2__abc_44228_n14873), .Y(u2__abc_44228_n14874) );
  INVX1 INVX1_3112 ( .A(u2__abc_44228_n14881), .Y(u2__abc_44228_n14882) );
  INVX1 INVX1_3113 ( .A(u2__abc_44228_n7005), .Y(u2__abc_44228_n14890) );
  INVX1 INVX1_3114 ( .A(u2__abc_44228_n14888), .Y(u2__abc_44228_n14891_1) );
  INVX1 INVX1_3115 ( .A(u2__abc_44228_n14898), .Y(u2__abc_44228_n14899) );
  INVX1 INVX1_3116 ( .A(u2__abc_44228_n14906), .Y(u2__abc_44228_n14907) );
  INVX1 INVX1_3117 ( .A(u2__abc_44228_n14908_1), .Y(u2__abc_44228_n14909) );
  INVX1 INVX1_3118 ( .A(u2__abc_44228_n14916), .Y(u2__abc_44228_n14917) );
  INVX1 INVX1_3119 ( .A(u2__abc_44228_n6991), .Y(u2__abc_44228_n14923) );
  INVX1 INVX1_312 ( .A(u2__abc_44228_n3396), .Y(u2__abc_44228_n3397) );
  INVX1 INVX1_3120 ( .A(u2__abc_44228_n14924), .Y(u2__abc_44228_n14925) );
  INVX1 INVX1_3121 ( .A(u2__abc_44228_n14933), .Y(u2__abc_44228_n14934) );
  INVX1 INVX1_3122 ( .A(u2__abc_44228_n14943_1), .Y(u2__abc_44228_n14944) );
  INVX1 INVX1_3123 ( .A(u2__abc_44228_n14950), .Y(u2__abc_44228_n14951) );
  INVX1 INVX1_3124 ( .A(u2__abc_44228_n6960), .Y(u2__abc_44228_n14957) );
  INVX1 INVX1_3125 ( .A(u2__abc_44228_n14958), .Y(u2__abc_44228_n14960) );
  INVX1 INVX1_3126 ( .A(u2__abc_44228_n14967), .Y(u2__abc_44228_n14968) );
  INVX1 INVX1_3127 ( .A(u2__abc_44228_n14976), .Y(u2__abc_44228_n14977) );
  INVX1 INVX1_3128 ( .A(u2__abc_44228_n14984), .Y(u2__abc_44228_n14985) );
  INVX1 INVX1_3129 ( .A(u2__abc_44228_n6974), .Y(u2__abc_44228_n14991) );
  INVX1 INVX1_313 ( .A(sqrto_54_), .Y(u2__abc_44228_n3399) );
  INVX1 INVX1_3130 ( .A(u2__abc_44228_n14992), .Y(u2__abc_44228_n14994) );
  INVX1 INVX1_3131 ( .A(u2__abc_44228_n15001), .Y(u2__abc_44228_n15002) );
  INVX1 INVX1_3132 ( .A(u2__abc_44228_n15009), .Y(u2__abc_44228_n15010) );
  INVX1 INVX1_3133 ( .A(u2__abc_44228_n15012), .Y(u2__abc_44228_n15013) );
  INVX1 INVX1_3134 ( .A(u2__abc_44228_n15019), .Y(u2__abc_44228_n15020) );
  INVX1 INVX1_3135 ( .A(u2__abc_44228_n15026_1), .Y(u2__abc_44228_n15027) );
  INVX1 INVX1_3136 ( .A(u2__abc_44228_n6951), .Y(u2__abc_44228_n15029) );
  INVX1 INVX1_3137 ( .A(u2__abc_44228_n15036), .Y(u2__abc_44228_n15037) );
  INVX1 INVX1_3138 ( .A(u2__abc_44228_n15044), .Y(u2__abc_44228_n15045) );
  INVX1 INVX1_3139 ( .A(u2__abc_44228_n15046), .Y(u2__abc_44228_n15047) );
  INVX1 INVX1_314 ( .A(u2_remHi_54_), .Y(u2__abc_44228_n3401) );
  INVX1 INVX1_3140 ( .A(u2__abc_44228_n15054), .Y(u2__abc_44228_n15055) );
  INVX1 INVX1_3141 ( .A(u2__abc_44228_n6931), .Y(u2__abc_44228_n15061_1) );
  INVX1 INVX1_3142 ( .A(u2__abc_44228_n15062), .Y(u2__abc_44228_n15063) );
  INVX1 INVX1_3143 ( .A(u2__abc_44228_n15071), .Y(u2__abc_44228_n15072) );
  INVX1 INVX1_3144 ( .A(u2__abc_44228_n15080), .Y(u2__abc_44228_n15081) );
  INVX1 INVX1_3145 ( .A(u2__abc_44228_n15088), .Y(u2__abc_44228_n15089) );
  INVX1 INVX1_3146 ( .A(u2__abc_44228_n6915_1), .Y(u2__abc_44228_n15097_1) );
  INVX1 INVX1_3147 ( .A(u2__abc_44228_n15095), .Y(u2__abc_44228_n15098) );
  INVX1 INVX1_3148 ( .A(u2__abc_44228_n15105_1), .Y(u2__abc_44228_n15106) );
  INVX1 INVX1_3149 ( .A(u2__abc_44228_n15113), .Y(u2__abc_44228_n15114_1) );
  INVX1 INVX1_315 ( .A(u2__abc_44228_n3403), .Y(u2__abc_44228_n3404) );
  INVX1 INVX1_3150 ( .A(u2__abc_44228_n15115), .Y(u2__abc_44228_n15116) );
  INVX1 INVX1_3151 ( .A(u2__abc_44228_n15123), .Y(u2__abc_44228_n15124) );
  INVX1 INVX1_3152 ( .A(u2__abc_44228_n6901), .Y(u2__abc_44228_n15130) );
  INVX1 INVX1_3153 ( .A(u2__abc_44228_n15131), .Y(u2__abc_44228_n15132_1) );
  INVX1 INVX1_3154 ( .A(u2__abc_44228_n15140_1), .Y(u2__abc_44228_n15141) );
  INVX1 INVX1_3155 ( .A(u2__abc_44228_n15150), .Y(u2__abc_44228_n15151) );
  INVX1 INVX1_3156 ( .A(u2__abc_44228_n15157_1), .Y(u2__abc_44228_n15158) );
  INVX1 INVX1_3157 ( .A(u2__abc_44228_n6886), .Y(u2__abc_44228_n15164) );
  INVX1 INVX1_3158 ( .A(u2__abc_44228_n15165), .Y(u2__abc_44228_n15167) );
  INVX1 INVX1_3159 ( .A(u2__abc_44228_n15174), .Y(u2__abc_44228_n15175) );
  INVX1 INVX1_316 ( .A(sqrto_53_), .Y(u2__abc_44228_n3408) );
  INVX1 INVX1_3160 ( .A(u2__abc_44228_n15183), .Y(u2__abc_44228_n15184) );
  INVX1 INVX1_3161 ( .A(u2__abc_44228_n15191), .Y(u2__abc_44228_n15192) );
  INVX1 INVX1_3162 ( .A(u2__abc_44228_n6872), .Y(u2__abc_44228_n15198) );
  INVX1 INVX1_3163 ( .A(u2__abc_44228_n15199), .Y(u2__abc_44228_n15200) );
  INVX1 INVX1_3164 ( .A(u2__abc_44228_n15208), .Y(u2__abc_44228_n15209) );
  INVX1 INVX1_3165 ( .A(u2__abc_44228_n15216), .Y(u2__abc_44228_n15217) );
  INVX1 INVX1_3166 ( .A(u2__abc_44228_n15223), .Y(u2__abc_44228_n15224) );
  INVX1 INVX1_3167 ( .A(u2__abc_44228_n7535), .Y(u2__abc_44228_n15230_1) );
  INVX1 INVX1_3168 ( .A(u2__abc_44228_n15231), .Y(u2__abc_44228_n15233) );
  INVX1 INVX1_3169 ( .A(u2__abc_44228_n15240), .Y(u2__abc_44228_n15241_1) );
  INVX1 INVX1_317 ( .A(u2__abc_44228_n3409), .Y(u2__abc_44228_n3410) );
  INVX1 INVX1_3170 ( .A(u2__abc_44228_n17776), .Y(u2__abc_44228_n17777) );
  INVX1 INVX1_3171 ( .A(u2__abc_44228_n17781), .Y(u2__abc_44228_n17782) );
  INVX1 INVX1_3172 ( .A(u2__abc_44228_n17789), .Y(u2__abc_44228_n17790) );
  INVX1 INVX1_3173 ( .A(u2__abc_44228_n17793), .Y(u2__abc_44228_n17794) );
  INVX1 INVX1_3174 ( .A(u2__abc_44228_n17801), .Y(u2__abc_44228_n17802) );
  INVX1 INVX1_3175 ( .A(u2__abc_44228_n17805), .Y(u2__abc_44228_n17806) );
  INVX1 INVX1_3176 ( .A(u2__abc_44228_n17813), .Y(u2__abc_44228_n17814) );
  INVX1 INVX1_3177 ( .A(u2__abc_44228_n17817), .Y(u2__abc_44228_n17818) );
  INVX1 INVX1_3178 ( .A(u2__abc_44228_n17825), .Y(u2__abc_44228_n17826) );
  INVX1 INVX1_3179 ( .A(u2__abc_44228_n17829), .Y(u2__abc_44228_n17830) );
  INVX1 INVX1_318 ( .A(u2_remHi_53_), .Y(u2__abc_44228_n3411) );
  INVX1 INVX1_3180 ( .A(u2__abc_44228_n17837), .Y(u2__abc_44228_n17838) );
  INVX1 INVX1_3181 ( .A(u2__abc_44228_n17841), .Y(u2__abc_44228_n17842) );
  INVX1 INVX1_3182 ( .A(u2__abc_44228_n17849), .Y(u2__abc_44228_n17850) );
  INVX1 INVX1_3183 ( .A(u2__abc_44228_n17853), .Y(u2__abc_44228_n17854) );
  INVX1 INVX1_3184 ( .A(u2__abc_44228_n17861), .Y(u2__abc_44228_n17862) );
  INVX1 INVX1_3185 ( .A(u2__abc_44228_n17865), .Y(u2__abc_44228_n17866) );
  INVX1 INVX1_3186 ( .A(u2__abc_44228_n17873), .Y(u2__abc_44228_n17874) );
  INVX1 INVX1_3187 ( .A(u2__abc_44228_n17877), .Y(u2__abc_44228_n17878) );
  INVX1 INVX1_3188 ( .A(u2__abc_44228_n17885), .Y(u2__abc_44228_n17886) );
  INVX1 INVX1_3189 ( .A(u2__abc_44228_n17889), .Y(u2__abc_44228_n17890) );
  INVX1 INVX1_319 ( .A(u2__abc_44228_n3412), .Y(u2__abc_44228_n3413) );
  INVX1 INVX1_3190 ( .A(u2__abc_44228_n17897), .Y(u2__abc_44228_n17898) );
  INVX1 INVX1_3191 ( .A(u2__abc_44228_n17901), .Y(u2__abc_44228_n17902) );
  INVX1 INVX1_3192 ( .A(u2__abc_44228_n17909), .Y(u2__abc_44228_n17910) );
  INVX1 INVX1_3193 ( .A(u2__abc_44228_n17913), .Y(u2__abc_44228_n17914) );
  INVX1 INVX1_3194 ( .A(u2__abc_44228_n17921), .Y(u2__abc_44228_n17922) );
  INVX1 INVX1_3195 ( .A(u2__abc_44228_n17925), .Y(u2__abc_44228_n17926) );
  INVX1 INVX1_3196 ( .A(u2__abc_44228_n17933), .Y(u2__abc_44228_n17934) );
  INVX1 INVX1_3197 ( .A(u2__abc_44228_n17937), .Y(u2__abc_44228_n17938) );
  INVX1 INVX1_3198 ( .A(u2__abc_44228_n17945), .Y(u2__abc_44228_n17946) );
  INVX1 INVX1_3199 ( .A(u2__abc_44228_n17949), .Y(u2__abc_44228_n17950) );
  INVX1 INVX1_32 ( .A(_abc_64468_n1616), .Y(_abc_64468_n1622) );
  INVX1 INVX1_320 ( .A(sqrto_52_), .Y(u2__abc_44228_n3415) );
  INVX1 INVX1_3200 ( .A(u2__abc_44228_n17957), .Y(u2__abc_44228_n17958) );
  INVX1 INVX1_3201 ( .A(u2__abc_44228_n17961), .Y(u2__abc_44228_n17962) );
  INVX1 INVX1_3202 ( .A(u2__abc_44228_n17969), .Y(u2__abc_44228_n17970) );
  INVX1 INVX1_3203 ( .A(u2__abc_44228_n17973), .Y(u2__abc_44228_n17974) );
  INVX1 INVX1_3204 ( .A(u2__abc_44228_n17981), .Y(u2__abc_44228_n17982) );
  INVX1 INVX1_3205 ( .A(u2__abc_44228_n17985), .Y(u2__abc_44228_n17986) );
  INVX1 INVX1_3206 ( .A(u2__abc_44228_n17993), .Y(u2__abc_44228_n17994) );
  INVX1 INVX1_3207 ( .A(u2__abc_44228_n17997), .Y(u2__abc_44228_n17998) );
  INVX1 INVX1_3208 ( .A(u2__abc_44228_n18005), .Y(u2__abc_44228_n18006) );
  INVX1 INVX1_3209 ( .A(u2__abc_44228_n18009), .Y(u2__abc_44228_n18010) );
  INVX1 INVX1_321 ( .A(u2_remHi_52_), .Y(u2__abc_44228_n3417) );
  INVX1 INVX1_3210 ( .A(u2__abc_44228_n18017), .Y(u2__abc_44228_n18018) );
  INVX1 INVX1_3211 ( .A(u2__abc_44228_n18021), .Y(u2__abc_44228_n18022) );
  INVX1 INVX1_3212 ( .A(u2__abc_44228_n18029), .Y(u2__abc_44228_n18030) );
  INVX1 INVX1_3213 ( .A(u2__abc_44228_n18033), .Y(u2__abc_44228_n18034) );
  INVX1 INVX1_3214 ( .A(u2__abc_44228_n18041), .Y(u2__abc_44228_n18042) );
  INVX1 INVX1_3215 ( .A(u2__abc_44228_n18045), .Y(u2__abc_44228_n18046) );
  INVX1 INVX1_3216 ( .A(u2__abc_44228_n18053), .Y(u2__abc_44228_n18054) );
  INVX1 INVX1_3217 ( .A(u2__abc_44228_n18057), .Y(u2__abc_44228_n18058) );
  INVX1 INVX1_3218 ( .A(u2__abc_44228_n18065), .Y(u2__abc_44228_n18066) );
  INVX1 INVX1_3219 ( .A(u2__abc_44228_n18069), .Y(u2__abc_44228_n18070) );
  INVX1 INVX1_322 ( .A(u2__abc_44228_n3419), .Y(u2__abc_44228_n3420) );
  INVX1 INVX1_3220 ( .A(u2__abc_44228_n18077), .Y(u2__abc_44228_n18078) );
  INVX1 INVX1_3221 ( .A(u2__abc_44228_n18081), .Y(u2__abc_44228_n18082) );
  INVX1 INVX1_3222 ( .A(u2__abc_44228_n18089), .Y(u2__abc_44228_n18090) );
  INVX1 INVX1_3223 ( .A(u2__abc_44228_n18093), .Y(u2__abc_44228_n18094) );
  INVX1 INVX1_3224 ( .A(u2__abc_44228_n18101), .Y(u2__abc_44228_n18102) );
  INVX1 INVX1_3225 ( .A(u2__abc_44228_n18105), .Y(u2__abc_44228_n18106) );
  INVX1 INVX1_3226 ( .A(u2__abc_44228_n18113), .Y(u2__abc_44228_n18114) );
  INVX1 INVX1_3227 ( .A(u2__abc_44228_n18117), .Y(u2__abc_44228_n18118) );
  INVX1 INVX1_3228 ( .A(u2__abc_44228_n18125), .Y(u2__abc_44228_n18126) );
  INVX1 INVX1_3229 ( .A(u2__abc_44228_n18129), .Y(u2__abc_44228_n18130) );
  INVX1 INVX1_323 ( .A(sqrto_50_), .Y(u2__abc_44228_n3422) );
  INVX1 INVX1_3230 ( .A(u2__abc_44228_n18137), .Y(u2__abc_44228_n18138) );
  INVX1 INVX1_3231 ( .A(u2__abc_44228_n18141), .Y(u2__abc_44228_n18142) );
  INVX1 INVX1_3232 ( .A(u2__abc_44228_n18149), .Y(u2__abc_44228_n18150) );
  INVX1 INVX1_3233 ( .A(u2__abc_44228_n18153), .Y(u2__abc_44228_n18154) );
  INVX1 INVX1_3234 ( .A(u2__abc_44228_n18161), .Y(u2__abc_44228_n18162) );
  INVX1 INVX1_3235 ( .A(u2__abc_44228_n18165), .Y(u2__abc_44228_n18166) );
  INVX1 INVX1_3236 ( .A(u2__abc_44228_n18173), .Y(u2__abc_44228_n18174) );
  INVX1 INVX1_3237 ( .A(u2__abc_44228_n18177), .Y(u2__abc_44228_n18178) );
  INVX1 INVX1_3238 ( .A(u2__abc_44228_n18185), .Y(u2__abc_44228_n18186) );
  INVX1 INVX1_3239 ( .A(u2__abc_44228_n18189), .Y(u2__abc_44228_n18190) );
  INVX1 INVX1_324 ( .A(u2_remHi_50_), .Y(u2__abc_44228_n3424) );
  INVX1 INVX1_3240 ( .A(u2__abc_44228_n18197), .Y(u2__abc_44228_n18198) );
  INVX1 INVX1_3241 ( .A(u2__abc_44228_n18201), .Y(u2__abc_44228_n18202) );
  INVX1 INVX1_3242 ( .A(u2__abc_44228_n18209), .Y(u2__abc_44228_n18210) );
  INVX1 INVX1_3243 ( .A(u2__abc_44228_n18213), .Y(u2__abc_44228_n18214) );
  INVX1 INVX1_3244 ( .A(u2__abc_44228_n18221), .Y(u2__abc_44228_n18222) );
  INVX1 INVX1_3245 ( .A(u2__abc_44228_n18225), .Y(u2__abc_44228_n18226) );
  INVX1 INVX1_3246 ( .A(u2__abc_44228_n18233), .Y(u2__abc_44228_n18234) );
  INVX1 INVX1_3247 ( .A(u2__abc_44228_n18237), .Y(u2__abc_44228_n18238) );
  INVX1 INVX1_3248 ( .A(u2__abc_44228_n18245), .Y(u2__abc_44228_n18246) );
  INVX1 INVX1_3249 ( .A(u2__abc_44228_n18249), .Y(u2__abc_44228_n18250) );
  INVX1 INVX1_325 ( .A(u2__abc_44228_n3426), .Y(u2__abc_44228_n3427) );
  INVX1 INVX1_3250 ( .A(u2__abc_44228_n18257), .Y(u2__abc_44228_n18258) );
  INVX1 INVX1_3251 ( .A(u2__abc_44228_n18261), .Y(u2__abc_44228_n18262) );
  INVX1 INVX1_3252 ( .A(u2__abc_44228_n18269), .Y(u2__abc_44228_n18270) );
  INVX1 INVX1_3253 ( .A(u2__abc_44228_n18273), .Y(u2__abc_44228_n18274) );
  INVX1 INVX1_3254 ( .A(u2__abc_44228_n18281), .Y(u2__abc_44228_n18282) );
  INVX1 INVX1_3255 ( .A(u2__abc_44228_n18285), .Y(u2__abc_44228_n18286) );
  INVX1 INVX1_3256 ( .A(u2__abc_44228_n18293), .Y(u2__abc_44228_n18294) );
  INVX1 INVX1_3257 ( .A(u2__abc_44228_n18297), .Y(u2__abc_44228_n18298) );
  INVX1 INVX1_3258 ( .A(u2__abc_44228_n18305), .Y(u2__abc_44228_n18306) );
  INVX1 INVX1_3259 ( .A(u2__abc_44228_n18309), .Y(u2__abc_44228_n18310) );
  INVX1 INVX1_326 ( .A(sqrto_51_), .Y(u2__abc_44228_n3428) );
  INVX1 INVX1_3260 ( .A(u2__abc_44228_n18317), .Y(u2__abc_44228_n18318) );
  INVX1 INVX1_3261 ( .A(u2__abc_44228_n18321), .Y(u2__abc_44228_n18322) );
  INVX1 INVX1_3262 ( .A(u2__abc_44228_n18329), .Y(u2__abc_44228_n18330) );
  INVX1 INVX1_3263 ( .A(u2__abc_44228_n18333), .Y(u2__abc_44228_n18334) );
  INVX1 INVX1_3264 ( .A(u2__abc_44228_n18341), .Y(u2__abc_44228_n18342) );
  INVX1 INVX1_3265 ( .A(u2__abc_44228_n18345), .Y(u2__abc_44228_n18346) );
  INVX1 INVX1_3266 ( .A(u2__abc_44228_n18353), .Y(u2__abc_44228_n18354) );
  INVX1 INVX1_3267 ( .A(u2__abc_44228_n18357), .Y(u2__abc_44228_n18358) );
  INVX1 INVX1_3268 ( .A(u2__abc_44228_n18365), .Y(u2__abc_44228_n18366) );
  INVX1 INVX1_3269 ( .A(u2__abc_44228_n18369), .Y(u2__abc_44228_n18370) );
  INVX1 INVX1_327 ( .A(u2__abc_44228_n3429), .Y(u2__abc_44228_n3430) );
  INVX1 INVX1_3270 ( .A(u2__abc_44228_n18377), .Y(u2__abc_44228_n18378) );
  INVX1 INVX1_3271 ( .A(u2__abc_44228_n18381), .Y(u2__abc_44228_n18382) );
  INVX1 INVX1_3272 ( .A(u2__abc_44228_n18389), .Y(u2__abc_44228_n18390) );
  INVX1 INVX1_3273 ( .A(u2__abc_44228_n18393), .Y(u2__abc_44228_n18394) );
  INVX1 INVX1_3274 ( .A(u2__abc_44228_n18401), .Y(u2__abc_44228_n18402) );
  INVX1 INVX1_3275 ( .A(u2__abc_44228_n18405), .Y(u2__abc_44228_n18406) );
  INVX1 INVX1_3276 ( .A(u2__abc_44228_n18413), .Y(u2__abc_44228_n18414) );
  INVX1 INVX1_3277 ( .A(u2__abc_44228_n18417), .Y(u2__abc_44228_n18418) );
  INVX1 INVX1_3278 ( .A(u2__abc_44228_n18425), .Y(u2__abc_44228_n18426) );
  INVX1 INVX1_3279 ( .A(u2__abc_44228_n18429), .Y(u2__abc_44228_n18430) );
  INVX1 INVX1_328 ( .A(u2_remHi_51_), .Y(u2__abc_44228_n3431) );
  INVX1 INVX1_3280 ( .A(u2__abc_44228_n18437), .Y(u2__abc_44228_n18438) );
  INVX1 INVX1_3281 ( .A(u2__abc_44228_n18441), .Y(u2__abc_44228_n18442) );
  INVX1 INVX1_3282 ( .A(u2__abc_44228_n18449), .Y(u2__abc_44228_n18450) );
  INVX1 INVX1_3283 ( .A(u2__abc_44228_n18453), .Y(u2__abc_44228_n18454) );
  INVX1 INVX1_3284 ( .A(u2__abc_44228_n18461), .Y(u2__abc_44228_n18462) );
  INVX1 INVX1_3285 ( .A(u2__abc_44228_n18465), .Y(u2__abc_44228_n18466) );
  INVX1 INVX1_3286 ( .A(u2__abc_44228_n18473), .Y(u2__abc_44228_n18474) );
  INVX1 INVX1_3287 ( .A(u2__abc_44228_n18477), .Y(u2__abc_44228_n18478) );
  INVX1 INVX1_3288 ( .A(u2__abc_44228_n18485), .Y(u2__abc_44228_n18486) );
  INVX1 INVX1_3289 ( .A(u2__abc_44228_n18489), .Y(u2__abc_44228_n18490) );
  INVX1 INVX1_329 ( .A(u2__abc_44228_n3432), .Y(u2__abc_44228_n3433) );
  INVX1 INVX1_3290 ( .A(u2__abc_44228_n18497), .Y(u2__abc_44228_n18498) );
  INVX1 INVX1_3291 ( .A(u2__abc_44228_n18501), .Y(u2__abc_44228_n18502) );
  INVX1 INVX1_3292 ( .A(u2__abc_44228_n18509), .Y(u2__abc_44228_n18510) );
  INVX1 INVX1_3293 ( .A(u2__abc_44228_n18513), .Y(u2__abc_44228_n18514) );
  INVX1 INVX1_3294 ( .A(u2__abc_44228_n18521), .Y(u2__abc_44228_n18522) );
  INVX1 INVX1_3295 ( .A(u2__abc_44228_n18525), .Y(u2__abc_44228_n18526) );
  INVX1 INVX1_3296 ( .A(u2__abc_44228_n18533), .Y(u2__abc_44228_n18534) );
  INVX1 INVX1_3297 ( .A(u2__abc_44228_n18537), .Y(u2__abc_44228_n18538) );
  INVX1 INVX1_3298 ( .A(u2__abc_44228_n18545), .Y(u2__abc_44228_n18546) );
  INVX1 INVX1_3299 ( .A(u2__abc_44228_n18549), .Y(u2__abc_44228_n18550) );
  INVX1 INVX1_33 ( .A(\a[122] ), .Y(_abc_64468_n1623) );
  INVX1 INVX1_330 ( .A(sqrto_49_), .Y(u2__abc_44228_n3437) );
  INVX1 INVX1_3300 ( .A(u2__abc_44228_n18557), .Y(u2__abc_44228_n18558) );
  INVX1 INVX1_3301 ( .A(u2__abc_44228_n18561), .Y(u2__abc_44228_n18562) );
  INVX1 INVX1_3302 ( .A(u2__abc_44228_n18569), .Y(u2__abc_44228_n18570) );
  INVX1 INVX1_3303 ( .A(u2__abc_44228_n18573), .Y(u2__abc_44228_n18574) );
  INVX1 INVX1_3304 ( .A(u2__abc_44228_n18581), .Y(u2__abc_44228_n18582) );
  INVX1 INVX1_3305 ( .A(u2__abc_44228_n18585), .Y(u2__abc_44228_n18586) );
  INVX1 INVX1_3306 ( .A(u2__abc_44228_n18593), .Y(u2__abc_44228_n18594) );
  INVX1 INVX1_3307 ( .A(u2__abc_44228_n18597), .Y(u2__abc_44228_n18598) );
  INVX1 INVX1_3308 ( .A(u2__abc_44228_n18605), .Y(u2__abc_44228_n18606) );
  INVX1 INVX1_3309 ( .A(u2__abc_44228_n18609), .Y(u2__abc_44228_n18610) );
  INVX1 INVX1_331 ( .A(u2__abc_44228_n3438), .Y(u2__abc_44228_n3439_1) );
  INVX1 INVX1_3310 ( .A(u2__abc_44228_n18617), .Y(u2__abc_44228_n18618) );
  INVX1 INVX1_3311 ( .A(u2__abc_44228_n18621), .Y(u2__abc_44228_n18622) );
  INVX1 INVX1_3312 ( .A(u2__abc_44228_n18629), .Y(u2__abc_44228_n18630) );
  INVX1 INVX1_3313 ( .A(u2__abc_44228_n18633), .Y(u2__abc_44228_n18634) );
  INVX1 INVX1_3314 ( .A(u2__abc_44228_n18641), .Y(u2__abc_44228_n18642) );
  INVX1 INVX1_3315 ( .A(u2__abc_44228_n18645), .Y(u2__abc_44228_n18646) );
  INVX1 INVX1_3316 ( .A(u2__abc_44228_n18653), .Y(u2__abc_44228_n18654) );
  INVX1 INVX1_3317 ( .A(u2__abc_44228_n18657), .Y(u2__abc_44228_n18658) );
  INVX1 INVX1_3318 ( .A(u2__abc_44228_n18665), .Y(u2__abc_44228_n18666) );
  INVX1 INVX1_3319 ( .A(u2__abc_44228_n18669), .Y(u2__abc_44228_n18670) );
  INVX1 INVX1_332 ( .A(u2_remHi_49_), .Y(u2__abc_44228_n3440) );
  INVX1 INVX1_3320 ( .A(u2__abc_44228_n18677), .Y(u2__abc_44228_n18678) );
  INVX1 INVX1_3321 ( .A(u2__abc_44228_n18681), .Y(u2__abc_44228_n18682) );
  INVX1 INVX1_3322 ( .A(u2__abc_44228_n18689), .Y(u2__abc_44228_n18690) );
  INVX1 INVX1_3323 ( .A(u2__abc_44228_n18693), .Y(u2__abc_44228_n18694) );
  INVX1 INVX1_3324 ( .A(u2__abc_44228_n18701), .Y(u2__abc_44228_n18702) );
  INVX1 INVX1_3325 ( .A(u2__abc_44228_n18705), .Y(u2__abc_44228_n18706) );
  INVX1 INVX1_3326 ( .A(u2__abc_44228_n18713), .Y(u2__abc_44228_n18714) );
  INVX1 INVX1_3327 ( .A(u2__abc_44228_n18717), .Y(u2__abc_44228_n18718) );
  INVX1 INVX1_3328 ( .A(u2__abc_44228_n18725), .Y(u2__abc_44228_n18726) );
  INVX1 INVX1_3329 ( .A(u2__abc_44228_n18729), .Y(u2__abc_44228_n18730) );
  INVX1 INVX1_333 ( .A(u2__abc_44228_n3441), .Y(u2__abc_44228_n3442) );
  INVX1 INVX1_3330 ( .A(u2__abc_44228_n18737), .Y(u2__abc_44228_n18738) );
  INVX1 INVX1_3331 ( .A(u2__abc_44228_n18741), .Y(u2__abc_44228_n18742) );
  INVX1 INVX1_3332 ( .A(u2__abc_44228_n18749), .Y(u2__abc_44228_n18750) );
  INVX1 INVX1_3333 ( .A(u2__abc_44228_n18753), .Y(u2__abc_44228_n18754) );
  INVX1 INVX1_3334 ( .A(u2__abc_44228_n18761), .Y(u2__abc_44228_n18762) );
  INVX1 INVX1_3335 ( .A(u2__abc_44228_n18765), .Y(u2__abc_44228_n18766) );
  INVX1 INVX1_3336 ( .A(u2__abc_44228_n18773), .Y(u2__abc_44228_n18774) );
  INVX1 INVX1_3337 ( .A(u2__abc_44228_n18777), .Y(u2__abc_44228_n18778) );
  INVX1 INVX1_3338 ( .A(u2__abc_44228_n18785), .Y(u2__abc_44228_n18786) );
  INVX1 INVX1_3339 ( .A(u2__abc_44228_n18789), .Y(u2__abc_44228_n18790) );
  INVX1 INVX1_334 ( .A(sqrto_48_), .Y(u2__abc_44228_n3444) );
  INVX1 INVX1_3340 ( .A(u2__abc_44228_n18797), .Y(u2__abc_44228_n18798) );
  INVX1 INVX1_3341 ( .A(u2__abc_44228_n18801), .Y(u2__abc_44228_n18802) );
  INVX1 INVX1_3342 ( .A(u2__abc_44228_n18809), .Y(u2__abc_44228_n18810) );
  INVX1 INVX1_3343 ( .A(u2__abc_44228_n18813), .Y(u2__abc_44228_n18814) );
  INVX1 INVX1_3344 ( .A(u2__abc_44228_n18821), .Y(u2__abc_44228_n18822) );
  INVX1 INVX1_3345 ( .A(u2__abc_44228_n18825), .Y(u2__abc_44228_n18826) );
  INVX1 INVX1_3346 ( .A(u2__abc_44228_n18833), .Y(u2__abc_44228_n18834) );
  INVX1 INVX1_3347 ( .A(u2__abc_44228_n18837), .Y(u2__abc_44228_n18838) );
  INVX1 INVX1_3348 ( .A(u2__abc_44228_n18845), .Y(u2__abc_44228_n18846) );
  INVX1 INVX1_3349 ( .A(u2__abc_44228_n18849), .Y(u2__abc_44228_n18850) );
  INVX1 INVX1_335 ( .A(u2_remHi_48_), .Y(u2__abc_44228_n3446) );
  INVX1 INVX1_3350 ( .A(u2__abc_44228_n18857), .Y(u2__abc_44228_n18858) );
  INVX1 INVX1_3351 ( .A(u2__abc_44228_n18861), .Y(u2__abc_44228_n18862) );
  INVX1 INVX1_3352 ( .A(u2__abc_44228_n18869), .Y(u2__abc_44228_n18870) );
  INVX1 INVX1_3353 ( .A(u2__abc_44228_n18873), .Y(u2__abc_44228_n18874) );
  INVX1 INVX1_3354 ( .A(u2__abc_44228_n18881), .Y(u2__abc_44228_n18882) );
  INVX1 INVX1_3355 ( .A(u2__abc_44228_n18885), .Y(u2__abc_44228_n18886) );
  INVX1 INVX1_3356 ( .A(u2__abc_44228_n18893), .Y(u2__abc_44228_n18894) );
  INVX1 INVX1_3357 ( .A(u2__abc_44228_n18897), .Y(u2__abc_44228_n18898) );
  INVX1 INVX1_3358 ( .A(u2__abc_44228_n18905), .Y(u2__abc_44228_n18906) );
  INVX1 INVX1_3359 ( .A(u2__abc_44228_n18909), .Y(u2__abc_44228_n18910) );
  INVX1 INVX1_336 ( .A(u2__abc_44228_n3448), .Y(u2__abc_44228_n3449_1) );
  INVX1 INVX1_3360 ( .A(u2__abc_44228_n18917), .Y(u2__abc_44228_n18918) );
  INVX1 INVX1_3361 ( .A(u2__abc_44228_n18921), .Y(u2__abc_44228_n18922) );
  INVX1 INVX1_3362 ( .A(u2__abc_44228_n18929), .Y(u2__abc_44228_n18930) );
  INVX1 INVX1_3363 ( .A(u2__abc_44228_n18933), .Y(u2__abc_44228_n18934) );
  INVX1 INVX1_3364 ( .A(u2__abc_44228_n18941), .Y(u2__abc_44228_n18942) );
  INVX1 INVX1_3365 ( .A(u2__abc_44228_n18945), .Y(u2__abc_44228_n18946) );
  INVX1 INVX1_3366 ( .A(u2__abc_44228_n18953), .Y(u2__abc_44228_n18954) );
  INVX1 INVX1_3367 ( .A(u2__abc_44228_n18957), .Y(u2__abc_44228_n18958) );
  INVX1 INVX1_3368 ( .A(u2__abc_44228_n18965), .Y(u2__abc_44228_n18966) );
  INVX1 INVX1_3369 ( .A(u2__abc_44228_n18969), .Y(u2__abc_44228_n18970) );
  INVX1 INVX1_337 ( .A(sqrto_47_), .Y(u2__abc_44228_n3451) );
  INVX1 INVX1_3370 ( .A(u2__abc_44228_n18977), .Y(u2__abc_44228_n18978) );
  INVX1 INVX1_3371 ( .A(u2__abc_44228_n18981), .Y(u2__abc_44228_n18982) );
  INVX1 INVX1_3372 ( .A(u2__abc_44228_n18989), .Y(u2__abc_44228_n18990) );
  INVX1 INVX1_3373 ( .A(u2__abc_44228_n18993), .Y(u2__abc_44228_n18994) );
  INVX1 INVX1_3374 ( .A(u2__abc_44228_n19001), .Y(u2__abc_44228_n19002) );
  INVX1 INVX1_3375 ( .A(u2__abc_44228_n19005), .Y(u2__abc_44228_n19006) );
  INVX1 INVX1_3376 ( .A(u2__abc_44228_n19013), .Y(u2__abc_44228_n19014) );
  INVX1 INVX1_3377 ( .A(u2__abc_44228_n19017), .Y(u2__abc_44228_n19018) );
  INVX1 INVX1_3378 ( .A(u2__abc_44228_n19025), .Y(u2__abc_44228_n19026) );
  INVX1 INVX1_3379 ( .A(u2__abc_44228_n19029), .Y(u2__abc_44228_n19030) );
  INVX1 INVX1_338 ( .A(u2__abc_44228_n3452), .Y(u2__abc_44228_n3453) );
  INVX1 INVX1_3380 ( .A(u2__abc_44228_n19037), .Y(u2__abc_44228_n19038) );
  INVX1 INVX1_3381 ( .A(u2__abc_44228_n19041), .Y(u2__abc_44228_n19042) );
  INVX1 INVX1_3382 ( .A(u2__abc_44228_n19049), .Y(u2__abc_44228_n19050) );
  INVX1 INVX1_3383 ( .A(u2__abc_44228_n19053), .Y(u2__abc_44228_n19054) );
  INVX1 INVX1_3384 ( .A(u2__abc_44228_n19061), .Y(u2__abc_44228_n19062) );
  INVX1 INVX1_3385 ( .A(u2__abc_44228_n19065), .Y(u2__abc_44228_n19066) );
  INVX1 INVX1_3386 ( .A(u2__abc_44228_n19073), .Y(u2__abc_44228_n19074) );
  INVX1 INVX1_3387 ( .A(u2__abc_44228_n19077), .Y(u2__abc_44228_n19078) );
  INVX1 INVX1_3388 ( .A(u2__abc_44228_n19085), .Y(u2__abc_44228_n19086) );
  INVX1 INVX1_3389 ( .A(u2__abc_44228_n19089), .Y(u2__abc_44228_n19090) );
  INVX1 INVX1_339 ( .A(u2_remHi_47_), .Y(u2__abc_44228_n3454) );
  INVX1 INVX1_3390 ( .A(u2__abc_44228_n19097), .Y(u2__abc_44228_n19098) );
  INVX1 INVX1_3391 ( .A(u2__abc_44228_n19101), .Y(u2__abc_44228_n19102) );
  INVX1 INVX1_3392 ( .A(u2__abc_44228_n19109), .Y(u2__abc_44228_n19110) );
  INVX1 INVX1_3393 ( .A(u2__abc_44228_n19113), .Y(u2__abc_44228_n19114) );
  INVX1 INVX1_3394 ( .A(u2__abc_44228_n19121), .Y(u2__abc_44228_n19122) );
  INVX1 INVX1_3395 ( .A(u2__abc_44228_n19125), .Y(u2__abc_44228_n19126) );
  INVX1 INVX1_3396 ( .A(u2__abc_44228_n19133), .Y(u2__abc_44228_n19134) );
  INVX1 INVX1_3397 ( .A(u2__abc_44228_n19137), .Y(u2__abc_44228_n19138) );
  INVX1 INVX1_3398 ( .A(u2__abc_44228_n19145), .Y(u2__abc_44228_n19146) );
  INVX1 INVX1_3399 ( .A(u2__abc_44228_n19149), .Y(u2__abc_44228_n19150) );
  INVX1 INVX1_34 ( .A(_abc_64468_n1626), .Y(_abc_64468_n1627) );
  INVX1 INVX1_340 ( .A(u2__abc_44228_n3455), .Y(u2__abc_44228_n3456) );
  INVX1 INVX1_3400 ( .A(u2__abc_44228_n19157), .Y(u2__abc_44228_n19158) );
  INVX1 INVX1_3401 ( .A(u2__abc_44228_n19161), .Y(u2__abc_44228_n19162) );
  INVX1 INVX1_3402 ( .A(u2__abc_44228_n19169), .Y(u2__abc_44228_n19170) );
  INVX1 INVX1_3403 ( .A(u2__abc_44228_n19173), .Y(u2__abc_44228_n19174) );
  INVX1 INVX1_3404 ( .A(u2__abc_44228_n19181), .Y(u2__abc_44228_n19182) );
  INVX1 INVX1_3405 ( .A(u2__abc_44228_n19185), .Y(u2__abc_44228_n19186) );
  INVX1 INVX1_3406 ( .A(u2__abc_44228_n19193), .Y(u2__abc_44228_n19194) );
  INVX1 INVX1_3407 ( .A(u2__abc_44228_n19197), .Y(u2__abc_44228_n19198) );
  INVX1 INVX1_3408 ( .A(u2__abc_44228_n19205), .Y(u2__abc_44228_n19206) );
  INVX1 INVX1_3409 ( .A(u2__abc_44228_n19209), .Y(u2__abc_44228_n19210) );
  INVX1 INVX1_341 ( .A(sqrto_46_), .Y(u2__abc_44228_n3458) );
  INVX1 INVX1_3410 ( .A(u2__abc_44228_n19217), .Y(u2__abc_44228_n19218) );
  INVX1 INVX1_3411 ( .A(u2__abc_44228_n19221), .Y(u2__abc_44228_n19222) );
  INVX1 INVX1_3412 ( .A(u2__abc_44228_n19229), .Y(u2__abc_44228_n19230) );
  INVX1 INVX1_3413 ( .A(u2__abc_44228_n19233), .Y(u2__abc_44228_n19234) );
  INVX1 INVX1_3414 ( .A(u2__abc_44228_n19241), .Y(u2__abc_44228_n19242) );
  INVX1 INVX1_3415 ( .A(u2__abc_44228_n19245), .Y(u2__abc_44228_n19246) );
  INVX1 INVX1_3416 ( .A(u2__abc_44228_n19253), .Y(u2__abc_44228_n19254) );
  INVX1 INVX1_3417 ( .A(u2__abc_44228_n19257), .Y(u2__abc_44228_n19258) );
  INVX1 INVX1_3418 ( .A(u2__abc_44228_n19265), .Y(u2__abc_44228_n19266) );
  INVX1 INVX1_3419 ( .A(u2__abc_44228_n19269), .Y(u2__abc_44228_n19270) );
  INVX1 INVX1_342 ( .A(u2_remHi_46_), .Y(u2__abc_44228_n3460) );
  INVX1 INVX1_3420 ( .A(u2__abc_44228_n19277), .Y(u2__abc_44228_n19278) );
  INVX1 INVX1_3421 ( .A(u2__abc_44228_n19281), .Y(u2__abc_44228_n19282) );
  INVX1 INVX1_3422 ( .A(u2__abc_44228_n19289), .Y(u2__abc_44228_n19290) );
  INVX1 INVX1_3423 ( .A(u2__abc_44228_n19293), .Y(u2__abc_44228_n19294) );
  INVX1 INVX1_3424 ( .A(u2__abc_44228_n19301), .Y(u2__abc_44228_n19302) );
  INVX1 INVX1_3425 ( .A(u2__abc_44228_n19305), .Y(u2__abc_44228_n19306) );
  INVX1 INVX1_3426 ( .A(u2__abc_44228_n19313), .Y(u2__abc_44228_n19314) );
  INVX1 INVX1_3427 ( .A(u2__abc_44228_n19317), .Y(u2__abc_44228_n19318) );
  INVX1 INVX1_3428 ( .A(u2__abc_44228_n19325), .Y(u2__abc_44228_n19326) );
  INVX1 INVX1_3429 ( .A(u2__abc_44228_n19329), .Y(u2__abc_44228_n19330) );
  INVX1 INVX1_343 ( .A(u2__abc_44228_n3462), .Y(u2__abc_44228_n3463) );
  INVX1 INVX1_3430 ( .A(u2__abc_44228_n19337), .Y(u2__abc_44228_n19338) );
  INVX1 INVX1_3431 ( .A(u2__abc_44228_n19341), .Y(u2__abc_44228_n19342) );
  INVX1 INVX1_3432 ( .A(u2__abc_44228_n19349), .Y(u2__abc_44228_n19350) );
  INVX1 INVX1_3433 ( .A(u2__abc_44228_n19353), .Y(u2__abc_44228_n19354) );
  INVX1 INVX1_3434 ( .A(u2__abc_44228_n19361), .Y(u2__abc_44228_n19362) );
  INVX1 INVX1_3435 ( .A(u2__abc_44228_n19365), .Y(u2__abc_44228_n19366) );
  INVX1 INVX1_3436 ( .A(u2__abc_44228_n19373), .Y(u2__abc_44228_n19374) );
  INVX1 INVX1_3437 ( .A(u2__abc_44228_n19377), .Y(u2__abc_44228_n19378) );
  INVX1 INVX1_3438 ( .A(u2__abc_44228_n19385), .Y(u2__abc_44228_n19386) );
  INVX1 INVX1_3439 ( .A(u2__abc_44228_n19389), .Y(u2__abc_44228_n19390) );
  INVX1 INVX1_344 ( .A(sqrto_45_), .Y(u2__abc_44228_n3468) );
  INVX1 INVX1_3440 ( .A(u2__abc_44228_n19397), .Y(u2__abc_44228_n19398) );
  INVX1 INVX1_3441 ( .A(u2__abc_44228_n19401), .Y(u2__abc_44228_n19402) );
  INVX1 INVX1_3442 ( .A(u2__abc_44228_n19409), .Y(u2__abc_44228_n19410) );
  INVX1 INVX1_3443 ( .A(u2__abc_44228_n19413), .Y(u2__abc_44228_n19414) );
  INVX1 INVX1_3444 ( .A(u2__abc_44228_n19421), .Y(u2__abc_44228_n19422) );
  INVX1 INVX1_3445 ( .A(u2__abc_44228_n19425), .Y(u2__abc_44228_n19426) );
  INVX1 INVX1_3446 ( .A(u2__abc_44228_n19433), .Y(u2__abc_44228_n19434) );
  INVX1 INVX1_3447 ( .A(u2__abc_44228_n19437), .Y(u2__abc_44228_n19438) );
  INVX1 INVX1_3448 ( .A(u2__abc_44228_n19445), .Y(u2__abc_44228_n19446) );
  INVX1 INVX1_3449 ( .A(u2__abc_44228_n19449), .Y(u2__abc_44228_n19450) );
  INVX1 INVX1_345 ( .A(u2__abc_44228_n3469), .Y(u2__abc_44228_n3470) );
  INVX1 INVX1_3450 ( .A(u2__abc_44228_n19457), .Y(u2__abc_44228_n19458) );
  INVX1 INVX1_3451 ( .A(u2__abc_44228_n19461), .Y(u2__abc_44228_n19462) );
  INVX1 INVX1_3452 ( .A(u2__abc_44228_n19469), .Y(u2__abc_44228_n19470) );
  INVX1 INVX1_3453 ( .A(u2__abc_44228_n19473), .Y(u2__abc_44228_n19474) );
  INVX1 INVX1_3454 ( .A(u2__abc_44228_n19481), .Y(u2__abc_44228_n19482) );
  INVX1 INVX1_3455 ( .A(u2__abc_44228_n19485), .Y(u2__abc_44228_n19486) );
  INVX1 INVX1_3456 ( .A(u2__abc_44228_n19493), .Y(u2__abc_44228_n19494) );
  INVX1 INVX1_3457 ( .A(u2__abc_44228_n19497), .Y(u2__abc_44228_n19498) );
  INVX1 INVX1_3458 ( .A(u2__abc_44228_n19505), .Y(u2__abc_44228_n19506) );
  INVX1 INVX1_3459 ( .A(u2__abc_44228_n19509), .Y(u2__abc_44228_n19510) );
  INVX1 INVX1_346 ( .A(u2_remHi_45_), .Y(u2__abc_44228_n3471) );
  INVX1 INVX1_3460 ( .A(u2__abc_44228_n19517), .Y(u2__abc_44228_n19518) );
  INVX1 INVX1_3461 ( .A(u2__abc_44228_n19521), .Y(u2__abc_44228_n19522) );
  INVX1 INVX1_3462 ( .A(u2__abc_44228_n19529), .Y(u2__abc_44228_n19530) );
  INVX1 INVX1_3463 ( .A(u2__abc_44228_n19533), .Y(u2__abc_44228_n19534) );
  INVX1 INVX1_3464 ( .A(u2__abc_44228_n19541), .Y(u2__abc_44228_n19542) );
  INVX1 INVX1_3465 ( .A(u2__abc_44228_n19545), .Y(u2__abc_44228_n19546) );
  INVX1 INVX1_3466 ( .A(u2__abc_44228_n19553), .Y(u2__abc_44228_n19554) );
  INVX1 INVX1_3467 ( .A(u2__abc_44228_n19557), .Y(u2__abc_44228_n19558) );
  INVX1 INVX1_3468 ( .A(u2__abc_44228_n19565), .Y(u2__abc_44228_n19566) );
  INVX1 INVX1_3469 ( .A(u2__abc_44228_n19569), .Y(u2__abc_44228_n19570) );
  INVX1 INVX1_347 ( .A(u2__abc_44228_n3472), .Y(u2__abc_44228_n3473) );
  INVX1 INVX1_3470 ( .A(u2__abc_44228_n19577), .Y(u2__abc_44228_n19578) );
  INVX1 INVX1_3471 ( .A(u2__abc_44228_n19581), .Y(u2__abc_44228_n19582) );
  INVX1 INVX1_3472 ( .A(u2__abc_44228_n19589), .Y(u2__abc_44228_n19590) );
  INVX1 INVX1_3473 ( .A(u2__abc_44228_n19593), .Y(u2__abc_44228_n19594) );
  INVX1 INVX1_3474 ( .A(u2__abc_44228_n19601), .Y(u2__abc_44228_n19602) );
  INVX1 INVX1_3475 ( .A(u2__abc_44228_n19605), .Y(u2__abc_44228_n19606) );
  INVX1 INVX1_3476 ( .A(u2__abc_44228_n19613), .Y(u2__abc_44228_n19614) );
  INVX1 INVX1_3477 ( .A(u2__abc_44228_n19617), .Y(u2__abc_44228_n19618) );
  INVX1 INVX1_3478 ( .A(u2__abc_44228_n19625), .Y(u2__abc_44228_n19626) );
  INVX1 INVX1_3479 ( .A(u2__abc_44228_n19629), .Y(u2__abc_44228_n19630) );
  INVX1 INVX1_348 ( .A(sqrto_44_), .Y(u2__abc_44228_n3475_1) );
  INVX1 INVX1_3480 ( .A(u2__abc_44228_n19637), .Y(u2__abc_44228_n19638) );
  INVX1 INVX1_3481 ( .A(u2__abc_44228_n19641), .Y(u2__abc_44228_n19642) );
  INVX1 INVX1_3482 ( .A(u2__abc_44228_n19649), .Y(u2__abc_44228_n19650) );
  INVX1 INVX1_3483 ( .A(u2__abc_44228_n19653), .Y(u2__abc_44228_n19654) );
  INVX1 INVX1_3484 ( .A(u2__abc_44228_n19661), .Y(u2__abc_44228_n19662) );
  INVX1 INVX1_3485 ( .A(u2__abc_44228_n19665), .Y(u2__abc_44228_n19666) );
  INVX1 INVX1_3486 ( .A(u2__abc_44228_n19673), .Y(u2__abc_44228_n19674) );
  INVX1 INVX1_3487 ( .A(u2__abc_44228_n19677), .Y(u2__abc_44228_n19678) );
  INVX1 INVX1_3488 ( .A(u2__abc_44228_n19685), .Y(u2__abc_44228_n19686) );
  INVX1 INVX1_3489 ( .A(u2__abc_44228_n19689), .Y(u2__abc_44228_n19690) );
  INVX1 INVX1_349 ( .A(u2_remHi_44_), .Y(u2__abc_44228_n3477) );
  INVX1 INVX1_3490 ( .A(u2__abc_44228_n19697), .Y(u2__abc_44228_n19698) );
  INVX1 INVX1_3491 ( .A(u2__abc_44228_n19701), .Y(u2__abc_44228_n19702) );
  INVX1 INVX1_3492 ( .A(u2__abc_44228_n19709), .Y(u2__abc_44228_n19710) );
  INVX1 INVX1_3493 ( .A(u2__abc_44228_n19713), .Y(u2__abc_44228_n19714) );
  INVX1 INVX1_3494 ( .A(u2__abc_44228_n19721), .Y(u2__abc_44228_n19722) );
  INVX1 INVX1_3495 ( .A(u2__abc_44228_n19725), .Y(u2__abc_44228_n19726) );
  INVX1 INVX1_3496 ( .A(u2__abc_44228_n19733), .Y(u2__abc_44228_n19734) );
  INVX1 INVX1_3497 ( .A(u2__abc_44228_n19737), .Y(u2__abc_44228_n19738) );
  INVX1 INVX1_3498 ( .A(u2__abc_44228_n19745), .Y(u2__abc_44228_n19746) );
  INVX1 INVX1_3499 ( .A(u2__abc_44228_n19749), .Y(u2__abc_44228_n19750) );
  INVX1 INVX1_35 ( .A(_abc_64468_n1628), .Y(_abc_64468_n1629) );
  INVX1 INVX1_350 ( .A(u2__abc_44228_n3479), .Y(u2__abc_44228_n3480) );
  INVX1 INVX1_3500 ( .A(u2__abc_44228_n19757), .Y(u2__abc_44228_n19758) );
  INVX1 INVX1_3501 ( .A(u2__abc_44228_n19761), .Y(u2__abc_44228_n19762) );
  INVX1 INVX1_3502 ( .A(u2__abc_44228_n19769), .Y(u2__abc_44228_n19770) );
  INVX1 INVX1_3503 ( .A(u2__abc_44228_n19773), .Y(u2__abc_44228_n19774) );
  INVX1 INVX1_3504 ( .A(u2__abc_44228_n19781), .Y(u2__abc_44228_n19782) );
  INVX1 INVX1_3505 ( .A(u2__abc_44228_n19785), .Y(u2__abc_44228_n19786) );
  INVX1 INVX1_3506 ( .A(u2__abc_44228_n19793), .Y(u2__abc_44228_n19794) );
  INVX1 INVX1_3507 ( .A(u2__abc_44228_n19797), .Y(u2__abc_44228_n19798) );
  INVX1 INVX1_3508 ( .A(u2__abc_44228_n19805), .Y(u2__abc_44228_n19806) );
  INVX1 INVX1_3509 ( .A(u2__abc_44228_n19809), .Y(u2__abc_44228_n19810) );
  INVX1 INVX1_351 ( .A(sqrto_42_), .Y(u2__abc_44228_n3482) );
  INVX1 INVX1_3510 ( .A(u2__abc_44228_n19817), .Y(u2__abc_44228_n19818) );
  INVX1 INVX1_3511 ( .A(u2__abc_44228_n19821), .Y(u2__abc_44228_n19822) );
  INVX1 INVX1_3512 ( .A(u2__abc_44228_n19829), .Y(u2__abc_44228_n19830) );
  INVX1 INVX1_3513 ( .A(u2__abc_44228_n19833), .Y(u2__abc_44228_n19834) );
  INVX1 INVX1_3514 ( .A(u2__abc_44228_n19841), .Y(u2__abc_44228_n19842) );
  INVX1 INVX1_3515 ( .A(u2__abc_44228_n19845), .Y(u2__abc_44228_n19846) );
  INVX1 INVX1_3516 ( .A(u2__abc_44228_n19853), .Y(u2__abc_44228_n19854) );
  INVX1 INVX1_3517 ( .A(u2__abc_44228_n19857), .Y(u2__abc_44228_n19858) );
  INVX1 INVX1_3518 ( .A(u2__abc_44228_n19865), .Y(u2__abc_44228_n19866) );
  INVX1 INVX1_3519 ( .A(u2__abc_44228_n19869), .Y(u2__abc_44228_n19870) );
  INVX1 INVX1_352 ( .A(u2_remHi_42_), .Y(u2__abc_44228_n3484_1) );
  INVX1 INVX1_3520 ( .A(u2__abc_44228_n19877), .Y(u2__abc_44228_n19878) );
  INVX1 INVX1_3521 ( .A(u2__abc_44228_n19881), .Y(u2__abc_44228_n19882) );
  INVX1 INVX1_3522 ( .A(u2__abc_44228_n19889), .Y(u2__abc_44228_n19890) );
  INVX1 INVX1_3523 ( .A(u2__abc_44228_n19893), .Y(u2__abc_44228_n19894) );
  INVX1 INVX1_3524 ( .A(u2__abc_44228_n19901), .Y(u2__abc_44228_n19902) );
  INVX1 INVX1_3525 ( .A(u2__abc_44228_n19905), .Y(u2__abc_44228_n19906) );
  INVX1 INVX1_3526 ( .A(u2__abc_44228_n19913), .Y(u2__abc_44228_n19914) );
  INVX1 INVX1_3527 ( .A(u2__abc_44228_n19917), .Y(u2__abc_44228_n19918) );
  INVX1 INVX1_3528 ( .A(u2__abc_44228_n19925), .Y(u2__abc_44228_n19926) );
  INVX1 INVX1_3529 ( .A(u2__abc_44228_n19929), .Y(u2__abc_44228_n19930) );
  INVX1 INVX1_353 ( .A(u2__abc_44228_n3486), .Y(u2__abc_44228_n3487) );
  INVX1 INVX1_3530 ( .A(u2__abc_44228_n19937), .Y(u2__abc_44228_n19938) );
  INVX1 INVX1_3531 ( .A(u2__abc_44228_n19941), .Y(u2__abc_44228_n19942) );
  INVX1 INVX1_3532 ( .A(u2__abc_44228_n19949), .Y(u2__abc_44228_n19950) );
  INVX1 INVX1_3533 ( .A(u2__abc_44228_n19953), .Y(u2__abc_44228_n19954) );
  INVX1 INVX1_3534 ( .A(u2__abc_44228_n19961), .Y(u2__abc_44228_n19962) );
  INVX1 INVX1_3535 ( .A(u2__abc_44228_n19965), .Y(u2__abc_44228_n19966) );
  INVX1 INVX1_3536 ( .A(u2__abc_44228_n19973), .Y(u2__abc_44228_n19974) );
  INVX1 INVX1_3537 ( .A(u2__abc_44228_n19977), .Y(u2__abc_44228_n19978) );
  INVX1 INVX1_3538 ( .A(u2__abc_44228_n19985), .Y(u2__abc_44228_n19986) );
  INVX1 INVX1_3539 ( .A(u2__abc_44228_n19989), .Y(u2__abc_44228_n19990) );
  INVX1 INVX1_354 ( .A(sqrto_43_), .Y(u2__abc_44228_n3488) );
  INVX1 INVX1_3540 ( .A(u2__abc_44228_n19997), .Y(u2__abc_44228_n19998) );
  INVX1 INVX1_3541 ( .A(u2__abc_44228_n20001), .Y(u2__abc_44228_n20002) );
  INVX1 INVX1_3542 ( .A(u2__abc_44228_n20009), .Y(u2__abc_44228_n20010) );
  INVX1 INVX1_3543 ( .A(u2__abc_44228_n20013), .Y(u2__abc_44228_n20014) );
  INVX1 INVX1_3544 ( .A(u2__abc_44228_n20021), .Y(u2__abc_44228_n20022) );
  INVX1 INVX1_3545 ( .A(u2__abc_44228_n20025), .Y(u2__abc_44228_n20026) );
  INVX1 INVX1_3546 ( .A(u2__abc_44228_n20033), .Y(u2__abc_44228_n20034) );
  INVX1 INVX1_3547 ( .A(u2__abc_44228_n20037), .Y(u2__abc_44228_n20038) );
  INVX1 INVX1_3548 ( .A(u2__abc_44228_n20045), .Y(u2__abc_44228_n20046) );
  INVX1 INVX1_3549 ( .A(u2__abc_44228_n20049), .Y(u2__abc_44228_n20050) );
  INVX1 INVX1_355 ( .A(u2__abc_44228_n3489), .Y(u2__abc_44228_n3490) );
  INVX1 INVX1_3550 ( .A(u2__abc_44228_n20057), .Y(u2__abc_44228_n20058) );
  INVX1 INVX1_3551 ( .A(u2__abc_44228_n20061), .Y(u2__abc_44228_n20062) );
  INVX1 INVX1_3552 ( .A(u2__abc_44228_n20069), .Y(u2__abc_44228_n20070) );
  INVX1 INVX1_3553 ( .A(u2__abc_44228_n20073), .Y(u2__abc_44228_n20074) );
  INVX1 INVX1_3554 ( .A(u2__abc_44228_n20081), .Y(u2__abc_44228_n20082) );
  INVX1 INVX1_3555 ( .A(u2__abc_44228_n20085), .Y(u2__abc_44228_n20086) );
  INVX1 INVX1_3556 ( .A(u2__abc_44228_n20093), .Y(u2__abc_44228_n20094) );
  INVX1 INVX1_3557 ( .A(u2__abc_44228_n20097), .Y(u2__abc_44228_n20098) );
  INVX1 INVX1_3558 ( .A(u2__abc_44228_n20105), .Y(u2__abc_44228_n20106) );
  INVX1 INVX1_3559 ( .A(u2__abc_44228_n20109), .Y(u2__abc_44228_n20110) );
  INVX1 INVX1_356 ( .A(u2_remHi_43_), .Y(u2__abc_44228_n3491) );
  INVX1 INVX1_3560 ( .A(u2__abc_44228_n20117), .Y(u2__abc_44228_n20118) );
  INVX1 INVX1_3561 ( .A(u2__abc_44228_n20121), .Y(u2__abc_44228_n20122) );
  INVX1 INVX1_3562 ( .A(u2__abc_44228_n20129), .Y(u2__abc_44228_n20130) );
  INVX1 INVX1_3563 ( .A(u2__abc_44228_n20133), .Y(u2__abc_44228_n20134) );
  INVX1 INVX1_3564 ( .A(u2__abc_44228_n20141), .Y(u2__abc_44228_n20142) );
  INVX1 INVX1_3565 ( .A(u2__abc_44228_n20145), .Y(u2__abc_44228_n20146) );
  INVX1 INVX1_3566 ( .A(u2__abc_44228_n20153), .Y(u2__abc_44228_n20154) );
  INVX1 INVX1_3567 ( .A(u2__abc_44228_n20157), .Y(u2__abc_44228_n20158) );
  INVX1 INVX1_3568 ( .A(u2__abc_44228_n20165), .Y(u2__abc_44228_n20166) );
  INVX1 INVX1_3569 ( .A(u2__abc_44228_n20169), .Y(u2__abc_44228_n20170) );
  INVX1 INVX1_357 ( .A(u2__abc_44228_n3492), .Y(u2__abc_44228_n3493) );
  INVX1 INVX1_3570 ( .A(u2__abc_44228_n20177), .Y(u2__abc_44228_n20178) );
  INVX1 INVX1_3571 ( .A(u2__abc_44228_n20181), .Y(u2__abc_44228_n20182) );
  INVX1 INVX1_3572 ( .A(u2__abc_44228_n20189), .Y(u2__abc_44228_n20190) );
  INVX1 INVX1_3573 ( .A(u2__abc_44228_n20193), .Y(u2__abc_44228_n20194) );
  INVX1 INVX1_3574 ( .A(u2__abc_44228_n20201), .Y(u2__abc_44228_n20202) );
  INVX1 INVX1_3575 ( .A(u2__abc_44228_n20205), .Y(u2__abc_44228_n20206) );
  INVX1 INVX1_3576 ( .A(u2__abc_44228_n20213), .Y(u2__abc_44228_n20214) );
  INVX1 INVX1_3577 ( .A(u2__abc_44228_n20217), .Y(u2__abc_44228_n20218) );
  INVX1 INVX1_3578 ( .A(u2__abc_44228_n20225), .Y(u2__abc_44228_n20226) );
  INVX1 INVX1_3579 ( .A(u2__abc_44228_n20229), .Y(u2__abc_44228_n20230) );
  INVX1 INVX1_358 ( .A(sqrto_39_), .Y(u2__abc_44228_n3497) );
  INVX1 INVX1_3580 ( .A(u2__abc_44228_n20237), .Y(u2__abc_44228_n20238) );
  INVX1 INVX1_3581 ( .A(u2__abc_44228_n20241), .Y(u2__abc_44228_n20242) );
  INVX1 INVX1_3582 ( .A(u2__abc_44228_n20249), .Y(u2__abc_44228_n20250) );
  INVX1 INVX1_3583 ( .A(u2__abc_44228_n20253), .Y(u2__abc_44228_n20254) );
  INVX1 INVX1_3584 ( .A(u2__abc_44228_n20261), .Y(u2__abc_44228_n20262) );
  INVX1 INVX1_3585 ( .A(u2__abc_44228_n20265), .Y(u2__abc_44228_n20266) );
  INVX1 INVX1_3586 ( .A(u2__abc_44228_n20273), .Y(u2__abc_44228_n20274) );
  INVX1 INVX1_3587 ( .A(u2__abc_44228_n20277), .Y(u2__abc_44228_n20278) );
  INVX1 INVX1_3588 ( .A(u2__abc_44228_n20285), .Y(u2__abc_44228_n20286) );
  INVX1 INVX1_3589 ( .A(u2__abc_44228_n20289), .Y(u2__abc_44228_n20290) );
  INVX1 INVX1_359 ( .A(u2__abc_44228_n3498), .Y(u2__abc_44228_n3499) );
  INVX1 INVX1_3590 ( .A(u2__abc_44228_n20297), .Y(u2__abc_44228_n20298) );
  INVX1 INVX1_3591 ( .A(u2__abc_44228_n20301), .Y(u2__abc_44228_n20302) );
  INVX1 INVX1_3592 ( .A(u2__abc_44228_n20309), .Y(u2__abc_44228_n20310) );
  INVX1 INVX1_3593 ( .A(u2__abc_44228_n20313), .Y(u2__abc_44228_n20314) );
  INVX1 INVX1_3594 ( .A(u2__abc_44228_n20321), .Y(u2__abc_44228_n20322) );
  INVX1 INVX1_3595 ( .A(u2__abc_44228_n20325), .Y(u2__abc_44228_n20326) );
  INVX1 INVX1_3596 ( .A(u2__abc_44228_n20333), .Y(u2__abc_44228_n20334) );
  INVX1 INVX1_3597 ( .A(u2__abc_44228_n20337), .Y(u2__abc_44228_n20338) );
  INVX1 INVX1_3598 ( .A(u2__abc_44228_n20345), .Y(u2__abc_44228_n20346) );
  INVX1 INVX1_3599 ( .A(u2__abc_44228_n20349), .Y(u2__abc_44228_n20350) );
  INVX1 INVX1_36 ( .A(_abc_64468_n1631), .Y(_abc_64468_n1635) );
  INVX1 INVX1_360 ( .A(u2_remHi_39_), .Y(u2__abc_44228_n3500) );
  INVX1 INVX1_3600 ( .A(u2__abc_44228_n20357), .Y(u2__abc_44228_n20358) );
  INVX1 INVX1_3601 ( .A(u2__abc_44228_n20361), .Y(u2__abc_44228_n20362) );
  INVX1 INVX1_3602 ( .A(u2__abc_44228_n20369), .Y(u2__abc_44228_n20370) );
  INVX1 INVX1_3603 ( .A(u2__abc_44228_n20373), .Y(u2__abc_44228_n20374) );
  INVX1 INVX1_3604 ( .A(u2__abc_44228_n20381), .Y(u2__abc_44228_n20382) );
  INVX1 INVX1_3605 ( .A(u2__abc_44228_n20385), .Y(u2__abc_44228_n20386) );
  INVX1 INVX1_3606 ( .A(u2__abc_44228_n20393), .Y(u2__abc_44228_n20394) );
  INVX1 INVX1_3607 ( .A(u2__abc_44228_n20397), .Y(u2__abc_44228_n20398) );
  INVX1 INVX1_3608 ( .A(u2__abc_44228_n20405), .Y(u2__abc_44228_n20406) );
  INVX1 INVX1_3609 ( .A(u2__abc_44228_n20409), .Y(u2__abc_44228_n20410) );
  INVX1 INVX1_361 ( .A(u2__abc_44228_n3501), .Y(u2__abc_44228_n3502) );
  INVX1 INVX1_3610 ( .A(u2__abc_44228_n20417), .Y(u2__abc_44228_n20418) );
  INVX1 INVX1_3611 ( .A(u2__abc_44228_n20421), .Y(u2__abc_44228_n20422) );
  INVX1 INVX1_3612 ( .A(u2__abc_44228_n20429), .Y(u2__abc_44228_n20430) );
  INVX1 INVX1_3613 ( .A(u2__abc_44228_n20433), .Y(u2__abc_44228_n20434) );
  INVX1 INVX1_3614 ( .A(u2__abc_44228_n20441), .Y(u2__abc_44228_n20442) );
  INVX1 INVX1_3615 ( .A(u2__abc_44228_n20445), .Y(u2__abc_44228_n20446) );
  INVX1 INVX1_3616 ( .A(u2__abc_44228_n20453), .Y(u2__abc_44228_n20454) );
  INVX1 INVX1_3617 ( .A(u2__abc_44228_n20457), .Y(u2__abc_44228_n20458) );
  INVX1 INVX1_3618 ( .A(u2__abc_44228_n20465), .Y(u2__abc_44228_n20466) );
  INVX1 INVX1_3619 ( .A(u2__abc_44228_n20469), .Y(u2__abc_44228_n20470) );
  INVX1 INVX1_362 ( .A(sqrto_38_), .Y(u2__abc_44228_n3504) );
  INVX1 INVX1_3620 ( .A(u2__abc_44228_n20477), .Y(u2__abc_44228_n20478) );
  INVX1 INVX1_3621 ( .A(u2__abc_44228_n20481), .Y(u2__abc_44228_n20482) );
  INVX1 INVX1_3622 ( .A(u2__abc_44228_n20489), .Y(u2__abc_44228_n20490) );
  INVX1 INVX1_3623 ( .A(u2__abc_44228_n20493), .Y(u2__abc_44228_n20494) );
  INVX1 INVX1_3624 ( .A(u2__abc_44228_n20501), .Y(u2__abc_44228_n20502) );
  INVX1 INVX1_3625 ( .A(u2__abc_44228_n20505), .Y(u2__abc_44228_n20506) );
  INVX1 INVX1_3626 ( .A(u2__abc_44228_n20513), .Y(u2__abc_44228_n20514) );
  INVX1 INVX1_3627 ( .A(u2__abc_44228_n20517), .Y(u2__abc_44228_n20518) );
  INVX1 INVX1_3628 ( .A(u2__abc_44228_n20525), .Y(u2__abc_44228_n20526) );
  INVX1 INVX1_3629 ( .A(u2__abc_44228_n20529), .Y(u2__abc_44228_n20530) );
  INVX1 INVX1_363 ( .A(u2_remHi_38_), .Y(u2__abc_44228_n3506) );
  INVX1 INVX1_3630 ( .A(u2__abc_44228_n20537), .Y(u2__abc_44228_n20538) );
  INVX1 INVX1_3631 ( .A(u2__abc_44228_n20541), .Y(u2__abc_44228_n20542) );
  INVX1 INVX1_3632 ( .A(u2__abc_44228_n20549), .Y(u2__abc_44228_n20550) );
  INVX1 INVX1_3633 ( .A(u2__abc_44228_n20553), .Y(u2__abc_44228_n20554) );
  INVX1 INVX1_3634 ( .A(u2__abc_44228_n20561), .Y(u2__abc_44228_n20562) );
  INVX1 INVX1_3635 ( .A(u2__abc_44228_n20565), .Y(u2__abc_44228_n20566) );
  INVX1 INVX1_3636 ( .A(u2__abc_44228_n20573), .Y(u2__abc_44228_n20574) );
  INVX1 INVX1_3637 ( .A(u2__abc_44228_n20577), .Y(u2__abc_44228_n20578) );
  INVX1 INVX1_3638 ( .A(u2__abc_44228_n20585), .Y(u2__abc_44228_n20586) );
  INVX1 INVX1_3639 ( .A(u2__abc_44228_n20589), .Y(u2__abc_44228_n20590) );
  INVX1 INVX1_364 ( .A(u2__abc_44228_n3508), .Y(u2__abc_44228_n3509) );
  INVX1 INVX1_3640 ( .A(u2__abc_44228_n20597), .Y(u2__abc_44228_n20598) );
  INVX1 INVX1_3641 ( .A(u2__abc_44228_n20601), .Y(u2__abc_44228_n20602) );
  INVX1 INVX1_3642 ( .A(u2__abc_44228_n20609), .Y(u2__abc_44228_n20610) );
  INVX1 INVX1_3643 ( .A(u2__abc_44228_n20613), .Y(u2__abc_44228_n20614) );
  INVX1 INVX1_3644 ( .A(u2__abc_44228_n20621), .Y(u2__abc_44228_n20622) );
  INVX1 INVX1_3645 ( .A(u2__abc_44228_n20625), .Y(u2__abc_44228_n20626) );
  INVX1 INVX1_3646 ( .A(u2__abc_44228_n20633), .Y(u2__abc_44228_n20634) );
  INVX1 INVX1_3647 ( .A(u2__abc_44228_n20637), .Y(u2__abc_44228_n20638) );
  INVX1 INVX1_3648 ( .A(u2__abc_44228_n20645), .Y(u2__abc_44228_n20646) );
  INVX1 INVX1_3649 ( .A(u2__abc_44228_n20649), .Y(u2__abc_44228_n20650) );
  INVX1 INVX1_365 ( .A(sqrto_41_), .Y(u2__abc_44228_n3511) );
  INVX1 INVX1_3650 ( .A(u2__abc_44228_n20657), .Y(u2__abc_44228_n20658) );
  INVX1 INVX1_3651 ( .A(u2__abc_44228_n20661), .Y(u2__abc_44228_n20662) );
  INVX1 INVX1_3652 ( .A(u2__abc_44228_n20669), .Y(u2__abc_44228_n20670) );
  INVX1 INVX1_3653 ( .A(u2__abc_44228_n20673), .Y(u2__abc_44228_n20674) );
  INVX1 INVX1_3654 ( .A(u2__abc_44228_n20681), .Y(u2__abc_44228_n20682) );
  INVX1 INVX1_3655 ( .A(u2__abc_44228_n20685), .Y(u2__abc_44228_n20686) );
  INVX1 INVX1_3656 ( .A(u2__abc_44228_n20693), .Y(u2__abc_44228_n20694) );
  INVX1 INVX1_3657 ( .A(u2__abc_44228_n20697), .Y(u2__abc_44228_n20698) );
  INVX1 INVX1_3658 ( .A(u2__abc_44228_n20705), .Y(u2__abc_44228_n20706) );
  INVX1 INVX1_3659 ( .A(u2__abc_44228_n20709), .Y(u2__abc_44228_n20710) );
  INVX1 INVX1_366 ( .A(u2__abc_44228_n3512), .Y(u2__abc_44228_n3513_1) );
  INVX1 INVX1_3660 ( .A(u2__abc_44228_n20717), .Y(u2__abc_44228_n20718) );
  INVX1 INVX1_3661 ( .A(u2__abc_44228_n20721), .Y(u2__abc_44228_n20722) );
  INVX1 INVX1_3662 ( .A(u2__abc_44228_n20729), .Y(u2__abc_44228_n20730) );
  INVX1 INVX1_3663 ( .A(u2__abc_44228_n20733), .Y(u2__abc_44228_n20734) );
  INVX1 INVX1_3664 ( .A(u2__abc_44228_n20741), .Y(u2__abc_44228_n20742) );
  INVX1 INVX1_3665 ( .A(u2__abc_44228_n20745), .Y(u2__abc_44228_n20746) );
  INVX1 INVX1_3666 ( .A(u2__abc_44228_n20753), .Y(u2__abc_44228_n20754) );
  INVX1 INVX1_3667 ( .A(u2__abc_44228_n20757), .Y(u2__abc_44228_n20758) );
  INVX1 INVX1_3668 ( .A(u2__abc_44228_n20765), .Y(u2__abc_44228_n20766) );
  INVX1 INVX1_3669 ( .A(u2__abc_44228_n20769), .Y(u2__abc_44228_n20770) );
  INVX1 INVX1_367 ( .A(u2_remHi_41_), .Y(u2__abc_44228_n3514) );
  INVX1 INVX1_3670 ( .A(u2__abc_44228_n20777), .Y(u2__abc_44228_n20778) );
  INVX1 INVX1_3671 ( .A(u2__abc_44228_n20781), .Y(u2__abc_44228_n20782) );
  INVX1 INVX1_3672 ( .A(u2__abc_44228_n20789), .Y(u2__abc_44228_n20790) );
  INVX1 INVX1_3673 ( .A(u2__abc_44228_n20793), .Y(u2__abc_44228_n20794) );
  INVX1 INVX1_3674 ( .A(u2__abc_44228_n20801), .Y(u2__abc_44228_n20802) );
  INVX1 INVX1_3675 ( .A(u2__abc_44228_n20805), .Y(u2__abc_44228_n20806) );
  INVX1 INVX1_3676 ( .A(u2__abc_44228_n20813), .Y(u2__abc_44228_n20814) );
  INVX1 INVX1_3677 ( .A(u2__abc_44228_n20817), .Y(u2__abc_44228_n20818) );
  INVX1 INVX1_3678 ( .A(u2__abc_44228_n20825), .Y(u2__abc_44228_n20826) );
  INVX1 INVX1_3679 ( .A(u2__abc_44228_n20829), .Y(u2__abc_44228_n20830) );
  INVX1 INVX1_368 ( .A(u2__abc_44228_n3515), .Y(u2__abc_44228_n3516) );
  INVX1 INVX1_3680 ( .A(u2__abc_44228_n20837), .Y(u2__abc_44228_n20838) );
  INVX1 INVX1_3681 ( .A(u2__abc_44228_n20841), .Y(u2__abc_44228_n20842) );
  INVX1 INVX1_3682 ( .A(u2__abc_44228_n20849), .Y(u2__abc_44228_n20850) );
  INVX1 INVX1_3683 ( .A(u2__abc_44228_n20853), .Y(u2__abc_44228_n20854) );
  INVX1 INVX1_3684 ( .A(u2__abc_44228_n20861), .Y(u2__abc_44228_n20862) );
  INVX1 INVX1_3685 ( .A(u2__abc_44228_n20865), .Y(u2__abc_44228_n20866) );
  INVX1 INVX1_3686 ( .A(u2__abc_44228_n20873), .Y(u2__abc_44228_n20874) );
  INVX1 INVX1_3687 ( .A(u2__abc_44228_n20877), .Y(u2__abc_44228_n20878) );
  INVX1 INVX1_3688 ( .A(u2__abc_44228_n20885), .Y(u2__abc_44228_n20886) );
  INVX1 INVX1_3689 ( .A(u2__abc_44228_n20889), .Y(u2__abc_44228_n20890) );
  INVX1 INVX1_369 ( .A(sqrto_40_), .Y(u2__abc_44228_n3518) );
  INVX1 INVX1_3690 ( .A(u2__abc_44228_n20897), .Y(u2__abc_44228_n20898) );
  INVX1 INVX1_3691 ( .A(u2__abc_44228_n20901), .Y(u2__abc_44228_n20902) );
  INVX1 INVX1_3692 ( .A(u2__abc_44228_n20909), .Y(u2__abc_44228_n20910) );
  INVX1 INVX1_3693 ( .A(u2__abc_44228_n20913), .Y(u2__abc_44228_n20914) );
  INVX1 INVX1_3694 ( .A(u2__abc_44228_n20921), .Y(u2__abc_44228_n20922) );
  INVX1 INVX1_3695 ( .A(u2__abc_44228_n20925), .Y(u2__abc_44228_n20926) );
  INVX1 INVX1_3696 ( .A(u2__abc_44228_n20933), .Y(u2__abc_44228_n20934) );
  INVX1 INVX1_3697 ( .A(u2__abc_44228_n20937), .Y(u2__abc_44228_n20938) );
  INVX1 INVX1_3698 ( .A(u2__abc_44228_n20945), .Y(u2__abc_44228_n20946) );
  INVX1 INVX1_3699 ( .A(u2__abc_44228_n20949), .Y(u2__abc_44228_n20950) );
  INVX1 INVX1_37 ( .A(\a[123] ), .Y(_abc_64468_n1636) );
  INVX1 INVX1_370 ( .A(u2_remHi_40_), .Y(u2__abc_44228_n3520) );
  INVX1 INVX1_3700 ( .A(u2__abc_44228_n20957), .Y(u2__abc_44228_n20958) );
  INVX1 INVX1_3701 ( .A(u2__abc_44228_n20961), .Y(u2__abc_44228_n20962) );
  INVX1 INVX1_3702 ( .A(u2__abc_44228_n20969), .Y(u2__abc_44228_n20970) );
  INVX1 INVX1_3703 ( .A(u2__abc_44228_n20973), .Y(u2__abc_44228_n20974) );
  INVX1 INVX1_3704 ( .A(u2__abc_44228_n20981), .Y(u2__abc_44228_n20982) );
  INVX1 INVX1_3705 ( .A(u2__abc_44228_n20985), .Y(u2__abc_44228_n20986) );
  INVX1 INVX1_3706 ( .A(u2__abc_44228_n20993), .Y(u2__abc_44228_n20994) );
  INVX1 INVX1_3707 ( .A(u2__abc_44228_n20997), .Y(u2__abc_44228_n20998) );
  INVX1 INVX1_3708 ( .A(u2__abc_44228_n21005), .Y(u2__abc_44228_n21006) );
  INVX1 INVX1_3709 ( .A(u2__abc_44228_n21009), .Y(u2__abc_44228_n21010) );
  INVX1 INVX1_371 ( .A(u2__abc_44228_n3522), .Y(u2__abc_44228_n3523_1) );
  INVX1 INVX1_3710 ( .A(u2__abc_44228_n21017), .Y(u2__abc_44228_n21018) );
  INVX1 INVX1_3711 ( .A(u2__abc_44228_n21021), .Y(u2__abc_44228_n21022) );
  INVX1 INVX1_3712 ( .A(u2__abc_44228_n21029), .Y(u2__abc_44228_n21030) );
  INVX1 INVX1_3713 ( .A(u2__abc_44228_n21033), .Y(u2__abc_44228_n21034) );
  INVX1 INVX1_3714 ( .A(u2__abc_44228_n21041), .Y(u2__abc_44228_n21042) );
  INVX1 INVX1_3715 ( .A(u2__abc_44228_n21045), .Y(u2__abc_44228_n21046) );
  INVX1 INVX1_3716 ( .A(u2__abc_44228_n21053), .Y(u2__abc_44228_n21054) );
  INVX1 INVX1_3717 ( .A(u2__abc_44228_n21057), .Y(u2__abc_44228_n21058) );
  INVX1 INVX1_3718 ( .A(u2__abc_44228_n21065), .Y(u2__abc_44228_n21066) );
  INVX1 INVX1_3719 ( .A(u2__abc_44228_n21069), .Y(u2__abc_44228_n21070) );
  INVX1 INVX1_372 ( .A(sqrto_37_), .Y(u2__abc_44228_n3527) );
  INVX1 INVX1_3720 ( .A(u2__abc_44228_n21077), .Y(u2__abc_44228_n21078) );
  INVX1 INVX1_3721 ( .A(u2__abc_44228_n21081), .Y(u2__abc_44228_n21082) );
  INVX1 INVX1_3722 ( .A(u2__abc_44228_n21089), .Y(u2__abc_44228_n21090) );
  INVX1 INVX1_3723 ( .A(u2__abc_44228_n21093), .Y(u2__abc_44228_n21094) );
  INVX1 INVX1_3724 ( .A(u2__abc_44228_n21101), .Y(u2__abc_44228_n21102) );
  INVX1 INVX1_3725 ( .A(u2__abc_44228_n21105), .Y(u2__abc_44228_n21106) );
  INVX1 INVX1_3726 ( .A(u2__abc_44228_n21113), .Y(u2__abc_44228_n21114) );
  INVX1 INVX1_3727 ( .A(u2__abc_44228_n21117), .Y(u2__abc_44228_n21118) );
  INVX1 INVX1_3728 ( .A(u2__abc_44228_n21125), .Y(u2__abc_44228_n21126) );
  INVX1 INVX1_3729 ( .A(u2__abc_44228_n21129), .Y(u2__abc_44228_n21130) );
  INVX1 INVX1_373 ( .A(u2__abc_44228_n3528), .Y(u2__abc_44228_n3529) );
  INVX1 INVX1_3730 ( .A(u2__abc_44228_n21137), .Y(u2__abc_44228_n21138) );
  INVX1 INVX1_3731 ( .A(u2__abc_44228_n21141), .Y(u2__abc_44228_n21142) );
  INVX1 INVX1_3732 ( .A(u2__abc_44228_n21149), .Y(u2__abc_44228_n21150) );
  INVX1 INVX1_3733 ( .A(u2__abc_44228_n21153), .Y(u2__abc_44228_n21154) );
  INVX1 INVX1_3734 ( .A(u2__abc_44228_n21161), .Y(u2__abc_44228_n21162) );
  INVX1 INVX1_3735 ( .A(u2__abc_44228_n21165), .Y(u2__abc_44228_n21166) );
  INVX1 INVX1_3736 ( .A(u2__abc_44228_n21173), .Y(u2__abc_44228_n21174) );
  INVX1 INVX1_3737 ( .A(u2__abc_44228_n21177), .Y(u2__abc_44228_n21178) );
  INVX1 INVX1_3738 ( .A(u2__abc_44228_n21185), .Y(u2__abc_44228_n21186) );
  INVX1 INVX1_3739 ( .A(u2__abc_44228_n21189), .Y(u2__abc_44228_n21190) );
  INVX1 INVX1_374 ( .A(u2_remHi_37_), .Y(u2__abc_44228_n3530) );
  INVX1 INVX1_3740 ( .A(u2__abc_44228_n21197), .Y(u2__abc_44228_n21198) );
  INVX1 INVX1_3741 ( .A(u2__abc_44228_n21201), .Y(u2__abc_44228_n21202) );
  INVX1 INVX1_3742 ( .A(u2__abc_44228_n21209), .Y(u2__abc_44228_n21210) );
  INVX1 INVX1_3743 ( .A(u2__abc_44228_n21213), .Y(u2__abc_44228_n21214) );
  INVX1 INVX1_3744 ( .A(u2__abc_44228_n21221), .Y(u2__abc_44228_n21222) );
  INVX1 INVX1_3745 ( .A(u2__abc_44228_n21225), .Y(u2__abc_44228_n21226) );
  INVX1 INVX1_3746 ( .A(u2__abc_44228_n21233), .Y(u2__abc_44228_n21234) );
  INVX1 INVX1_3747 ( .A(u2__abc_44228_n21237), .Y(u2__abc_44228_n21238) );
  INVX1 INVX1_3748 ( .A(u2__abc_44228_n21245), .Y(u2__abc_44228_n21246) );
  INVX1 INVX1_3749 ( .A(u2__abc_44228_n21249), .Y(u2__abc_44228_n21250) );
  INVX1 INVX1_375 ( .A(u2__abc_44228_n3531), .Y(u2__abc_44228_n3532_1) );
  INVX1 INVX1_3750 ( .A(u2__abc_44228_n21257), .Y(u2__abc_44228_n21258) );
  INVX1 INVX1_3751 ( .A(u2__abc_44228_n21261), .Y(u2__abc_44228_n21262) );
  INVX1 INVX1_3752 ( .A(u2__abc_44228_n21269), .Y(u2__abc_44228_n21270) );
  INVX1 INVX1_3753 ( .A(u2__abc_44228_n21273), .Y(u2__abc_44228_n21274) );
  INVX1 INVX1_3754 ( .A(u2__abc_44228_n21281), .Y(u2__abc_44228_n21282) );
  INVX1 INVX1_3755 ( .A(u2__abc_44228_n21285), .Y(u2__abc_44228_n21286) );
  INVX1 INVX1_3756 ( .A(u2__abc_44228_n21293), .Y(u2__abc_44228_n21294) );
  INVX1 INVX1_3757 ( .A(u2__abc_44228_n21297), .Y(u2__abc_44228_n21298) );
  INVX1 INVX1_3758 ( .A(u2__abc_44228_n21305), .Y(u2__abc_44228_n21306) );
  INVX1 INVX1_3759 ( .A(u2__abc_44228_n21309), .Y(u2__abc_44228_n21310) );
  INVX1 INVX1_376 ( .A(sqrto_36_), .Y(u2__abc_44228_n3534) );
  INVX1 INVX1_3760 ( .A(u2__abc_44228_n21317), .Y(u2__abc_44228_n21318) );
  INVX1 INVX1_3761 ( .A(u2__abc_44228_n21321), .Y(u2__abc_44228_n21322) );
  INVX1 INVX1_3762 ( .A(u2__abc_44228_n21329), .Y(u2__abc_44228_n21330) );
  INVX1 INVX1_3763 ( .A(u2__abc_44228_n21333), .Y(u2__abc_44228_n21334) );
  INVX1 INVX1_3764 ( .A(u2__abc_44228_n21341), .Y(u2__abc_44228_n21342) );
  INVX1 INVX1_3765 ( .A(u2__abc_44228_n21345), .Y(u2__abc_44228_n21346) );
  INVX1 INVX1_3766 ( .A(u2__abc_44228_n21353), .Y(u2__abc_44228_n21354) );
  INVX1 INVX1_3767 ( .A(u2__abc_44228_n21357), .Y(u2__abc_44228_n21358) );
  INVX1 INVX1_3768 ( .A(u2__abc_44228_n21365), .Y(u2__abc_44228_n21366) );
  INVX1 INVX1_3769 ( .A(u2__abc_44228_n21369), .Y(u2__abc_44228_n21370) );
  INVX1 INVX1_377 ( .A(u2_remHi_36_), .Y(u2__abc_44228_n3536) );
  INVX1 INVX1_3770 ( .A(u2__abc_44228_n21377), .Y(u2__abc_44228_n21378) );
  INVX1 INVX1_3771 ( .A(u2__abc_44228_n21381), .Y(u2__abc_44228_n21382) );
  INVX1 INVX1_3772 ( .A(u2__abc_44228_n21389), .Y(u2__abc_44228_n21390) );
  INVX1 INVX1_3773 ( .A(u2__abc_44228_n21393), .Y(u2__abc_44228_n21394) );
  INVX1 INVX1_3774 ( .A(u2__abc_44228_n21401), .Y(u2__abc_44228_n21402) );
  INVX1 INVX1_3775 ( .A(u2__abc_44228_n21405), .Y(u2__abc_44228_n21406) );
  INVX1 INVX1_3776 ( .A(u2__abc_44228_n21413), .Y(u2__abc_44228_n21414) );
  INVX1 INVX1_3777 ( .A(u2__abc_44228_n21417), .Y(u2__abc_44228_n21418) );
  INVX1 INVX1_3778 ( .A(u2__abc_44228_n21425), .Y(u2__abc_44228_n21426) );
  INVX1 INVX1_3779 ( .A(u2__abc_44228_n21429), .Y(u2__abc_44228_n21430) );
  INVX1 INVX1_378 ( .A(u2__abc_44228_n3538), .Y(u2__abc_44228_n3539) );
  INVX1 INVX1_3780 ( .A(u2__abc_44228_n21437), .Y(u2__abc_44228_n21438) );
  INVX1 INVX1_3781 ( .A(u2__abc_44228_n21441), .Y(u2__abc_44228_n21442) );
  INVX1 INVX1_3782 ( .A(u2__abc_44228_n21449), .Y(u2__abc_44228_n21450) );
  INVX1 INVX1_3783 ( .A(u2__abc_44228_n21453), .Y(u2__abc_44228_n21454) );
  INVX1 INVX1_3784 ( .A(u2__abc_44228_n21461), .Y(u2__abc_44228_n21462) );
  INVX1 INVX1_3785 ( .A(u2__abc_44228_n21465), .Y(u2__abc_44228_n21466) );
  INVX1 INVX1_3786 ( .A(u2__abc_44228_n21473), .Y(u2__abc_44228_n21474) );
  INVX1 INVX1_3787 ( .A(u2__abc_44228_n21477), .Y(u2__abc_44228_n21478) );
  INVX1 INVX1_3788 ( .A(u2__abc_44228_n21485), .Y(u2__abc_44228_n21486) );
  INVX1 INVX1_3789 ( .A(u2__abc_44228_n21489), .Y(u2__abc_44228_n21490) );
  INVX1 INVX1_379 ( .A(sqrto_34_), .Y(u2__abc_44228_n3541_1) );
  INVX1 INVX1_3790 ( .A(u2__abc_44228_n21497), .Y(u2__abc_44228_n21498) );
  INVX1 INVX1_3791 ( .A(u2__abc_44228_n21501), .Y(u2__abc_44228_n21502) );
  INVX1 INVX1_3792 ( .A(u2__abc_44228_n21509), .Y(u2__abc_44228_n21510) );
  INVX1 INVX1_3793 ( .A(u2__abc_44228_n21513), .Y(u2__abc_44228_n21514) );
  INVX1 INVX1_3794 ( .A(u2__abc_44228_n21521), .Y(u2__abc_44228_n21522) );
  INVX1 INVX1_3795 ( .A(u2__abc_44228_n21525), .Y(u2__abc_44228_n21526) );
  INVX1 INVX1_3796 ( .A(u2__abc_44228_n21533), .Y(u2__abc_44228_n21534) );
  INVX1 INVX1_3797 ( .A(u2__abc_44228_n21537), .Y(u2__abc_44228_n21538) );
  INVX1 INVX1_3798 ( .A(u2__abc_44228_n21545), .Y(u2__abc_44228_n21546) );
  INVX1 INVX1_3799 ( .A(u2__abc_44228_n21549), .Y(u2__abc_44228_n21550) );
  INVX1 INVX1_38 ( .A(_abc_64468_n1639), .Y(_abc_64468_n1640) );
  INVX1 INVX1_380 ( .A(u2_remHi_34_), .Y(u2__abc_44228_n3543) );
  INVX1 INVX1_3800 ( .A(u2__abc_44228_n21557), .Y(u2__abc_44228_n21558) );
  INVX1 INVX1_3801 ( .A(u2__abc_44228_n21561), .Y(u2__abc_44228_n21562) );
  INVX1 INVX1_3802 ( .A(u2__abc_44228_n21569), .Y(u2__abc_44228_n21570) );
  INVX1 INVX1_3803 ( .A(u2__abc_44228_n21573), .Y(u2__abc_44228_n21574) );
  INVX1 INVX1_3804 ( .A(u2__abc_44228_n21581), .Y(u2__abc_44228_n21582) );
  INVX1 INVX1_3805 ( .A(u2__abc_44228_n21585), .Y(u2__abc_44228_n21586) );
  INVX1 INVX1_3806 ( .A(u2__abc_44228_n21593), .Y(u2__abc_44228_n21594) );
  INVX1 INVX1_3807 ( .A(u2__abc_44228_n21597), .Y(u2__abc_44228_n21598) );
  INVX1 INVX1_3808 ( .A(u2__abc_44228_n21605), .Y(u2__abc_44228_n21606) );
  INVX1 INVX1_3809 ( .A(u2__abc_44228_n21609), .Y(u2__abc_44228_n21610) );
  INVX1 INVX1_381 ( .A(u2__abc_44228_n3545), .Y(u2__abc_44228_n3546) );
  INVX1 INVX1_3810 ( .A(u2__abc_44228_n21617), .Y(u2__abc_44228_n21618) );
  INVX1 INVX1_3811 ( .A(u2__abc_44228_n21621), .Y(u2__abc_44228_n21622) );
  INVX1 INVX1_3812 ( .A(u2__abc_44228_n21629), .Y(u2__abc_44228_n21630) );
  INVX1 INVX1_3813 ( .A(u2__abc_44228_n21633), .Y(u2__abc_44228_n21634) );
  INVX1 INVX1_3814 ( .A(u2__abc_44228_n21641), .Y(u2__abc_44228_n21642) );
  INVX1 INVX1_3815 ( .A(u2__abc_44228_n21645), .Y(u2__abc_44228_n21646) );
  INVX1 INVX1_3816 ( .A(u2__abc_44228_n21653), .Y(u2__abc_44228_n21654) );
  INVX1 INVX1_3817 ( .A(u2__abc_44228_n21657), .Y(u2__abc_44228_n21658) );
  INVX1 INVX1_3818 ( .A(u2__abc_44228_n21665), .Y(u2__abc_44228_n21666) );
  INVX1 INVX1_3819 ( .A(u2__abc_44228_n21669), .Y(u2__abc_44228_n21670) );
  INVX1 INVX1_382 ( .A(sqrto_35_), .Y(u2__abc_44228_n3547) );
  INVX1 INVX1_3820 ( .A(u2__abc_44228_n21677), .Y(u2__abc_44228_n21678) );
  INVX1 INVX1_3821 ( .A(u2__abc_44228_n21681), .Y(u2__abc_44228_n21682) );
  INVX1 INVX1_3822 ( .A(u2__abc_44228_n21689), .Y(u2__abc_44228_n21690) );
  INVX1 INVX1_3823 ( .A(u2__abc_44228_n21693), .Y(u2__abc_44228_n21694) );
  INVX1 INVX1_3824 ( .A(u2__abc_44228_n21701), .Y(u2__abc_44228_n21702) );
  INVX1 INVX1_3825 ( .A(u2__abc_44228_n21705), .Y(u2__abc_44228_n21706) );
  INVX1 INVX1_3826 ( .A(u2__abc_44228_n21713), .Y(u2__abc_44228_n21714) );
  INVX1 INVX1_3827 ( .A(u2__abc_44228_n21717), .Y(u2__abc_44228_n21718) );
  INVX1 INVX1_3828 ( .A(u2__abc_44228_n21725), .Y(u2__abc_44228_n21726) );
  INVX1 INVX1_3829 ( .A(u2__abc_44228_n21729), .Y(u2__abc_44228_n21730) );
  INVX1 INVX1_383 ( .A(u2__abc_44228_n3548), .Y(u2__abc_44228_n3549) );
  INVX1 INVX1_3830 ( .A(u2__abc_44228_n21737), .Y(u2__abc_44228_n21738) );
  INVX1 INVX1_3831 ( .A(u2__abc_44228_n21741), .Y(u2__abc_44228_n21742) );
  INVX1 INVX1_3832 ( .A(u2__abc_44228_n21749), .Y(u2__abc_44228_n21750) );
  INVX1 INVX1_3833 ( .A(u2__abc_44228_n21753), .Y(u2__abc_44228_n21754) );
  INVX1 INVX1_3834 ( .A(u2__abc_44228_n21761), .Y(u2__abc_44228_n21762) );
  INVX1 INVX1_3835 ( .A(u2__abc_44228_n21765), .Y(u2__abc_44228_n21766) );
  INVX1 INVX1_3836 ( .A(u2__abc_44228_n21773), .Y(u2__abc_44228_n21774) );
  INVX1 INVX1_3837 ( .A(u2__abc_44228_n21777), .Y(u2__abc_44228_n21778) );
  INVX1 INVX1_3838 ( .A(u2__abc_44228_n21785), .Y(u2__abc_44228_n21786) );
  INVX1 INVX1_3839 ( .A(u2__abc_44228_n21789), .Y(u2__abc_44228_n21790) );
  INVX1 INVX1_384 ( .A(u2_remHi_35_), .Y(u2__abc_44228_n3550) );
  INVX1 INVX1_3840 ( .A(u2__abc_44228_n21797), .Y(u2__abc_44228_n21798) );
  INVX1 INVX1_3841 ( .A(u2__abc_44228_n21801), .Y(u2__abc_44228_n21802) );
  INVX1 INVX1_3842 ( .A(u2__abc_44228_n21809), .Y(u2__abc_44228_n21810) );
  INVX1 INVX1_3843 ( .A(u2__abc_44228_n21813), .Y(u2__abc_44228_n21814) );
  INVX1 INVX1_3844 ( .A(u2__abc_44228_n21821), .Y(u2__abc_44228_n21822) );
  INVX1 INVX1_3845 ( .A(u2__abc_44228_n21825), .Y(u2__abc_44228_n21826) );
  INVX1 INVX1_3846 ( .A(u2__abc_44228_n21833), .Y(u2__abc_44228_n21834) );
  INVX1 INVX1_3847 ( .A(u2__abc_44228_n21837), .Y(u2__abc_44228_n21838) );
  INVX1 INVX1_3848 ( .A(u2__abc_44228_n21845), .Y(u2__abc_44228_n21846) );
  INVX1 INVX1_3849 ( .A(u2__abc_44228_n21849), .Y(u2__abc_44228_n21850) );
  INVX1 INVX1_385 ( .A(u2__abc_44228_n3551), .Y(u2__abc_44228_n3552_1) );
  INVX1 INVX1_3850 ( .A(u2__abc_44228_n21857), .Y(u2__abc_44228_n21858) );
  INVX1 INVX1_3851 ( .A(u2__abc_44228_n21861), .Y(u2__abc_44228_n21862) );
  INVX1 INVX1_3852 ( .A(u2__abc_44228_n21869), .Y(u2__abc_44228_n21870) );
  INVX1 INVX1_3853 ( .A(u2__abc_44228_n21873), .Y(u2__abc_44228_n21874) );
  INVX1 INVX1_3854 ( .A(u2__abc_44228_n21881), .Y(u2__abc_44228_n21882) );
  INVX1 INVX1_3855 ( .A(u2__abc_44228_n21885), .Y(u2__abc_44228_n21886) );
  INVX1 INVX1_3856 ( .A(u2__abc_44228_n21893), .Y(u2__abc_44228_n21894) );
  INVX1 INVX1_3857 ( .A(u2__abc_44228_n21897), .Y(u2__abc_44228_n21898) );
  INVX1 INVX1_3858 ( .A(u2__abc_44228_n21905), .Y(u2__abc_44228_n21906) );
  INVX1 INVX1_3859 ( .A(u2__abc_44228_n21909), .Y(u2__abc_44228_n21910) );
  INVX1 INVX1_386 ( .A(u2_remHi_33_), .Y(u2__abc_44228_n3556) );
  INVX1 INVX1_3860 ( .A(u2__abc_44228_n21917), .Y(u2__abc_44228_n21918) );
  INVX1 INVX1_3861 ( .A(u2__abc_44228_n21921), .Y(u2__abc_44228_n21922) );
  INVX1 INVX1_3862 ( .A(u2__abc_44228_n21929), .Y(u2__abc_44228_n21930) );
  INVX1 INVX1_3863 ( .A(u2__abc_44228_n21933), .Y(u2__abc_44228_n21934) );
  INVX1 INVX1_3864 ( .A(u2__abc_44228_n21941), .Y(u2__abc_44228_n21942) );
  INVX1 INVX1_3865 ( .A(u2__abc_44228_n21945), .Y(u2__abc_44228_n21946) );
  INVX1 INVX1_3866 ( .A(u2__abc_44228_n21953), .Y(u2__abc_44228_n21954) );
  INVX1 INVX1_3867 ( .A(u2__abc_44228_n21957), .Y(u2__abc_44228_n21958) );
  INVX1 INVX1_3868 ( .A(u2__abc_44228_n21965), .Y(u2__abc_44228_n21966) );
  INVX1 INVX1_3869 ( .A(u2__abc_44228_n21969), .Y(u2__abc_44228_n21970) );
  INVX1 INVX1_387 ( .A(sqrto_33_), .Y(u2__abc_44228_n3558) );
  INVX1 INVX1_3870 ( .A(u2__abc_44228_n21977), .Y(u2__abc_44228_n21978) );
  INVX1 INVX1_3871 ( .A(u2__abc_44228_n21981), .Y(u2__abc_44228_n21982) );
  INVX1 INVX1_3872 ( .A(u2__abc_44228_n21989), .Y(u2__abc_44228_n21990) );
  INVX1 INVX1_3873 ( .A(u2__abc_44228_n21993), .Y(u2__abc_44228_n21994) );
  INVX1 INVX1_3874 ( .A(u2__abc_44228_n22001), .Y(u2__abc_44228_n22002) );
  INVX1 INVX1_3875 ( .A(u2__abc_44228_n22005), .Y(u2__abc_44228_n22006) );
  INVX1 INVX1_3876 ( .A(u2__abc_44228_n22013), .Y(u2__abc_44228_n22014) );
  INVX1 INVX1_3877 ( .A(u2__abc_44228_n22017), .Y(u2__abc_44228_n22018) );
  INVX1 INVX1_3878 ( .A(u2__abc_44228_n22025), .Y(u2__abc_44228_n22026) );
  INVX1 INVX1_3879 ( .A(u2__abc_44228_n22029), .Y(u2__abc_44228_n22030) );
  INVX1 INVX1_388 ( .A(u2_remHi_32_), .Y(u2__abc_44228_n3561) );
  INVX1 INVX1_3880 ( .A(u2__abc_44228_n22037), .Y(u2__abc_44228_n22038) );
  INVX1 INVX1_3881 ( .A(u2__abc_44228_n22041), .Y(u2__abc_44228_n22042) );
  INVX1 INVX1_3882 ( .A(u2__abc_44228_n22049), .Y(u2__abc_44228_n22050) );
  INVX1 INVX1_3883 ( .A(u2__abc_44228_n22053), .Y(u2__abc_44228_n22054) );
  INVX1 INVX1_3884 ( .A(u2__abc_44228_n22061), .Y(u2__abc_44228_n22062) );
  INVX1 INVX1_3885 ( .A(u2__abc_44228_n22065), .Y(u2__abc_44228_n22066) );
  INVX1 INVX1_3886 ( .A(u2__abc_44228_n22073), .Y(u2__abc_44228_n22074) );
  INVX1 INVX1_3887 ( .A(u2__abc_44228_n22077), .Y(u2__abc_44228_n22078) );
  INVX1 INVX1_3888 ( .A(u2__abc_44228_n22085), .Y(u2__abc_44228_n22086) );
  INVX1 INVX1_3889 ( .A(u2__abc_44228_n22089), .Y(u2__abc_44228_n22090) );
  INVX1 INVX1_389 ( .A(sqrto_32_), .Y(u2__abc_44228_n3563) );
  INVX1 INVX1_3890 ( .A(u2__abc_44228_n22097), .Y(u2__abc_44228_n22098) );
  INVX1 INVX1_3891 ( .A(u2__abc_44228_n22101), .Y(u2__abc_44228_n22102) );
  INVX1 INVX1_3892 ( .A(u2__abc_44228_n22109), .Y(u2__abc_44228_n22110) );
  INVX1 INVX1_3893 ( .A(u2__abc_44228_n22113), .Y(u2__abc_44228_n22114) );
  INVX1 INVX1_3894 ( .A(u2__abc_44228_n22121), .Y(u2__abc_44228_n22122) );
  INVX1 INVX1_3895 ( .A(u2__abc_44228_n22125), .Y(u2__abc_44228_n22126) );
  INVX1 INVX1_3896 ( .A(u2__abc_44228_n22133), .Y(u2__abc_44228_n22134) );
  INVX1 INVX1_3897 ( .A(u2__abc_44228_n22137), .Y(u2__abc_44228_n22138) );
  INVX1 INVX1_3898 ( .A(u2__abc_44228_n22145), .Y(u2__abc_44228_n22146) );
  INVX1 INVX1_3899 ( .A(u2__abc_44228_n22149), .Y(u2__abc_44228_n22150) );
  INVX1 INVX1_39 ( .A(_abc_64468_n1641), .Y(_abc_64468_n1642) );
  INVX1 INVX1_390 ( .A(sqrto_30_), .Y(u2__abc_44228_n3567) );
  INVX1 INVX1_3900 ( .A(u2__abc_44228_n22157), .Y(u2__abc_44228_n22158) );
  INVX1 INVX1_3901 ( .A(u2__abc_44228_n22161), .Y(u2__abc_44228_n22162) );
  INVX1 INVX1_3902 ( .A(u2__abc_44228_n22169), .Y(u2__abc_44228_n22170) );
  INVX1 INVX1_3903 ( .A(u2__abc_44228_n22173), .Y(u2__abc_44228_n22174) );
  INVX1 INVX1_3904 ( .A(u2__abc_44228_n22181), .Y(u2__abc_44228_n22182) );
  INVX1 INVX1_3905 ( .A(u2__abc_44228_n22185), .Y(u2__abc_44228_n22186) );
  INVX1 INVX1_3906 ( .A(u2__abc_44228_n22193), .Y(u2__abc_44228_n22194) );
  INVX1 INVX1_3907 ( .A(u2__abc_44228_n22197), .Y(u2__abc_44228_n22198) );
  INVX1 INVX1_3908 ( .A(u2__abc_44228_n22205), .Y(u2__abc_44228_n22206) );
  INVX1 INVX1_3909 ( .A(u2__abc_44228_n22209), .Y(u2__abc_44228_n22210) );
  INVX1 INVX1_391 ( .A(u2_remHi_30_), .Y(u2__abc_44228_n3569) );
  INVX1 INVX1_3910 ( .A(u2__abc_44228_n22217), .Y(u2__abc_44228_n22218) );
  INVX1 INVX1_3911 ( .A(u2__abc_44228_n22221), .Y(u2__abc_44228_n22222) );
  INVX1 INVX1_3912 ( .A(u2__abc_44228_n22229), .Y(u2__abc_44228_n22230) );
  INVX1 INVX1_3913 ( .A(u2__abc_44228_n22233), .Y(u2__abc_44228_n22234) );
  INVX1 INVX1_3914 ( .A(u2__abc_44228_n22241), .Y(u2__abc_44228_n22242) );
  INVX1 INVX1_3915 ( .A(u2__abc_44228_n22245), .Y(u2__abc_44228_n22246) );
  INVX1 INVX1_3916 ( .A(u2__abc_44228_n22253), .Y(u2__abc_44228_n22254) );
  INVX1 INVX1_3917 ( .A(u2__abc_44228_n22257), .Y(u2__abc_44228_n22258) );
  INVX1 INVX1_3918 ( .A(u2__abc_44228_n22265), .Y(u2__abc_44228_n22266) );
  INVX1 INVX1_3919 ( .A(u2__abc_44228_n22269), .Y(u2__abc_44228_n22270) );
  INVX1 INVX1_392 ( .A(u2__abc_44228_n3571_1), .Y(u2__abc_44228_n3572) );
  INVX1 INVX1_3920 ( .A(u2__abc_44228_n22277), .Y(u2__abc_44228_n22278) );
  INVX1 INVX1_3921 ( .A(u2__abc_44228_n22281), .Y(u2__abc_44228_n22282) );
  INVX1 INVX1_3922 ( .A(u2__abc_44228_n22289), .Y(u2__abc_44228_n22290) );
  INVX1 INVX1_3923 ( .A(u2__abc_44228_n22293), .Y(u2__abc_44228_n22294) );
  INVX1 INVX1_3924 ( .A(u2__abc_44228_n22301), .Y(u2__abc_44228_n22302) );
  INVX1 INVX1_3925 ( .A(u2__abc_44228_n22305), .Y(u2__abc_44228_n22306) );
  INVX1 INVX1_3926 ( .A(u2__abc_44228_n22313), .Y(u2__abc_44228_n22314) );
  INVX1 INVX1_3927 ( .A(u2__abc_44228_n22317), .Y(u2__abc_44228_n22318) );
  INVX1 INVX1_3928 ( .A(u2__abc_44228_n22325), .Y(u2__abc_44228_n22326) );
  INVX1 INVX1_3929 ( .A(u2__abc_44228_n22329), .Y(u2__abc_44228_n22330) );
  INVX1 INVX1_393 ( .A(sqrto_31_), .Y(u2__abc_44228_n3573) );
  INVX1 INVX1_3930 ( .A(u2__abc_44228_n22337), .Y(u2__abc_44228_n22338) );
  INVX1 INVX1_3931 ( .A(u2__abc_44228_n22341), .Y(u2__abc_44228_n22342) );
  INVX1 INVX1_3932 ( .A(u2__abc_44228_n22349), .Y(u2__abc_44228_n22350) );
  INVX1 INVX1_3933 ( .A(u2__abc_44228_n22353), .Y(u2__abc_44228_n22354) );
  INVX1 INVX1_3934 ( .A(u2__abc_44228_n22361), .Y(u2__abc_44228_n22362) );
  INVX1 INVX1_3935 ( .A(u2__abc_44228_n22365), .Y(u2__abc_44228_n22366) );
  INVX1 INVX1_3936 ( .A(u2__abc_44228_n22373), .Y(u2__abc_44228_n22374) );
  INVX1 INVX1_3937 ( .A(u2__abc_44228_n22377), .Y(u2__abc_44228_n22378) );
  INVX1 INVX1_3938 ( .A(u2__abc_44228_n22385), .Y(u2__abc_44228_n22386) );
  INVX1 INVX1_3939 ( .A(u2__abc_44228_n22389), .Y(u2__abc_44228_n22390) );
  INVX1 INVX1_394 ( .A(u2__abc_44228_n3574), .Y(u2__abc_44228_n3575) );
  INVX1 INVX1_3940 ( .A(u2__abc_44228_n22397), .Y(u2__abc_44228_n22398) );
  INVX1 INVX1_3941 ( .A(u2__abc_44228_n22401), .Y(u2__abc_44228_n22402) );
  INVX1 INVX1_3942 ( .A(u2__abc_44228_n22409), .Y(u2__abc_44228_n22410) );
  INVX1 INVX1_3943 ( .A(u2__abc_44228_n22413), .Y(u2__abc_44228_n22414) );
  INVX1 INVX1_3944 ( .A(u2__abc_44228_n22421), .Y(u2__abc_44228_n22422) );
  INVX1 INVX1_3945 ( .A(u2__abc_44228_n22425), .Y(u2__abc_44228_n22426) );
  INVX1 INVX1_3946 ( .A(u2__abc_44228_n22433), .Y(u2__abc_44228_n22434) );
  INVX1 INVX1_3947 ( .A(u2__abc_44228_n22437), .Y(u2__abc_44228_n22438) );
  INVX1 INVX1_3948 ( .A(u2__abc_44228_n22445), .Y(u2__abc_44228_n22446) );
  INVX1 INVX1_3949 ( .A(u2__abc_44228_n22449), .Y(u2__abc_44228_n22450) );
  INVX1 INVX1_395 ( .A(u2_remHi_31_), .Y(u2__abc_44228_n3576) );
  INVX1 INVX1_3950 ( .A(u2__abc_44228_n22457), .Y(u2__abc_44228_n22458) );
  INVX1 INVX1_3951 ( .A(u2__abc_44228_n22461), .Y(u2__abc_44228_n22462) );
  INVX1 INVX1_3952 ( .A(u2__abc_44228_n22469), .Y(u2__abc_44228_n22470) );
  INVX1 INVX1_3953 ( .A(u2__abc_44228_n22473), .Y(u2__abc_44228_n22474) );
  INVX1 INVX1_3954 ( .A(u2__abc_44228_n22481), .Y(u2__abc_44228_n22482) );
  INVX1 INVX1_3955 ( .A(u2__abc_44228_n22485), .Y(u2__abc_44228_n22486) );
  INVX1 INVX1_3956 ( .A(u2__abc_44228_n22493), .Y(u2__abc_44228_n22494) );
  INVX1 INVX1_3957 ( .A(u2__abc_44228_n22497), .Y(u2__abc_44228_n22498) );
  INVX1 INVX1_3958 ( .A(u2__abc_44228_n22505), .Y(u2__abc_44228_n22506) );
  INVX1 INVX1_3959 ( .A(u2__abc_44228_n22509), .Y(u2__abc_44228_n22510) );
  INVX1 INVX1_396 ( .A(u2__abc_44228_n3577), .Y(u2__abc_44228_n3578) );
  INVX1 INVX1_3960 ( .A(u2__abc_44228_n22517), .Y(u2__abc_44228_n22518) );
  INVX1 INVX1_3961 ( .A(u2__abc_44228_n22521), .Y(u2__abc_44228_n22522) );
  INVX1 INVX1_3962 ( .A(u2__abc_44228_n22529), .Y(u2__abc_44228_n22530) );
  INVX1 INVX1_3963 ( .A(u2__abc_44228_n22533), .Y(u2__abc_44228_n22534) );
  INVX1 INVX1_3964 ( .A(u2__abc_44228_n22541), .Y(u2__abc_44228_n22542) );
  INVX1 INVX1_3965 ( .A(u2__abc_44228_n22545), .Y(u2__abc_44228_n22546) );
  INVX1 INVX1_3966 ( .A(u2__abc_44228_n22553), .Y(u2__abc_44228_n22554) );
  INVX1 INVX1_3967 ( .A(u2__abc_44228_n22557), .Y(u2__abc_44228_n22558) );
  INVX1 INVX1_3968 ( .A(u2__abc_44228_n22565), .Y(u2__abc_44228_n22566) );
  INVX1 INVX1_3969 ( .A(u2__abc_44228_n22569), .Y(u2__abc_44228_n22570) );
  INVX1 INVX1_397 ( .A(u2__abc_44228_n3557), .Y(u2__abc_44228_n3589) );
  INVX1 INVX1_3970 ( .A(u2__abc_44228_n22577), .Y(u2__abc_44228_n22578) );
  INVX1 INVX1_3971 ( .A(u2__abc_44228_n22581), .Y(u2__abc_44228_n22582) );
  INVX1 INVX1_3972 ( .A(u2__abc_44228_n22589), .Y(u2__abc_44228_n22590) );
  INVX1 INVX1_3973 ( .A(u2__abc_44228_n22593), .Y(u2__abc_44228_n22594) );
  INVX1 INVX1_3974 ( .A(u2__abc_44228_n22601), .Y(u2__abc_44228_n22602) );
  INVX1 INVX1_3975 ( .A(u2__abc_44228_n22605), .Y(u2__abc_44228_n22606) );
  INVX1 INVX1_3976 ( .A(u2__abc_44228_n22613), .Y(u2__abc_44228_n22614) );
  INVX1 INVX1_3977 ( .A(u2__abc_44228_n22617), .Y(u2__abc_44228_n22618) );
  INVX1 INVX1_3978 ( .A(u2__abc_44228_n22625), .Y(u2__abc_44228_n22626) );
  INVX1 INVX1_3979 ( .A(u2__abc_44228_n22629), .Y(u2__abc_44228_n22630) );
  INVX1 INVX1_398 ( .A(u2__abc_44228_n3562_1), .Y(u2__abc_44228_n3590) );
  INVX1 INVX1_3980 ( .A(u2__abc_44228_n22637), .Y(u2__abc_44228_n22638) );
  INVX1 INVX1_3981 ( .A(u2__abc_44228_n22641), .Y(u2__abc_44228_n22642) );
  INVX1 INVX1_3982 ( .A(u2__abc_44228_n22649), .Y(u2__abc_44228_n22650) );
  INVX1 INVX1_3983 ( .A(u2__abc_44228_n22653), .Y(u2__abc_44228_n22654) );
  INVX1 INVX1_3984 ( .A(u2__abc_44228_n22661), .Y(u2__abc_44228_n22662) );
  INVX1 INVX1_3985 ( .A(u2__abc_44228_n22665), .Y(u2__abc_44228_n22666) );
  INVX1 INVX1_3986 ( .A(u2__abc_44228_n22673), .Y(u2__abc_44228_n22674) );
  INVX1 INVX1_3987 ( .A(u2__abc_44228_n22677), .Y(u2__abc_44228_n22678) );
  INVX1 INVX1_3988 ( .A(u2__abc_44228_n22685), .Y(u2__abc_44228_n22686) );
  INVX1 INVX1_3989 ( .A(u2__abc_44228_n22689), .Y(u2__abc_44228_n22690) );
  INVX1 INVX1_399 ( .A(u2__abc_44228_n3542), .Y(u2__abc_44228_n3595) );
  INVX1 INVX1_3990 ( .A(u2__abc_44228_n22697), .Y(u2__abc_44228_n22698) );
  INVX1 INVX1_3991 ( .A(u2__abc_44228_n22701), .Y(u2__abc_44228_n22702) );
  INVX1 INVX1_3992 ( .A(u2__abc_44228_n22709), .Y(u2__abc_44228_n22710) );
  INVX1 INVX1_3993 ( .A(u2__abc_44228_n22713), .Y(u2__abc_44228_n22714) );
  INVX1 INVX1_3994 ( .A(u2__abc_44228_n22721), .Y(u2__abc_44228_n22722) );
  INVX1 INVX1_3995 ( .A(u2__abc_44228_n22725), .Y(u2__abc_44228_n22726) );
  INVX1 INVX1_3996 ( .A(u2__abc_44228_n22733), .Y(u2__abc_44228_n22734) );
  INVX1 INVX1_3997 ( .A(u2__abc_44228_n22737), .Y(u2__abc_44228_n22738) );
  INVX1 INVX1_3998 ( .A(u2__abc_44228_n22745), .Y(u2__abc_44228_n22746) );
  INVX1 INVX1_3999 ( .A(u2__abc_44228_n22749), .Y(u2__abc_44228_n22750) );
  INVX1 INVX1_4 ( .A(\a[114] ), .Y(_abc_64468_n1518) );
  INVX1 INVX1_40 ( .A(_abc_64468_n1644), .Y(_abc_64468_n1650) );
  INVX1 INVX1_400 ( .A(u2__abc_44228_n3596), .Y(u2__abc_44228_n3597_1) );
  INVX1 INVX1_4000 ( .A(u2__abc_44228_n22757), .Y(u2__abc_44228_n22758) );
  INVX1 INVX1_4001 ( .A(u2__abc_44228_n22761), .Y(u2__abc_44228_n22762) );
  INVX1 INVX1_4002 ( .A(u2__abc_44228_n22769), .Y(u2__abc_44228_n22770) );
  INVX1 INVX1_4003 ( .A(u2__abc_44228_n22773), .Y(u2__abc_44228_n22774) );
  INVX1 INVX1_4004 ( .A(u2__abc_44228_n22781), .Y(u2__abc_44228_n22782) );
  INVX1 INVX1_4005 ( .A(u2__abc_44228_n22785), .Y(u2__abc_44228_n22786) );
  INVX1 INVX1_4006 ( .A(u2__abc_44228_n22793), .Y(u2__abc_44228_n22794) );
  INVX1 INVX1_4007 ( .A(u2__abc_44228_n22797), .Y(u2__abc_44228_n22798) );
  INVX1 INVX1_4008 ( .A(u2__abc_44228_n22805), .Y(u2__abc_44228_n22806) );
  INVX1 INVX1_4009 ( .A(u2__abc_44228_n22809), .Y(u2__abc_44228_n22810) );
  INVX1 INVX1_401 ( .A(u2__abc_44228_n3519), .Y(u2__abc_44228_n3608_1) );
  INVX1 INVX1_4010 ( .A(u2__abc_44228_n22817), .Y(u2__abc_44228_n22818) );
  INVX1 INVX1_4011 ( .A(u2__abc_44228_n22821), .Y(u2__abc_44228_n22822) );
  INVX1 INVX1_4012 ( .A(u2__abc_44228_n22829), .Y(u2__abc_44228_n22830) );
  INVX1 INVX1_4013 ( .A(u2__abc_44228_n22833), .Y(u2__abc_44228_n22834) );
  INVX1 INVX1_4014 ( .A(u2__abc_44228_n22841), .Y(u2__abc_44228_n22842) );
  INVX1 INVX1_4015 ( .A(u2__abc_44228_n22845), .Y(u2__abc_44228_n22846) );
  INVX1 INVX1_4016 ( .A(u2__abc_44228_n22853), .Y(u2__abc_44228_n22854) );
  INVX1 INVX1_4017 ( .A(u2__abc_44228_n22857), .Y(u2__abc_44228_n22858) );
  INVX1 INVX1_4018 ( .A(u2__abc_44228_n22865), .Y(u2__abc_44228_n22866) );
  INVX1 INVX1_4019 ( .A(u2__abc_44228_n22869), .Y(u2__abc_44228_n22870) );
  INVX1 INVX1_402 ( .A(u2__abc_44228_n3609), .Y(u2__abc_44228_n3610) );
  INVX1 INVX1_4020 ( .A(u2__abc_44228_n22877), .Y(u2__abc_44228_n22878) );
  INVX1 INVX1_4021 ( .A(u2__abc_44228_n22881), .Y(u2__abc_44228_n22882) );
  INVX1 INVX1_4022 ( .A(u2__abc_44228_n22889), .Y(u2__abc_44228_n22890) );
  INVX1 INVX1_4023 ( .A(u2__abc_44228_n22893), .Y(u2__abc_44228_n22894) );
  INVX1 INVX1_4024 ( .A(u2__abc_44228_n22901), .Y(u2__abc_44228_n22902) );
  INVX1 INVX1_4025 ( .A(u2__abc_44228_n22905), .Y(u2__abc_44228_n22906) );
  INVX1 INVX1_4026 ( .A(u2__abc_44228_n22913), .Y(u2__abc_44228_n22914) );
  INVX1 INVX1_4027 ( .A(u2__abc_44228_n22917), .Y(u2__abc_44228_n22918) );
  INVX1 INVX1_4028 ( .A(u2__abc_44228_n22925), .Y(u2__abc_44228_n22926) );
  INVX1 INVX1_4029 ( .A(u2__abc_44228_n22929), .Y(u2__abc_44228_n22930) );
  INVX1 INVX1_403 ( .A(u2__abc_44228_n3483), .Y(u2__abc_44228_n3616) );
  INVX1 INVX1_4030 ( .A(u2__abc_44228_n22937), .Y(u2__abc_44228_n22938) );
  INVX1 INVX1_4031 ( .A(u2__abc_44228_n22941), .Y(u2__abc_44228_n22942) );
  INVX1 INVX1_4032 ( .A(u2__abc_44228_n22949), .Y(u2__abc_44228_n22950) );
  INVX1 INVX1_4033 ( .A(u2__abc_44228_n22953), .Y(u2__abc_44228_n22954) );
  INVX1 INVX1_4034 ( .A(u2__abc_44228_n22961), .Y(u2__abc_44228_n22962) );
  INVX1 INVX1_4035 ( .A(u2__abc_44228_n22965), .Y(u2__abc_44228_n22966) );
  INVX1 INVX1_4036 ( .A(u2__abc_44228_n22973), .Y(u2__abc_44228_n22974) );
  INVX1 INVX1_4037 ( .A(u2__abc_44228_n22977), .Y(u2__abc_44228_n22978) );
  INVX1 INVX1_4038 ( .A(u2__abc_44228_n22985), .Y(u2__abc_44228_n22986) );
  INVX1 INVX1_4039 ( .A(u2__abc_44228_n22989), .Y(u2__abc_44228_n22990) );
  INVX1 INVX1_404 ( .A(u2__abc_44228_n3617_1), .Y(u2__abc_44228_n3618) );
  INVX1 INVX1_4040 ( .A(u2__abc_44228_n22997), .Y(u2__abc_44228_n22998) );
  INVX1 INVX1_4041 ( .A(u2__abc_44228_n23001), .Y(u2__abc_44228_n23002) );
  INVX1 INVX1_4042 ( .A(u2__abc_44228_n23009), .Y(u2__abc_44228_n23010) );
  INVX1 INVX1_4043 ( .A(u2__abc_44228_n23013), .Y(u2__abc_44228_n23014) );
  INVX1 INVX1_4044 ( .A(u2__abc_44228_n23021), .Y(u2__abc_44228_n23022) );
  INVX1 INVX1_4045 ( .A(u2__abc_44228_n23025), .Y(u2__abc_44228_n23026) );
  INVX1 INVX1_4046 ( .A(u2__abc_44228_n23033), .Y(u2__abc_44228_n23034) );
  INVX1 INVX1_4047 ( .A(u2__abc_44228_n23037), .Y(u2__abc_44228_n23038) );
  INVX1 INVX1_4048 ( .A(u2__abc_44228_n23045), .Y(u2__abc_44228_n23046) );
  INVX1 INVX1_4049 ( .A(u2__abc_44228_n23049), .Y(u2__abc_44228_n23050) );
  INVX1 INVX1_405 ( .A(u2__abc_44228_n3423), .Y(u2__abc_44228_n3632) );
  INVX1 INVX1_4050 ( .A(u2__abc_44228_n23057), .Y(u2__abc_44228_n23058) );
  INVX1 INVX1_4051 ( .A(u2__abc_44228_n23061), .Y(u2__abc_44228_n23062) );
  INVX1 INVX1_4052 ( .A(u2__abc_44228_n23069), .Y(u2__abc_44228_n23070) );
  INVX1 INVX1_4053 ( .A(u2__abc_44228_n23073), .Y(u2__abc_44228_n23074) );
  INVX1 INVX1_4054 ( .A(u2__abc_44228_n23081), .Y(u2__abc_44228_n23082) );
  INVX1 INVX1_4055 ( .A(u2__abc_44228_n23085), .Y(u2__abc_44228_n23086) );
  INVX1 INVX1_4056 ( .A(u2__abc_44228_n23093), .Y(u2__abc_44228_n23094) );
  INVX1 INVX1_4057 ( .A(u2__abc_44228_n23097), .Y(u2__abc_44228_n23098) );
  INVX1 INVX1_4058 ( .A(u2__abc_44228_n23105), .Y(u2__abc_44228_n23106) );
  INVX1 INVX1_4059 ( .A(u2__abc_44228_n23109), .Y(u2__abc_44228_n23110) );
  INVX1 INVX1_406 ( .A(u2__abc_44228_n3633), .Y(u2__abc_44228_n3634) );
  INVX1 INVX1_4060 ( .A(u2__abc_44228_n23117), .Y(u2__abc_44228_n23118) );
  INVX1 INVX1_4061 ( .A(u2__abc_44228_n23121), .Y(u2__abc_44228_n23122) );
  INVX1 INVX1_4062 ( .A(u2__abc_44228_n23129), .Y(u2__abc_44228_n23130) );
  INVX1 INVX1_4063 ( .A(u2__abc_44228_n23133), .Y(u2__abc_44228_n23134) );
  INVX1 INVX1_4064 ( .A(u2__abc_44228_n23141), .Y(u2__abc_44228_n23142) );
  INVX1 INVX1_4065 ( .A(u2__abc_44228_n23145), .Y(u2__abc_44228_n23146) );
  INVX1 INVX1_4066 ( .A(u2__abc_44228_n23153), .Y(u2__abc_44228_n23154) );
  INVX1 INVX1_4067 ( .A(u2__abc_44228_n23157), .Y(u2__abc_44228_n23158) );
  INVX1 INVX1_4068 ( .A(u2__abc_44228_n23165), .Y(u2__abc_44228_n23166) );
  INVX1 INVX1_4069 ( .A(u2__abc_44228_n23169), .Y(u2__abc_44228_n23170) );
  INVX1 INVX1_407 ( .A(u2__abc_44228_n3400), .Y(u2__abc_44228_n3642) );
  INVX1 INVX1_408 ( .A(u2__abc_44228_n3644), .Y(u2__abc_44228_n3645) );
  INVX1 INVX1_409 ( .A(u2__abc_44228_n3386), .Y(u2__abc_44228_n3647_1) );
  INVX1 INVX1_41 ( .A(\a[124] ), .Y(_abc_64468_n1651) );
  INVX1 INVX1_410 ( .A(u2__abc_44228_n3648), .Y(u2__abc_44228_n3649) );
  INVX1 INVX1_411 ( .A(u2__abc_44228_n3364), .Y(u2__abc_44228_n3655) );
  INVX1 INVX1_412 ( .A(u2__abc_44228_n3656_1), .Y(u2__abc_44228_n3657) );
  INVX1 INVX1_413 ( .A(sqrto_125_), .Y(u2__abc_44228_n3665) );
  INVX1 INVX1_414 ( .A(u2__abc_44228_n3666_1), .Y(u2__abc_44228_n3667) );
  INVX1 INVX1_415 ( .A(u2_remHi_125_), .Y(u2__abc_44228_n3668) );
  INVX1 INVX1_416 ( .A(u2__abc_44228_n3669), .Y(u2__abc_44228_n3670) );
  INVX1 INVX1_417 ( .A(sqrto_124_), .Y(u2__abc_44228_n3672) );
  INVX1 INVX1_418 ( .A(u2_remHi_124_), .Y(u2__abc_44228_n3674) );
  INVX1 INVX1_419 ( .A(u2__abc_44228_n3676), .Y(u2__abc_44228_n3677) );
  INVX1 INVX1_42 ( .A(_abc_64468_n1654), .Y(_abc_64468_n1655) );
  INVX1 INVX1_420 ( .A(sqrto_122_), .Y(u2__abc_44228_n3679) );
  INVX1 INVX1_421 ( .A(u2_remHi_122_), .Y(u2__abc_44228_n3681) );
  INVX1 INVX1_422 ( .A(u2__abc_44228_n3683), .Y(u2__abc_44228_n3684) );
  INVX1 INVX1_423 ( .A(sqrto_123_), .Y(u2__abc_44228_n3685_1) );
  INVX1 INVX1_424 ( .A(u2__abc_44228_n3686), .Y(u2__abc_44228_n3687) );
  INVX1 INVX1_425 ( .A(u2_remHi_123_), .Y(u2__abc_44228_n3688) );
  INVX1 INVX1_426 ( .A(u2__abc_44228_n3689), .Y(u2__abc_44228_n3690) );
  INVX1 INVX1_427 ( .A(sqrto_119_), .Y(u2__abc_44228_n3694_1) );
  INVX1 INVX1_428 ( .A(u2__abc_44228_n3695), .Y(u2__abc_44228_n3696) );
  INVX1 INVX1_429 ( .A(u2_remHi_119_), .Y(u2__abc_44228_n3697) );
  INVX1 INVX1_43 ( .A(_abc_64468_n1656), .Y(_abc_64468_n1657) );
  INVX1 INVX1_430 ( .A(u2__abc_44228_n3698), .Y(u2__abc_44228_n3699) );
  INVX1 INVX1_431 ( .A(sqrto_118_), .Y(u2__abc_44228_n3701) );
  INVX1 INVX1_432 ( .A(u2_remHi_118_), .Y(u2__abc_44228_n3703) );
  INVX1 INVX1_433 ( .A(u2__abc_44228_n3705), .Y(u2__abc_44228_n3706) );
  INVX1 INVX1_434 ( .A(sqrto_121_), .Y(u2__abc_44228_n3708) );
  INVX1 INVX1_435 ( .A(u2__abc_44228_n3709), .Y(u2__abc_44228_n3710) );
  INVX1 INVX1_436 ( .A(u2_remHi_121_), .Y(u2__abc_44228_n3711) );
  INVX1 INVX1_437 ( .A(u2__abc_44228_n3712), .Y(u2__abc_44228_n3713) );
  INVX1 INVX1_438 ( .A(sqrto_120_), .Y(u2__abc_44228_n3715) );
  INVX1 INVX1_439 ( .A(u2_remHi_120_), .Y(u2__abc_44228_n3717) );
  INVX1 INVX1_44 ( .A(_abc_64468_n1659), .Y(_abc_64468_n1663) );
  INVX1 INVX1_440 ( .A(u2__abc_44228_n3719), .Y(u2__abc_44228_n3720) );
  INVX1 INVX1_441 ( .A(sqrto_117_), .Y(u2__abc_44228_n3724) );
  INVX1 INVX1_442 ( .A(u2__abc_44228_n3725), .Y(u2__abc_44228_n3726) );
  INVX1 INVX1_443 ( .A(u2_remHi_117_), .Y(u2__abc_44228_n3727) );
  INVX1 INVX1_444 ( .A(u2__abc_44228_n3728), .Y(u2__abc_44228_n3729) );
  INVX1 INVX1_445 ( .A(sqrto_116_), .Y(u2__abc_44228_n3731) );
  INVX1 INVX1_446 ( .A(u2_remHi_116_), .Y(u2__abc_44228_n3733) );
  INVX1 INVX1_447 ( .A(u2__abc_44228_n3735), .Y(u2__abc_44228_n3736) );
  INVX1 INVX1_448 ( .A(sqrto_115_), .Y(u2__abc_44228_n3738) );
  INVX1 INVX1_449 ( .A(u2__abc_44228_n3739), .Y(u2__abc_44228_n3740_1) );
  INVX1 INVX1_45 ( .A(\a[125] ), .Y(_abc_64468_n1664) );
  INVX1 INVX1_450 ( .A(u2_remHi_115_), .Y(u2__abc_44228_n3741) );
  INVX1 INVX1_451 ( .A(u2__abc_44228_n3742), .Y(u2__abc_44228_n3743) );
  INVX1 INVX1_452 ( .A(sqrto_114_), .Y(u2__abc_44228_n3745) );
  INVX1 INVX1_453 ( .A(u2_remHi_114_), .Y(u2__abc_44228_n3747) );
  INVX1 INVX1_454 ( .A(u2__abc_44228_n3749), .Y(u2__abc_44228_n3750_1) );
  INVX1 INVX1_455 ( .A(sqrto_113_), .Y(u2__abc_44228_n3753) );
  INVX1 INVX1_456 ( .A(u2__abc_44228_n3754), .Y(u2__abc_44228_n3755) );
  INVX1 INVX1_457 ( .A(u2_remHi_113_), .Y(u2__abc_44228_n3756) );
  INVX1 INVX1_458 ( .A(u2__abc_44228_n3757), .Y(u2__abc_44228_n3758) );
  INVX1 INVX1_459 ( .A(sqrto_112_), .Y(u2__abc_44228_n3760) );
  INVX1 INVX1_46 ( .A(_abc_64468_n1667), .Y(_abc_64468_n1668) );
  INVX1 INVX1_460 ( .A(u2_remHi_112_), .Y(u2__abc_44228_n3762) );
  INVX1 INVX1_461 ( .A(u2__abc_44228_n3764), .Y(u2__abc_44228_n3765) );
  INVX1 INVX1_462 ( .A(sqrto_110_), .Y(u2__abc_44228_n3767) );
  INVX1 INVX1_463 ( .A(u2_remHi_110_), .Y(u2__abc_44228_n3769) );
  INVX1 INVX1_464 ( .A(u2__abc_44228_n3771), .Y(u2__abc_44228_n3772) );
  INVX1 INVX1_465 ( .A(sqrto_111_), .Y(u2__abc_44228_n3773) );
  INVX1 INVX1_466 ( .A(u2__abc_44228_n3774), .Y(u2__abc_44228_n3775) );
  INVX1 INVX1_467 ( .A(u2_remHi_111_), .Y(u2__abc_44228_n3776) );
  INVX1 INVX1_468 ( .A(u2__abc_44228_n3777), .Y(u2__abc_44228_n3778) );
  INVX1 INVX1_469 ( .A(sqrto_109_), .Y(u2__abc_44228_n3784) );
  INVX1 INVX1_47 ( .A(_abc_64468_n1669), .Y(_abc_64468_n1670) );
  INVX1 INVX1_470 ( .A(u2__abc_44228_n3785), .Y(u2__abc_44228_n3786) );
  INVX1 INVX1_471 ( .A(u2_remHi_109_), .Y(u2__abc_44228_n3787) );
  INVX1 INVX1_472 ( .A(u2__abc_44228_n3788), .Y(u2__abc_44228_n3789_1) );
  INVX1 INVX1_473 ( .A(sqrto_108_), .Y(u2__abc_44228_n3791) );
  INVX1 INVX1_474 ( .A(u2_remHi_108_), .Y(u2__abc_44228_n3793) );
  INVX1 INVX1_475 ( .A(u2__abc_44228_n3795), .Y(u2__abc_44228_n3796) );
  INVX1 INVX1_476 ( .A(sqrto_106_), .Y(u2__abc_44228_n3798_1) );
  INVX1 INVX1_477 ( .A(u2_remHi_106_), .Y(u2__abc_44228_n3800) );
  INVX1 INVX1_478 ( .A(u2__abc_44228_n3802), .Y(u2__abc_44228_n3803) );
  INVX1 INVX1_479 ( .A(sqrto_107_), .Y(u2__abc_44228_n3804) );
  INVX1 INVX1_48 ( .A(\a[126] ), .Y(_abc_64468_n1678) );
  INVX1 INVX1_480 ( .A(u2__abc_44228_n3805), .Y(u2__abc_44228_n3806) );
  INVX1 INVX1_481 ( .A(u2_remHi_107_), .Y(u2__abc_44228_n3807_1) );
  INVX1 INVX1_482 ( .A(u2__abc_44228_n3808), .Y(u2__abc_44228_n3809) );
  INVX1 INVX1_483 ( .A(sqrto_103_), .Y(u2__abc_44228_n3813) );
  INVX1 INVX1_484 ( .A(u2__abc_44228_n3814), .Y(u2__abc_44228_n3815) );
  INVX1 INVX1_485 ( .A(u2_remHi_103_), .Y(u2__abc_44228_n3816_1) );
  INVX1 INVX1_486 ( .A(u2__abc_44228_n3817), .Y(u2__abc_44228_n3818) );
  INVX1 INVX1_487 ( .A(sqrto_102_), .Y(u2__abc_44228_n3820) );
  INVX1 INVX1_488 ( .A(u2_remHi_102_), .Y(u2__abc_44228_n3822) );
  INVX1 INVX1_489 ( .A(u2__abc_44228_n3824), .Y(u2__abc_44228_n3825_1) );
  INVX1 INVX1_49 ( .A(_abc_64468_n1681), .Y(_abc_64468_n1682) );
  INVX1 INVX1_490 ( .A(sqrto_105_), .Y(u2__abc_44228_n3827) );
  INVX1 INVX1_491 ( .A(u2__abc_44228_n3828), .Y(u2__abc_44228_n3829) );
  INVX1 INVX1_492 ( .A(u2_remHi_105_), .Y(u2__abc_44228_n3830) );
  INVX1 INVX1_493 ( .A(u2__abc_44228_n3831), .Y(u2__abc_44228_n3832) );
  INVX1 INVX1_494 ( .A(sqrto_104_), .Y(u2__abc_44228_n3834) );
  INVX1 INVX1_495 ( .A(u2_remHi_104_), .Y(u2__abc_44228_n3836) );
  INVX1 INVX1_496 ( .A(u2__abc_44228_n3838), .Y(u2__abc_44228_n3839) );
  INVX1 INVX1_497 ( .A(sqrto_101_), .Y(u2__abc_44228_n3843) );
  INVX1 INVX1_498 ( .A(u2__abc_44228_n3844_1), .Y(u2__abc_44228_n3845) );
  INVX1 INVX1_499 ( .A(u2_remHi_101_), .Y(u2__abc_44228_n3846) );
  INVX1 INVX1_5 ( .A(\a[115] ), .Y(_abc_64468_n1525) );
  INVX1 INVX1_50 ( .A(_abc_64468_n1685), .Y(_abc_64468_n1686) );
  INVX1 INVX1_500 ( .A(u2__abc_44228_n3847), .Y(u2__abc_44228_n3848) );
  INVX1 INVX1_501 ( .A(sqrto_100_), .Y(u2__abc_44228_n3850) );
  INVX1 INVX1_502 ( .A(u2_remHi_100_), .Y(u2__abc_44228_n3852) );
  INVX1 INVX1_503 ( .A(u2__abc_44228_n3854_1), .Y(u2__abc_44228_n3855) );
  INVX1 INVX1_504 ( .A(sqrto_98_), .Y(u2__abc_44228_n3857) );
  INVX1 INVX1_505 ( .A(u2_remHi_98_), .Y(u2__abc_44228_n3859) );
  INVX1 INVX1_506 ( .A(u2__abc_44228_n3861), .Y(u2__abc_44228_n3862) );
  INVX1 INVX1_507 ( .A(sqrto_99_), .Y(u2__abc_44228_n3863) );
  INVX1 INVX1_508 ( .A(u2__abc_44228_n3864_1), .Y(u2__abc_44228_n3865) );
  INVX1 INVX1_509 ( .A(u2_remHi_99_), .Y(u2__abc_44228_n3866) );
  INVX1 INVX1_51 ( .A(_abc_64468_n1684), .Y(_abc_64468_n1692) );
  INVX1 INVX1_510 ( .A(u2__abc_44228_n3867), .Y(u2__abc_44228_n3868) );
  INVX1 INVX1_511 ( .A(sqrto_97_), .Y(u2__abc_44228_n3872) );
  INVX1 INVX1_512 ( .A(u2__abc_44228_n3873_1), .Y(u2__abc_44228_n3874) );
  INVX1 INVX1_513 ( .A(u2_remHi_97_), .Y(u2__abc_44228_n3875) );
  INVX1 INVX1_514 ( .A(u2__abc_44228_n3876), .Y(u2__abc_44228_n3877) );
  INVX1 INVX1_515 ( .A(sqrto_96_), .Y(u2__abc_44228_n3879) );
  INVX1 INVX1_516 ( .A(u2_remHi_96_), .Y(u2__abc_44228_n3881) );
  INVX1 INVX1_517 ( .A(u2__abc_44228_n3883), .Y(u2__abc_44228_n3884) );
  INVX1 INVX1_518 ( .A(sqrto_94_), .Y(u2__abc_44228_n3886) );
  INVX1 INVX1_519 ( .A(u2_remHi_94_), .Y(u2__abc_44228_n3888) );
  INVX1 INVX1_52 ( .A(\a[78] ), .Y(u1__abc_43968_n166) );
  INVX1 INVX1_520 ( .A(u2__abc_44228_n3890), .Y(u2__abc_44228_n3891) );
  INVX1 INVX1_521 ( .A(sqrto_95_), .Y(u2__abc_44228_n3892) );
  INVX1 INVX1_522 ( .A(u2__abc_44228_n3893_1), .Y(u2__abc_44228_n3894) );
  INVX1 INVX1_523 ( .A(u2_remHi_95_), .Y(u2__abc_44228_n3895) );
  INVX1 INVX1_524 ( .A(u2__abc_44228_n3896), .Y(u2__abc_44228_n3897) );
  INVX1 INVX1_525 ( .A(sqrto_93_), .Y(u2__abc_44228_n3904) );
  INVX1 INVX1_526 ( .A(u2__abc_44228_n3905), .Y(u2__abc_44228_n3906) );
  INVX1 INVX1_527 ( .A(u2_remHi_93_), .Y(u2__abc_44228_n3907) );
  INVX1 INVX1_528 ( .A(u2__abc_44228_n3908), .Y(u2__abc_44228_n3909) );
  INVX1 INVX1_529 ( .A(sqrto_92_), .Y(u2__abc_44228_n3911) );
  INVX1 INVX1_53 ( .A(\a[79] ), .Y(u1__abc_43968_n167) );
  INVX1 INVX1_530 ( .A(u2_remHi_92_), .Y(u2__abc_44228_n3913) );
  INVX1 INVX1_531 ( .A(u2__abc_44228_n3915), .Y(u2__abc_44228_n3916) );
  INVX1 INVX1_532 ( .A(sqrto_90_), .Y(u2__abc_44228_n3918) );
  INVX1 INVX1_533 ( .A(u2_remHi_90_), .Y(u2__abc_44228_n3920) );
  INVX1 INVX1_534 ( .A(u2__abc_44228_n3922), .Y(u2__abc_44228_n3923) );
  INVX1 INVX1_535 ( .A(sqrto_91_), .Y(u2__abc_44228_n3924) );
  INVX1 INVX1_536 ( .A(u2__abc_44228_n3925), .Y(u2__abc_44228_n3926) );
  INVX1 INVX1_537 ( .A(u2_remHi_91_), .Y(u2__abc_44228_n3927) );
  INVX1 INVX1_538 ( .A(u2__abc_44228_n3928), .Y(u2__abc_44228_n3929) );
  INVX1 INVX1_539 ( .A(sqrto_89_), .Y(u2__abc_44228_n3933) );
  INVX1 INVX1_54 ( .A(\a[76] ), .Y(u1__abc_43968_n169) );
  INVX1 INVX1_540 ( .A(u2__abc_44228_n3934), .Y(u2__abc_44228_n3935) );
  INVX1 INVX1_541 ( .A(u2_remHi_89_), .Y(u2__abc_44228_n3936) );
  INVX1 INVX1_542 ( .A(u2__abc_44228_n3937), .Y(u2__abc_44228_n3938) );
  INVX1 INVX1_543 ( .A(sqrto_88_), .Y(u2__abc_44228_n3940_1) );
  INVX1 INVX1_544 ( .A(u2_remHi_88_), .Y(u2__abc_44228_n3942) );
  INVX1 INVX1_545 ( .A(u2__abc_44228_n3944), .Y(u2__abc_44228_n3945) );
  INVX1 INVX1_546 ( .A(sqrto_86_), .Y(u2__abc_44228_n3947) );
  INVX1 INVX1_547 ( .A(u2_remHi_86_), .Y(u2__abc_44228_n3949_1) );
  INVX1 INVX1_548 ( .A(u2__abc_44228_n3951), .Y(u2__abc_44228_n3952) );
  INVX1 INVX1_549 ( .A(sqrto_87_), .Y(u2__abc_44228_n3953) );
  INVX1 INVX1_55 ( .A(\a[77] ), .Y(u1__abc_43968_n170_1) );
  INVX1 INVX1_550 ( .A(u2__abc_44228_n3954), .Y(u2__abc_44228_n3955) );
  INVX1 INVX1_551 ( .A(u2_remHi_87_), .Y(u2__abc_44228_n3956) );
  INVX1 INVX1_552 ( .A(u2__abc_44228_n3957), .Y(u2__abc_44228_n3958_1) );
  INVX1 INVX1_553 ( .A(sqrto_85_), .Y(u2__abc_44228_n3963) );
  INVX1 INVX1_554 ( .A(u2__abc_44228_n3964), .Y(u2__abc_44228_n3965) );
  INVX1 INVX1_555 ( .A(u2_remHi_85_), .Y(u2__abc_44228_n3966) );
  INVX1 INVX1_556 ( .A(u2__abc_44228_n3967_1), .Y(u2__abc_44228_n3968) );
  INVX1 INVX1_557 ( .A(sqrto_84_), .Y(u2__abc_44228_n3970) );
  INVX1 INVX1_558 ( .A(u2_remHi_84_), .Y(u2__abc_44228_n3972) );
  INVX1 INVX1_559 ( .A(u2__abc_44228_n3974), .Y(u2__abc_44228_n3975) );
  INVX1 INVX1_56 ( .A(\a[74] ), .Y(u1__abc_43968_n173_1) );
  INVX1 INVX1_560 ( .A(sqrto_82_), .Y(u2__abc_44228_n3977) );
  INVX1 INVX1_561 ( .A(u2_remHi_82_), .Y(u2__abc_44228_n3979) );
  INVX1 INVX1_562 ( .A(u2__abc_44228_n3981), .Y(u2__abc_44228_n3982) );
  INVX1 INVX1_563 ( .A(sqrto_83_), .Y(u2__abc_44228_n3983) );
  INVX1 INVX1_564 ( .A(u2__abc_44228_n3984), .Y(u2__abc_44228_n3985) );
  INVX1 INVX1_565 ( .A(u2_remHi_83_), .Y(u2__abc_44228_n3986_1) );
  INVX1 INVX1_566 ( .A(u2__abc_44228_n3987), .Y(u2__abc_44228_n3988) );
  INVX1 INVX1_567 ( .A(sqrto_81_), .Y(u2__abc_44228_n3992) );
  INVX1 INVX1_568 ( .A(u2__abc_44228_n3993), .Y(u2__abc_44228_n3994) );
  INVX1 INVX1_569 ( .A(u2_remHi_81_), .Y(u2__abc_44228_n3995_1) );
  INVX1 INVX1_57 ( .A(\a[75] ), .Y(u1__abc_43968_n174_1) );
  INVX1 INVX1_570 ( .A(u2__abc_44228_n3996), .Y(u2__abc_44228_n3997) );
  INVX1 INVX1_571 ( .A(sqrto_80_), .Y(u2__abc_44228_n3999) );
  INVX1 INVX1_572 ( .A(u2_remHi_80_), .Y(u2__abc_44228_n4001) );
  INVX1 INVX1_573 ( .A(u2__abc_44228_n4003), .Y(u2__abc_44228_n4004) );
  INVX1 INVX1_574 ( .A(sqrto_78_), .Y(u2__abc_44228_n4006) );
  INVX1 INVX1_575 ( .A(u2_remHi_78_), .Y(u2__abc_44228_n4008) );
  INVX1 INVX1_576 ( .A(u2__abc_44228_n4010), .Y(u2__abc_44228_n4011) );
  INVX1 INVX1_577 ( .A(sqrto_79_), .Y(u2__abc_44228_n4012) );
  INVX1 INVX1_578 ( .A(u2__abc_44228_n4013), .Y(u2__abc_44228_n4014) );
  INVX1 INVX1_579 ( .A(u2_remHi_79_), .Y(u2__abc_44228_n4015_1) );
  INVX1 INVX1_58 ( .A(\a[72] ), .Y(u1__abc_43968_n176) );
  INVX1 INVX1_580 ( .A(u2__abc_44228_n4016), .Y(u2__abc_44228_n4017) );
  INVX1 INVX1_581 ( .A(sqrto_77_), .Y(u2__abc_44228_n4023) );
  INVX1 INVX1_582 ( .A(u2__abc_44228_n4024_1), .Y(u2__abc_44228_n4025) );
  INVX1 INVX1_583 ( .A(u2_remHi_77_), .Y(u2__abc_44228_n4026) );
  INVX1 INVX1_584 ( .A(u2__abc_44228_n4027), .Y(u2__abc_44228_n4028) );
  INVX1 INVX1_585 ( .A(sqrto_76_), .Y(u2__abc_44228_n4030) );
  INVX1 INVX1_586 ( .A(u2_remHi_76_), .Y(u2__abc_44228_n4032) );
  INVX1 INVX1_587 ( .A(u2__abc_44228_n4034), .Y(u2__abc_44228_n4035) );
  INVX1 INVX1_588 ( .A(sqrto_74_), .Y(u2__abc_44228_n4037) );
  INVX1 INVX1_589 ( .A(u2_remHi_74_), .Y(u2__abc_44228_n4039) );
  INVX1 INVX1_59 ( .A(\a[73] ), .Y(u1__abc_43968_n177_1) );
  INVX1 INVX1_590 ( .A(u2__abc_44228_n4041_1), .Y(u2__abc_44228_n4042) );
  INVX1 INVX1_591 ( .A(sqrto_75_), .Y(u2__abc_44228_n4043) );
  INVX1 INVX1_592 ( .A(u2__abc_44228_n4044), .Y(u2__abc_44228_n4045) );
  INVX1 INVX1_593 ( .A(u2_remHi_75_), .Y(u2__abc_44228_n4046) );
  INVX1 INVX1_594 ( .A(u2__abc_44228_n4047), .Y(u2__abc_44228_n4048) );
  INVX1 INVX1_595 ( .A(sqrto_71_), .Y(u2__abc_44228_n4052) );
  INVX1 INVX1_596 ( .A(u2__abc_44228_n4053), .Y(u2__abc_44228_n4054) );
  INVX1 INVX1_597 ( .A(u2_remHi_71_), .Y(u2__abc_44228_n4055) );
  INVX1 INVX1_598 ( .A(u2__abc_44228_n4056), .Y(u2__abc_44228_n4057) );
  INVX1 INVX1_599 ( .A(sqrto_70_), .Y(u2__abc_44228_n4059) );
  INVX1 INVX1_6 ( .A(_abc_64468_n1528), .Y(_abc_64468_n1529) );
  INVX1 INVX1_60 ( .A(\a[70] ), .Y(u1__abc_43968_n181_1) );
  INVX1 INVX1_600 ( .A(u2_remHi_70_), .Y(u2__abc_44228_n4061_1) );
  INVX1 INVX1_601 ( .A(u2__abc_44228_n4063), .Y(u2__abc_44228_n4064) );
  INVX1 INVX1_602 ( .A(sqrto_73_), .Y(u2__abc_44228_n4066) );
  INVX1 INVX1_603 ( .A(u2__abc_44228_n4067), .Y(u2__abc_44228_n4068) );
  INVX1 INVX1_604 ( .A(u2_remHi_73_), .Y(u2__abc_44228_n4069) );
  INVX1 INVX1_605 ( .A(u2__abc_44228_n4070_1), .Y(u2__abc_44228_n4071) );
  INVX1 INVX1_606 ( .A(sqrto_72_), .Y(u2__abc_44228_n4073) );
  INVX1 INVX1_607 ( .A(u2_remHi_72_), .Y(u2__abc_44228_n4075) );
  INVX1 INVX1_608 ( .A(u2__abc_44228_n4077), .Y(u2__abc_44228_n4078) );
  INVX1 INVX1_609 ( .A(sqrto_69_), .Y(u2__abc_44228_n4082) );
  INVX1 INVX1_61 ( .A(\a[71] ), .Y(u1__abc_43968_n182) );
  INVX1 INVX1_610 ( .A(u2__abc_44228_n4083), .Y(u2__abc_44228_n4084) );
  INVX1 INVX1_611 ( .A(u2_remHi_69_), .Y(u2__abc_44228_n4085) );
  INVX1 INVX1_612 ( .A(u2__abc_44228_n4086), .Y(u2__abc_44228_n4087) );
  INVX1 INVX1_613 ( .A(sqrto_68_), .Y(u2__abc_44228_n4089) );
  INVX1 INVX1_614 ( .A(u2_remHi_68_), .Y(u2__abc_44228_n4091) );
  INVX1 INVX1_615 ( .A(u2__abc_44228_n4093), .Y(u2__abc_44228_n4094) );
  INVX1 INVX1_616 ( .A(sqrto_67_), .Y(u2__abc_44228_n4096) );
  INVX1 INVX1_617 ( .A(u2__abc_44228_n4097), .Y(u2__abc_44228_n4098) );
  INVX1 INVX1_618 ( .A(u2_remHi_67_), .Y(u2__abc_44228_n4099) );
  INVX1 INVX1_619 ( .A(u2__abc_44228_n4100_1), .Y(u2__abc_44228_n4101) );
  INVX1 INVX1_62 ( .A(\a[68] ), .Y(u1__abc_43968_n184) );
  INVX1 INVX1_620 ( .A(sqrto_66_), .Y(u2__abc_44228_n4103) );
  INVX1 INVX1_621 ( .A(u2_remHi_66_), .Y(u2__abc_44228_n4105) );
  INVX1 INVX1_622 ( .A(u2__abc_44228_n4107), .Y(u2__abc_44228_n4108) );
  INVX1 INVX1_623 ( .A(u2_remHi_65_), .Y(u2__abc_44228_n4111) );
  INVX1 INVX1_624 ( .A(sqrto_65_), .Y(u2__abc_44228_n4113) );
  INVX1 INVX1_625 ( .A(u2_remHi_64_), .Y(u2__abc_44228_n4116) );
  INVX1 INVX1_626 ( .A(sqrto_64_), .Y(u2__abc_44228_n4118) );
  INVX1 INVX1_627 ( .A(sqrto_63_), .Y(u2__abc_44228_n4122) );
  INVX1 INVX1_628 ( .A(u2__abc_44228_n4123), .Y(u2__abc_44228_n4124) );
  INVX1 INVX1_629 ( .A(u2_remHi_63_), .Y(u2__abc_44228_n4125) );
  INVX1 INVX1_63 ( .A(\a[69] ), .Y(u1__abc_43968_n185_1) );
  INVX1 INVX1_630 ( .A(u2__abc_44228_n4126), .Y(u2__abc_44228_n4127) );
  INVX1 INVX1_631 ( .A(sqrto_62_), .Y(u2__abc_44228_n4129) );
  INVX1 INVX1_632 ( .A(u2_remHi_62_), .Y(u2__abc_44228_n4131) );
  INVX1 INVX1_633 ( .A(u2__abc_44228_n4133), .Y(u2__abc_44228_n4134) );
  INVX1 INVX1_634 ( .A(u2__abc_44228_n4112), .Y(u2__abc_44228_n4145) );
  INVX1 INVX1_635 ( .A(u2__abc_44228_n4117), .Y(u2__abc_44228_n4146) );
  INVX1 INVX1_636 ( .A(u2__abc_44228_n4074), .Y(u2__abc_44228_n4162) );
  INVX1 INVX1_637 ( .A(u2__abc_44228_n4163), .Y(u2__abc_44228_n4164) );
  INVX1 INVX1_638 ( .A(u2__abc_44228_n4038), .Y(u2__abc_44228_n4169) );
  INVX1 INVX1_639 ( .A(u2__abc_44228_n4170), .Y(u2__abc_44228_n4171) );
  INVX1 INVX1_64 ( .A(\a[66] ), .Y(u1__abc_43968_n188_1) );
  INVX1 INVX1_640 ( .A(u2__abc_44228_n4007), .Y(u2__abc_44228_n4179) );
  INVX1 INVX1_641 ( .A(u2__abc_44228_n4180), .Y(u2__abc_44228_n4181) );
  INVX1 INVX1_642 ( .A(u2__abc_44228_n3978), .Y(u2__abc_44228_n4188) );
  INVX1 INVX1_643 ( .A(u2__abc_44228_n4190), .Y(u2__abc_44228_n4191) );
  INVX1 INVX1_644 ( .A(u2__abc_44228_n3948), .Y(u2__abc_44228_n4198) );
  INVX1 INVX1_645 ( .A(u2__abc_44228_n4199), .Y(u2__abc_44228_n4200) );
  INVX1 INVX1_646 ( .A(u2__abc_44228_n3919), .Y(u2__abc_44228_n4207) );
  INVX1 INVX1_647 ( .A(u2__abc_44228_n4208), .Y(u2__abc_44228_n4209) );
  INVX1 INVX1_648 ( .A(u2__abc_44228_n3887), .Y(u2__abc_44228_n4219) );
  INVX1 INVX1_649 ( .A(u2__abc_44228_n4220), .Y(u2__abc_44228_n4221) );
  INVX1 INVX1_65 ( .A(\a[67] ), .Y(u1__abc_43968_n189_1) );
  INVX1 INVX1_650 ( .A(u2__abc_44228_n3858), .Y(u2__abc_44228_n4228) );
  INVX1 INVX1_651 ( .A(u2__abc_44228_n4230), .Y(u2__abc_44228_n4231) );
  INVX1 INVX1_652 ( .A(u2__abc_44228_n3821), .Y(u2__abc_44228_n4238) );
  INVX1 INVX1_653 ( .A(u2__abc_44228_n4240), .Y(u2__abc_44228_n4241) );
  INVX1 INVX1_654 ( .A(u2__abc_44228_n3835_1), .Y(u2__abc_44228_n4243_1) );
  INVX1 INVX1_655 ( .A(u2__abc_44228_n4244), .Y(u2__abc_44228_n4245) );
  INVX1 INVX1_656 ( .A(u2__abc_44228_n3799), .Y(u2__abc_44228_n4249) );
  INVX1 INVX1_657 ( .A(u2__abc_44228_n4250), .Y(u2__abc_44228_n4251) );
  INVX1 INVX1_658 ( .A(u2__abc_44228_n3702), .Y(u2__abc_44228_n4260) );
  INVX1 INVX1_659 ( .A(u2__abc_44228_n4262_1), .Y(u2__abc_44228_n4263) );
  INVX1 INVX1_66 ( .A(\a[64] ), .Y(u1__abc_43968_n191) );
  INVX1 INVX1_660 ( .A(u2__abc_44228_n3680), .Y(u2__abc_44228_n4269) );
  INVX1 INVX1_661 ( .A(u2__abc_44228_n4270), .Y(u2__abc_44228_n4271) );
  INVX1 INVX1_662 ( .A(u2__abc_44228_n3768_1), .Y(u2__abc_44228_n4278) );
  INVX1 INVX1_663 ( .A(u2__abc_44228_n4279), .Y(u2__abc_44228_n4280) );
  INVX1 INVX1_664 ( .A(u2__abc_44228_n3746), .Y(u2__abc_44228_n4287) );
  INVX1 INVX1_665 ( .A(u2__abc_44228_n4289), .Y(u2__abc_44228_n4290) );
  INVX1 INVX1_666 ( .A(u2_o_253_), .Y(u2__abc_44228_n4301) );
  INVX1 INVX1_667 ( .A(u2__abc_44228_n4302), .Y(u2__abc_44228_n4303) );
  INVX1 INVX1_668 ( .A(u2_remHi_253_), .Y(u2__abc_44228_n4304) );
  INVX1 INVX1_669 ( .A(u2__abc_44228_n4305), .Y(u2__abc_44228_n4306) );
  INVX1 INVX1_67 ( .A(\a[65] ), .Y(u1__abc_43968_n192_1) );
  INVX1 INVX1_670 ( .A(u2_o_252_), .Y(u2__abc_44228_n4308) );
  INVX1 INVX1_671 ( .A(u2_remHi_252_), .Y(u2__abc_44228_n4310_1) );
  INVX1 INVX1_672 ( .A(u2__abc_44228_n4312), .Y(u2__abc_44228_n4313) );
  INVX1 INVX1_673 ( .A(u2_o_250_), .Y(u2__abc_44228_n4315) );
  INVX1 INVX1_674 ( .A(u2_remHi_250_), .Y(u2__abc_44228_n4317) );
  INVX1 INVX1_675 ( .A(u2__abc_44228_n4319), .Y(u2__abc_44228_n4320_1) );
  INVX1 INVX1_676 ( .A(u2_o_251_), .Y(u2__abc_44228_n4321) );
  INVX1 INVX1_677 ( .A(u2__abc_44228_n4322), .Y(u2__abc_44228_n4323) );
  INVX1 INVX1_678 ( .A(u2_remHi_251_), .Y(u2__abc_44228_n4324) );
  INVX1 INVX1_679 ( .A(u2__abc_44228_n4325), .Y(u2__abc_44228_n4326) );
  INVX1 INVX1_68 ( .A(\a[62] ), .Y(u1__abc_43968_n197) );
  INVX1 INVX1_680 ( .A(u2_o_249_), .Y(u2__abc_44228_n4330) );
  INVX1 INVX1_681 ( .A(u2__abc_44228_n4331), .Y(u2__abc_44228_n4332) );
  INVX1 INVX1_682 ( .A(u2_remHi_249_), .Y(u2__abc_44228_n4333) );
  INVX1 INVX1_683 ( .A(u2__abc_44228_n4334), .Y(u2__abc_44228_n4335) );
  INVX1 INVX1_684 ( .A(u2_o_248_), .Y(u2__abc_44228_n4337) );
  INVX1 INVX1_685 ( .A(u2_remHi_248_), .Y(u2__abc_44228_n4339) );
  INVX1 INVX1_686 ( .A(u2__abc_44228_n4341), .Y(u2__abc_44228_n4342) );
  INVX1 INVX1_687 ( .A(u2_o_246_), .Y(u2__abc_44228_n4344) );
  INVX1 INVX1_688 ( .A(u2_remHi_246_), .Y(u2__abc_44228_n4346) );
  INVX1 INVX1_689 ( .A(u2__abc_44228_n4348), .Y(u2__abc_44228_n4349_1) );
  INVX1 INVX1_69 ( .A(\a[63] ), .Y(u1__abc_43968_n198) );
  INVX1 INVX1_690 ( .A(u2_o_247_), .Y(u2__abc_44228_n4350) );
  INVX1 INVX1_691 ( .A(u2__abc_44228_n4351), .Y(u2__abc_44228_n4352) );
  INVX1 INVX1_692 ( .A(u2_remHi_247_), .Y(u2__abc_44228_n4353) );
  INVX1 INVX1_693 ( .A(u2__abc_44228_n4354), .Y(u2__abc_44228_n4355) );
  INVX1 INVX1_694 ( .A(u2_o_245_), .Y(u2__abc_44228_n4360) );
  INVX1 INVX1_695 ( .A(u2__abc_44228_n4361), .Y(u2__abc_44228_n4362) );
  INVX1 INVX1_696 ( .A(u2_remHi_245_), .Y(u2__abc_44228_n4363) );
  INVX1 INVX1_697 ( .A(u2__abc_44228_n4364), .Y(u2__abc_44228_n4365) );
  INVX1 INVX1_698 ( .A(u2_o_244_), .Y(u2__abc_44228_n4367) );
  INVX1 INVX1_699 ( .A(u2_remHi_244_), .Y(u2__abc_44228_n4369) );
  INVX1 INVX1_7 ( .A(_abc_64468_n1524), .Y(_abc_64468_n1532) );
  INVX1 INVX1_70 ( .A(\a[60] ), .Y(u1__abc_43968_n200) );
  INVX1 INVX1_700 ( .A(u2__abc_44228_n4371), .Y(u2__abc_44228_n4372) );
  INVX1 INVX1_701 ( .A(u2_o_242_), .Y(u2__abc_44228_n4374) );
  INVX1 INVX1_702 ( .A(u2_remHi_242_), .Y(u2__abc_44228_n4376) );
  INVX1 INVX1_703 ( .A(u2__abc_44228_n4378), .Y(u2__abc_44228_n4379) );
  INVX1 INVX1_704 ( .A(u2_o_243_), .Y(u2__abc_44228_n4380) );
  INVX1 INVX1_705 ( .A(u2__abc_44228_n4381), .Y(u2__abc_44228_n4382) );
  INVX1 INVX1_706 ( .A(u2_remHi_243_), .Y(u2__abc_44228_n4383) );
  INVX1 INVX1_707 ( .A(u2__abc_44228_n4384), .Y(u2__abc_44228_n4385) );
  INVX1 INVX1_708 ( .A(u2_o_241_), .Y(u2__abc_44228_n4389) );
  INVX1 INVX1_709 ( .A(u2__abc_44228_n4390), .Y(u2__abc_44228_n4391) );
  INVX1 INVX1_71 ( .A(\a[61] ), .Y(u1__abc_43968_n201) );
  INVX1 INVX1_710 ( .A(u2_remHi_241_), .Y(u2__abc_44228_n4392) );
  INVX1 INVX1_711 ( .A(u2__abc_44228_n4393), .Y(u2__abc_44228_n4394) );
  INVX1 INVX1_712 ( .A(u2_o_240_), .Y(u2__abc_44228_n4396_1) );
  INVX1 INVX1_713 ( .A(u2_remHi_240_), .Y(u2__abc_44228_n4398) );
  INVX1 INVX1_714 ( .A(u2__abc_44228_n4400), .Y(u2__abc_44228_n4401) );
  INVX1 INVX1_715 ( .A(u2_o_238_), .Y(u2__abc_44228_n4403) );
  INVX1 INVX1_716 ( .A(u2_remHi_238_), .Y(u2__abc_44228_n4405_1) );
  INVX1 INVX1_717 ( .A(u2__abc_44228_n4407), .Y(u2__abc_44228_n4408) );
  INVX1 INVX1_718 ( .A(u2_o_239_), .Y(u2__abc_44228_n4409) );
  INVX1 INVX1_719 ( .A(u2__abc_44228_n4410), .Y(u2__abc_44228_n4411) );
  INVX1 INVX1_72 ( .A(\a[58] ), .Y(u1__abc_43968_n204) );
  INVX1 INVX1_720 ( .A(u2_remHi_239_), .Y(u2__abc_44228_n4412) );
  INVX1 INVX1_721 ( .A(u2__abc_44228_n4413), .Y(u2__abc_44228_n4414_1) );
  INVX1 INVX1_722 ( .A(u2_o_237_), .Y(u2__abc_44228_n4420) );
  INVX1 INVX1_723 ( .A(u2__abc_44228_n4421), .Y(u2__abc_44228_n4422) );
  INVX1 INVX1_724 ( .A(u2_remHi_237_), .Y(u2__abc_44228_n4423_1) );
  INVX1 INVX1_725 ( .A(u2__abc_44228_n4424), .Y(u2__abc_44228_n4425) );
  INVX1 INVX1_726 ( .A(u2_o_236_), .Y(u2__abc_44228_n4427) );
  INVX1 INVX1_727 ( .A(u2_remHi_236_), .Y(u2__abc_44228_n4429) );
  INVX1 INVX1_728 ( .A(u2__abc_44228_n4431), .Y(u2__abc_44228_n4432_1) );
  INVX1 INVX1_729 ( .A(u2_o_234_), .Y(u2__abc_44228_n4434) );
  INVX1 INVX1_73 ( .A(\a[59] ), .Y(u1__abc_43968_n205_1) );
  INVX1 INVX1_730 ( .A(u2_remHi_234_), .Y(u2__abc_44228_n4436) );
  INVX1 INVX1_731 ( .A(u2__abc_44228_n4438), .Y(u2__abc_44228_n4439) );
  INVX1 INVX1_732 ( .A(u2_o_235_), .Y(u2__abc_44228_n4440) );
  INVX1 INVX1_733 ( .A(u2__abc_44228_n4441), .Y(u2__abc_44228_n4442_1) );
  INVX1 INVX1_734 ( .A(u2_remHi_235_), .Y(u2__abc_44228_n4443) );
  INVX1 INVX1_735 ( .A(u2__abc_44228_n4444), .Y(u2__abc_44228_n4445) );
  INVX1 INVX1_736 ( .A(u2_o_231_), .Y(u2__abc_44228_n4449) );
  INVX1 INVX1_737 ( .A(u2__abc_44228_n4450), .Y(u2__abc_44228_n4451_1) );
  INVX1 INVX1_738 ( .A(u2_remHi_231_), .Y(u2__abc_44228_n4452) );
  INVX1 INVX1_739 ( .A(u2__abc_44228_n4453), .Y(u2__abc_44228_n4454) );
  INVX1 INVX1_74 ( .A(\a[56] ), .Y(u1__abc_43968_n207) );
  INVX1 INVX1_740 ( .A(u2_o_230_), .Y(u2__abc_44228_n4456) );
  INVX1 INVX1_741 ( .A(u2_remHi_230_), .Y(u2__abc_44228_n4458) );
  INVX1 INVX1_742 ( .A(u2__abc_44228_n4460), .Y(u2__abc_44228_n4461_1) );
  INVX1 INVX1_743 ( .A(u2_o_233_), .Y(u2__abc_44228_n4463) );
  INVX1 INVX1_744 ( .A(u2__abc_44228_n4464), .Y(u2__abc_44228_n4465) );
  INVX1 INVX1_745 ( .A(u2_remHi_233_), .Y(u2__abc_44228_n4466) );
  INVX1 INVX1_746 ( .A(u2__abc_44228_n4467), .Y(u2__abc_44228_n4468) );
  INVX1 INVX1_747 ( .A(u2_o_232_), .Y(u2__abc_44228_n4470) );
  INVX1 INVX1_748 ( .A(u2_remHi_232_), .Y(u2__abc_44228_n4472) );
  INVX1 INVX1_749 ( .A(u2__abc_44228_n4474), .Y(u2__abc_44228_n4475) );
  INVX1 INVX1_75 ( .A(\a[57] ), .Y(u1__abc_43968_n208) );
  INVX1 INVX1_750 ( .A(u2_o_229_), .Y(u2__abc_44228_n4479) );
  INVX1 INVX1_751 ( .A(u2__abc_44228_n4480_1), .Y(u2__abc_44228_n4481) );
  INVX1 INVX1_752 ( .A(u2_remHi_229_), .Y(u2__abc_44228_n4482) );
  INVX1 INVX1_753 ( .A(u2__abc_44228_n4483), .Y(u2__abc_44228_n4484) );
  INVX1 INVX1_754 ( .A(u2_o_228_), .Y(u2__abc_44228_n4486) );
  INVX1 INVX1_755 ( .A(u2_remHi_228_), .Y(u2__abc_44228_n4488) );
  INVX1 INVX1_756 ( .A(u2__abc_44228_n4490), .Y(u2__abc_44228_n4491) );
  INVX1 INVX1_757 ( .A(u2_o_226_), .Y(u2__abc_44228_n4493) );
  INVX1 INVX1_758 ( .A(u2_remHi_226_), .Y(u2__abc_44228_n4495) );
  INVX1 INVX1_759 ( .A(u2__abc_44228_n4497), .Y(u2__abc_44228_n4498_1) );
  INVX1 INVX1_76 ( .A(\a[54] ), .Y(u1__abc_43968_n212_1) );
  INVX1 INVX1_760 ( .A(u2_o_227_), .Y(u2__abc_44228_n4499) );
  INVX1 INVX1_761 ( .A(u2__abc_44228_n4500), .Y(u2__abc_44228_n4501) );
  INVX1 INVX1_762 ( .A(u2_remHi_227_), .Y(u2__abc_44228_n4502) );
  INVX1 INVX1_763 ( .A(u2__abc_44228_n4503), .Y(u2__abc_44228_n4504) );
  INVX1 INVX1_764 ( .A(sqrto_225_), .Y(u2__abc_44228_n4508_1) );
  INVX1 INVX1_765 ( .A(u2__abc_44228_n4509), .Y(u2__abc_44228_n4510) );
  INVX1 INVX1_766 ( .A(u2_remHi_225_), .Y(u2__abc_44228_n4511) );
  INVX1 INVX1_767 ( .A(u2__abc_44228_n4512), .Y(u2__abc_44228_n4513) );
  INVX1 INVX1_768 ( .A(sqrto_224_), .Y(u2__abc_44228_n4515) );
  INVX1 INVX1_769 ( .A(u2_remHi_224_), .Y(u2__abc_44228_n4517_1) );
  INVX1 INVX1_77 ( .A(\a[55] ), .Y(u1__abc_43968_n213_1) );
  INVX1 INVX1_770 ( .A(u2__abc_44228_n4519), .Y(u2__abc_44228_n4520) );
  INVX1 INVX1_771 ( .A(sqrto_222_), .Y(u2__abc_44228_n4522) );
  INVX1 INVX1_772 ( .A(u2_remHi_222_), .Y(u2__abc_44228_n4524) );
  INVX1 INVX1_773 ( .A(u2__abc_44228_n4526_1), .Y(u2__abc_44228_n4527) );
  INVX1 INVX1_774 ( .A(sqrto_223_), .Y(u2__abc_44228_n4528) );
  INVX1 INVX1_775 ( .A(u2__abc_44228_n4529), .Y(u2__abc_44228_n4530) );
  INVX1 INVX1_776 ( .A(u2_remHi_223_), .Y(u2__abc_44228_n4531) );
  INVX1 INVX1_777 ( .A(u2__abc_44228_n4532), .Y(u2__abc_44228_n4533) );
  INVX1 INVX1_778 ( .A(sqrto_221_), .Y(u2__abc_44228_n4540) );
  INVX1 INVX1_779 ( .A(u2__abc_44228_n4541), .Y(u2__abc_44228_n4542) );
  INVX1 INVX1_78 ( .A(\a[52] ), .Y(u1__abc_43968_n215) );
  INVX1 INVX1_780 ( .A(u2_remHi_221_), .Y(u2__abc_44228_n4543) );
  INVX1 INVX1_781 ( .A(u2__abc_44228_n4544), .Y(u2__abc_44228_n4545_1) );
  INVX1 INVX1_782 ( .A(sqrto_220_), .Y(u2__abc_44228_n4547) );
  INVX1 INVX1_783 ( .A(u2_remHi_220_), .Y(u2__abc_44228_n4549) );
  INVX1 INVX1_784 ( .A(u2__abc_44228_n4551), .Y(u2__abc_44228_n4552) );
  INVX1 INVX1_785 ( .A(sqrto_218_), .Y(u2__abc_44228_n4554_1) );
  INVX1 INVX1_786 ( .A(u2_remHi_218_), .Y(u2__abc_44228_n4556) );
  INVX1 INVX1_787 ( .A(u2__abc_44228_n4558), .Y(u2__abc_44228_n4559) );
  INVX1 INVX1_788 ( .A(sqrto_219_), .Y(u2__abc_44228_n4560) );
  INVX1 INVX1_789 ( .A(u2__abc_44228_n4561), .Y(u2__abc_44228_n4562) );
  INVX1 INVX1_79 ( .A(\a[53] ), .Y(u1__abc_43968_n216) );
  INVX1 INVX1_790 ( .A(u2_remHi_219_), .Y(u2__abc_44228_n4563_1) );
  INVX1 INVX1_791 ( .A(u2__abc_44228_n4564), .Y(u2__abc_44228_n4565) );
  INVX1 INVX1_792 ( .A(sqrto_217_), .Y(u2__abc_44228_n4569) );
  INVX1 INVX1_793 ( .A(u2__abc_44228_n4570), .Y(u2__abc_44228_n4571) );
  INVX1 INVX1_794 ( .A(u2_remHi_217_), .Y(u2__abc_44228_n4572_1) );
  INVX1 INVX1_795 ( .A(u2__abc_44228_n4573), .Y(u2__abc_44228_n4574) );
  INVX1 INVX1_796 ( .A(sqrto_216_), .Y(u2__abc_44228_n4576) );
  INVX1 INVX1_797 ( .A(u2_remHi_216_), .Y(u2__abc_44228_n4578) );
  INVX1 INVX1_798 ( .A(u2__abc_44228_n4580), .Y(u2__abc_44228_n4581_1) );
  INVX1 INVX1_799 ( .A(sqrto_214_), .Y(u2__abc_44228_n4583) );
  INVX1 INVX1_8 ( .A(\a[116] ), .Y(_abc_64468_n1538) );
  INVX1 INVX1_80 ( .A(\a[50] ), .Y(u1__abc_43968_n219) );
  INVX1 INVX1_800 ( .A(u2_remHi_214_), .Y(u2__abc_44228_n4585) );
  INVX1 INVX1_801 ( .A(u2__abc_44228_n4587), .Y(u2__abc_44228_n4588) );
  INVX1 INVX1_802 ( .A(sqrto_215_), .Y(u2__abc_44228_n4589) );
  INVX1 INVX1_803 ( .A(u2__abc_44228_n4590), .Y(u2__abc_44228_n4591_1) );
  INVX1 INVX1_804 ( .A(u2_remHi_215_), .Y(u2__abc_44228_n4592) );
  INVX1 INVX1_805 ( .A(u2__abc_44228_n4593), .Y(u2__abc_44228_n4594) );
  INVX1 INVX1_806 ( .A(sqrto_213_), .Y(u2__abc_44228_n4599) );
  INVX1 INVX1_807 ( .A(u2__abc_44228_n4600_1), .Y(u2__abc_44228_n4601) );
  INVX1 INVX1_808 ( .A(u2_remHi_213_), .Y(u2__abc_44228_n4602) );
  INVX1 INVX1_809 ( .A(u2__abc_44228_n4603), .Y(u2__abc_44228_n4604) );
  INVX1 INVX1_81 ( .A(\a[51] ), .Y(u1__abc_43968_n220_1) );
  INVX1 INVX1_810 ( .A(sqrto_212_), .Y(u2__abc_44228_n4606) );
  INVX1 INVX1_811 ( .A(u2_remHi_212_), .Y(u2__abc_44228_n4608) );
  INVX1 INVX1_812 ( .A(u2__abc_44228_n4610_1), .Y(u2__abc_44228_n4611) );
  INVX1 INVX1_813 ( .A(sqrto_210_), .Y(u2__abc_44228_n4613) );
  INVX1 INVX1_814 ( .A(u2_remHi_210_), .Y(u2__abc_44228_n4615) );
  INVX1 INVX1_815 ( .A(u2__abc_44228_n4617), .Y(u2__abc_44228_n4618) );
  INVX1 INVX1_816 ( .A(sqrto_211_), .Y(u2__abc_44228_n4619) );
  INVX1 INVX1_817 ( .A(u2__abc_44228_n4620_1), .Y(u2__abc_44228_n4621) );
  INVX1 INVX1_818 ( .A(u2_remHi_211_), .Y(u2__abc_44228_n4622) );
  INVX1 INVX1_819 ( .A(u2__abc_44228_n4623), .Y(u2__abc_44228_n4624) );
  INVX1 INVX1_82 ( .A(\a[48] ), .Y(u1__abc_43968_n222) );
  INVX1 INVX1_820 ( .A(sqrto_209_), .Y(u2__abc_44228_n4628) );
  INVX1 INVX1_821 ( .A(u2__abc_44228_n4629_1), .Y(u2__abc_44228_n4630) );
  INVX1 INVX1_822 ( .A(u2_remHi_209_), .Y(u2__abc_44228_n4631) );
  INVX1 INVX1_823 ( .A(u2__abc_44228_n4632), .Y(u2__abc_44228_n4633) );
  INVX1 INVX1_824 ( .A(sqrto_208_), .Y(u2__abc_44228_n4635) );
  INVX1 INVX1_825 ( .A(u2_remHi_208_), .Y(u2__abc_44228_n4637) );
  INVX1 INVX1_826 ( .A(u2__abc_44228_n4639), .Y(u2__abc_44228_n4640) );
  INVX1 INVX1_827 ( .A(sqrto_207_), .Y(u2__abc_44228_n4642) );
  INVX1 INVX1_828 ( .A(u2__abc_44228_n4643), .Y(u2__abc_44228_n4644) );
  INVX1 INVX1_829 ( .A(u2_remHi_207_), .Y(u2__abc_44228_n4645) );
  INVX1 INVX1_83 ( .A(\a[49] ), .Y(u1__abc_43968_n223) );
  INVX1 INVX1_830 ( .A(u2__abc_44228_n4646_1), .Y(u2__abc_44228_n4647) );
  INVX1 INVX1_831 ( .A(sqrto_206_), .Y(u2__abc_44228_n4649) );
  INVX1 INVX1_832 ( .A(u2_remHi_206_), .Y(u2__abc_44228_n4651) );
  INVX1 INVX1_833 ( .A(u2__abc_44228_n4653), .Y(u2__abc_44228_n4654) );
  INVX1 INVX1_834 ( .A(sqrto_205_), .Y(u2__abc_44228_n4659) );
  INVX1 INVX1_835 ( .A(u2__abc_44228_n4660), .Y(u2__abc_44228_n4661) );
  INVX1 INVX1_836 ( .A(u2_remHi_205_), .Y(u2__abc_44228_n4662) );
  INVX1 INVX1_837 ( .A(u2__abc_44228_n4663), .Y(u2__abc_44228_n4664) );
  INVX1 INVX1_838 ( .A(sqrto_204_), .Y(u2__abc_44228_n4666) );
  INVX1 INVX1_839 ( .A(u2_remHi_204_), .Y(u2__abc_44228_n4668) );
  INVX1 INVX1_84 ( .A(\a[110] ), .Y(u1__abc_43968_n228_1) );
  INVX1 INVX1_840 ( .A(u2__abc_44228_n4670), .Y(u2__abc_44228_n4671) );
  INVX1 INVX1_841 ( .A(sqrto_203_), .Y(u2__abc_44228_n4673) );
  INVX1 INVX1_842 ( .A(u2__abc_44228_n4674_1), .Y(u2__abc_44228_n4675) );
  INVX1 INVX1_843 ( .A(u2_remHi_203_), .Y(u2__abc_44228_n4676) );
  INVX1 INVX1_844 ( .A(u2__abc_44228_n4677), .Y(u2__abc_44228_n4678) );
  INVX1 INVX1_845 ( .A(sqrto_202_), .Y(u2__abc_44228_n4680) );
  INVX1 INVX1_846 ( .A(u2_remHi_202_), .Y(u2__abc_44228_n4682) );
  INVX1 INVX1_847 ( .A(u2__abc_44228_n4684), .Y(u2__abc_44228_n4685_1) );
  INVX1 INVX1_848 ( .A(sqrto_201_), .Y(u2__abc_44228_n4688) );
  INVX1 INVX1_849 ( .A(u2__abc_44228_n4689), .Y(u2__abc_44228_n4690) );
  INVX1 INVX1_85 ( .A(\a[111] ), .Y(u1__abc_43968_n229) );
  INVX1 INVX1_850 ( .A(u2_remHi_201_), .Y(u2__abc_44228_n4691) );
  INVX1 INVX1_851 ( .A(u2__abc_44228_n4692), .Y(u2__abc_44228_n4693) );
  INVX1 INVX1_852 ( .A(sqrto_200_), .Y(u2__abc_44228_n4695_1) );
  INVX1 INVX1_853 ( .A(u2_remHi_200_), .Y(u2__abc_44228_n4697) );
  INVX1 INVX1_854 ( .A(u2__abc_44228_n4699), .Y(u2__abc_44228_n4700) );
  INVX1 INVX1_855 ( .A(sqrto_198_), .Y(u2__abc_44228_n4702) );
  INVX1 INVX1_856 ( .A(u2_remHi_198_), .Y(u2__abc_44228_n4704_1) );
  INVX1 INVX1_857 ( .A(u2__abc_44228_n4706), .Y(u2__abc_44228_n4707) );
  INVX1 INVX1_858 ( .A(sqrto_199_), .Y(u2__abc_44228_n4708) );
  INVX1 INVX1_859 ( .A(u2__abc_44228_n4709), .Y(u2__abc_44228_n4710) );
  INVX1 INVX1_86 ( .A(\a[108] ), .Y(u1__abc_43968_n231) );
  INVX1 INVX1_860 ( .A(u2_remHi_199_), .Y(u2__abc_44228_n4711) );
  INVX1 INVX1_861 ( .A(u2__abc_44228_n4712), .Y(u2__abc_44228_n4713_1) );
  INVX1 INVX1_862 ( .A(sqrto_197_), .Y(u2__abc_44228_n4718) );
  INVX1 INVX1_863 ( .A(u2__abc_44228_n4719), .Y(u2__abc_44228_n4720) );
  INVX1 INVX1_864 ( .A(u2_remHi_197_), .Y(u2__abc_44228_n4721) );
  INVX1 INVX1_865 ( .A(u2__abc_44228_n4722_1), .Y(u2__abc_44228_n4723) );
  INVX1 INVX1_866 ( .A(sqrto_196_), .Y(u2__abc_44228_n4725) );
  INVX1 INVX1_867 ( .A(u2_remHi_196_), .Y(u2__abc_44228_n4727) );
  INVX1 INVX1_868 ( .A(u2__abc_44228_n4729), .Y(u2__abc_44228_n4730) );
  INVX1 INVX1_869 ( .A(sqrto_195_), .Y(u2__abc_44228_n4732) );
  INVX1 INVX1_87 ( .A(\a[109] ), .Y(u1__abc_43968_n232) );
  INVX1 INVX1_870 ( .A(u2__abc_44228_n4733), .Y(u2__abc_44228_n4734) );
  INVX1 INVX1_871 ( .A(u2_remHi_195_), .Y(u2__abc_44228_n4735) );
  INVX1 INVX1_872 ( .A(u2__abc_44228_n4736), .Y(u2__abc_44228_n4737) );
  INVX1 INVX1_873 ( .A(sqrto_194_), .Y(u2__abc_44228_n4739) );
  INVX1 INVX1_874 ( .A(u2_remHi_194_), .Y(u2__abc_44228_n4741_1) );
  INVX1 INVX1_875 ( .A(u2__abc_44228_n4743), .Y(u2__abc_44228_n4744) );
  INVX1 INVX1_876 ( .A(sqrto_193_), .Y(u2__abc_44228_n4747) );
  INVX1 INVX1_877 ( .A(u2__abc_44228_n4748), .Y(u2__abc_44228_n4749) );
  INVX1 INVX1_878 ( .A(u2_remHi_193_), .Y(u2__abc_44228_n4750_1) );
  INVX1 INVX1_879 ( .A(u2__abc_44228_n4751), .Y(u2__abc_44228_n4752) );
  INVX1 INVX1_88 ( .A(\a[106] ), .Y(u1__abc_43968_n235) );
  INVX1 INVX1_880 ( .A(sqrto_192_), .Y(u2__abc_44228_n4754) );
  INVX1 INVX1_881 ( .A(u2_remHi_192_), .Y(u2__abc_44228_n4756) );
  INVX1 INVX1_882 ( .A(u2__abc_44228_n4758), .Y(u2__abc_44228_n4759) );
  INVX1 INVX1_883 ( .A(sqrto_190_), .Y(u2__abc_44228_n4761) );
  INVX1 INVX1_884 ( .A(u2_remHi_190_), .Y(u2__abc_44228_n4763) );
  INVX1 INVX1_885 ( .A(u2__abc_44228_n4765), .Y(u2__abc_44228_n4766) );
  INVX1 INVX1_886 ( .A(sqrto_191_), .Y(u2__abc_44228_n4767) );
  INVX1 INVX1_887 ( .A(u2__abc_44228_n4768), .Y(u2__abc_44228_n4769) );
  INVX1 INVX1_888 ( .A(u2_remHi_191_), .Y(u2__abc_44228_n4770_1) );
  INVX1 INVX1_889 ( .A(u2__abc_44228_n4771), .Y(u2__abc_44228_n4772) );
  INVX1 INVX1_89 ( .A(\a[107] ), .Y(u1__abc_43968_n236_1) );
  INVX1 INVX1_890 ( .A(sqrto_189_), .Y(u2__abc_44228_n4780) );
  INVX1 INVX1_891 ( .A(u2__abc_44228_n4781), .Y(u2__abc_44228_n4782) );
  INVX1 INVX1_892 ( .A(u2_remHi_189_), .Y(u2__abc_44228_n4783) );
  INVX1 INVX1_893 ( .A(u2__abc_44228_n4784), .Y(u2__abc_44228_n4785) );
  INVX1 INVX1_894 ( .A(sqrto_188_), .Y(u2__abc_44228_n4787) );
  INVX1 INVX1_895 ( .A(u2_remHi_188_), .Y(u2__abc_44228_n4789) );
  INVX1 INVX1_896 ( .A(u2__abc_44228_n4791), .Y(u2__abc_44228_n4792) );
  INVX1 INVX1_897 ( .A(sqrto_187_), .Y(u2__abc_44228_n4794) );
  INVX1 INVX1_898 ( .A(u2__abc_44228_n4795), .Y(u2__abc_44228_n4796) );
  INVX1 INVX1_899 ( .A(u2_remHi_187_), .Y(u2__abc_44228_n4797) );
  INVX1 INVX1_9 ( .A(_abc_64468_n1541), .Y(_abc_64468_n1542) );
  INVX1 INVX1_90 ( .A(\a[104] ), .Y(u1__abc_43968_n238) );
  INVX1 INVX1_900 ( .A(u2__abc_44228_n4798), .Y(u2__abc_44228_n4799_1) );
  INVX1 INVX1_901 ( .A(sqrto_186_), .Y(u2__abc_44228_n4801) );
  INVX1 INVX1_902 ( .A(u2_remHi_186_), .Y(u2__abc_44228_n4803) );
  INVX1 INVX1_903 ( .A(u2__abc_44228_n4805), .Y(u2__abc_44228_n4806) );
  INVX1 INVX1_904 ( .A(sqrto_183_), .Y(u2__abc_44228_n4809_1) );
  INVX1 INVX1_905 ( .A(u2__abc_44228_n4810), .Y(u2__abc_44228_n4811) );
  INVX1 INVX1_906 ( .A(u2_remHi_183_), .Y(u2__abc_44228_n4812) );
  INVX1 INVX1_907 ( .A(u2__abc_44228_n4813), .Y(u2__abc_44228_n4814) );
  INVX1 INVX1_908 ( .A(sqrto_182_), .Y(u2__abc_44228_n4816) );
  INVX1 INVX1_909 ( .A(u2_remHi_182_), .Y(u2__abc_44228_n4818_1) );
  INVX1 INVX1_91 ( .A(\a[105] ), .Y(u1__abc_43968_n239) );
  INVX1 INVX1_910 ( .A(u2__abc_44228_n4820), .Y(u2__abc_44228_n4821) );
  INVX1 INVX1_911 ( .A(sqrto_185_), .Y(u2__abc_44228_n4823) );
  INVX1 INVX1_912 ( .A(u2__abc_44228_n4824), .Y(u2__abc_44228_n4825) );
  INVX1 INVX1_913 ( .A(u2_remHi_185_), .Y(u2__abc_44228_n4826) );
  INVX1 INVX1_914 ( .A(u2__abc_44228_n4827_1), .Y(u2__abc_44228_n4828) );
  INVX1 INVX1_915 ( .A(sqrto_184_), .Y(u2__abc_44228_n4830) );
  INVX1 INVX1_916 ( .A(u2_remHi_184_), .Y(u2__abc_44228_n4832) );
  INVX1 INVX1_917 ( .A(u2__abc_44228_n4834), .Y(u2__abc_44228_n4835) );
  INVX1 INVX1_918 ( .A(sqrto_181_), .Y(u2__abc_44228_n4839) );
  INVX1 INVX1_919 ( .A(u2__abc_44228_n4840), .Y(u2__abc_44228_n4841) );
  INVX1 INVX1_92 ( .A(\a[102] ), .Y(u1__abc_43968_n243_1) );
  INVX1 INVX1_920 ( .A(u2_remHi_181_), .Y(u2__abc_44228_n4842) );
  INVX1 INVX1_921 ( .A(u2__abc_44228_n4843), .Y(u2__abc_44228_n4844) );
  INVX1 INVX1_922 ( .A(sqrto_180_), .Y(u2__abc_44228_n4846_1) );
  INVX1 INVX1_923 ( .A(u2_remHi_180_), .Y(u2__abc_44228_n4848) );
  INVX1 INVX1_924 ( .A(u2__abc_44228_n4850), .Y(u2__abc_44228_n4851) );
  INVX1 INVX1_925 ( .A(sqrto_179_), .Y(u2__abc_44228_n4853) );
  INVX1 INVX1_926 ( .A(u2__abc_44228_n4854), .Y(u2__abc_44228_n4855_1) );
  INVX1 INVX1_927 ( .A(u2_remHi_179_), .Y(u2__abc_44228_n4856) );
  INVX1 INVX1_928 ( .A(u2__abc_44228_n4857), .Y(u2__abc_44228_n4858) );
  INVX1 INVX1_929 ( .A(sqrto_178_), .Y(u2__abc_44228_n4860) );
  INVX1 INVX1_93 ( .A(\a[103] ), .Y(u1__abc_43968_n244_1) );
  INVX1 INVX1_930 ( .A(u2_remHi_178_), .Y(u2__abc_44228_n4862) );
  INVX1 INVX1_931 ( .A(u2__abc_44228_n4864_1), .Y(u2__abc_44228_n4865) );
  INVX1 INVX1_932 ( .A(sqrto_177_), .Y(u2__abc_44228_n4868) );
  INVX1 INVX1_933 ( .A(u2__abc_44228_n4869), .Y(u2__abc_44228_n4870) );
  INVX1 INVX1_934 ( .A(u2_remHi_177_), .Y(u2__abc_44228_n4871) );
  INVX1 INVX1_935 ( .A(u2__abc_44228_n4872), .Y(u2__abc_44228_n4873_1) );
  INVX1 INVX1_936 ( .A(sqrto_176_), .Y(u2__abc_44228_n4875) );
  INVX1 INVX1_937 ( .A(u2_remHi_176_), .Y(u2__abc_44228_n4877) );
  INVX1 INVX1_938 ( .A(u2__abc_44228_n4879), .Y(u2__abc_44228_n4880) );
  INVX1 INVX1_939 ( .A(sqrto_175_), .Y(u2__abc_44228_n4882_1) );
  INVX1 INVX1_94 ( .A(\a[100] ), .Y(u1__abc_43968_n246) );
  INVX1 INVX1_940 ( .A(u2__abc_44228_n4883), .Y(u2__abc_44228_n4884) );
  INVX1 INVX1_941 ( .A(u2_remHi_175_), .Y(u2__abc_44228_n4885) );
  INVX1 INVX1_942 ( .A(u2__abc_44228_n4886), .Y(u2__abc_44228_n4887) );
  INVX1 INVX1_943 ( .A(sqrto_174_), .Y(u2__abc_44228_n4889) );
  INVX1 INVX1_944 ( .A(u2_remHi_174_), .Y(u2__abc_44228_n4891) );
  INVX1 INVX1_945 ( .A(u2__abc_44228_n4893), .Y(u2__abc_44228_n4894) );
  INVX1 INVX1_946 ( .A(sqrto_173_), .Y(u2__abc_44228_n4899) );
  INVX1 INVX1_947 ( .A(u2__abc_44228_n4900), .Y(u2__abc_44228_n4901_1) );
  INVX1 INVX1_948 ( .A(u2_remHi_173_), .Y(u2__abc_44228_n4902) );
  INVX1 INVX1_949 ( .A(u2__abc_44228_n4903), .Y(u2__abc_44228_n4904) );
  INVX1 INVX1_95 ( .A(\a[101] ), .Y(u1__abc_43968_n247) );
  INVX1 INVX1_950 ( .A(sqrto_172_), .Y(u2__abc_44228_n4906) );
  INVX1 INVX1_951 ( .A(u2_remHi_172_), .Y(u2__abc_44228_n4908) );
  INVX1 INVX1_952 ( .A(u2__abc_44228_n4910), .Y(u2__abc_44228_n4911_1) );
  INVX1 INVX1_953 ( .A(sqrto_170_), .Y(u2__abc_44228_n4913) );
  INVX1 INVX1_954 ( .A(u2_remHi_170_), .Y(u2__abc_44228_n4915) );
  INVX1 INVX1_955 ( .A(u2__abc_44228_n4917), .Y(u2__abc_44228_n4918) );
  INVX1 INVX1_956 ( .A(sqrto_171_), .Y(u2__abc_44228_n4919) );
  INVX1 INVX1_957 ( .A(u2__abc_44228_n4920), .Y(u2__abc_44228_n4921_1) );
  INVX1 INVX1_958 ( .A(u2_remHi_171_), .Y(u2__abc_44228_n4922) );
  INVX1 INVX1_959 ( .A(u2__abc_44228_n4923), .Y(u2__abc_44228_n4924) );
  INVX1 INVX1_96 ( .A(\a[98] ), .Y(u1__abc_43968_n250) );
  INVX1 INVX1_960 ( .A(sqrto_169_), .Y(u2__abc_44228_n4928) );
  INVX1 INVX1_961 ( .A(u2__abc_44228_n4929), .Y(u2__abc_44228_n4930_1) );
  INVX1 INVX1_962 ( .A(u2_remHi_169_), .Y(u2__abc_44228_n4931) );
  INVX1 INVX1_963 ( .A(u2__abc_44228_n4932), .Y(u2__abc_44228_n4933) );
  INVX1 INVX1_964 ( .A(sqrto_168_), .Y(u2__abc_44228_n4935) );
  INVX1 INVX1_965 ( .A(u2_remHi_168_), .Y(u2__abc_44228_n4937) );
  INVX1 INVX1_966 ( .A(u2__abc_44228_n4939_1), .Y(u2__abc_44228_n4940) );
  INVX1 INVX1_967 ( .A(sqrto_166_), .Y(u2__abc_44228_n4942) );
  INVX1 INVX1_968 ( .A(u2_remHi_166_), .Y(u2__abc_44228_n4944) );
  INVX1 INVX1_969 ( .A(u2__abc_44228_n4946), .Y(u2__abc_44228_n4947) );
  INVX1 INVX1_97 ( .A(\a[99] ), .Y(u1__abc_43968_n251_1) );
  INVX1 INVX1_970 ( .A(sqrto_167_), .Y(u2__abc_44228_n4948_1) );
  INVX1 INVX1_971 ( .A(u2__abc_44228_n4949), .Y(u2__abc_44228_n4950) );
  INVX1 INVX1_972 ( .A(u2_remHi_167_), .Y(u2__abc_44228_n4951) );
  INVX1 INVX1_973 ( .A(u2__abc_44228_n4952), .Y(u2__abc_44228_n4953) );
  INVX1 INVX1_974 ( .A(sqrto_165_), .Y(u2__abc_44228_n4958) );
  INVX1 INVX1_975 ( .A(u2__abc_44228_n4959), .Y(u2__abc_44228_n4960) );
  INVX1 INVX1_976 ( .A(u2_remHi_165_), .Y(u2__abc_44228_n4961) );
  INVX1 INVX1_977 ( .A(u2__abc_44228_n4962), .Y(u2__abc_44228_n4963) );
  INVX1 INVX1_978 ( .A(sqrto_164_), .Y(u2__abc_44228_n4965) );
  INVX1 INVX1_979 ( .A(u2_remHi_164_), .Y(u2__abc_44228_n4967_1) );
  INVX1 INVX1_98 ( .A(\a[96] ), .Y(u1__abc_43968_n253) );
  INVX1 INVX1_980 ( .A(u2__abc_44228_n4969), .Y(u2__abc_44228_n4970) );
  INVX1 INVX1_981 ( .A(sqrto_162_), .Y(u2__abc_44228_n4972) );
  INVX1 INVX1_982 ( .A(u2_remHi_162_), .Y(u2__abc_44228_n4974) );
  INVX1 INVX1_983 ( .A(u2__abc_44228_n4976_1), .Y(u2__abc_44228_n4977) );
  INVX1 INVX1_984 ( .A(sqrto_163_), .Y(u2__abc_44228_n4978) );
  INVX1 INVX1_985 ( .A(u2__abc_44228_n4979), .Y(u2__abc_44228_n4980) );
  INVX1 INVX1_986 ( .A(u2_remHi_163_), .Y(u2__abc_44228_n4981) );
  INVX1 INVX1_987 ( .A(u2__abc_44228_n4982), .Y(u2__abc_44228_n4983) );
  INVX1 INVX1_988 ( .A(sqrto_161_), .Y(u2__abc_44228_n4987) );
  INVX1 INVX1_989 ( .A(u2__abc_44228_n4988), .Y(u2__abc_44228_n4989) );
  INVX1 INVX1_99 ( .A(\a[97] ), .Y(u1__abc_43968_n254) );
  INVX1 INVX1_990 ( .A(u2_remHi_161_), .Y(u2__abc_44228_n4990) );
  INVX1 INVX1_991 ( .A(u2__abc_44228_n4991), .Y(u2__abc_44228_n4992) );
  INVX1 INVX1_992 ( .A(sqrto_160_), .Y(u2__abc_44228_n4994) );
  INVX1 INVX1_993 ( .A(u2_remHi_160_), .Y(u2__abc_44228_n4996_1) );
  INVX1 INVX1_994 ( .A(u2__abc_44228_n4998), .Y(u2__abc_44228_n4999) );
  INVX1 INVX1_995 ( .A(sqrto_158_), .Y(u2__abc_44228_n5001) );
  INVX1 INVX1_996 ( .A(u2_remHi_158_), .Y(u2__abc_44228_n5003) );
  INVX1 INVX1_997 ( .A(u2__abc_44228_n5005_1), .Y(u2__abc_44228_n5006) );
  INVX1 INVX1_998 ( .A(sqrto_159_), .Y(u2__abc_44228_n5007) );
  INVX1 INVX1_999 ( .A(u2__abc_44228_n5008), .Y(u2__abc_44228_n5009) );
  INVX8 INVX8_1 ( .A(aNan_bF_buf10), .Y(_abc_64468_n753) );
  INVX8 INVX8_2 ( .A(a_112_bF_buf7), .Y(_abc_64468_n1170) );
  INVX8 INVX8_3 ( .A(rst), .Y(u2__abc_44228_n2966) );
  INVX8 INVX8_4 ( .A(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n2984) );
  INVX8 INVX8_5 ( .A(u2__abc_44228_n7547_bF_buf57), .Y(u2__abc_44228_n7548_1) );
  OR2X2 OR2X2_1 ( .A(aNan_bF_buf9), .B(sqrto_76_), .Y(_abc_64468_n830) );
  OR2X2 OR2X2_10 ( .A(_abc_64468_n753_bF_buf3), .B(\a[4] ), .Y(_abc_64468_n843) );
  OR2X2 OR2X2_100 ( .A(_abc_64468_n753_bF_buf0), .B(\a[49] ), .Y(_abc_64468_n978) );
  OR2X2 OR2X2_1000 ( .A(u2__abc_44228_n6623), .B(u2__abc_44228_n6248), .Y(u2__abc_44228_n6624) );
  OR2X2 OR2X2_1001 ( .A(u2__abc_44228_n6628), .B(u2__abc_44228_n6231), .Y(u2__abc_44228_n6629) );
  OR2X2 OR2X2_1002 ( .A(u2__abc_44228_n6627), .B(u2__abc_44228_n6629), .Y(u2__abc_44228_n6630) );
  OR2X2 OR2X2_1003 ( .A(u2__abc_44228_n6622), .B(u2__abc_44228_n6630), .Y(u2__abc_44228_n6631) );
  OR2X2 OR2X2_1004 ( .A(u2__abc_44228_n6633), .B(u2__abc_44228_n6204), .Y(u2__abc_44228_n6634_1) );
  OR2X2 OR2X2_1005 ( .A(u2__abc_44228_n6637), .B(u2__abc_44228_n6641), .Y(u2__abc_44228_n6642) );
  OR2X2 OR2X2_1006 ( .A(u2__abc_44228_n6649), .B(u2__abc_44228_n6172), .Y(u2__abc_44228_n6650) );
  OR2X2 OR2X2_1007 ( .A(u2__abc_44228_n6648), .B(u2__abc_44228_n6650), .Y(u2__abc_44228_n6651) );
  OR2X2 OR2X2_1008 ( .A(u2__abc_44228_n6643), .B(u2__abc_44228_n6651), .Y(u2__abc_44228_n6652) );
  OR2X2 OR2X2_1009 ( .A(u2__abc_44228_n6632), .B(u2__abc_44228_n6652), .Y(u2__abc_44228_n6653_1) );
  OR2X2 OR2X2_101 ( .A(aNan_bF_buf3), .B(sqrto_126_), .Y(_abc_64468_n980) );
  OR2X2 OR2X2_1010 ( .A(u2__abc_44228_n6655), .B(u2__abc_44228_n6164), .Y(u2__abc_44228_n6656) );
  OR2X2 OR2X2_1011 ( .A(u2__abc_44228_n6660), .B(u2__abc_44228_n6141_1), .Y(u2__abc_44228_n6661) );
  OR2X2 OR2X2_1012 ( .A(u2__abc_44228_n6659), .B(u2__abc_44228_n6661), .Y(u2__abc_44228_n6662) );
  OR2X2 OR2X2_1013 ( .A(u2__abc_44228_n6664), .B(u2__abc_44228_n6135), .Y(u2__abc_44228_n6665) );
  OR2X2 OR2X2_1014 ( .A(u2__abc_44228_n6669), .B(u2__abc_44228_n6112), .Y(u2__abc_44228_n6670) );
  OR2X2 OR2X2_1015 ( .A(u2__abc_44228_n6668), .B(u2__abc_44228_n6670), .Y(u2__abc_44228_n6671_1) );
  OR2X2 OR2X2_1016 ( .A(u2__abc_44228_n6663_1), .B(u2__abc_44228_n6671_1), .Y(u2__abc_44228_n6672) );
  OR2X2 OR2X2_1017 ( .A(u2__abc_44228_n6674), .B(u2__abc_44228_n6099), .Y(u2__abc_44228_n6675) );
  OR2X2 OR2X2_1018 ( .A(u2__abc_44228_n6678), .B(u2__abc_44228_n6682), .Y(u2__abc_44228_n6683) );
  OR2X2 OR2X2_1019 ( .A(u2__abc_44228_n6685), .B(u2__abc_44228_n6053), .Y(u2__abc_44228_n6686) );
  OR2X2 OR2X2_102 ( .A(_abc_64468_n753_bF_buf13), .B(\a[50] ), .Y(_abc_64468_n981) );
  OR2X2 OR2X2_1020 ( .A(u2__abc_44228_n6687), .B(u2__abc_44228_n6070), .Y(u2__abc_44228_n6688) );
  OR2X2 OR2X2_1021 ( .A(u2__abc_44228_n6691), .B(u2__abc_44228_n6686), .Y(u2__abc_44228_n6692) );
  OR2X2 OR2X2_1022 ( .A(u2__abc_44228_n6684), .B(u2__abc_44228_n6692), .Y(u2__abc_44228_n6693) );
  OR2X2 OR2X2_1023 ( .A(u2__abc_44228_n6673), .B(u2__abc_44228_n6693), .Y(u2__abc_44228_n6694) );
  OR2X2 OR2X2_1024 ( .A(u2__abc_44228_n6654), .B(u2__abc_44228_n6694), .Y(u2__abc_44228_n6695) );
  OR2X2 OR2X2_1025 ( .A(u2__abc_44228_n6613), .B(u2__abc_44228_n6695), .Y(u2__abc_44228_n6696) );
  OR2X2 OR2X2_1026 ( .A(u2__abc_44228_n6703), .B(u2__abc_44228_n6020), .Y(u2__abc_44228_n6704) );
  OR2X2 OR2X2_1027 ( .A(u2__abc_44228_n6702), .B(u2__abc_44228_n6704), .Y(u2__abc_44228_n6705) );
  OR2X2 OR2X2_1028 ( .A(u2__abc_44228_n6712), .B(u2__abc_44228_n5991), .Y(u2__abc_44228_n6713) );
  OR2X2 OR2X2_1029 ( .A(u2__abc_44228_n6711), .B(u2__abc_44228_n6713), .Y(u2__abc_44228_n6714) );
  OR2X2 OR2X2_103 ( .A(aNan_bF_buf2), .B(sqrto_127_), .Y(_abc_64468_n983) );
  OR2X2 OR2X2_1030 ( .A(u2__abc_44228_n6706), .B(u2__abc_44228_n6714), .Y(u2__abc_44228_n6715) );
  OR2X2 OR2X2_1031 ( .A(u2__abc_44228_n5961), .B(u2__abc_44228_n5968), .Y(u2__abc_44228_n6717_1) );
  OR2X2 OR2X2_1032 ( .A(u2__abc_44228_n6723), .B(u2__abc_44228_n6718), .Y(u2__abc_44228_n6724) );
  OR2X2 OR2X2_1033 ( .A(u2__abc_44228_n6731), .B(u2__abc_44228_n5932), .Y(u2__abc_44228_n6732) );
  OR2X2 OR2X2_1034 ( .A(u2__abc_44228_n6730), .B(u2__abc_44228_n6732), .Y(u2__abc_44228_n6733) );
  OR2X2 OR2X2_1035 ( .A(u2__abc_44228_n6725_1), .B(u2__abc_44228_n6733), .Y(u2__abc_44228_n6734) );
  OR2X2 OR2X2_1036 ( .A(u2__abc_44228_n6716), .B(u2__abc_44228_n6734), .Y(u2__abc_44228_n6735_1) );
  OR2X2 OR2X2_1037 ( .A(u2__abc_44228_n6737), .B(u2__abc_44228_n5918), .Y(u2__abc_44228_n6738) );
  OR2X2 OR2X2_1038 ( .A(u2__abc_44228_n6742), .B(u2__abc_44228_n5901_1), .Y(u2__abc_44228_n6743_1) );
  OR2X2 OR2X2_1039 ( .A(u2__abc_44228_n6741), .B(u2__abc_44228_n6743_1), .Y(u2__abc_44228_n6744) );
  OR2X2 OR2X2_104 ( .A(_abc_64468_n753_bF_buf12), .B(\a[51] ), .Y(_abc_64468_n984) );
  OR2X2 OR2X2_1040 ( .A(u2__abc_44228_n6751), .B(u2__abc_44228_n5872), .Y(u2__abc_44228_n6752) );
  OR2X2 OR2X2_1041 ( .A(u2__abc_44228_n6750), .B(u2__abc_44228_n6752), .Y(u2__abc_44228_n6753_1) );
  OR2X2 OR2X2_1042 ( .A(u2__abc_44228_n6745), .B(u2__abc_44228_n6753_1), .Y(u2__abc_44228_n6754) );
  OR2X2 OR2X2_1043 ( .A(u2__abc_44228_n6756), .B(u2__abc_44228_n5845_1), .Y(u2__abc_44228_n6757) );
  OR2X2 OR2X2_1044 ( .A(u2__abc_44228_n6760), .B(u2__abc_44228_n6764), .Y(u2__abc_44228_n6765) );
  OR2X2 OR2X2_1045 ( .A(u2__abc_44228_n6767), .B(u2__abc_44228_n5813), .Y(u2__abc_44228_n6768) );
  OR2X2 OR2X2_1046 ( .A(u2__abc_44228_n6773), .B(u2__abc_44228_n6768), .Y(u2__abc_44228_n6774) );
  OR2X2 OR2X2_1047 ( .A(u2__abc_44228_n6766), .B(u2__abc_44228_n6774), .Y(u2__abc_44228_n6775) );
  OR2X2 OR2X2_1048 ( .A(u2__abc_44228_n6755), .B(u2__abc_44228_n6775), .Y(u2__abc_44228_n6776) );
  OR2X2 OR2X2_1049 ( .A(u2__abc_44228_n6736), .B(u2__abc_44228_n6776), .Y(u2__abc_44228_n6777) );
  OR2X2 OR2X2_105 ( .A(aNan_bF_buf1), .B(sqrto_128_), .Y(_abc_64468_n986) );
  OR2X2 OR2X2_1050 ( .A(u2__abc_44228_n6779_1), .B(u2__abc_44228_n5798), .Y(u2__abc_44228_n6780) );
  OR2X2 OR2X2_1051 ( .A(u2__abc_44228_n6784), .B(u2__abc_44228_n5781), .Y(u2__abc_44228_n6785) );
  OR2X2 OR2X2_1052 ( .A(u2__abc_44228_n6783), .B(u2__abc_44228_n6785), .Y(u2__abc_44228_n6786) );
  OR2X2 OR2X2_1053 ( .A(u2__abc_44228_n6793), .B(u2__abc_44228_n5752), .Y(u2__abc_44228_n6794) );
  OR2X2 OR2X2_1054 ( .A(u2__abc_44228_n6792), .B(u2__abc_44228_n6794), .Y(u2__abc_44228_n6795) );
  OR2X2 OR2X2_1055 ( .A(u2__abc_44228_n6787), .B(u2__abc_44228_n6795), .Y(u2__abc_44228_n6796) );
  OR2X2 OR2X2_1056 ( .A(u2__abc_44228_n6798), .B(u2__abc_44228_n5725), .Y(u2__abc_44228_n6799) );
  OR2X2 OR2X2_1057 ( .A(u2__abc_44228_n6802), .B(u2__abc_44228_n6806), .Y(u2__abc_44228_n6807_1) );
  OR2X2 OR2X2_1058 ( .A(u2__abc_44228_n6809), .B(u2__abc_44228_n5693), .Y(u2__abc_44228_n6810) );
  OR2X2 OR2X2_1059 ( .A(u2__abc_44228_n6811), .B(u2__abc_44228_n5710_1), .Y(u2__abc_44228_n6812) );
  OR2X2 OR2X2_106 ( .A(_abc_64468_n753_bF_buf11), .B(\a[52] ), .Y(_abc_64468_n987) );
  OR2X2 OR2X2_1060 ( .A(u2__abc_44228_n6815_1), .B(u2__abc_44228_n6810), .Y(u2__abc_44228_n6816) );
  OR2X2 OR2X2_1061 ( .A(u2__abc_44228_n6808), .B(u2__abc_44228_n6816), .Y(u2__abc_44228_n6817) );
  OR2X2 OR2X2_1062 ( .A(u2__abc_44228_n6797_1), .B(u2__abc_44228_n6817), .Y(u2__abc_44228_n6818) );
  OR2X2 OR2X2_1063 ( .A(u2__abc_44228_n6820), .B(u2__abc_44228_n5665), .Y(u2__abc_44228_n6821) );
  OR2X2 OR2X2_1064 ( .A(u2__abc_44228_n6824), .B(u2__abc_44228_n6828), .Y(u2__abc_44228_n6829) );
  OR2X2 OR2X2_1065 ( .A(u2__abc_44228_n6836), .B(u2__abc_44228_n5633_1), .Y(u2__abc_44228_n6837) );
  OR2X2 OR2X2_1066 ( .A(u2__abc_44228_n6835), .B(u2__abc_44228_n6837), .Y(u2__abc_44228_n6838) );
  OR2X2 OR2X2_1067 ( .A(u2__abc_44228_n6830), .B(u2__abc_44228_n6838), .Y(u2__abc_44228_n6839) );
  OR2X2 OR2X2_1068 ( .A(u2__abc_44228_n6841), .B(u2__abc_44228_n5606_1), .Y(u2__abc_44228_n6842_1) );
  OR2X2 OR2X2_1069 ( .A(u2__abc_44228_n6845), .B(u2__abc_44228_n6849), .Y(u2__abc_44228_n6850) );
  OR2X2 OR2X2_107 ( .A(aNan_bF_buf0), .B(sqrto_129_), .Y(_abc_64468_n989) );
  OR2X2 OR2X2_1070 ( .A(u2__abc_44228_n6852), .B(u2__abc_44228_n5574), .Y(u2__abc_44228_n6853) );
  OR2X2 OR2X2_1071 ( .A(u2__abc_44228_n6858), .B(u2__abc_44228_n6853), .Y(u2__abc_44228_n6859) );
  OR2X2 OR2X2_1072 ( .A(u2__abc_44228_n6851_1), .B(u2__abc_44228_n6859), .Y(u2__abc_44228_n6860) );
  OR2X2 OR2X2_1073 ( .A(u2__abc_44228_n6840), .B(u2__abc_44228_n6860), .Y(u2__abc_44228_n6861_1) );
  OR2X2 OR2X2_1074 ( .A(u2__abc_44228_n6819), .B(u2__abc_44228_n6861_1), .Y(u2__abc_44228_n6862) );
  OR2X2 OR2X2_1075 ( .A(u2__abc_44228_n6778), .B(u2__abc_44228_n6862), .Y(u2__abc_44228_n6863) );
  OR2X2 OR2X2_1076 ( .A(u2__abc_44228_n6697), .B(u2__abc_44228_n6863), .Y(u2__abc_44228_n6864) );
  OR2X2 OR2X2_1077 ( .A(u2__abc_44228_n6532), .B(u2__abc_44228_n6864), .Y(u2__abc_44228_n6865) );
  OR2X2 OR2X2_1078 ( .A(u2__abc_44228_n6874), .B(u2__abc_44228_n6876), .Y(u2__abc_44228_n6877) );
  OR2X2 OR2X2_1079 ( .A(u2__abc_44228_n6888), .B(u2__abc_44228_n6890), .Y(u2__abc_44228_n6891) );
  OR2X2 OR2X2_108 ( .A(_abc_64468_n753_bF_buf10), .B(\a[53] ), .Y(_abc_64468_n990) );
  OR2X2 OR2X2_1080 ( .A(u2__abc_44228_n6903), .B(u2__abc_44228_n6905), .Y(u2__abc_44228_n6906_1) );
  OR2X2 OR2X2_1081 ( .A(u2__abc_44228_n6917), .B(u2__abc_44228_n6919), .Y(u2__abc_44228_n6920) );
  OR2X2 OR2X2_1082 ( .A(u2__abc_44228_n6933), .B(u2__abc_44228_n6935), .Y(u2__abc_44228_n6936) );
  OR2X2 OR2X2_1083 ( .A(u2__abc_44228_n6940), .B(u2__abc_44228_n6942), .Y(u2__abc_44228_n6943_1) );
  OR2X2 OR2X2_1084 ( .A(u2__abc_44228_n6962), .B(u2__abc_44228_n6964), .Y(u2__abc_44228_n6965) );
  OR2X2 OR2X2_1085 ( .A(u2__abc_44228_n6976), .B(u2__abc_44228_n6978), .Y(u2__abc_44228_n6979_1) );
  OR2X2 OR2X2_1086 ( .A(u2__abc_44228_n6993), .B(u2__abc_44228_n6995), .Y(u2__abc_44228_n6996) );
  OR2X2 OR2X2_1087 ( .A(u2__abc_44228_n7007_1), .B(u2__abc_44228_n7009), .Y(u2__abc_44228_n7010) );
  OR2X2 OR2X2_1088 ( .A(u2__abc_44228_n7022_1), .B(u2__abc_44228_n7024), .Y(u2__abc_44228_n7025) );
  OR2X2 OR2X2_1089 ( .A(u2__abc_44228_n7036), .B(u2__abc_44228_n7038), .Y(u2__abc_44228_n7039) );
  OR2X2 OR2X2_109 ( .A(aNan_bF_buf10), .B(sqrto_130_), .Y(_abc_64468_n992) );
  OR2X2 OR2X2_1090 ( .A(u2__abc_44228_n7052), .B(u2__abc_44228_n7054), .Y(u2__abc_44228_n7055) );
  OR2X2 OR2X2_1091 ( .A(u2__abc_44228_n7066), .B(u2__abc_44228_n7068_1), .Y(u2__abc_44228_n7069) );
  OR2X2 OR2X2_1092 ( .A(u2__abc_44228_n7081), .B(u2__abc_44228_n7083), .Y(u2__abc_44228_n7084) );
  OR2X2 OR2X2_1093 ( .A(u2__abc_44228_n7088_1), .B(u2__abc_44228_n7090), .Y(u2__abc_44228_n7091) );
  OR2X2 OR2X2_1094 ( .A(u2__abc_44228_n7113), .B(u2__abc_44228_n7115), .Y(u2__abc_44228_n7116_1) );
  OR2X2 OR2X2_1095 ( .A(u2__abc_44228_n7127), .B(u2__abc_44228_n7129), .Y(u2__abc_44228_n7130) );
  OR2X2 OR2X2_1096 ( .A(u2__abc_44228_n7142), .B(u2__abc_44228_n7144), .Y(u2__abc_44228_n7145) );
  OR2X2 OR2X2_1097 ( .A(u2__abc_44228_n7156), .B(u2__abc_44228_n7158), .Y(u2__abc_44228_n7159) );
  OR2X2 OR2X2_1098 ( .A(u2__abc_44228_n7172), .B(u2__abc_44228_n7174), .Y(u2__abc_44228_n7175) );
  OR2X2 OR2X2_1099 ( .A(u2__abc_44228_n7186), .B(u2__abc_44228_n7188), .Y(u2__abc_44228_n7189_1) );
  OR2X2 OR2X2_11 ( .A(aNan_bF_buf4), .B(sqrto_81_), .Y(_abc_64468_n845) );
  OR2X2 OR2X2_110 ( .A(_abc_64468_n753_bF_buf9), .B(\a[54] ), .Y(_abc_64468_n993) );
  OR2X2 OR2X2_1100 ( .A(u2__abc_44228_n7201), .B(u2__abc_44228_n7203), .Y(u2__abc_44228_n7204) );
  OR2X2 OR2X2_1101 ( .A(u2__abc_44228_n7208), .B(u2__abc_44228_n7210), .Y(u2__abc_44228_n7211) );
  OR2X2 OR2X2_1102 ( .A(u2__abc_44228_n7232), .B(u2__abc_44228_n7234_1), .Y(u2__abc_44228_n7235) );
  OR2X2 OR2X2_1103 ( .A(u2__abc_44228_n7239), .B(u2__abc_44228_n7241), .Y(u2__abc_44228_n7242) );
  OR2X2 OR2X2_1104 ( .A(u2__abc_44228_n7261), .B(u2__abc_44228_n7263), .Y(u2__abc_44228_n7264) );
  OR2X2 OR2X2_1105 ( .A(u2__abc_44228_n7268), .B(u2__abc_44228_n7270), .Y(u2__abc_44228_n7271_1) );
  OR2X2 OR2X2_1106 ( .A(u2__abc_44228_n7291), .B(u2__abc_44228_n7293), .Y(u2__abc_44228_n7294) );
  OR2X2 OR2X2_1107 ( .A(u2__abc_44228_n7298), .B(u2__abc_44228_n7300), .Y(u2__abc_44228_n7301) );
  OR2X2 OR2X2_1108 ( .A(u2__abc_44228_n7320), .B(u2__abc_44228_n7322), .Y(u2__abc_44228_n7323) );
  OR2X2 OR2X2_1109 ( .A(u2__abc_44228_n7334), .B(u2__abc_44228_n7336), .Y(u2__abc_44228_n7337_1) );
  OR2X2 OR2X2_111 ( .A(aNan_bF_buf9), .B(sqrto_131_), .Y(_abc_64468_n995) );
  OR2X2 OR2X2_1110 ( .A(u2__abc_44228_n7346_1), .B(u2__abc_44228_n7330), .Y(u2__abc_44228_n7347) );
  OR2X2 OR2X2_1111 ( .A(u2__abc_44228_n7351), .B(u2__abc_44228_n7313), .Y(u2__abc_44228_n7352) );
  OR2X2 OR2X2_1112 ( .A(u2__abc_44228_n7350), .B(u2__abc_44228_n7352), .Y(u2__abc_44228_n7353) );
  OR2X2 OR2X2_1113 ( .A(u2__abc_44228_n7360), .B(u2__abc_44228_n7284), .Y(u2__abc_44228_n7361) );
  OR2X2 OR2X2_1114 ( .A(u2__abc_44228_n7359), .B(u2__abc_44228_n7361), .Y(u2__abc_44228_n7362) );
  OR2X2 OR2X2_1115 ( .A(u2__abc_44228_n7354), .B(u2__abc_44228_n7362), .Y(u2__abc_44228_n7363) );
  OR2X2 OR2X2_1116 ( .A(u2__abc_44228_n7370), .B(u2__abc_44228_n7254), .Y(u2__abc_44228_n7371) );
  OR2X2 OR2X2_1117 ( .A(u2__abc_44228_n7369), .B(u2__abc_44228_n7371), .Y(u2__abc_44228_n7372) );
  OR2X2 OR2X2_1118 ( .A(u2__abc_44228_n7374_1), .B(u2__abc_44228_n7225_1), .Y(u2__abc_44228_n7375) );
  OR2X2 OR2X2_1119 ( .A(u2__abc_44228_n7380), .B(u2__abc_44228_n7375), .Y(u2__abc_44228_n7381) );
  OR2X2 OR2X2_112 ( .A(_abc_64468_n753_bF_buf8), .B(\a[55] ), .Y(_abc_64468_n996) );
  OR2X2 OR2X2_1120 ( .A(u2__abc_44228_n7373), .B(u2__abc_44228_n7381), .Y(u2__abc_44228_n7382_1) );
  OR2X2 OR2X2_1121 ( .A(u2__abc_44228_n7364_1), .B(u2__abc_44228_n7382_1), .Y(u2__abc_44228_n7383) );
  OR2X2 OR2X2_1122 ( .A(u2__abc_44228_n7390), .B(u2__abc_44228_n7194), .Y(u2__abc_44228_n7391) );
  OR2X2 OR2X2_1123 ( .A(u2__abc_44228_n7389), .B(u2__abc_44228_n7391), .Y(u2__abc_44228_n7392_1) );
  OR2X2 OR2X2_1124 ( .A(u2__abc_44228_n7394), .B(u2__abc_44228_n7182), .Y(u2__abc_44228_n7395) );
  OR2X2 OR2X2_1125 ( .A(u2__abc_44228_n7399), .B(u2__abc_44228_n7165), .Y(u2__abc_44228_n7400_1) );
  OR2X2 OR2X2_1126 ( .A(u2__abc_44228_n7398), .B(u2__abc_44228_n7400_1), .Y(u2__abc_44228_n7401) );
  OR2X2 OR2X2_1127 ( .A(u2__abc_44228_n7393), .B(u2__abc_44228_n7401), .Y(u2__abc_44228_n7402) );
  OR2X2 OR2X2_1128 ( .A(u2__abc_44228_n7135), .B(u2__abc_44228_n7142), .Y(u2__abc_44228_n7404) );
  OR2X2 OR2X2_1129 ( .A(u2__abc_44228_n7410_1), .B(u2__abc_44228_n7405), .Y(u2__abc_44228_n7411) );
  OR2X2 OR2X2_113 ( .A(aNan_bF_buf8), .B(sqrto_132_), .Y(_abc_64468_n998) );
  OR2X2 OR2X2_1130 ( .A(u2__abc_44228_n7418), .B(u2__abc_44228_n7106_1), .Y(u2__abc_44228_n7419_1) );
  OR2X2 OR2X2_1131 ( .A(u2__abc_44228_n7417), .B(u2__abc_44228_n7419_1), .Y(u2__abc_44228_n7420) );
  OR2X2 OR2X2_1132 ( .A(u2__abc_44228_n7412), .B(u2__abc_44228_n7420), .Y(u2__abc_44228_n7421) );
  OR2X2 OR2X2_1133 ( .A(u2__abc_44228_n7403), .B(u2__abc_44228_n7421), .Y(u2__abc_44228_n7422) );
  OR2X2 OR2X2_1134 ( .A(u2__abc_44228_n7384), .B(u2__abc_44228_n7422), .Y(u2__abc_44228_n7423) );
  OR2X2 OR2X2_1135 ( .A(u2__abc_44228_n7430), .B(u2__abc_44228_n7074), .Y(u2__abc_44228_n7431) );
  OR2X2 OR2X2_1136 ( .A(u2__abc_44228_n7429), .B(u2__abc_44228_n7431), .Y(u2__abc_44228_n7432) );
  OR2X2 OR2X2_1137 ( .A(u2__abc_44228_n7434), .B(u2__abc_44228_n7062), .Y(u2__abc_44228_n7435) );
  OR2X2 OR2X2_1138 ( .A(u2__abc_44228_n7439), .B(u2__abc_44228_n7045), .Y(u2__abc_44228_n7440) );
  OR2X2 OR2X2_1139 ( .A(u2__abc_44228_n7438), .B(u2__abc_44228_n7440), .Y(u2__abc_44228_n7441) );
  OR2X2 OR2X2_114 ( .A(_abc_64468_n753_bF_buf7), .B(\a[56] ), .Y(_abc_64468_n999) );
  OR2X2 OR2X2_1140 ( .A(u2__abc_44228_n7433), .B(u2__abc_44228_n7441), .Y(u2__abc_44228_n7442) );
  OR2X2 OR2X2_1141 ( .A(u2__abc_44228_n7444), .B(u2__abc_44228_n7032_1), .Y(u2__abc_44228_n7445) );
  OR2X2 OR2X2_1142 ( .A(u2__abc_44228_n7448), .B(u2__abc_44228_n7452), .Y(u2__abc_44228_n7453) );
  OR2X2 OR2X2_1143 ( .A(u2__abc_44228_n7455_1), .B(u2__abc_44228_n6986), .Y(u2__abc_44228_n7456) );
  OR2X2 OR2X2_1144 ( .A(u2__abc_44228_n7461), .B(u2__abc_44228_n7456), .Y(u2__abc_44228_n7462) );
  OR2X2 OR2X2_1145 ( .A(u2__abc_44228_n7454), .B(u2__abc_44228_n7462), .Y(u2__abc_44228_n7463) );
  OR2X2 OR2X2_1146 ( .A(u2__abc_44228_n7443), .B(u2__abc_44228_n7463), .Y(u2__abc_44228_n7464_1) );
  OR2X2 OR2X2_1147 ( .A(u2__abc_44228_n7466), .B(u2__abc_44228_n6958), .Y(u2__abc_44228_n7467) );
  OR2X2 OR2X2_1148 ( .A(u2__abc_44228_n7470), .B(u2__abc_44228_n7474), .Y(u2__abc_44228_n7475) );
  OR2X2 OR2X2_1149 ( .A(u2__abc_44228_n7482), .B(u2__abc_44228_n6926), .Y(u2__abc_44228_n7483_1) );
  OR2X2 OR2X2_115 ( .A(aNan_bF_buf7), .B(sqrto_133_), .Y(_abc_64468_n1001) );
  OR2X2 OR2X2_1150 ( .A(u2__abc_44228_n7481), .B(u2__abc_44228_n7483_1), .Y(u2__abc_44228_n7484) );
  OR2X2 OR2X2_1151 ( .A(u2__abc_44228_n7476), .B(u2__abc_44228_n7484), .Y(u2__abc_44228_n7485) );
  OR2X2 OR2X2_1152 ( .A(u2__abc_44228_n6896), .B(u2__abc_44228_n6903), .Y(u2__abc_44228_n7487) );
  OR2X2 OR2X2_1153 ( .A(u2__abc_44228_n7493_1), .B(u2__abc_44228_n7488), .Y(u2__abc_44228_n7494) );
  OR2X2 OR2X2_1154 ( .A(u2__abc_44228_n7496), .B(u2__abc_44228_n6884), .Y(u2__abc_44228_n7497) );
  OR2X2 OR2X2_1155 ( .A(u2__abc_44228_n7501), .B(u2__abc_44228_n6867), .Y(u2__abc_44228_n7502_1) );
  OR2X2 OR2X2_1156 ( .A(u2__abc_44228_n7500), .B(u2__abc_44228_n7502_1), .Y(u2__abc_44228_n7503) );
  OR2X2 OR2X2_1157 ( .A(u2__abc_44228_n7495), .B(u2__abc_44228_n7503), .Y(u2__abc_44228_n7504) );
  OR2X2 OR2X2_1158 ( .A(u2__abc_44228_n7486), .B(u2__abc_44228_n7504), .Y(u2__abc_44228_n7505) );
  OR2X2 OR2X2_1159 ( .A(u2__abc_44228_n7465), .B(u2__abc_44228_n7505), .Y(u2__abc_44228_n7506) );
  OR2X2 OR2X2_116 ( .A(_abc_64468_n753_bF_buf6), .B(\a[57] ), .Y(_abc_64468_n1002) );
  OR2X2 OR2X2_1160 ( .A(u2__abc_44228_n7424), .B(u2__abc_44228_n7506), .Y(u2__abc_44228_n7507) );
  OR2X2 OR2X2_1161 ( .A(u2__abc_44228_n7345), .B(u2__abc_44228_n7507), .Y(u2__abc_44228_n7508) );
  OR2X2 OR2X2_1162 ( .A(u2__abc_44228_n7517), .B(u2__abc_44228_n7519), .Y(u2__abc_44228_n7520) );
  OR2X2 OR2X2_1163 ( .A(u2__abc_44228_n7524), .B(u2__abc_44228_n7526), .Y(u2__abc_44228_n7527) );
  OR2X2 OR2X2_1164 ( .A(u2__abc_44228_n7540_1), .B(u2__abc_44228_n7533), .Y(u2__abc_44228_n7541) );
  OR2X2 OR2X2_1165 ( .A(u2__abc_44228_n7544), .B(u2__abc_44228_n7510), .Y(u2__abc_44228_n7545) );
  OR2X2 OR2X2_1166 ( .A(u2__abc_44228_n7543), .B(u2__abc_44228_n7545), .Y(u2__abc_44228_n7546) );
  OR2X2 OR2X2_1167 ( .A(u2__abc_44228_n7538), .B(u2__abc_44228_n7546), .Y(u2__abc_44228_n7547) );
  OR2X2 OR2X2_1168 ( .A(u2__abc_44228_n7551), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n7552) );
  OR2X2 OR2X2_1169 ( .A(u2__abc_44228_n7552), .B(u2__abc_44228_n7549), .Y(u2__abc_44228_n7553) );
  OR2X2 OR2X2_117 ( .A(aNan_bF_buf6), .B(sqrto_134_), .Y(_abc_64468_n1004) );
  OR2X2 OR2X2_1170 ( .A(u2__abc_44228_n7558_1), .B(u2__abc_44228_n3063), .Y(u2__abc_44228_n7559) );
  OR2X2 OR2X2_1171 ( .A(u2__abc_44228_n3069), .B(u2_remHiShift_0_), .Y(u2__abc_44228_n7563) );
  OR2X2 OR2X2_1172 ( .A(u2__abc_44228_n7566), .B(u2__abc_44228_n7565), .Y(u2__abc_44228_n7567_1) );
  OR2X2 OR2X2_1173 ( .A(u2__abc_44228_n7567_1), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n7568) );
  OR2X2 OR2X2_1174 ( .A(u2__abc_44228_n7572), .B(u2__abc_44228_n7561), .Y(u2__abc_44228_n7573) );
  OR2X2 OR2X2_1175 ( .A(u2__abc_44228_n3071), .B(u2__abc_44228_n3081), .Y(u2__abc_44228_n7578) );
  OR2X2 OR2X2_1176 ( .A(u2__abc_44228_n7581), .B(u2__abc_44228_n7580), .Y(u2__abc_44228_n7582) );
  OR2X2 OR2X2_1177 ( .A(u2__abc_44228_n7582), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n7583) );
  OR2X2 OR2X2_1178 ( .A(u2__abc_44228_n7588), .B(u2__abc_44228_n7575), .Y(u2__abc_44228_n7589) );
  OR2X2 OR2X2_1179 ( .A(u2__abc_44228_n7593), .B(u2__abc_44228_n3076), .Y(u2__abc_44228_n7594) );
  OR2X2 OR2X2_118 ( .A(_abc_64468_n753_bF_buf5), .B(\a[58] ), .Y(_abc_64468_n1005) );
  OR2X2 OR2X2_1180 ( .A(u2__abc_44228_n7592), .B(u2__abc_44228_n7595), .Y(u2__abc_44228_n7596) );
  OR2X2 OR2X2_1181 ( .A(u2__abc_44228_n7599), .B(u2__abc_44228_n7598), .Y(u2__abc_44228_n7600) );
  OR2X2 OR2X2_1182 ( .A(u2__abc_44228_n7600), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n7601) );
  OR2X2 OR2X2_1183 ( .A(u2__abc_44228_n7606), .B(u2__abc_44228_n7591), .Y(u2__abc_44228_n7607) );
  OR2X2 OR2X2_1184 ( .A(u2__abc_44228_n3087), .B(u2__abc_44228_n3108), .Y(u2__abc_44228_n7610) );
  OR2X2 OR2X2_1185 ( .A(u2__abc_44228_n7615_1), .B(u2__abc_44228_n7614), .Y(u2__abc_44228_n7616_1) );
  OR2X2 OR2X2_1186 ( .A(u2__abc_44228_n7616_1), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n7617) );
  OR2X2 OR2X2_1187 ( .A(u2__abc_44228_n7621), .B(u2__abc_44228_n7609), .Y(u2__abc_44228_n7622_1) );
  OR2X2 OR2X2_1188 ( .A(u2__abc_44228_n7626), .B(u2__abc_44228_n7625), .Y(u2__abc_44228_n7627) );
  OR2X2 OR2X2_1189 ( .A(u2__abc_44228_n7628), .B(u2__abc_44228_n3103), .Y(u2__abc_44228_n7629_1) );
  OR2X2 OR2X2_119 ( .A(aNan_bF_buf5), .B(sqrto_135_), .Y(_abc_64468_n1007) );
  OR2X2 OR2X2_1190 ( .A(u2__abc_44228_n7632), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n7633) );
  OR2X2 OR2X2_1191 ( .A(u2__abc_44228_n7633), .B(u2__abc_44228_n7631), .Y(u2__abc_44228_n7634) );
  OR2X2 OR2X2_1192 ( .A(u2__abc_44228_n7638), .B(u2__abc_44228_n7624), .Y(u2__abc_44228_n7639) );
  OR2X2 OR2X2_1193 ( .A(u2__abc_44228_n7642), .B(u2__abc_44228_n3113), .Y(u2__abc_44228_n7643_1) );
  OR2X2 OR2X2_1194 ( .A(u2__abc_44228_n7643_1), .B(u2__abc_44228_n3097), .Y(u2__abc_44228_n7646) );
  OR2X2 OR2X2_1195 ( .A(u2__abc_44228_n7649), .B(u2__abc_44228_n7648), .Y(u2__abc_44228_n7650_1) );
  OR2X2 OR2X2_1196 ( .A(u2__abc_44228_n7650_1), .B(u2__abc_44228_n2983_bF_buf127), .Y(u2__abc_44228_n7651_1) );
  OR2X2 OR2X2_1197 ( .A(u2__abc_44228_n7655), .B(u2__abc_44228_n7641), .Y(u2__abc_44228_n7656) );
  OR2X2 OR2X2_1198 ( .A(u2__abc_44228_n7660), .B(u2__abc_44228_n3092), .Y(u2__abc_44228_n7661) );
  OR2X2 OR2X2_1199 ( .A(u2__abc_44228_n7659), .B(u2__abc_44228_n7662), .Y(u2__abc_44228_n7663) );
  OR2X2 OR2X2_12 ( .A(_abc_64468_n753_bF_buf2), .B(\a[5] ), .Y(_abc_64468_n846) );
  OR2X2 OR2X2_120 ( .A(_abc_64468_n753_bF_buf4), .B(\a[59] ), .Y(_abc_64468_n1008) );
  OR2X2 OR2X2_1200 ( .A(u2__abc_44228_n7666), .B(u2__abc_44228_n7665_1), .Y(u2__abc_44228_n7667) );
  OR2X2 OR2X2_1201 ( .A(u2__abc_44228_n7667), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n7668) );
  OR2X2 OR2X2_1202 ( .A(u2__abc_44228_n7672_1), .B(u2__abc_44228_n7658_1), .Y(u2__abc_44228_n7673) );
  OR2X2 OR2X2_1203 ( .A(u2__abc_44228_n3120), .B(u2__abc_44228_n3166), .Y(u2__abc_44228_n7678_1) );
  OR2X2 OR2X2_1204 ( .A(u2__abc_44228_n7681), .B(u2__abc_44228_n7680), .Y(u2__abc_44228_n7682) );
  OR2X2 OR2X2_1205 ( .A(u2__abc_44228_n7682), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n7683) );
  OR2X2 OR2X2_1206 ( .A(u2__abc_44228_n7687), .B(u2__abc_44228_n7675), .Y(u2__abc_44228_n7688) );
  OR2X2 OR2X2_1207 ( .A(u2__abc_44228_n7676), .B(u2__abc_44228_n3162), .Y(u2__abc_44228_n7692_1) );
  OR2X2 OR2X2_1208 ( .A(u2__abc_44228_n7695), .B(u2__abc_44228_n7693_1), .Y(u2__abc_44228_n7696) );
  OR2X2 OR2X2_1209 ( .A(u2__abc_44228_n7698), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n7699_1) );
  OR2X2 OR2X2_121 ( .A(aNan_bF_buf4), .B(sqrto_136_), .Y(_abc_64468_n1010) );
  OR2X2 OR2X2_1210 ( .A(u2__abc_44228_n7699_1), .B(u2__abc_44228_n7697), .Y(u2__abc_44228_n7700_1) );
  OR2X2 OR2X2_1211 ( .A(u2__abc_44228_n7704), .B(u2__abc_44228_n7690), .Y(u2__abc_44228_n7705) );
  OR2X2 OR2X2_1212 ( .A(u2__abc_44228_n7708), .B(u2__abc_44228_n3179), .Y(u2__abc_44228_n7709) );
  OR2X2 OR2X2_1213 ( .A(u2__abc_44228_n7709), .B(u2__abc_44228_n3159), .Y(u2__abc_44228_n7710) );
  OR2X2 OR2X2_1214 ( .A(u2__abc_44228_n7715), .B(u2__abc_44228_n7714_1), .Y(u2__abc_44228_n7716) );
  OR2X2 OR2X2_1215 ( .A(u2__abc_44228_n7716), .B(u2__abc_44228_n2983_bF_buf119), .Y(u2__abc_44228_n7717) );
  OR2X2 OR2X2_1216 ( .A(u2__abc_44228_n7721_1), .B(u2__abc_44228_n7707_1), .Y(u2__abc_44228_n7722) );
  OR2X2 OR2X2_1217 ( .A(u2__abc_44228_n7726), .B(u2__abc_44228_n3154), .Y(u2__abc_44228_n7727_1) );
  OR2X2 OR2X2_1218 ( .A(u2__abc_44228_n7725), .B(u2__abc_44228_n7728_1), .Y(u2__abc_44228_n7729) );
  OR2X2 OR2X2_1219 ( .A(u2__abc_44228_n7732), .B(u2__abc_44228_n7731), .Y(u2__abc_44228_n7733) );
  OR2X2 OR2X2_122 ( .A(_abc_64468_n753_bF_buf3), .B(\a[60] ), .Y(_abc_64468_n1011) );
  OR2X2 OR2X2_1220 ( .A(u2__abc_44228_n7733), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n7734_1) );
  OR2X2 OR2X2_1221 ( .A(u2__abc_44228_n7738), .B(u2__abc_44228_n7724), .Y(u2__abc_44228_n7739) );
  OR2X2 OR2X2_1222 ( .A(u2__abc_44228_n7742_1), .B(u2__abc_44228_n3185), .Y(u2__abc_44228_n7743) );
  OR2X2 OR2X2_1223 ( .A(u2__abc_44228_n7743), .B(u2__abc_44228_n3147), .Y(u2__abc_44228_n7746) );
  OR2X2 OR2X2_1224 ( .A(u2__abc_44228_n7749_1), .B(u2__abc_44228_n7748_1), .Y(u2__abc_44228_n7750) );
  OR2X2 OR2X2_1225 ( .A(u2__abc_44228_n7750), .B(u2__abc_44228_n2983_bF_buf115), .Y(u2__abc_44228_n7751) );
  OR2X2 OR2X2_1226 ( .A(u2__abc_44228_n7755_1), .B(u2__abc_44228_n7741_1), .Y(u2__abc_44228_n7756_1) );
  OR2X2 OR2X2_1227 ( .A(u2__abc_44228_n7744), .B(u2__abc_44228_n3143), .Y(u2__abc_44228_n7759) );
  OR2X2 OR2X2_1228 ( .A(u2__abc_44228_n7759), .B(u2__abc_44228_n3141), .Y(u2__abc_44228_n7760) );
  OR2X2 OR2X2_1229 ( .A(u2__abc_44228_n7762_1), .B(u2__abc_44228_n7761), .Y(u2__abc_44228_n7763_1) );
  OR2X2 OR2X2_123 ( .A(aNan_bF_buf3), .B(sqrto_137_), .Y(_abc_64468_n1013) );
  OR2X2 OR2X2_1230 ( .A(u2__abc_44228_n7766), .B(u2__abc_44228_n7765), .Y(u2__abc_44228_n7767) );
  OR2X2 OR2X2_1231 ( .A(u2__abc_44228_n7767), .B(u2__abc_44228_n2983_bF_buf113), .Y(u2__abc_44228_n7768) );
  OR2X2 OR2X2_1232 ( .A(u2__abc_44228_n7772), .B(u2__abc_44228_n7758), .Y(u2__abc_44228_n7773) );
  OR2X2 OR2X2_1233 ( .A(u2__abc_44228_n7776_1), .B(u2__abc_44228_n3188), .Y(u2__abc_44228_n7777_1) );
  OR2X2 OR2X2_1234 ( .A(u2__abc_44228_n7777_1), .B(u2__abc_44228_n3133), .Y(u2__abc_44228_n7778) );
  OR2X2 OR2X2_1235 ( .A(u2__abc_44228_n7783_1), .B(u2__abc_44228_n7782), .Y(u2__abc_44228_n7784_1) );
  OR2X2 OR2X2_1236 ( .A(u2__abc_44228_n7784_1), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n7785) );
  OR2X2 OR2X2_1237 ( .A(u2__abc_44228_n7789), .B(u2__abc_44228_n7775), .Y(u2__abc_44228_n7790_1) );
  OR2X2 OR2X2_1238 ( .A(u2__abc_44228_n7779), .B(u2__abc_44228_n3129), .Y(u2__abc_44228_n7794) );
  OR2X2 OR2X2_1239 ( .A(u2__abc_44228_n7795), .B(u2__abc_44228_n7793), .Y(u2__abc_44228_n7796) );
  OR2X2 OR2X2_124 ( .A(_abc_64468_n753_bF_buf2), .B(\a[61] ), .Y(_abc_64468_n1014) );
  OR2X2 OR2X2_1240 ( .A(u2__abc_44228_n7794), .B(u2__abc_44228_n3127), .Y(u2__abc_44228_n7797_1) );
  OR2X2 OR2X2_1241 ( .A(u2__abc_44228_n7800), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n7801) );
  OR2X2 OR2X2_1242 ( .A(u2__abc_44228_n7801), .B(u2__abc_44228_n7799), .Y(u2__abc_44228_n7802) );
  OR2X2 OR2X2_1243 ( .A(u2__abc_44228_n7806), .B(u2__abc_44228_n7792), .Y(u2__abc_44228_n7807) );
  OR2X2 OR2X2_1244 ( .A(u2__abc_44228_n3194), .B(u2__abc_44228_n3306), .Y(u2__abc_44228_n7810) );
  OR2X2 OR2X2_1245 ( .A(u2__abc_44228_n7815), .B(u2__abc_44228_n7814), .Y(u2__abc_44228_n7816) );
  OR2X2 OR2X2_1246 ( .A(u2__abc_44228_n7816), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n7817) );
  OR2X2 OR2X2_1247 ( .A(u2__abc_44228_n7821), .B(u2__abc_44228_n7809), .Y(u2__abc_44228_n7822) );
  OR2X2 OR2X2_1248 ( .A(u2__abc_44228_n7811_1), .B(u2__abc_44228_n3302), .Y(u2__abc_44228_n7825_1) );
  OR2X2 OR2X2_1249 ( .A(u2__abc_44228_n7825_1), .B(u2__abc_44228_n3300), .Y(u2__abc_44228_n7826_1) );
  OR2X2 OR2X2_125 ( .A(aNan_bF_buf2), .B(sqrto_138_), .Y(_abc_64468_n1016) );
  OR2X2 OR2X2_1250 ( .A(u2__abc_44228_n7828), .B(u2__abc_44228_n7827), .Y(u2__abc_44228_n7829) );
  OR2X2 OR2X2_1251 ( .A(u2__abc_44228_n7832_1), .B(u2__abc_44228_n7831), .Y(u2__abc_44228_n7833_1) );
  OR2X2 OR2X2_1252 ( .A(u2__abc_44228_n7833_1), .B(u2__abc_44228_n2983_bF_buf105), .Y(u2__abc_44228_n7834) );
  OR2X2 OR2X2_1253 ( .A(u2__abc_44228_n7838), .B(u2__abc_44228_n7824), .Y(u2__abc_44228_n7839_1) );
  OR2X2 OR2X2_1254 ( .A(u2__abc_44228_n7842), .B(u2__abc_44228_n3313), .Y(u2__abc_44228_n7843) );
  OR2X2 OR2X2_1255 ( .A(u2__abc_44228_n7843), .B(u2__abc_44228_n3292), .Y(u2__abc_44228_n7844) );
  OR2X2 OR2X2_1256 ( .A(u2__abc_44228_n7849), .B(u2__abc_44228_n7848), .Y(u2__abc_44228_n7850_1) );
  OR2X2 OR2X2_1257 ( .A(u2__abc_44228_n7850_1), .B(u2__abc_44228_n2983_bF_buf103), .Y(u2__abc_44228_n7851_1) );
  OR2X2 OR2X2_1258 ( .A(u2__abc_44228_n7855), .B(u2__abc_44228_n7841), .Y(u2__abc_44228_n7856_1) );
  OR2X2 OR2X2_1259 ( .A(u2__abc_44228_n7860), .B(u2__abc_44228_n3287), .Y(u2__abc_44228_n7861_1) );
  OR2X2 OR2X2_126 ( .A(_abc_64468_n753_bF_buf1), .B(\a[62] ), .Y(_abc_64468_n1017) );
  OR2X2 OR2X2_1260 ( .A(u2__abc_44228_n7859), .B(u2__abc_44228_n7862_1), .Y(u2__abc_44228_n7863) );
  OR2X2 OR2X2_1261 ( .A(u2__abc_44228_n7866), .B(u2__abc_44228_n7865), .Y(u2__abc_44228_n7867_1) );
  OR2X2 OR2X2_1262 ( .A(u2__abc_44228_n7867_1), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n7868) );
  OR2X2 OR2X2_1263 ( .A(u2__abc_44228_n7872_1), .B(u2__abc_44228_n7858), .Y(u2__abc_44228_n7873_1) );
  OR2X2 OR2X2_1264 ( .A(u2__abc_44228_n7876), .B(u2__abc_44228_n3319), .Y(u2__abc_44228_n7877) );
  OR2X2 OR2X2_1265 ( .A(u2__abc_44228_n7877), .B(u2__abc_44228_n3273), .Y(u2__abc_44228_n7880) );
  OR2X2 OR2X2_1266 ( .A(u2__abc_44228_n7883_1), .B(u2__abc_44228_n7882), .Y(u2__abc_44228_n7884_1) );
  OR2X2 OR2X2_1267 ( .A(u2__abc_44228_n7884_1), .B(u2__abc_44228_n2983_bF_buf99), .Y(u2__abc_44228_n7885) );
  OR2X2 OR2X2_1268 ( .A(u2__abc_44228_n7889_1), .B(u2__abc_44228_n7875), .Y(u2__abc_44228_n7890) );
  OR2X2 OR2X2_1269 ( .A(u2__abc_44228_n7878_1), .B(u2__abc_44228_n3269), .Y(u2__abc_44228_n7894_1) );
  OR2X2 OR2X2_127 ( .A(aNan_bF_buf1), .B(sqrto_139_), .Y(_abc_64468_n1019) );
  OR2X2 OR2X2_1270 ( .A(u2__abc_44228_n7897), .B(u2__abc_44228_n7895_1), .Y(u2__abc_44228_n7898) );
  OR2X2 OR2X2_1271 ( .A(u2__abc_44228_n7900_1), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n7901) );
  OR2X2 OR2X2_1272 ( .A(u2__abc_44228_n7901), .B(u2__abc_44228_n7899), .Y(u2__abc_44228_n7902) );
  OR2X2 OR2X2_1273 ( .A(u2__abc_44228_n7906_1), .B(u2__abc_44228_n7892), .Y(u2__abc_44228_n7907) );
  OR2X2 OR2X2_1274 ( .A(u2__abc_44228_n7910), .B(u2__abc_44228_n3322), .Y(u2__abc_44228_n7911_1) );
  OR2X2 OR2X2_1275 ( .A(u2__abc_44228_n7911_1), .B(u2__abc_44228_n3266), .Y(u2__abc_44228_n7912) );
  OR2X2 OR2X2_1276 ( .A(u2__abc_44228_n7917_1), .B(u2__abc_44228_n7916_1), .Y(u2__abc_44228_n7918) );
  OR2X2 OR2X2_1277 ( .A(u2__abc_44228_n7918), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n7919) );
  OR2X2 OR2X2_1278 ( .A(u2__abc_44228_n7923), .B(u2__abc_44228_n7909), .Y(u2__abc_44228_n7924) );
  OR2X2 OR2X2_1279 ( .A(u2__abc_44228_n7913), .B(u2__abc_44228_n3262), .Y(u2__abc_44228_n7928_1) );
  OR2X2 OR2X2_128 ( .A(_abc_64468_n753_bF_buf0), .B(\a[63] ), .Y(_abc_64468_n1020) );
  OR2X2 OR2X2_1280 ( .A(u2__abc_44228_n7931), .B(u2__abc_44228_n7929), .Y(u2__abc_44228_n7932) );
  OR2X2 OR2X2_1281 ( .A(u2__abc_44228_n7934), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n7935) );
  OR2X2 OR2X2_1282 ( .A(u2__abc_44228_n7935), .B(u2__abc_44228_n7933_1), .Y(u2__abc_44228_n7936) );
  OR2X2 OR2X2_1283 ( .A(u2__abc_44228_n7940), .B(u2__abc_44228_n7926), .Y(u2__abc_44228_n7941) );
  OR2X2 OR2X2_1284 ( .A(u2__abc_44228_n7944_1), .B(u2__abc_44228_n3327), .Y(u2__abc_44228_n7945) );
  OR2X2 OR2X2_1285 ( .A(u2__abc_44228_n7945), .B(u2__abc_44228_n3236), .Y(u2__abc_44228_n7946) );
  OR2X2 OR2X2_1286 ( .A(u2__abc_44228_n7951), .B(u2__abc_44228_n7950_1), .Y(u2__abc_44228_n7952) );
  OR2X2 OR2X2_1287 ( .A(u2__abc_44228_n7952), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n7953) );
  OR2X2 OR2X2_1288 ( .A(u2__abc_44228_n7957), .B(u2__abc_44228_n7943), .Y(u2__abc_44228_n7958) );
  OR2X2 OR2X2_1289 ( .A(u2__abc_44228_n7947), .B(u2__abc_44228_n3232), .Y(u2__abc_44228_n7962) );
  OR2X2 OR2X2_129 ( .A(aNan_bF_buf0), .B(sqrto_140_), .Y(_abc_64468_n1022) );
  OR2X2 OR2X2_1290 ( .A(u2__abc_44228_n7963), .B(u2__abc_44228_n7961_1), .Y(u2__abc_44228_n7964) );
  OR2X2 OR2X2_1291 ( .A(u2__abc_44228_n7962), .B(u2__abc_44228_n3230), .Y(u2__abc_44228_n7965) );
  OR2X2 OR2X2_1292 ( .A(u2__abc_44228_n7968), .B(u2__abc_44228_n2983_bF_buf89), .Y(u2__abc_44228_n7969) );
  OR2X2 OR2X2_1293 ( .A(u2__abc_44228_n7969), .B(u2__abc_44228_n7967), .Y(u2__abc_44228_n7970) );
  OR2X2 OR2X2_1294 ( .A(u2__abc_44228_n7974), .B(u2__abc_44228_n7960_1), .Y(u2__abc_44228_n7975) );
  OR2X2 OR2X2_1295 ( .A(u2__abc_44228_n7978), .B(u2__abc_44228_n3330), .Y(u2__abc_44228_n7979) );
  OR2X2 OR2X2_1296 ( .A(u2__abc_44228_n7979), .B(u2__abc_44228_n3250), .Y(u2__abc_44228_n7980) );
  OR2X2 OR2X2_1297 ( .A(u2__abc_44228_n7985), .B(u2__abc_44228_n7984), .Y(u2__abc_44228_n7986) );
  OR2X2 OR2X2_1298 ( .A(u2__abc_44228_n7986), .B(u2__abc_44228_n2983_bF_buf87), .Y(u2__abc_44228_n7987) );
  OR2X2 OR2X2_1299 ( .A(u2__abc_44228_n7991), .B(u2__abc_44228_n7977_1), .Y(u2__abc_44228_n7992) );
  OR2X2 OR2X2_13 ( .A(aNan_bF_buf3), .B(sqrto_82_), .Y(_abc_64468_n848) );
  OR2X2 OR2X2_130 ( .A(_abc_64468_n753_bF_buf13), .B(\a[64] ), .Y(_abc_64468_n1023) );
  OR2X2 OR2X2_1300 ( .A(u2__abc_44228_n7996), .B(u2__abc_44228_n3244), .Y(u2__abc_44228_n7997) );
  OR2X2 OR2X2_1301 ( .A(u2__abc_44228_n7995), .B(u2__abc_44228_n7998), .Y(u2__abc_44228_n7999_1) );
  OR2X2 OR2X2_1302 ( .A(u2__abc_44228_n8002), .B(u2__abc_44228_n8001), .Y(u2__abc_44228_n8003) );
  OR2X2 OR2X2_1303 ( .A(u2__abc_44228_n8003), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n8004_1) );
  OR2X2 OR2X2_1304 ( .A(u2__abc_44228_n8008), .B(u2__abc_44228_n7994_1), .Y(u2__abc_44228_n8009) );
  OR2X2 OR2X2_1305 ( .A(u2__abc_44228_n8013), .B(u2__abc_44228_n3242), .Y(u2__abc_44228_n8014) );
  OR2X2 OR2X2_1306 ( .A(u2__abc_44228_n8015_1), .B(u2__abc_44228_n3214), .Y(u2__abc_44228_n8018) );
  OR2X2 OR2X2_1307 ( .A(u2__abc_44228_n8020), .B(u2__abc_44228_n2983_bF_buf83), .Y(u2__abc_44228_n8021_1) );
  OR2X2 OR2X2_1308 ( .A(u2__abc_44228_n8021_1), .B(u2__abc_44228_n8012), .Y(u2__abc_44228_n8022) );
  OR2X2 OR2X2_1309 ( .A(u2__abc_44228_n8026_1), .B(u2__abc_44228_n8011), .Y(u2__abc_44228_n8027_1) );
  OR2X2 OR2X2_131 ( .A(aNan_bF_buf10), .B(sqrto_141_), .Y(_abc_64468_n1025) );
  OR2X2 OR2X2_1310 ( .A(u2__abc_44228_n7547_bF_buf27), .B(u2_remHi_27_), .Y(u2__abc_44228_n8030) );
  OR2X2 OR2X2_1311 ( .A(u2__abc_44228_n8034), .B(u2__abc_44228_n8035), .Y(u2__abc_44228_n8036) );
  OR2X2 OR2X2_1312 ( .A(u2__abc_44228_n7548_1_bF_buf28), .B(u2__abc_44228_n8036), .Y(u2__abc_44228_n8037_1) );
  OR2X2 OR2X2_1313 ( .A(u2__abc_44228_n8038_1), .B(u2__abc_44228_n2983_bF_buf81), .Y(u2__abc_44228_n8039) );
  OR2X2 OR2X2_1314 ( .A(u2__abc_44228_n8043_1), .B(u2__abc_44228_n8029), .Y(u2__abc_44228_n8044) );
  OR2X2 OR2X2_1315 ( .A(u2__abc_44228_n8047), .B(u2__abc_44228_n3219), .Y(u2__abc_44228_n8048_1) );
  OR2X2 OR2X2_1316 ( .A(u2__abc_44228_n8049_1), .B(u2__abc_44228_n3207), .Y(u2__abc_44228_n8050) );
  OR2X2 OR2X2_1317 ( .A(u2__abc_44228_n7548_1_bF_buf27), .B(u2__abc_44228_n8053), .Y(u2__abc_44228_n8054_1) );
  OR2X2 OR2X2_1318 ( .A(u2__abc_44228_n7547_bF_buf26), .B(u2_remHi_28_), .Y(u2__abc_44228_n8055) );
  OR2X2 OR2X2_1319 ( .A(u2__abc_44228_n8056), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n8057) );
  OR2X2 OR2X2_132 ( .A(_abc_64468_n753_bF_buf12), .B(\a[65] ), .Y(_abc_64468_n1026) );
  OR2X2 OR2X2_1320 ( .A(u2__abc_44228_n8061), .B(u2__abc_44228_n8046), .Y(u2__abc_44228_n8062) );
  OR2X2 OR2X2_1321 ( .A(u2__abc_44228_n8051), .B(u2__abc_44228_n3203), .Y(u2__abc_44228_n8066) );
  OR2X2 OR2X2_1322 ( .A(u2__abc_44228_n8067), .B(u2__abc_44228_n8065_1), .Y(u2__abc_44228_n8068) );
  OR2X2 OR2X2_1323 ( .A(u2__abc_44228_n8066), .B(u2__abc_44228_n3201), .Y(u2__abc_44228_n8069) );
  OR2X2 OR2X2_1324 ( .A(u2__abc_44228_n8072), .B(u2__abc_44228_n2983_bF_buf77), .Y(u2__abc_44228_n8073) );
  OR2X2 OR2X2_1325 ( .A(u2__abc_44228_n8071_1), .B(u2__abc_44228_n8073), .Y(u2__abc_44228_n8074) );
  OR2X2 OR2X2_1326 ( .A(u2__abc_44228_n8078), .B(u2__abc_44228_n8064), .Y(u2__abc_44228_n8079) );
  OR2X2 OR2X2_1327 ( .A(u2__abc_44228_n3348), .B(u2__abc_44228_n3572), .Y(u2__abc_44228_n8084) );
  OR2X2 OR2X2_1328 ( .A(u2__abc_44228_n8087_1), .B(u2__abc_44228_n8086), .Y(u2__abc_44228_n8088) );
  OR2X2 OR2X2_1329 ( .A(u2__abc_44228_n8088), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n8089) );
  OR2X2 OR2X2_133 ( .A(aNan_bF_buf9), .B(sqrto_142_), .Y(_abc_64468_n1028) );
  OR2X2 OR2X2_1330 ( .A(u2__abc_44228_n8093_1), .B(u2__abc_44228_n8081_1), .Y(u2__abc_44228_n8094) );
  OR2X2 OR2X2_1331 ( .A(u2__abc_44228_n8082_1), .B(u2__abc_44228_n3568), .Y(u2__abc_44228_n8097) );
  OR2X2 OR2X2_1332 ( .A(u2__abc_44228_n8097), .B(u2__abc_44228_n3579), .Y(u2__abc_44228_n8098_1) );
  OR2X2 OR2X2_1333 ( .A(u2__abc_44228_n8100), .B(u2__abc_44228_n8099), .Y(u2__abc_44228_n8101) );
  OR2X2 OR2X2_1334 ( .A(u2__abc_44228_n8104_1), .B(u2__abc_44228_n8103_1), .Y(u2__abc_44228_n8105) );
  OR2X2 OR2X2_1335 ( .A(u2__abc_44228_n8105), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n8106) );
  OR2X2 OR2X2_1336 ( .A(u2__abc_44228_n8110), .B(u2__abc_44228_n8096), .Y(u2__abc_44228_n8111) );
  OR2X2 OR2X2_1337 ( .A(u2__abc_44228_n8114_1), .B(u2__abc_44228_n3587), .Y(u2__abc_44228_n8115_1) );
  OR2X2 OR2X2_1338 ( .A(u2__abc_44228_n8115_1), .B(u2__abc_44228_n3565), .Y(u2__abc_44228_n8116) );
  OR2X2 OR2X2_1339 ( .A(u2__abc_44228_n8121), .B(u2__abc_44228_n8120_1), .Y(u2__abc_44228_n8122) );
  OR2X2 OR2X2_134 ( .A(_abc_64468_n753_bF_buf11), .B(\a[66] ), .Y(_abc_64468_n1029) );
  OR2X2 OR2X2_1340 ( .A(u2__abc_44228_n8122), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n8123) );
  OR2X2 OR2X2_1341 ( .A(u2__abc_44228_n8127), .B(u2__abc_44228_n8113), .Y(u2__abc_44228_n8128) );
  OR2X2 OR2X2_1342 ( .A(u2__abc_44228_n8133), .B(u2__abc_44228_n8132), .Y(u2__abc_44228_n8134) );
  OR2X2 OR2X2_1343 ( .A(u2__abc_44228_n8135), .B(u2__abc_44228_n3560), .Y(u2__abc_44228_n8136_1) );
  OR2X2 OR2X2_1344 ( .A(u2__abc_44228_n8138), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n8139) );
  OR2X2 OR2X2_1345 ( .A(u2__abc_44228_n8139), .B(u2__abc_44228_n8131_1), .Y(u2__abc_44228_n8140) );
  OR2X2 OR2X2_1346 ( .A(u2__abc_44228_n8144), .B(u2__abc_44228_n8130), .Y(u2__abc_44228_n8145) );
  OR2X2 OR2X2_1347 ( .A(u2__abc_44228_n8148_1), .B(u2__abc_44228_n3593), .Y(u2__abc_44228_n8149) );
  OR2X2 OR2X2_1348 ( .A(u2__abc_44228_n8149), .B(u2__abc_44228_n3546), .Y(u2__abc_44228_n8152) );
  OR2X2 OR2X2_1349 ( .A(u2__abc_44228_n8155), .B(u2__abc_44228_n8154), .Y(u2__abc_44228_n8156) );
  OR2X2 OR2X2_135 ( .A(aNan_bF_buf8), .B(sqrto_143_), .Y(_abc_64468_n1031) );
  OR2X2 OR2X2_1350 ( .A(u2__abc_44228_n8156), .B(u2__abc_44228_n2983_bF_buf67), .Y(u2__abc_44228_n8157) );
  OR2X2 OR2X2_1351 ( .A(u2__abc_44228_n8161), .B(u2__abc_44228_n8147_1), .Y(u2__abc_44228_n8162) );
  OR2X2 OR2X2_1352 ( .A(u2__abc_44228_n8166), .B(u2__abc_44228_n8165), .Y(u2__abc_44228_n8167) );
  OR2X2 OR2X2_1353 ( .A(u2__abc_44228_n8168), .B(u2__abc_44228_n3553), .Y(u2__abc_44228_n8169_1) );
  OR2X2 OR2X2_1354 ( .A(u2__abc_44228_n8172), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n8173) );
  OR2X2 OR2X2_1355 ( .A(u2__abc_44228_n8173), .B(u2__abc_44228_n8171), .Y(u2__abc_44228_n8174) );
  OR2X2 OR2X2_1356 ( .A(u2__abc_44228_n8178), .B(u2__abc_44228_n8164_1), .Y(u2__abc_44228_n8179) );
  OR2X2 OR2X2_1357 ( .A(u2__abc_44228_n8183), .B(u2__abc_44228_n3551), .Y(u2__abc_44228_n8184) );
  OR2X2 OR2X2_1358 ( .A(u2__abc_44228_n8185), .B(u2__abc_44228_n3539), .Y(u2__abc_44228_n8186_1) );
  OR2X2 OR2X2_1359 ( .A(u2__abc_44228_n8190), .B(u2__abc_44228_n2983_bF_buf63), .Y(u2__abc_44228_n8191_1) );
  OR2X2 OR2X2_136 ( .A(_abc_64468_n753_bF_buf10), .B(\a[67] ), .Y(_abc_64468_n1032) );
  OR2X2 OR2X2_1360 ( .A(u2__abc_44228_n8191_1), .B(u2__abc_44228_n8182), .Y(u2__abc_44228_n8192_1) );
  OR2X2 OR2X2_1361 ( .A(u2__abc_44228_n8196), .B(u2__abc_44228_n8181_1), .Y(u2__abc_44228_n8197_1) );
  OR2X2 OR2X2_1362 ( .A(u2__abc_44228_n8187), .B(u2__abc_44228_n3535), .Y(u2__abc_44228_n8201) );
  OR2X2 OR2X2_1363 ( .A(u2__abc_44228_n8204), .B(u2__abc_44228_n8202_1), .Y(u2__abc_44228_n8205) );
  OR2X2 OR2X2_1364 ( .A(u2__abc_44228_n8210), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n8211) );
  OR2X2 OR2X2_1365 ( .A(u2__abc_44228_n8211), .B(u2__abc_44228_n8206), .Y(u2__abc_44228_n8212) );
  OR2X2 OR2X2_1366 ( .A(u2__abc_44228_n8216), .B(u2__abc_44228_n8199), .Y(u2__abc_44228_n8217) );
  OR2X2 OR2X2_1367 ( .A(u2__abc_44228_n8220), .B(u2__abc_44228_n3603), .Y(u2__abc_44228_n8221) );
  OR2X2 OR2X2_1368 ( .A(u2__abc_44228_n8221), .B(u2__abc_44228_n3509), .Y(u2__abc_44228_n8222) );
  OR2X2 OR2X2_1369 ( .A(u2__abc_44228_n8227), .B(u2__abc_44228_n8226), .Y(u2__abc_44228_n8228) );
  OR2X2 OR2X2_137 ( .A(aNan_bF_buf7), .B(sqrto_144_), .Y(_abc_64468_n1034) );
  OR2X2 OR2X2_1370 ( .A(u2__abc_44228_n8228), .B(u2__abc_44228_n2983_bF_buf60), .Y(u2__abc_44228_n8229) );
  OR2X2 OR2X2_1371 ( .A(u2__abc_44228_n8233), .B(u2__abc_44228_n8219_1), .Y(u2__abc_44228_n8234) );
  OR2X2 OR2X2_1372 ( .A(u2__abc_44228_n8223), .B(u2__abc_44228_n3505_1), .Y(u2__abc_44228_n8238) );
  OR2X2 OR2X2_1373 ( .A(u2__abc_44228_n8239), .B(u2__abc_44228_n8237), .Y(u2__abc_44228_n8240) );
  OR2X2 OR2X2_1374 ( .A(u2__abc_44228_n8238), .B(u2__abc_44228_n3503), .Y(u2__abc_44228_n8241_1) );
  OR2X2 OR2X2_1375 ( .A(u2__abc_44228_n8244), .B(u2__abc_44228_n2983_bF_buf58), .Y(u2__abc_44228_n8245) );
  OR2X2 OR2X2_1376 ( .A(u2__abc_44228_n8245), .B(u2__abc_44228_n8243), .Y(u2__abc_44228_n8246_1) );
  OR2X2 OR2X2_1377 ( .A(u2__abc_44228_n8250), .B(u2__abc_44228_n8236_1), .Y(u2__abc_44228_n8251) );
  OR2X2 OR2X2_1378 ( .A(u2__abc_44228_n8254), .B(u2__abc_44228_n3606), .Y(u2__abc_44228_n8255) );
  OR2X2 OR2X2_1379 ( .A(u2__abc_44228_n8255), .B(u2__abc_44228_n3523_1), .Y(u2__abc_44228_n8256) );
  OR2X2 OR2X2_138 ( .A(_abc_64468_n753_bF_buf9), .B(\a[68] ), .Y(_abc_64468_n1035) );
  OR2X2 OR2X2_1380 ( .A(u2__abc_44228_n8261), .B(u2__abc_44228_n8260), .Y(u2__abc_44228_n8262) );
  OR2X2 OR2X2_1381 ( .A(u2__abc_44228_n8262), .B(u2__abc_44228_n2983_bF_buf56), .Y(u2__abc_44228_n8263_1) );
  OR2X2 OR2X2_1382 ( .A(u2__abc_44228_n8267), .B(u2__abc_44228_n8253), .Y(u2__abc_44228_n8268_1) );
  OR2X2 OR2X2_1383 ( .A(u2__abc_44228_n8274_1), .B(u2__abc_44228_n8275), .Y(u2__abc_44228_n8276) );
  OR2X2 OR2X2_1384 ( .A(u2__abc_44228_n8278), .B(u2__abc_44228_n2983_bF_buf54), .Y(u2__abc_44228_n8279_1) );
  OR2X2 OR2X2_1385 ( .A(u2__abc_44228_n8279_1), .B(u2__abc_44228_n8277), .Y(u2__abc_44228_n8280_1) );
  OR2X2 OR2X2_1386 ( .A(u2__abc_44228_n8284), .B(u2__abc_44228_n8270), .Y(u2__abc_44228_n8285_1) );
  OR2X2 OR2X2_1387 ( .A(u2__abc_44228_n8288), .B(u2__abc_44228_n3515), .Y(u2__abc_44228_n8289) );
  OR2X2 OR2X2_1388 ( .A(u2__abc_44228_n8290_1), .B(u2__abc_44228_n3487), .Y(u2__abc_44228_n8293) );
  OR2X2 OR2X2_1389 ( .A(u2__abc_44228_n8296_1), .B(u2__abc_44228_n8295), .Y(u2__abc_44228_n8297) );
  OR2X2 OR2X2_139 ( .A(aNan_bF_buf6), .B(sqrto_145_), .Y(_abc_64468_n1037) );
  OR2X2 OR2X2_1390 ( .A(u2__abc_44228_n8297), .B(u2__abc_44228_n2983_bF_buf52), .Y(u2__abc_44228_n8298) );
  OR2X2 OR2X2_1391 ( .A(u2__abc_44228_n8302_1), .B(u2__abc_44228_n8287), .Y(u2__abc_44228_n8303) );
  OR2X2 OR2X2_1392 ( .A(u2__abc_44228_n8307_1), .B(u2__abc_44228_n8306), .Y(u2__abc_44228_n8308) );
  OR2X2 OR2X2_1393 ( .A(u2__abc_44228_n8309), .B(u2__abc_44228_n3494), .Y(u2__abc_44228_n8310) );
  OR2X2 OR2X2_1394 ( .A(u2__abc_44228_n8313_1), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n8314) );
  OR2X2 OR2X2_1395 ( .A(u2__abc_44228_n8314), .B(u2__abc_44228_n8312_1), .Y(u2__abc_44228_n8315) );
  OR2X2 OR2X2_1396 ( .A(u2__abc_44228_n8319), .B(u2__abc_44228_n8305), .Y(u2__abc_44228_n8320) );
  OR2X2 OR2X2_1397 ( .A(u2__abc_44228_n8323_1), .B(u2__abc_44228_n3492), .Y(u2__abc_44228_n8324_1) );
  OR2X2 OR2X2_1398 ( .A(u2__abc_44228_n8325), .B(u2__abc_44228_n3480), .Y(u2__abc_44228_n8326) );
  OR2X2 OR2X2_1399 ( .A(u2__abc_44228_n8329_1), .B(u2__abc_44228_n7548_1_bF_buf11), .Y(u2__abc_44228_n8330) );
  OR2X2 OR2X2_14 ( .A(_abc_64468_n753_bF_buf1), .B(\a[6] ), .Y(_abc_64468_n849) );
  OR2X2 OR2X2_140 ( .A(_abc_64468_n753_bF_buf8), .B(\a[69] ), .Y(_abc_64468_n1038) );
  OR2X2 OR2X2_1400 ( .A(u2__abc_44228_n7547_bF_buf10), .B(u2_remHi_44_), .Y(u2__abc_44228_n8331) );
  OR2X2 OR2X2_1401 ( .A(u2__abc_44228_n8332), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n8333) );
  OR2X2 OR2X2_1402 ( .A(u2__abc_44228_n8337), .B(u2__abc_44228_n8322), .Y(u2__abc_44228_n8338) );
  OR2X2 OR2X2_1403 ( .A(u2__abc_44228_n8327), .B(u2__abc_44228_n3476), .Y(u2__abc_44228_n8342) );
  OR2X2 OR2X2_1404 ( .A(u2__abc_44228_n8343), .B(u2__abc_44228_n8341), .Y(u2__abc_44228_n8344) );
  OR2X2 OR2X2_1405 ( .A(u2__abc_44228_n8342), .B(u2__abc_44228_n3474), .Y(u2__abc_44228_n8345_1) );
  OR2X2 OR2X2_1406 ( .A(u2__abc_44228_n8348), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n8349) );
  OR2X2 OR2X2_1407 ( .A(u2__abc_44228_n8347), .B(u2__abc_44228_n8349), .Y(u2__abc_44228_n8350) );
  OR2X2 OR2X2_1408 ( .A(u2__abc_44228_n8354), .B(u2__abc_44228_n8340_1), .Y(u2__abc_44228_n8355) );
  OR2X2 OR2X2_1409 ( .A(u2__abc_44228_n8358), .B(u2__abc_44228_n3623), .Y(u2__abc_44228_n8359) );
  OR2X2 OR2X2_141 ( .A(aNan_bF_buf5), .B(sqrto_146_), .Y(_abc_64468_n1040) );
  OR2X2 OR2X2_1410 ( .A(u2__abc_44228_n8359), .B(u2__abc_44228_n3463), .Y(u2__abc_44228_n8362_1) );
  OR2X2 OR2X2_1411 ( .A(u2__abc_44228_n8365), .B(u2__abc_44228_n8364), .Y(u2__abc_44228_n8366) );
  OR2X2 OR2X2_1412 ( .A(u2__abc_44228_n8366), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n8367_1) );
  OR2X2 OR2X2_1413 ( .A(u2__abc_44228_n8371), .B(u2__abc_44228_n8357_1), .Y(u2__abc_44228_n8372) );
  OR2X2 OR2X2_1414 ( .A(u2__abc_44228_n8360), .B(u2__abc_44228_n3459), .Y(u2__abc_44228_n8376) );
  OR2X2 OR2X2_1415 ( .A(u2__abc_44228_n8377), .B(u2__abc_44228_n8375), .Y(u2__abc_44228_n8378_1) );
  OR2X2 OR2X2_1416 ( .A(u2__abc_44228_n8376), .B(u2__abc_44228_n3457_1), .Y(u2__abc_44228_n8379_1) );
  OR2X2 OR2X2_1417 ( .A(u2__abc_44228_n8382), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n8383) );
  OR2X2 OR2X2_1418 ( .A(u2__abc_44228_n8383), .B(u2__abc_44228_n8381), .Y(u2__abc_44228_n8384_1) );
  OR2X2 OR2X2_1419 ( .A(u2__abc_44228_n8388), .B(u2__abc_44228_n8374), .Y(u2__abc_44228_n8389_1) );
  OR2X2 OR2X2_142 ( .A(_abc_64468_n753_bF_buf7), .B(\a[70] ), .Y(_abc_64468_n1041) );
  OR2X2 OR2X2_1420 ( .A(u2__abc_44228_n8392), .B(u2__abc_44228_n3626), .Y(u2__abc_44228_n8393) );
  OR2X2 OR2X2_1421 ( .A(u2__abc_44228_n8393), .B(u2__abc_44228_n3449_1), .Y(u2__abc_44228_n8394) );
  OR2X2 OR2X2_1422 ( .A(u2__abc_44228_n8399), .B(u2__abc_44228_n8398), .Y(u2__abc_44228_n8400_1) );
  OR2X2 OR2X2_1423 ( .A(u2__abc_44228_n8400_1), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n8401_1) );
  OR2X2 OR2X2_1424 ( .A(u2__abc_44228_n8405), .B(u2__abc_44228_n8391), .Y(u2__abc_44228_n8406_1) );
  OR2X2 OR2X2_1425 ( .A(u2__abc_44228_n8395_1), .B(u2__abc_44228_n3445), .Y(u2__abc_44228_n8410) );
  OR2X2 OR2X2_1426 ( .A(u2__abc_44228_n8413), .B(u2__abc_44228_n8411_1), .Y(u2__abc_44228_n8414) );
  OR2X2 OR2X2_1427 ( .A(u2__abc_44228_n8416), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n8417_1) );
  OR2X2 OR2X2_1428 ( .A(u2__abc_44228_n8417_1), .B(u2__abc_44228_n8415), .Y(u2__abc_44228_n8418) );
  OR2X2 OR2X2_1429 ( .A(u2__abc_44228_n8422_1), .B(u2__abc_44228_n8408), .Y(u2__abc_44228_n8423_1) );
  OR2X2 OR2X2_143 ( .A(aNan_bF_buf4), .B(sqrto_147_), .Y(_abc_64468_n1043) );
  OR2X2 OR2X2_1430 ( .A(u2__abc_44228_n8426), .B(u2__abc_44228_n3630), .Y(u2__abc_44228_n8427) );
  OR2X2 OR2X2_1431 ( .A(u2__abc_44228_n8427), .B(u2__abc_44228_n3427), .Y(u2__abc_44228_n8430) );
  OR2X2 OR2X2_1432 ( .A(u2__abc_44228_n8433_1), .B(u2__abc_44228_n8432), .Y(u2__abc_44228_n8434_1) );
  OR2X2 OR2X2_1433 ( .A(u2__abc_44228_n8434_1), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n8435) );
  OR2X2 OR2X2_1434 ( .A(u2__abc_44228_n8439_1), .B(u2__abc_44228_n8425), .Y(u2__abc_44228_n8440) );
  OR2X2 OR2X2_1435 ( .A(u2__abc_44228_n8447), .B(u2__abc_44228_n8444_1), .Y(u2__abc_44228_n8448) );
  OR2X2 OR2X2_1436 ( .A(u2__abc_44228_n8450_1), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n8451) );
  OR2X2 OR2X2_1437 ( .A(u2__abc_44228_n8451), .B(u2__abc_44228_n8449), .Y(u2__abc_44228_n8452) );
  OR2X2 OR2X2_1438 ( .A(u2__abc_44228_n8456_1), .B(u2__abc_44228_n8442), .Y(u2__abc_44228_n8457) );
  OR2X2 OR2X2_1439 ( .A(u2__abc_44228_n8460), .B(u2__abc_44228_n3432), .Y(u2__abc_44228_n8461_1) );
  OR2X2 OR2X2_144 ( .A(_abc_64468_n753_bF_buf6), .B(\a[71] ), .Y(_abc_64468_n1044) );
  OR2X2 OR2X2_1440 ( .A(u2__abc_44228_n8462), .B(u2__abc_44228_n3420), .Y(u2__abc_44228_n8463) );
  OR2X2 OR2X2_1441 ( .A(u2__abc_44228_n8468), .B(u2__abc_44228_n8467_1), .Y(u2__abc_44228_n8469) );
  OR2X2 OR2X2_1442 ( .A(u2__abc_44228_n8469), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n8470) );
  OR2X2 OR2X2_1443 ( .A(u2__abc_44228_n8474), .B(u2__abc_44228_n8459), .Y(u2__abc_44228_n8475) );
  OR2X2 OR2X2_1444 ( .A(u2__abc_44228_n8464), .B(u2__abc_44228_n3416), .Y(u2__abc_44228_n8479) );
  OR2X2 OR2X2_1445 ( .A(u2__abc_44228_n8480), .B(u2__abc_44228_n8478_1), .Y(u2__abc_44228_n8481) );
  OR2X2 OR2X2_1446 ( .A(u2__abc_44228_n8479), .B(u2__abc_44228_n3414), .Y(u2__abc_44228_n8482) );
  OR2X2 OR2X2_1447 ( .A(u2__abc_44228_n8485), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n8486) );
  OR2X2 OR2X2_1448 ( .A(u2__abc_44228_n8486), .B(u2__abc_44228_n8484), .Y(u2__abc_44228_n8487) );
  OR2X2 OR2X2_1449 ( .A(u2__abc_44228_n8491), .B(u2__abc_44228_n8477_1), .Y(u2__abc_44228_n8492) );
  OR2X2 OR2X2_145 ( .A(aNan_bF_buf3), .B(sqrto_148_), .Y(_abc_64468_n1046) );
  OR2X2 OR2X2_1450 ( .A(u2__abc_44228_n8495), .B(u2__abc_44228_n3640), .Y(u2__abc_44228_n8496) );
  OR2X2 OR2X2_1451 ( .A(u2__abc_44228_n8496), .B(u2__abc_44228_n3404), .Y(u2__abc_44228_n8497) );
  OR2X2 OR2X2_1452 ( .A(u2__abc_44228_n8502), .B(u2__abc_44228_n8501), .Y(u2__abc_44228_n8503) );
  OR2X2 OR2X2_1453 ( .A(u2__abc_44228_n8503), .B(u2__abc_44228_n2983_bF_buf30), .Y(u2__abc_44228_n8504) );
  OR2X2 OR2X2_1454 ( .A(u2__abc_44228_n8508), .B(u2__abc_44228_n8494_1), .Y(u2__abc_44228_n8509) );
  OR2X2 OR2X2_1455 ( .A(u2__abc_44228_n8514), .B(u2__abc_44228_n8513), .Y(u2__abc_44228_n8515) );
  OR2X2 OR2X2_1456 ( .A(u2__abc_44228_n8516_1), .B(u2__abc_44228_n3398), .Y(u2__abc_44228_n8517) );
  OR2X2 OR2X2_1457 ( .A(u2__abc_44228_n8519), .B(u2__abc_44228_n2983_bF_buf28), .Y(u2__abc_44228_n8520) );
  OR2X2 OR2X2_1458 ( .A(u2__abc_44228_n8520), .B(u2__abc_44228_n8512), .Y(u2__abc_44228_n8521_1) );
  OR2X2 OR2X2_1459 ( .A(u2__abc_44228_n8525), .B(u2__abc_44228_n8511_1), .Y(u2__abc_44228_n8526) );
  OR2X2 OR2X2_146 ( .A(_abc_64468_n753_bF_buf5), .B(\a[72] ), .Y(_abc_64468_n1047) );
  OR2X2 OR2X2_1460 ( .A(u2__abc_44228_n8529), .B(u2__abc_44228_n3645), .Y(u2__abc_44228_n8530) );
  OR2X2 OR2X2_1461 ( .A(u2__abc_44228_n8530), .B(u2__abc_44228_n3390), .Y(u2__abc_44228_n8531) );
  OR2X2 OR2X2_1462 ( .A(u2__abc_44228_n7548_1_bF_buf57), .B(u2__abc_44228_n8534), .Y(u2__abc_44228_n8535) );
  OR2X2 OR2X2_1463 ( .A(u2__abc_44228_n7547_bF_buf56), .B(u2_remHi_56_), .Y(u2__abc_44228_n8536) );
  OR2X2 OR2X2_1464 ( .A(u2__abc_44228_n8537), .B(u2__abc_44228_n2983_bF_buf26), .Y(u2__abc_44228_n8538_1) );
  OR2X2 OR2X2_1465 ( .A(u2__abc_44228_n8542), .B(u2__abc_44228_n8528), .Y(u2__abc_44228_n8543_1) );
  OR2X2 OR2X2_1466 ( .A(u2__abc_44228_n8547), .B(u2__abc_44228_n3384), .Y(u2__abc_44228_n8548) );
  OR2X2 OR2X2_1467 ( .A(u2__abc_44228_n8546), .B(u2__abc_44228_n8549_1), .Y(u2__abc_44228_n8550) );
  OR2X2 OR2X2_1468 ( .A(u2__abc_44228_n8553), .B(u2__abc_44228_n2983_bF_buf24), .Y(u2__abc_44228_n8554_1) );
  OR2X2 OR2X2_1469 ( .A(u2__abc_44228_n8554_1), .B(u2__abc_44228_n8552), .Y(u2__abc_44228_n8555_1) );
  OR2X2 OR2X2_147 ( .A(aNan_bF_buf2), .B(sqrto_149_), .Y(_abc_64468_n1049) );
  OR2X2 OR2X2_1470 ( .A(u2__abc_44228_n8559), .B(u2__abc_44228_n8545), .Y(u2__abc_44228_n8560_1) );
  OR2X2 OR2X2_1471 ( .A(u2__abc_44228_n8563), .B(u2__abc_44228_n3382), .Y(u2__abc_44228_n8564) );
  OR2X2 OR2X2_1472 ( .A(u2__abc_44228_n8565_1), .B(u2__abc_44228_n3368), .Y(u2__abc_44228_n8568) );
  OR2X2 OR2X2_1473 ( .A(u2__abc_44228_n7548_1_bF_buf55), .B(u2__abc_44228_n8569), .Y(u2__abc_44228_n8570) );
  OR2X2 OR2X2_1474 ( .A(u2__abc_44228_n7547_bF_buf54), .B(u2_remHi_58_), .Y(u2__abc_44228_n8571_1) );
  OR2X2 OR2X2_1475 ( .A(u2__abc_44228_n8572), .B(u2__abc_44228_n2983_bF_buf22), .Y(u2__abc_44228_n8573) );
  OR2X2 OR2X2_1476 ( .A(u2__abc_44228_n8577_1), .B(u2__abc_44228_n8562), .Y(u2__abc_44228_n8578) );
  OR2X2 OR2X2_1477 ( .A(u2__abc_44228_n8582_1), .B(u2__abc_44228_n3375), .Y(u2__abc_44228_n8583) );
  OR2X2 OR2X2_1478 ( .A(u2__abc_44228_n8581), .B(u2__abc_44228_n8584), .Y(u2__abc_44228_n8585) );
  OR2X2 OR2X2_1479 ( .A(u2__abc_44228_n8588_1), .B(u2__abc_44228_n2983_bF_buf20), .Y(u2__abc_44228_n8589) );
  OR2X2 OR2X2_148 ( .A(_abc_64468_n753_bF_buf4), .B(\a[73] ), .Y(_abc_64468_n1050) );
  OR2X2 OR2X2_1480 ( .A(u2__abc_44228_n8587_1), .B(u2__abc_44228_n8589), .Y(u2__abc_44228_n8590) );
  OR2X2 OR2X2_1481 ( .A(u2__abc_44228_n8594), .B(u2__abc_44228_n8580), .Y(u2__abc_44228_n8595) );
  OR2X2 OR2X2_1482 ( .A(u2__abc_44228_n8598_1), .B(u2__abc_44228_n3373), .Y(u2__abc_44228_n8599_1) );
  OR2X2 OR2X2_1483 ( .A(u2__abc_44228_n8600), .B(u2__abc_44228_n3361), .Y(u2__abc_44228_n8601) );
  OR2X2 OR2X2_1484 ( .A(u2__abc_44228_n8606), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n8607) );
  OR2X2 OR2X2_1485 ( .A(u2__abc_44228_n8605), .B(u2__abc_44228_n8607), .Y(u2__abc_44228_n8608) );
  OR2X2 OR2X2_1486 ( .A(u2__abc_44228_n8612), .B(u2__abc_44228_n8597), .Y(u2__abc_44228_n8613) );
  OR2X2 OR2X2_1487 ( .A(u2__abc_44228_n8602), .B(u2__abc_44228_n3357), .Y(u2__abc_44228_n8617) );
  OR2X2 OR2X2_1488 ( .A(u2__abc_44228_n8618), .B(u2__abc_44228_n8616), .Y(u2__abc_44228_n8619) );
  OR2X2 OR2X2_1489 ( .A(u2__abc_44228_n8617), .B(u2__abc_44228_n3355), .Y(u2__abc_44228_n8620_1) );
  OR2X2 OR2X2_149 ( .A(aNan_bF_buf1), .B(sqrto_150_), .Y(_abc_64468_n1052) );
  OR2X2 OR2X2_1490 ( .A(u2__abc_44228_n8623), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n8624) );
  OR2X2 OR2X2_1491 ( .A(u2__abc_44228_n8622), .B(u2__abc_44228_n8624), .Y(u2__abc_44228_n8625) );
  OR2X2 OR2X2_1492 ( .A(u2__abc_44228_n8629), .B(u2__abc_44228_n8615_1), .Y(u2__abc_44228_n8630) );
  OR2X2 OR2X2_1493 ( .A(u2__abc_44228_n3664), .B(u2__abc_44228_n4134), .Y(u2__abc_44228_n8633) );
  OR2X2 OR2X2_1494 ( .A(u2__abc_44228_n8638), .B(u2__abc_44228_n8637_1), .Y(u2__abc_44228_n8639) );
  OR2X2 OR2X2_1495 ( .A(u2__abc_44228_n8639), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n8640) );
  OR2X2 OR2X2_1496 ( .A(u2__abc_44228_n8644), .B(u2__abc_44228_n8632_1), .Y(u2__abc_44228_n8645) );
  OR2X2 OR2X2_1497 ( .A(u2__abc_44228_n8634), .B(u2__abc_44228_n4130), .Y(u2__abc_44228_n8649) );
  OR2X2 OR2X2_1498 ( .A(u2__abc_44228_n8650), .B(u2__abc_44228_n8648_1), .Y(u2__abc_44228_n8651) );
  OR2X2 OR2X2_1499 ( .A(u2__abc_44228_n8649), .B(u2__abc_44228_n4128_1), .Y(u2__abc_44228_n8652) );
  OR2X2 OR2X2_15 ( .A(aNan_bF_buf2), .B(sqrto_83_), .Y(_abc_64468_n851) );
  OR2X2 OR2X2_150 ( .A(_abc_64468_n753_bF_buf3), .B(\a[74] ), .Y(_abc_64468_n1053) );
  OR2X2 OR2X2_1500 ( .A(u2__abc_44228_n8655), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n8656) );
  OR2X2 OR2X2_1501 ( .A(u2__abc_44228_n8656), .B(u2__abc_44228_n8654_1), .Y(u2__abc_44228_n8657) );
  OR2X2 OR2X2_1502 ( .A(u2__abc_44228_n8661), .B(u2__abc_44228_n8647), .Y(u2__abc_44228_n8662) );
  OR2X2 OR2X2_1503 ( .A(u2__abc_44228_n8665_1), .B(u2__abc_44228_n4143), .Y(u2__abc_44228_n8666) );
  OR2X2 OR2X2_1504 ( .A(u2__abc_44228_n8666), .B(u2__abc_44228_n4120), .Y(u2__abc_44228_n8667) );
  OR2X2 OR2X2_1505 ( .A(u2__abc_44228_n8672), .B(u2__abc_44228_n8671), .Y(u2__abc_44228_n8673) );
  OR2X2 OR2X2_1506 ( .A(u2__abc_44228_n8673), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n8674) );
  OR2X2 OR2X2_1507 ( .A(u2__abc_44228_n8678), .B(u2__abc_44228_n8664_1), .Y(u2__abc_44228_n8679) );
  OR2X2 OR2X2_1508 ( .A(u2__abc_44228_n8685), .B(u2__abc_44228_n8686_1), .Y(u2__abc_44228_n8687_1) );
  OR2X2 OR2X2_1509 ( .A(u2__abc_44228_n8689), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n8690) );
  OR2X2 OR2X2_151 ( .A(aNan_bF_buf0), .B(sqrto_151_), .Y(_abc_64468_n1055) );
  OR2X2 OR2X2_1510 ( .A(u2__abc_44228_n8690), .B(u2__abc_44228_n8688), .Y(u2__abc_44228_n8691) );
  OR2X2 OR2X2_1511 ( .A(u2__abc_44228_n8695), .B(u2__abc_44228_n8681_1), .Y(u2__abc_44228_n8696) );
  OR2X2 OR2X2_1512 ( .A(u2__abc_44228_n8699), .B(u2__abc_44228_n4149), .Y(u2__abc_44228_n8700) );
  OR2X2 OR2X2_1513 ( .A(u2__abc_44228_n8700), .B(u2__abc_44228_n4108), .Y(u2__abc_44228_n8703_1) );
  OR2X2 OR2X2_1514 ( .A(u2__abc_44228_n8706), .B(u2__abc_44228_n8705), .Y(u2__abc_44228_n8707) );
  OR2X2 OR2X2_1515 ( .A(u2__abc_44228_n8707), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n8708_1) );
  OR2X2 OR2X2_1516 ( .A(u2__abc_44228_n8712), .B(u2__abc_44228_n8698_1), .Y(u2__abc_44228_n8713) );
  OR2X2 OR2X2_1517 ( .A(u2__abc_44228_n8701), .B(u2__abc_44228_n4104), .Y(u2__abc_44228_n8717) );
  OR2X2 OR2X2_1518 ( .A(u2__abc_44228_n8720_1), .B(u2__abc_44228_n8718), .Y(u2__abc_44228_n8721) );
  OR2X2 OR2X2_1519 ( .A(u2__abc_44228_n8723), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n8724) );
  OR2X2 OR2X2_152 ( .A(_abc_64468_n753_bF_buf2), .B(\a[75] ), .Y(_abc_64468_n1056) );
  OR2X2 OR2X2_1520 ( .A(u2__abc_44228_n8724), .B(u2__abc_44228_n8722), .Y(u2__abc_44228_n8725_1) );
  OR2X2 OR2X2_1521 ( .A(u2__abc_44228_n8729), .B(u2__abc_44228_n8715), .Y(u2__abc_44228_n8730_1) );
  OR2X2 OR2X2_1522 ( .A(u2__abc_44228_n8734), .B(u2__abc_44228_n4152), .Y(u2__abc_44228_n8735) );
  OR2X2 OR2X2_1523 ( .A(u2__abc_44228_n8735), .B(u2__abc_44228_n4094), .Y(u2__abc_44228_n8736_1) );
  OR2X2 OR2X2_1524 ( .A(u2__abc_44228_n8740), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n8741_1) );
  OR2X2 OR2X2_1525 ( .A(u2__abc_44228_n8741_1), .B(u2__abc_44228_n8733), .Y(u2__abc_44228_n8742_1) );
  OR2X2 OR2X2_1526 ( .A(u2__abc_44228_n8746), .B(u2__abc_44228_n8732), .Y(u2__abc_44228_n8747_1) );
  OR2X2 OR2X2_1527 ( .A(u2__abc_44228_n8737), .B(u2__abc_44228_n4090_1), .Y(u2__abc_44228_n8752_1) );
  OR2X2 OR2X2_1528 ( .A(u2__abc_44228_n8755), .B(u2__abc_44228_n8753_1), .Y(u2__abc_44228_n8756) );
  OR2X2 OR2X2_1529 ( .A(u2__abc_44228_n8757), .B(u2__abc_44228_n2983_bF_buf1), .Y(u2__abc_44228_n8758_1) );
  OR2X2 OR2X2_153 ( .A(aNan_bF_buf10), .B(sqrto_152_), .Y(_abc_64468_n1058) );
  OR2X2 OR2X2_1530 ( .A(u2__abc_44228_n8758_1), .B(u2__abc_44228_n8750), .Y(u2__abc_44228_n8759) );
  OR2X2 OR2X2_1531 ( .A(u2__abc_44228_n8763_1), .B(u2__abc_44228_n8749), .Y(u2__abc_44228_n8764_1) );
  OR2X2 OR2X2_1532 ( .A(u2__abc_44228_n8767), .B(u2__abc_44228_n4157_1), .Y(u2__abc_44228_n8768) );
  OR2X2 OR2X2_1533 ( .A(u2__abc_44228_n8768), .B(u2__abc_44228_n4064), .Y(u2__abc_44228_n8769_1) );
  OR2X2 OR2X2_1534 ( .A(u2__abc_44228_n8774_1), .B(u2__abc_44228_n8773), .Y(u2__abc_44228_n8775_1) );
  OR2X2 OR2X2_1535 ( .A(u2__abc_44228_n8775_1), .B(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n8776) );
  OR2X2 OR2X2_1536 ( .A(u2__abc_44228_n8780_1), .B(u2__abc_44228_n8766), .Y(u2__abc_44228_n8781) );
  OR2X2 OR2X2_1537 ( .A(u2__abc_44228_n8770), .B(u2__abc_44228_n4060), .Y(u2__abc_44228_n8785_1) );
  OR2X2 OR2X2_1538 ( .A(u2__abc_44228_n8788), .B(u2__abc_44228_n8786_1), .Y(u2__abc_44228_n8789) );
  OR2X2 OR2X2_1539 ( .A(u2__abc_44228_n8791_1), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n8792) );
  OR2X2 OR2X2_154 ( .A(_abc_64468_n753_bF_buf1), .B(\a[76] ), .Y(_abc_64468_n1059) );
  OR2X2 OR2X2_1540 ( .A(u2__abc_44228_n8792), .B(u2__abc_44228_n8790), .Y(u2__abc_44228_n8793) );
  OR2X2 OR2X2_1541 ( .A(u2__abc_44228_n8797_1), .B(u2__abc_44228_n8783), .Y(u2__abc_44228_n8798) );
  OR2X2 OR2X2_1542 ( .A(u2__abc_44228_n8802_1), .B(u2__abc_44228_n4160), .Y(u2__abc_44228_n8803) );
  OR2X2 OR2X2_1543 ( .A(u2__abc_44228_n8803), .B(u2__abc_44228_n4078), .Y(u2__abc_44228_n8804) );
  OR2X2 OR2X2_1544 ( .A(u2__abc_44228_n8808_1), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n8809) );
  OR2X2 OR2X2_1545 ( .A(u2__abc_44228_n8809), .B(u2__abc_44228_n8801), .Y(u2__abc_44228_n8810) );
  OR2X2 OR2X2_1546 ( .A(u2__abc_44228_n8814), .B(u2__abc_44228_n8800), .Y(u2__abc_44228_n8815) );
  OR2X2 OR2X2_1547 ( .A(u2__abc_44228_n8822), .B(u2__abc_44228_n8823), .Y(u2__abc_44228_n8824_1) );
  OR2X2 OR2X2_1548 ( .A(u2__abc_44228_n8825), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n8826) );
  OR2X2 OR2X2_1549 ( .A(u2__abc_44228_n8826), .B(u2__abc_44228_n8818_1), .Y(u2__abc_44228_n8827) );
  OR2X2 OR2X2_155 ( .A(aNan_bF_buf9), .B(sqrto_153_), .Y(_abc_64468_n1061) );
  OR2X2 OR2X2_1550 ( .A(u2__abc_44228_n8831), .B(u2__abc_44228_n8817), .Y(u2__abc_44228_n8832) );
  OR2X2 OR2X2_1551 ( .A(u2__abc_44228_n8835_1), .B(u2__abc_44228_n4070_1), .Y(u2__abc_44228_n8836) );
  OR2X2 OR2X2_1552 ( .A(u2__abc_44228_n8837), .B(u2__abc_44228_n4042), .Y(u2__abc_44228_n8840_1) );
  OR2X2 OR2X2_1553 ( .A(u2__abc_44228_n7548_1_bF_buf39), .B(u2__abc_44228_n8841_1), .Y(u2__abc_44228_n8842) );
  OR2X2 OR2X2_1554 ( .A(u2__abc_44228_n7547_bF_buf38), .B(u2_remHi_74_), .Y(u2__abc_44228_n8843) );
  OR2X2 OR2X2_1555 ( .A(u2__abc_44228_n8844), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n8845) );
  OR2X2 OR2X2_1556 ( .A(u2__abc_44228_n8849), .B(u2__abc_44228_n8834), .Y(u2__abc_44228_n8850) );
  OR2X2 OR2X2_1557 ( .A(u2__abc_44228_n8854), .B(u2__abc_44228_n4049), .Y(u2__abc_44228_n8855) );
  OR2X2 OR2X2_1558 ( .A(u2__abc_44228_n8853), .B(u2__abc_44228_n8856), .Y(u2__abc_44228_n8857_1) );
  OR2X2 OR2X2_1559 ( .A(u2__abc_44228_n8860), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n8861) );
  OR2X2 OR2X2_156 ( .A(_abc_64468_n753_bF_buf0), .B(\a[77] ), .Y(_abc_64468_n1062) );
  OR2X2 OR2X2_1560 ( .A(u2__abc_44228_n8859), .B(u2__abc_44228_n8861), .Y(u2__abc_44228_n8862_1) );
  OR2X2 OR2X2_1561 ( .A(u2__abc_44228_n8866), .B(u2__abc_44228_n8852_1), .Y(u2__abc_44228_n8867) );
  OR2X2 OR2X2_1562 ( .A(u2__abc_44228_n8870), .B(u2__abc_44228_n4047), .Y(u2__abc_44228_n8871) );
  OR2X2 OR2X2_1563 ( .A(u2__abc_44228_n8872), .B(u2__abc_44228_n4035), .Y(u2__abc_44228_n8873_1) );
  OR2X2 OR2X2_1564 ( .A(u2__abc_44228_n8878), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n8879_1) );
  OR2X2 OR2X2_1565 ( .A(u2__abc_44228_n8877), .B(u2__abc_44228_n8879_1), .Y(u2__abc_44228_n8880) );
  OR2X2 OR2X2_1566 ( .A(u2__abc_44228_n8884_1), .B(u2__abc_44228_n8869), .Y(u2__abc_44228_n8885_1) );
  OR2X2 OR2X2_1567 ( .A(u2__abc_44228_n8890_1), .B(u2__abc_44228_n8888), .Y(u2__abc_44228_n8891) );
  OR2X2 OR2X2_1568 ( .A(u2__abc_44228_n8892), .B(u2__abc_44228_n4029), .Y(u2__abc_44228_n8893) );
  OR2X2 OR2X2_1569 ( .A(u2__abc_44228_n8896_1), .B(u2__abc_44228_n2983_bF_buf128), .Y(u2__abc_44228_n8897) );
  OR2X2 OR2X2_157 ( .A(aNan_bF_buf8), .B(sqrto_154_), .Y(_abc_64468_n1064) );
  OR2X2 OR2X2_1570 ( .A(u2__abc_44228_n8895_1), .B(u2__abc_44228_n8897), .Y(u2__abc_44228_n8898) );
  OR2X2 OR2X2_1571 ( .A(u2__abc_44228_n8902), .B(u2__abc_44228_n8887), .Y(u2__abc_44228_n8903) );
  OR2X2 OR2X2_1572 ( .A(u2__abc_44228_n8906_1), .B(u2__abc_44228_n4177), .Y(u2__abc_44228_n8907_1) );
  OR2X2 OR2X2_1573 ( .A(u2__abc_44228_n8907_1), .B(u2__abc_44228_n4011), .Y(u2__abc_44228_n8910) );
  OR2X2 OR2X2_1574 ( .A(u2__abc_44228_n8913), .B(u2__abc_44228_n8912_1), .Y(u2__abc_44228_n8914) );
  OR2X2 OR2X2_1575 ( .A(u2__abc_44228_n8914), .B(u2__abc_44228_n2983_bF_buf126), .Y(u2__abc_44228_n8915) );
  OR2X2 OR2X2_1576 ( .A(u2__abc_44228_n8919), .B(u2__abc_44228_n8905), .Y(u2__abc_44228_n8920) );
  OR2X2 OR2X2_1577 ( .A(u2__abc_44228_n8926), .B(u2__abc_44228_n8927), .Y(u2__abc_44228_n8928_1) );
  OR2X2 OR2X2_1578 ( .A(u2__abc_44228_n8930), .B(u2__abc_44228_n2983_bF_buf124), .Y(u2__abc_44228_n8931) );
  OR2X2 OR2X2_1579 ( .A(u2__abc_44228_n8931), .B(u2__abc_44228_n8929_1), .Y(u2__abc_44228_n8932) );
  OR2X2 OR2X2_158 ( .A(_abc_64468_n753_bF_buf13), .B(\a[78] ), .Y(_abc_64468_n1065) );
  OR2X2 OR2X2_1580 ( .A(u2__abc_44228_n8936), .B(u2__abc_44228_n8922), .Y(u2__abc_44228_n8937) );
  OR2X2 OR2X2_1581 ( .A(u2__abc_44228_n8940_1), .B(u2__abc_44228_n4016), .Y(u2__abc_44228_n8941) );
  OR2X2 OR2X2_1582 ( .A(u2__abc_44228_n8942), .B(u2__abc_44228_n4004), .Y(u2__abc_44228_n8943) );
  OR2X2 OR2X2_1583 ( .A(u2__abc_44228_n8948), .B(u2__abc_44228_n8947), .Y(u2__abc_44228_n8949) );
  OR2X2 OR2X2_1584 ( .A(u2__abc_44228_n8949), .B(u2__abc_44228_n2983_bF_buf122), .Y(u2__abc_44228_n8950_1) );
  OR2X2 OR2X2_1585 ( .A(u2__abc_44228_n8954), .B(u2__abc_44228_n8939_1), .Y(u2__abc_44228_n8955) );
  OR2X2 OR2X2_1586 ( .A(u2__abc_44228_n8944), .B(u2__abc_44228_n4000), .Y(u2__abc_44228_n8958) );
  OR2X2 OR2X2_1587 ( .A(u2__abc_44228_n8958), .B(u2__abc_44228_n3998), .Y(u2__abc_44228_n8959) );
  OR2X2 OR2X2_1588 ( .A(u2__abc_44228_n8961_1), .B(u2__abc_44228_n8960), .Y(u2__abc_44228_n8962_1) );
  OR2X2 OR2X2_1589 ( .A(u2__abc_44228_n8963), .B(u2__abc_44228_n7548_1_bF_buf32), .Y(u2__abc_44228_n8964) );
  OR2X2 OR2X2_159 ( .A(aNan_bF_buf7), .B(sqrto_155_), .Y(_abc_64468_n1067) );
  OR2X2 OR2X2_1590 ( .A(u2__abc_44228_n7547_bF_buf31), .B(u2_remHi_81_), .Y(u2__abc_44228_n8965) );
  OR2X2 OR2X2_1591 ( .A(u2__abc_44228_n8966), .B(u2__abc_44228_n2983_bF_buf120), .Y(u2__abc_44228_n8967_1) );
  OR2X2 OR2X2_1592 ( .A(u2__abc_44228_n8971), .B(u2__abc_44228_n8957), .Y(u2__abc_44228_n8972_1) );
  OR2X2 OR2X2_1593 ( .A(u2__abc_44228_n8976), .B(u2__abc_44228_n4186), .Y(u2__abc_44228_n8977) );
  OR2X2 OR2X2_1594 ( .A(u2__abc_44228_n8977), .B(u2__abc_44228_n3982), .Y(u2__abc_44228_n8980) );
  OR2X2 OR2X2_1595 ( .A(u2__abc_44228_n8982), .B(u2__abc_44228_n2983_bF_buf118), .Y(u2__abc_44228_n8983_1) );
  OR2X2 OR2X2_1596 ( .A(u2__abc_44228_n8983_1), .B(u2__abc_44228_n8975), .Y(u2__abc_44228_n8984_1) );
  OR2X2 OR2X2_1597 ( .A(u2__abc_44228_n8988), .B(u2__abc_44228_n8974), .Y(u2__abc_44228_n8989_1) );
  OR2X2 OR2X2_1598 ( .A(u2__abc_44228_n8993), .B(u2__abc_44228_n8992), .Y(u2__abc_44228_n8994_1) );
  OR2X2 OR2X2_1599 ( .A(u2__abc_44228_n8995_1), .B(u2__abc_44228_n3989), .Y(u2__abc_44228_n8996) );
  OR2X2 OR2X2_16 ( .A(_abc_64468_n753_bF_buf0), .B(\a[7] ), .Y(_abc_64468_n852) );
  OR2X2 OR2X2_160 ( .A(_abc_64468_n753_bF_buf12), .B(\a[79] ), .Y(_abc_64468_n1068) );
  OR2X2 OR2X2_1600 ( .A(u2__abc_44228_n7548_1_bF_buf30), .B(u2__abc_44228_n8997), .Y(u2__abc_44228_n8998) );
  OR2X2 OR2X2_1601 ( .A(u2__abc_44228_n7547_bF_buf29), .B(u2_remHi_83_), .Y(u2__abc_44228_n8999) );
  OR2X2 OR2X2_1602 ( .A(u2__abc_44228_n9000_1), .B(u2__abc_44228_n2983_bF_buf116), .Y(u2__abc_44228_n9001) );
  OR2X2 OR2X2_1603 ( .A(u2__abc_44228_n9005_1), .B(u2__abc_44228_n8991), .Y(u2__abc_44228_n9006_1) );
  OR2X2 OR2X2_1604 ( .A(u2__abc_44228_n9009), .B(u2__abc_44228_n4191), .Y(u2__abc_44228_n9010) );
  OR2X2 OR2X2_1605 ( .A(u2__abc_44228_n9010), .B(u2__abc_44228_n3975), .Y(u2__abc_44228_n9011_1) );
  OR2X2 OR2X2_1606 ( .A(u2__abc_44228_n7548_1_bF_buf29), .B(u2__abc_44228_n9014), .Y(u2__abc_44228_n9015) );
  OR2X2 OR2X2_1607 ( .A(u2__abc_44228_n7547_bF_buf28), .B(u2_remHi_84_), .Y(u2__abc_44228_n9016_1) );
  OR2X2 OR2X2_1608 ( .A(u2__abc_44228_n9017_1), .B(u2__abc_44228_n2983_bF_buf114), .Y(u2__abc_44228_n9018) );
  OR2X2 OR2X2_1609 ( .A(u2__abc_44228_n9022_1), .B(u2__abc_44228_n9008), .Y(u2__abc_44228_n9023) );
  OR2X2 OR2X2_161 ( .A(aNan_bF_buf6), .B(sqrto_156_), .Y(_abc_64468_n1070) );
  OR2X2 OR2X2_1610 ( .A(u2__abc_44228_n9012), .B(u2__abc_44228_n3971), .Y(u2__abc_44228_n9026) );
  OR2X2 OR2X2_1611 ( .A(u2__abc_44228_n9026), .B(u2__abc_44228_n3969), .Y(u2__abc_44228_n9027_1) );
  OR2X2 OR2X2_1612 ( .A(u2__abc_44228_n9029), .B(u2__abc_44228_n9028_1), .Y(u2__abc_44228_n9030) );
  OR2X2 OR2X2_1613 ( .A(u2__abc_44228_n9033_1), .B(u2__abc_44228_n2983_bF_buf112), .Y(u2__abc_44228_n9034) );
  OR2X2 OR2X2_1614 ( .A(u2__abc_44228_n9034), .B(u2__abc_44228_n9032), .Y(u2__abc_44228_n9035) );
  OR2X2 OR2X2_1615 ( .A(u2__abc_44228_n9039_1), .B(u2__abc_44228_n9025), .Y(u2__abc_44228_n9040) );
  OR2X2 OR2X2_1616 ( .A(u2__abc_44228_n9044_1), .B(u2__abc_44228_n4196), .Y(u2__abc_44228_n9045) );
  OR2X2 OR2X2_1617 ( .A(u2__abc_44228_n9045), .B(u2__abc_44228_n3952), .Y(u2__abc_44228_n9046) );
  OR2X2 OR2X2_1618 ( .A(u2__abc_44228_n9050_1), .B(u2__abc_44228_n2983_bF_buf110), .Y(u2__abc_44228_n9051) );
  OR2X2 OR2X2_1619 ( .A(u2__abc_44228_n9051), .B(u2__abc_44228_n9043), .Y(u2__abc_44228_n9052) );
  OR2X2 OR2X2_162 ( .A(_abc_64468_n753_bF_buf11), .B(\a[80] ), .Y(_abc_64468_n1071) );
  OR2X2 OR2X2_1620 ( .A(u2__abc_44228_n9056), .B(u2__abc_44228_n9042), .Y(u2__abc_44228_n9057) );
  OR2X2 OR2X2_1621 ( .A(u2__abc_44228_n9064), .B(u2__abc_44228_n9065), .Y(u2__abc_44228_n9066_1) );
  OR2X2 OR2X2_1622 ( .A(u2__abc_44228_n9067), .B(u2__abc_44228_n2983_bF_buf108), .Y(u2__abc_44228_n9068) );
  OR2X2 OR2X2_1623 ( .A(u2__abc_44228_n9068), .B(u2__abc_44228_n9060_1), .Y(u2__abc_44228_n9069) );
  OR2X2 OR2X2_1624 ( .A(u2__abc_44228_n9073), .B(u2__abc_44228_n9059), .Y(u2__abc_44228_n9074) );
  OR2X2 OR2X2_1625 ( .A(u2__abc_44228_n9077_1), .B(u2__abc_44228_n3957), .Y(u2__abc_44228_n9078) );
  OR2X2 OR2X2_1626 ( .A(u2__abc_44228_n9079), .B(u2__abc_44228_n3945), .Y(u2__abc_44228_n9080) );
  OR2X2 OR2X2_1627 ( .A(u2__abc_44228_n7548_1_bF_buf25), .B(u2__abc_44228_n9083_1), .Y(u2__abc_44228_n9084) );
  OR2X2 OR2X2_1628 ( .A(u2__abc_44228_n7547_bF_buf24), .B(u2_remHi_88_), .Y(u2__abc_44228_n9085) );
  OR2X2 OR2X2_1629 ( .A(u2__abc_44228_n9086), .B(u2__abc_44228_n2983_bF_buf106), .Y(u2__abc_44228_n9087) );
  OR2X2 OR2X2_163 ( .A(aNan_bF_buf5), .B(sqrto_157_), .Y(_abc_64468_n1073) );
  OR2X2 OR2X2_1630 ( .A(u2__abc_44228_n9091), .B(u2__abc_44228_n9076), .Y(u2__abc_44228_n9092) );
  OR2X2 OR2X2_1631 ( .A(u2__abc_44228_n9081), .B(u2__abc_44228_n3941), .Y(u2__abc_44228_n9096) );
  OR2X2 OR2X2_1632 ( .A(u2__abc_44228_n9097), .B(u2__abc_44228_n9095), .Y(u2__abc_44228_n9098) );
  OR2X2 OR2X2_1633 ( .A(u2__abc_44228_n9096), .B(u2__abc_44228_n3939), .Y(u2__abc_44228_n9099_1) );
  OR2X2 OR2X2_1634 ( .A(u2__abc_44228_n9102), .B(u2__abc_44228_n2983_bF_buf104), .Y(u2__abc_44228_n9103) );
  OR2X2 OR2X2_1635 ( .A(u2__abc_44228_n9101), .B(u2__abc_44228_n9103), .Y(u2__abc_44228_n9104_1) );
  OR2X2 OR2X2_1636 ( .A(u2__abc_44228_n9108), .B(u2__abc_44228_n9094_1), .Y(u2__abc_44228_n9109) );
  OR2X2 OR2X2_1637 ( .A(u2__abc_44228_n9112), .B(u2__abc_44228_n4205_1), .Y(u2__abc_44228_n9113) );
  OR2X2 OR2X2_1638 ( .A(u2__abc_44228_n9113), .B(u2__abc_44228_n3923), .Y(u2__abc_44228_n9116_1) );
  OR2X2 OR2X2_1639 ( .A(u2__abc_44228_n7548_1_bF_buf23), .B(u2__abc_44228_n9117), .Y(u2__abc_44228_n9118) );
  OR2X2 OR2X2_164 ( .A(_abc_64468_n753_bF_buf10), .B(\a[81] ), .Y(_abc_64468_n1074) );
  OR2X2 OR2X2_1640 ( .A(u2__abc_44228_n7547_bF_buf22), .B(u2_remHi_90_), .Y(u2__abc_44228_n9119) );
  OR2X2 OR2X2_1641 ( .A(u2__abc_44228_n9120), .B(u2__abc_44228_n2983_bF_buf102), .Y(u2__abc_44228_n9121_1) );
  OR2X2 OR2X2_1642 ( .A(u2__abc_44228_n9125), .B(u2__abc_44228_n9111), .Y(u2__abc_44228_n9126_1) );
  OR2X2 OR2X2_1643 ( .A(u2__abc_44228_n9133), .B(u2__abc_44228_n9130), .Y(u2__abc_44228_n9134) );
  OR2X2 OR2X2_1644 ( .A(u2__abc_44228_n9136), .B(u2__abc_44228_n2983_bF_buf100), .Y(u2__abc_44228_n9137_1) );
  OR2X2 OR2X2_1645 ( .A(u2__abc_44228_n9137_1), .B(u2__abc_44228_n9135), .Y(u2__abc_44228_n9138_1) );
  OR2X2 OR2X2_1646 ( .A(u2__abc_44228_n9142), .B(u2__abc_44228_n9128), .Y(u2__abc_44228_n9143_1) );
  OR2X2 OR2X2_1647 ( .A(u2__abc_44228_n9146), .B(u2__abc_44228_n3928), .Y(u2__abc_44228_n9147) );
  OR2X2 OR2X2_1648 ( .A(u2__abc_44228_n9148_1), .B(u2__abc_44228_n3916), .Y(u2__abc_44228_n9149_1) );
  OR2X2 OR2X2_1649 ( .A(u2__abc_44228_n9154_1), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n9155) );
  OR2X2 OR2X2_165 ( .A(aNan_bF_buf4), .B(sqrto_158_), .Y(_abc_64468_n1076) );
  OR2X2 OR2X2_1650 ( .A(u2__abc_44228_n9153), .B(u2__abc_44228_n9155), .Y(u2__abc_44228_n9156) );
  OR2X2 OR2X2_1651 ( .A(u2__abc_44228_n9160_1), .B(u2__abc_44228_n9145), .Y(u2__abc_44228_n9161) );
  OR2X2 OR2X2_1652 ( .A(u2__abc_44228_n9150), .B(u2__abc_44228_n3912_1), .Y(u2__abc_44228_n9165_1) );
  OR2X2 OR2X2_1653 ( .A(u2__abc_44228_n9166), .B(u2__abc_44228_n9164), .Y(u2__abc_44228_n9167) );
  OR2X2 OR2X2_1654 ( .A(u2__abc_44228_n9165_1), .B(u2__abc_44228_n3910), .Y(u2__abc_44228_n9168) );
  OR2X2 OR2X2_1655 ( .A(u2__abc_44228_n9171_1), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n9172) );
  OR2X2 OR2X2_1656 ( .A(u2__abc_44228_n9170_1), .B(u2__abc_44228_n9172), .Y(u2__abc_44228_n9173) );
  OR2X2 OR2X2_1657 ( .A(u2__abc_44228_n9177), .B(u2__abc_44228_n9163), .Y(u2__abc_44228_n9178) );
  OR2X2 OR2X2_1658 ( .A(u2__abc_44228_n9181_1), .B(u2__abc_44228_n4217), .Y(u2__abc_44228_n9182_1) );
  OR2X2 OR2X2_1659 ( .A(u2__abc_44228_n9182_1), .B(u2__abc_44228_n3891), .Y(u2__abc_44228_n9185) );
  OR2X2 OR2X2_166 ( .A(_abc_64468_n753_bF_buf9), .B(\a[82] ), .Y(_abc_64468_n1077) );
  OR2X2 OR2X2_1660 ( .A(u2__abc_44228_n9188), .B(u2__abc_44228_n9187_1), .Y(u2__abc_44228_n9189) );
  OR2X2 OR2X2_1661 ( .A(u2__abc_44228_n9189), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n9190) );
  OR2X2 OR2X2_1662 ( .A(u2__abc_44228_n9194), .B(u2__abc_44228_n9180), .Y(u2__abc_44228_n9195) );
  OR2X2 OR2X2_1663 ( .A(u2__abc_44228_n9202), .B(u2__abc_44228_n9199), .Y(u2__abc_44228_n9203_1) );
  OR2X2 OR2X2_1664 ( .A(u2__abc_44228_n9205), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n9206) );
  OR2X2 OR2X2_1665 ( .A(u2__abc_44228_n9206), .B(u2__abc_44228_n9204_1), .Y(u2__abc_44228_n9207) );
  OR2X2 OR2X2_1666 ( .A(u2__abc_44228_n9211), .B(u2__abc_44228_n9197), .Y(u2__abc_44228_n9212) );
  OR2X2 OR2X2_1667 ( .A(u2__abc_44228_n9215_1), .B(u2__abc_44228_n3896), .Y(u2__abc_44228_n9216) );
  OR2X2 OR2X2_1668 ( .A(u2__abc_44228_n9217), .B(u2__abc_44228_n3884), .Y(u2__abc_44228_n9218) );
  OR2X2 OR2X2_1669 ( .A(u2__abc_44228_n9223), .B(u2__abc_44228_n9222), .Y(u2__abc_44228_n9224) );
  OR2X2 OR2X2_167 ( .A(aNan_bF_buf3), .B(sqrto_159_), .Y(_abc_64468_n1079) );
  OR2X2 OR2X2_1670 ( .A(u2__abc_44228_n9224), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n9225_1) );
  OR2X2 OR2X2_1671 ( .A(u2__abc_44228_n9229), .B(u2__abc_44228_n9214_1), .Y(u2__abc_44228_n9230) );
  OR2X2 OR2X2_1672 ( .A(u2__abc_44228_n9219), .B(u2__abc_44228_n3880), .Y(u2__abc_44228_n9233) );
  OR2X2 OR2X2_1673 ( .A(u2__abc_44228_n9233), .B(u2__abc_44228_n3878), .Y(u2__abc_44228_n9234) );
  OR2X2 OR2X2_1674 ( .A(u2__abc_44228_n9236_1), .B(u2__abc_44228_n9235), .Y(u2__abc_44228_n9237_1) );
  OR2X2 OR2X2_1675 ( .A(u2__abc_44228_n9238), .B(u2__abc_44228_n7548_1_bF_buf16), .Y(u2__abc_44228_n9239) );
  OR2X2 OR2X2_1676 ( .A(u2__abc_44228_n7547_bF_buf15), .B(u2_remHi_97_), .Y(u2__abc_44228_n9240) );
  OR2X2 OR2X2_1677 ( .A(u2__abc_44228_n9241), .B(u2__abc_44228_n2983_bF_buf89), .Y(u2__abc_44228_n9242_1) );
  OR2X2 OR2X2_1678 ( .A(u2__abc_44228_n9246), .B(u2__abc_44228_n9232), .Y(u2__abc_44228_n9247_1) );
  OR2X2 OR2X2_1679 ( .A(u2__abc_44228_n9251), .B(u2__abc_44228_n4226), .Y(u2__abc_44228_n9252) );
  OR2X2 OR2X2_168 ( .A(_abc_64468_n753_bF_buf8), .B(\a[83] ), .Y(_abc_64468_n1080) );
  OR2X2 OR2X2_1680 ( .A(u2__abc_44228_n9252), .B(u2__abc_44228_n3862), .Y(u2__abc_44228_n9255) );
  OR2X2 OR2X2_1681 ( .A(u2__abc_44228_n9257), .B(u2__abc_44228_n2983_bF_buf87), .Y(u2__abc_44228_n9258_1) );
  OR2X2 OR2X2_1682 ( .A(u2__abc_44228_n9258_1), .B(u2__abc_44228_n9250), .Y(u2__abc_44228_n9259_1) );
  OR2X2 OR2X2_1683 ( .A(u2__abc_44228_n9263), .B(u2__abc_44228_n9249), .Y(u2__abc_44228_n9264_1) );
  OR2X2 OR2X2_1684 ( .A(u2__abc_44228_n9268), .B(u2__abc_44228_n9267), .Y(u2__abc_44228_n9269_1) );
  OR2X2 OR2X2_1685 ( .A(u2__abc_44228_n9270_1), .B(u2__abc_44228_n3869), .Y(u2__abc_44228_n9271) );
  OR2X2 OR2X2_1686 ( .A(u2__abc_44228_n7548_1_bF_buf14), .B(u2__abc_44228_n9272), .Y(u2__abc_44228_n9273) );
  OR2X2 OR2X2_1687 ( .A(u2__abc_44228_n7547_bF_buf13), .B(u2_remHi_99_), .Y(u2__abc_44228_n9274) );
  OR2X2 OR2X2_1688 ( .A(u2__abc_44228_n9275_1), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n9276) );
  OR2X2 OR2X2_1689 ( .A(u2__abc_44228_n9280_1), .B(u2__abc_44228_n9266), .Y(u2__abc_44228_n9281_1) );
  OR2X2 OR2X2_169 ( .A(aNan_bF_buf2), .B(sqrto_160_), .Y(_abc_64468_n1082) );
  OR2X2 OR2X2_1690 ( .A(u2__abc_44228_n9284), .B(u2__abc_44228_n4231), .Y(u2__abc_44228_n9285) );
  OR2X2 OR2X2_1691 ( .A(u2__abc_44228_n9285), .B(u2__abc_44228_n3855), .Y(u2__abc_44228_n9286_1) );
  OR2X2 OR2X2_1692 ( .A(u2__abc_44228_n7548_1_bF_buf13), .B(u2__abc_44228_n9289), .Y(u2__abc_44228_n9290) );
  OR2X2 OR2X2_1693 ( .A(u2__abc_44228_n7547_bF_buf12), .B(u2_remHi_100_), .Y(u2__abc_44228_n9291_1) );
  OR2X2 OR2X2_1694 ( .A(u2__abc_44228_n9292_1), .B(u2__abc_44228_n2983_bF_buf83), .Y(u2__abc_44228_n9293) );
  OR2X2 OR2X2_1695 ( .A(u2__abc_44228_n9297_1), .B(u2__abc_44228_n9283), .Y(u2__abc_44228_n9298) );
  OR2X2 OR2X2_1696 ( .A(u2__abc_44228_n9287), .B(u2__abc_44228_n3851), .Y(u2__abc_44228_n9301) );
  OR2X2 OR2X2_1697 ( .A(u2__abc_44228_n9301), .B(u2__abc_44228_n3849), .Y(u2__abc_44228_n9302_1) );
  OR2X2 OR2X2_1698 ( .A(u2__abc_44228_n9304), .B(u2__abc_44228_n9303_1), .Y(u2__abc_44228_n9305) );
  OR2X2 OR2X2_1699 ( .A(u2__abc_44228_n9308_1), .B(u2__abc_44228_n2983_bF_buf81), .Y(u2__abc_44228_n9309) );
  OR2X2 OR2X2_17 ( .A(aNan_bF_buf1), .B(sqrto_84_), .Y(_abc_64468_n854) );
  OR2X2 OR2X2_170 ( .A(_abc_64468_n753_bF_buf7), .B(\a[84] ), .Y(_abc_64468_n1083) );
  OR2X2 OR2X2_1700 ( .A(u2__abc_44228_n9309), .B(u2__abc_44228_n9307), .Y(u2__abc_44228_n9310) );
  OR2X2 OR2X2_1701 ( .A(u2__abc_44228_n9314_1), .B(u2__abc_44228_n9300), .Y(u2__abc_44228_n9315) );
  OR2X2 OR2X2_1702 ( .A(u2__abc_44228_n9319_1), .B(u2__abc_44228_n4236), .Y(u2__abc_44228_n9320) );
  OR2X2 OR2X2_1703 ( .A(u2__abc_44228_n9320), .B(u2__abc_44228_n3825_1), .Y(u2__abc_44228_n9321) );
  OR2X2 OR2X2_1704 ( .A(u2__abc_44228_n9325_1), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n9326) );
  OR2X2 OR2X2_1705 ( .A(u2__abc_44228_n9326), .B(u2__abc_44228_n9318), .Y(u2__abc_44228_n9327) );
  OR2X2 OR2X2_1706 ( .A(u2__abc_44228_n9331), .B(u2__abc_44228_n9317), .Y(u2__abc_44228_n9332) );
  OR2X2 OR2X2_1707 ( .A(u2__abc_44228_n9339), .B(u2__abc_44228_n9340), .Y(u2__abc_44228_n9341_1) );
  OR2X2 OR2X2_1708 ( .A(u2__abc_44228_n9342), .B(u2__abc_44228_n2983_bF_buf77), .Y(u2__abc_44228_n9343) );
  OR2X2 OR2X2_1709 ( .A(u2__abc_44228_n9343), .B(u2__abc_44228_n9335_1), .Y(u2__abc_44228_n9344) );
  OR2X2 OR2X2_171 ( .A(aNan_bF_buf1), .B(sqrto_161_), .Y(_abc_64468_n1085) );
  OR2X2 OR2X2_1710 ( .A(u2__abc_44228_n9348), .B(u2__abc_44228_n9334), .Y(u2__abc_44228_n9349) );
  OR2X2 OR2X2_1711 ( .A(u2__abc_44228_n9352_1), .B(u2__abc_44228_n4241), .Y(u2__abc_44228_n9353) );
  OR2X2 OR2X2_1712 ( .A(u2__abc_44228_n9353), .B(u2__abc_44228_n3839), .Y(u2__abc_44228_n9354) );
  OR2X2 OR2X2_1713 ( .A(u2__abc_44228_n7548_1_bF_buf9), .B(u2__abc_44228_n9357_1), .Y(u2__abc_44228_n9358_1) );
  OR2X2 OR2X2_1714 ( .A(u2__abc_44228_n7547_bF_buf8), .B(u2_remHi_104_), .Y(u2__abc_44228_n9359) );
  OR2X2 OR2X2_1715 ( .A(u2__abc_44228_n9360), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n9361) );
  OR2X2 OR2X2_1716 ( .A(u2__abc_44228_n9365), .B(u2__abc_44228_n9351), .Y(u2__abc_44228_n9366) );
  OR2X2 OR2X2_1717 ( .A(u2__abc_44228_n9370), .B(u2__abc_44228_n9369_1), .Y(u2__abc_44228_n9371) );
  OR2X2 OR2X2_1718 ( .A(u2__abc_44228_n9372), .B(u2__abc_44228_n3833), .Y(u2__abc_44228_n9373) );
  OR2X2 OR2X2_1719 ( .A(u2__abc_44228_n9376), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n9377) );
  OR2X2 OR2X2_172 ( .A(_abc_64468_n753_bF_buf6), .B(\a[85] ), .Y(_abc_64468_n1086) );
  OR2X2 OR2X2_1720 ( .A(u2__abc_44228_n9377), .B(u2__abc_44228_n9375), .Y(u2__abc_44228_n9378) );
  OR2X2 OR2X2_1721 ( .A(u2__abc_44228_n9382), .B(u2__abc_44228_n9368_1), .Y(u2__abc_44228_n9383) );
  OR2X2 OR2X2_1722 ( .A(u2__abc_44228_n9386), .B(u2__abc_44228_n3831), .Y(u2__abc_44228_n9387) );
  OR2X2 OR2X2_1723 ( .A(u2__abc_44228_n9388), .B(u2__abc_44228_n3803), .Y(u2__abc_44228_n9391_1) );
  OR2X2 OR2X2_1724 ( .A(u2__abc_44228_n9392), .B(u2__abc_44228_n7548_1_bF_buf7), .Y(u2__abc_44228_n9393) );
  OR2X2 OR2X2_1725 ( .A(u2__abc_44228_n7547_bF_buf6), .B(u2_remHi_106_), .Y(u2__abc_44228_n9394) );
  OR2X2 OR2X2_1726 ( .A(u2__abc_44228_n9395), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n9396_1) );
  OR2X2 OR2X2_1727 ( .A(u2__abc_44228_n9400), .B(u2__abc_44228_n9385_1), .Y(u2__abc_44228_n9401_1) );
  OR2X2 OR2X2_1728 ( .A(u2__abc_44228_n9408), .B(u2__abc_44228_n9405), .Y(u2__abc_44228_n9409) );
  OR2X2 OR2X2_1729 ( .A(u2__abc_44228_n9411), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n9412_1) );
  OR2X2 OR2X2_173 ( .A(aNan_bF_buf0), .B(sqrto_162_), .Y(_abc_64468_n1088) );
  OR2X2 OR2X2_1730 ( .A(u2__abc_44228_n9410), .B(u2__abc_44228_n9412_1), .Y(u2__abc_44228_n9413_1) );
  OR2X2 OR2X2_1731 ( .A(u2__abc_44228_n9417), .B(u2__abc_44228_n9403), .Y(u2__abc_44228_n9418_1) );
  OR2X2 OR2X2_1732 ( .A(u2__abc_44228_n9421), .B(u2__abc_44228_n3808), .Y(u2__abc_44228_n9422) );
  OR2X2 OR2X2_1733 ( .A(u2__abc_44228_n9423_1), .B(u2__abc_44228_n3796), .Y(u2__abc_44228_n9424_1) );
  OR2X2 OR2X2_1734 ( .A(u2__abc_44228_n9429_1), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n9430) );
  OR2X2 OR2X2_1735 ( .A(u2__abc_44228_n9428), .B(u2__abc_44228_n9430), .Y(u2__abc_44228_n9431) );
  OR2X2 OR2X2_1736 ( .A(u2__abc_44228_n9435_1), .B(u2__abc_44228_n9420), .Y(u2__abc_44228_n9436) );
  OR2X2 OR2X2_1737 ( .A(u2__abc_44228_n9425), .B(u2__abc_44228_n3792), .Y(u2__abc_44228_n9440_1) );
  OR2X2 OR2X2_1738 ( .A(u2__abc_44228_n9441), .B(u2__abc_44228_n9439), .Y(u2__abc_44228_n9442) );
  OR2X2 OR2X2_1739 ( .A(u2__abc_44228_n9440_1), .B(u2__abc_44228_n3790), .Y(u2__abc_44228_n9443) );
  OR2X2 OR2X2_174 ( .A(_abc_64468_n753_bF_buf5), .B(\a[86] ), .Y(_abc_64468_n1089) );
  OR2X2 OR2X2_1740 ( .A(u2__abc_44228_n9446_1), .B(u2__abc_44228_n2983_bF_buf66), .Y(u2__abc_44228_n9447) );
  OR2X2 OR2X2_1741 ( .A(u2__abc_44228_n9445_1), .B(u2__abc_44228_n9447), .Y(u2__abc_44228_n9448) );
  OR2X2 OR2X2_1742 ( .A(u2__abc_44228_n9452), .B(u2__abc_44228_n9438), .Y(u2__abc_44228_n9453) );
  OR2X2 OR2X2_1743 ( .A(u2__abc_44228_n9457_1), .B(u2__abc_44228_n4258), .Y(u2__abc_44228_n9458) );
  OR2X2 OR2X2_1744 ( .A(u2__abc_44228_n9458), .B(u2__abc_44228_n3772), .Y(u2__abc_44228_n9461) );
  OR2X2 OR2X2_1745 ( .A(u2__abc_44228_n9463), .B(u2__abc_44228_n2983_bF_buf64), .Y(u2__abc_44228_n9464) );
  OR2X2 OR2X2_1746 ( .A(u2__abc_44228_n9464), .B(u2__abc_44228_n9456_1), .Y(u2__abc_44228_n9465) );
  OR2X2 OR2X2_1747 ( .A(u2__abc_44228_n9469), .B(u2__abc_44228_n9455), .Y(u2__abc_44228_n9470) );
  OR2X2 OR2X2_1748 ( .A(u2__abc_44228_n9477), .B(u2__abc_44228_n9478_1), .Y(u2__abc_44228_n9479_1) );
  OR2X2 OR2X2_1749 ( .A(u2__abc_44228_n9480), .B(u2__abc_44228_n2983_bF_buf62), .Y(u2__abc_44228_n9481) );
  OR2X2 OR2X2_175 ( .A(aNan_bF_buf10), .B(sqrto_163_), .Y(_abc_64468_n1091) );
  OR2X2 OR2X2_1750 ( .A(u2__abc_44228_n9481), .B(u2__abc_44228_n9473_1), .Y(u2__abc_44228_n9482) );
  OR2X2 OR2X2_1751 ( .A(u2__abc_44228_n9486), .B(u2__abc_44228_n9472), .Y(u2__abc_44228_n9487) );
  OR2X2 OR2X2_1752 ( .A(u2__abc_44228_n9490_1), .B(u2__abc_44228_n3777), .Y(u2__abc_44228_n9491) );
  OR2X2 OR2X2_1753 ( .A(u2__abc_44228_n9492), .B(u2__abc_44228_n3765), .Y(u2__abc_44228_n9493) );
  OR2X2 OR2X2_1754 ( .A(u2__abc_44228_n7548_1_bF_buf1), .B(u2__abc_44228_n9496), .Y(u2__abc_44228_n9497) );
  OR2X2 OR2X2_1755 ( .A(u2__abc_44228_n7547_bF_buf0), .B(u2_remHi_112_), .Y(u2__abc_44228_n9498) );
  OR2X2 OR2X2_1756 ( .A(u2__abc_44228_n9499), .B(u2__abc_44228_n2983_bF_buf60), .Y(u2__abc_44228_n9500_1) );
  OR2X2 OR2X2_1757 ( .A(u2__abc_44228_n9504), .B(u2__abc_44228_n9489_1), .Y(u2__abc_44228_n9505) );
  OR2X2 OR2X2_1758 ( .A(u2__abc_44228_n9494), .B(u2__abc_44228_n3761), .Y(u2__abc_44228_n9509) );
  OR2X2 OR2X2_1759 ( .A(u2__abc_44228_n9510), .B(u2__abc_44228_n9508), .Y(u2__abc_44228_n9511_1) );
  OR2X2 OR2X2_176 ( .A(_abc_64468_n753_bF_buf4), .B(\a[87] ), .Y(_abc_64468_n1092) );
  OR2X2 OR2X2_1760 ( .A(u2__abc_44228_n9509), .B(u2__abc_44228_n3759_1), .Y(u2__abc_44228_n9512_1) );
  OR2X2 OR2X2_1761 ( .A(u2__abc_44228_n9515), .B(u2__abc_44228_n2983_bF_buf58), .Y(u2__abc_44228_n9516) );
  OR2X2 OR2X2_1762 ( .A(u2__abc_44228_n9514), .B(u2__abc_44228_n9516), .Y(u2__abc_44228_n9517_1) );
  OR2X2 OR2X2_1763 ( .A(u2__abc_44228_n9521), .B(u2__abc_44228_n9507), .Y(u2__abc_44228_n9522_1) );
  OR2X2 OR2X2_1764 ( .A(u2__abc_44228_n9525), .B(u2__abc_44228_n4285), .Y(u2__abc_44228_n9526) );
  OR2X2 OR2X2_1765 ( .A(u2__abc_44228_n9526), .B(u2__abc_44228_n3750_1), .Y(u2__abc_44228_n9529) );
  OR2X2 OR2X2_1766 ( .A(u2__abc_44228_n7548_1_bF_buf57), .B(u2__abc_44228_n9530), .Y(u2__abc_44228_n9531) );
  OR2X2 OR2X2_1767 ( .A(u2__abc_44228_n7547_bF_buf56), .B(u2_remHi_114_), .Y(u2__abc_44228_n9532) );
  OR2X2 OR2X2_1768 ( .A(u2__abc_44228_n9533_1), .B(u2__abc_44228_n2983_bF_buf56), .Y(u2__abc_44228_n9534_1) );
  OR2X2 OR2X2_1769 ( .A(u2__abc_44228_n9538), .B(u2__abc_44228_n9524), .Y(u2__abc_44228_n9539_1) );
  OR2X2 OR2X2_177 ( .A(aNan_bF_buf9), .B(sqrto_164_), .Y(_abc_64468_n1094) );
  OR2X2 OR2X2_1770 ( .A(u2__abc_44228_n9543), .B(u2__abc_44228_n3744), .Y(u2__abc_44228_n9544_1) );
  OR2X2 OR2X2_1771 ( .A(u2__abc_44228_n9542), .B(u2__abc_44228_n9545_1), .Y(u2__abc_44228_n9546) );
  OR2X2 OR2X2_1772 ( .A(u2__abc_44228_n9549), .B(u2__abc_44228_n2983_bF_buf54), .Y(u2__abc_44228_n9550_1) );
  OR2X2 OR2X2_1773 ( .A(u2__abc_44228_n9550_1), .B(u2__abc_44228_n9548), .Y(u2__abc_44228_n9551) );
  OR2X2 OR2X2_1774 ( .A(u2__abc_44228_n9555_1), .B(u2__abc_44228_n9541), .Y(u2__abc_44228_n9556_1) );
  OR2X2 OR2X2_1775 ( .A(u2__abc_44228_n9559), .B(u2__abc_44228_n4290), .Y(u2__abc_44228_n9560) );
  OR2X2 OR2X2_1776 ( .A(u2__abc_44228_n9560), .B(u2__abc_44228_n3736), .Y(u2__abc_44228_n9561_1) );
  OR2X2 OR2X2_1777 ( .A(u2__abc_44228_n7548_1_bF_buf55), .B(u2__abc_44228_n9564), .Y(u2__abc_44228_n9565) );
  OR2X2 OR2X2_1778 ( .A(u2__abc_44228_n7547_bF_buf54), .B(u2_remHi_116_), .Y(u2__abc_44228_n9566_1) );
  OR2X2 OR2X2_1779 ( .A(u2__abc_44228_n9567_1), .B(u2__abc_44228_n2983_bF_buf52), .Y(u2__abc_44228_n9568) );
  OR2X2 OR2X2_178 ( .A(_abc_64468_n753_bF_buf3), .B(\a[88] ), .Y(_abc_64468_n1095) );
  OR2X2 OR2X2_1780 ( .A(u2__abc_44228_n9572_1), .B(u2__abc_44228_n9558), .Y(u2__abc_44228_n9573) );
  OR2X2 OR2X2_1781 ( .A(u2__abc_44228_n9562), .B(u2__abc_44228_n3732_1), .Y(u2__abc_44228_n9577_1) );
  OR2X2 OR2X2_1782 ( .A(u2__abc_44228_n9578_1), .B(u2__abc_44228_n9576), .Y(u2__abc_44228_n9579) );
  OR2X2 OR2X2_1783 ( .A(u2__abc_44228_n9577_1), .B(u2__abc_44228_n3730), .Y(u2__abc_44228_n9580) );
  OR2X2 OR2X2_1784 ( .A(u2__abc_44228_n9583_1), .B(u2__abc_44228_n2983_bF_buf50), .Y(u2__abc_44228_n9584) );
  OR2X2 OR2X2_1785 ( .A(u2__abc_44228_n9582), .B(u2__abc_44228_n9584), .Y(u2__abc_44228_n9585) );
  OR2X2 OR2X2_1786 ( .A(u2__abc_44228_n9589_1), .B(u2__abc_44228_n9575), .Y(u2__abc_44228_n9590) );
  OR2X2 OR2X2_1787 ( .A(u2__abc_44228_n9593), .B(u2__abc_44228_n4295), .Y(u2__abc_44228_n9594_1) );
  OR2X2 OR2X2_1788 ( .A(u2__abc_44228_n9594_1), .B(u2__abc_44228_n3706), .Y(u2__abc_44228_n9595) );
  OR2X2 OR2X2_1789 ( .A(u2__abc_44228_n7548_1_bF_buf53), .B(u2__abc_44228_n9598), .Y(u2__abc_44228_n9599_1) );
  OR2X2 OR2X2_179 ( .A(aNan_bF_buf8), .B(sqrto_165_), .Y(_abc_64468_n1097) );
  OR2X2 OR2X2_1790 ( .A(u2__abc_44228_n7547_bF_buf52), .B(u2_remHi_118_), .Y(u2__abc_44228_n9600_1) );
  OR2X2 OR2X2_1791 ( .A(u2__abc_44228_n9601), .B(u2__abc_44228_n2983_bF_buf48), .Y(u2__abc_44228_n9602) );
  OR2X2 OR2X2_1792 ( .A(u2__abc_44228_n9606), .B(u2__abc_44228_n9592), .Y(u2__abc_44228_n9607) );
  OR2X2 OR2X2_1793 ( .A(u2__abc_44228_n9611_1), .B(u2__abc_44228_n9610_1), .Y(u2__abc_44228_n9612) );
  OR2X2 OR2X2_1794 ( .A(u2__abc_44228_n9613), .B(u2__abc_44228_n3700), .Y(u2__abc_44228_n9614) );
  OR2X2 OR2X2_1795 ( .A(u2__abc_44228_n9617), .B(u2__abc_44228_n2983_bF_buf46), .Y(u2__abc_44228_n9618) );
  OR2X2 OR2X2_1796 ( .A(u2__abc_44228_n9618), .B(u2__abc_44228_n9616_1), .Y(u2__abc_44228_n9619) );
  OR2X2 OR2X2_1797 ( .A(u2__abc_44228_n9623), .B(u2__abc_44228_n9609), .Y(u2__abc_44228_n9624) );
  OR2X2 OR2X2_1798 ( .A(u2__abc_44228_n9627_1), .B(u2__abc_44228_n4263), .Y(u2__abc_44228_n9628) );
  OR2X2 OR2X2_1799 ( .A(u2__abc_44228_n9628), .B(u2__abc_44228_n3720), .Y(u2__abc_44228_n9629) );
  OR2X2 OR2X2_18 ( .A(_abc_64468_n753_bF_buf13), .B(\a[8] ), .Y(_abc_64468_n855) );
  OR2X2 OR2X2_180 ( .A(_abc_64468_n753_bF_buf2), .B(\a[89] ), .Y(_abc_64468_n1098) );
  OR2X2 OR2X2_1800 ( .A(u2__abc_44228_n7548_1_bF_buf51), .B(u2__abc_44228_n9632_1), .Y(u2__abc_44228_n9633_1) );
  OR2X2 OR2X2_1801 ( .A(u2__abc_44228_n7547_bF_buf50), .B(u2_remHi_120_), .Y(u2__abc_44228_n9634) );
  OR2X2 OR2X2_1802 ( .A(u2__abc_44228_n9635), .B(u2__abc_44228_n2983_bF_buf44), .Y(u2__abc_44228_n9636) );
  OR2X2 OR2X2_1803 ( .A(u2__abc_44228_n9640), .B(u2__abc_44228_n9626), .Y(u2__abc_44228_n9641) );
  OR2X2 OR2X2_1804 ( .A(u2__abc_44228_n9630), .B(u2__abc_44228_n3716), .Y(u2__abc_44228_n9645) );
  OR2X2 OR2X2_1805 ( .A(u2__abc_44228_n9646), .B(u2__abc_44228_n9644_1), .Y(u2__abc_44228_n9647) );
  OR2X2 OR2X2_1806 ( .A(u2__abc_44228_n9645), .B(u2__abc_44228_n3714_1), .Y(u2__abc_44228_n9648) );
  OR2X2 OR2X2_1807 ( .A(u2__abc_44228_n9651), .B(u2__abc_44228_n2983_bF_buf42), .Y(u2__abc_44228_n9652) );
  OR2X2 OR2X2_1808 ( .A(u2__abc_44228_n9650), .B(u2__abc_44228_n9652), .Y(u2__abc_44228_n9653) );
  OR2X2 OR2X2_1809 ( .A(u2__abc_44228_n9657), .B(u2__abc_44228_n9643_1), .Y(u2__abc_44228_n9658) );
  OR2X2 OR2X2_181 ( .A(aNan_bF_buf7), .B(sqrto_166_), .Y(_abc_64468_n1100) );
  OR2X2 OR2X2_1810 ( .A(u2__abc_44228_n9661), .B(u2__abc_44228_n4267), .Y(u2__abc_44228_n9662) );
  OR2X2 OR2X2_1811 ( .A(u2__abc_44228_n9662), .B(u2__abc_44228_n3684), .Y(u2__abc_44228_n9665_1) );
  OR2X2 OR2X2_1812 ( .A(u2__abc_44228_n7548_1_bF_buf49), .B(u2__abc_44228_n9666_1), .Y(u2__abc_44228_n9667) );
  OR2X2 OR2X2_1813 ( .A(u2__abc_44228_n7547_bF_buf48), .B(u2_remHi_122_), .Y(u2__abc_44228_n9668) );
  OR2X2 OR2X2_1814 ( .A(u2__abc_44228_n9669), .B(u2__abc_44228_n2983_bF_buf40), .Y(u2__abc_44228_n9670) );
  OR2X2 OR2X2_1815 ( .A(u2__abc_44228_n9674), .B(u2__abc_44228_n9660_1), .Y(u2__abc_44228_n9675) );
  OR2X2 OR2X2_1816 ( .A(u2__abc_44228_n9682_1), .B(u2__abc_44228_n9679), .Y(u2__abc_44228_n9683) );
  OR2X2 OR2X2_1817 ( .A(u2__abc_44228_n9685), .B(u2__abc_44228_n2983_bF_buf38), .Y(u2__abc_44228_n9686) );
  OR2X2 OR2X2_1818 ( .A(u2__abc_44228_n9684), .B(u2__abc_44228_n9686), .Y(u2__abc_44228_n9687_1) );
  OR2X2 OR2X2_1819 ( .A(u2__abc_44228_n9691), .B(u2__abc_44228_n9677_1), .Y(u2__abc_44228_n9692) );
  OR2X2 OR2X2_182 ( .A(_abc_64468_n753_bF_buf1), .B(\a[90] ), .Y(_abc_64468_n1101) );
  OR2X2 OR2X2_1820 ( .A(u2__abc_44228_n9695), .B(u2__abc_44228_n3689), .Y(u2__abc_44228_n9696) );
  OR2X2 OR2X2_1821 ( .A(u2__abc_44228_n9697), .B(u2__abc_44228_n3677), .Y(u2__abc_44228_n9698_1) );
  OR2X2 OR2X2_1822 ( .A(u2__abc_44228_n9703), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n9704_1) );
  OR2X2 OR2X2_1823 ( .A(u2__abc_44228_n9702), .B(u2__abc_44228_n9704_1), .Y(u2__abc_44228_n9705) );
  OR2X2 OR2X2_1824 ( .A(u2__abc_44228_n9709_1), .B(u2__abc_44228_n9694), .Y(u2__abc_44228_n9710_1) );
  OR2X2 OR2X2_1825 ( .A(u2__abc_44228_n9699_1), .B(u2__abc_44228_n3673), .Y(u2__abc_44228_n9714) );
  OR2X2 OR2X2_1826 ( .A(u2__abc_44228_n9715_1), .B(u2__abc_44228_n9713), .Y(u2__abc_44228_n9716) );
  OR2X2 OR2X2_1827 ( .A(u2__abc_44228_n9714), .B(u2__abc_44228_n3671), .Y(u2__abc_44228_n9717) );
  OR2X2 OR2X2_1828 ( .A(u2__abc_44228_n9720_1), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n9721_1) );
  OR2X2 OR2X2_1829 ( .A(u2__abc_44228_n9719), .B(u2__abc_44228_n9721_1), .Y(u2__abc_44228_n9722) );
  OR2X2 OR2X2_183 ( .A(aNan_bF_buf6), .B(sqrto_167_), .Y(_abc_64468_n1103) );
  OR2X2 OR2X2_1830 ( .A(u2__abc_44228_n9726_1), .B(u2__abc_44228_n9712), .Y(u2__abc_44228_n9727) );
  OR2X2 OR2X2_1831 ( .A(u2__abc_44228_n4300_1), .B(u2__abc_44228_n5249), .Y(u2__abc_44228_n9732_1) );
  OR2X2 OR2X2_1832 ( .A(u2__abc_44228_n9735), .B(u2__abc_44228_n9734), .Y(u2__abc_44228_n9736) );
  OR2X2 OR2X2_1833 ( .A(u2__abc_44228_n9736), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n9737_1) );
  OR2X2 OR2X2_1834 ( .A(u2__abc_44228_n9741), .B(u2__abc_44228_n9729), .Y(u2__abc_44228_n9742_1) );
  OR2X2 OR2X2_1835 ( .A(u2__abc_44228_n9730), .B(u2__abc_44228_n5245), .Y(u2__abc_44228_n9746) );
  OR2X2 OR2X2_1836 ( .A(u2__abc_44228_n9749), .B(u2__abc_44228_n9747), .Y(u2__abc_44228_n9750) );
  OR2X2 OR2X2_1837 ( .A(u2__abc_44228_n9752), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n9753_1) );
  OR2X2 OR2X2_1838 ( .A(u2__abc_44228_n9753_1), .B(u2__abc_44228_n9751), .Y(u2__abc_44228_n9754_1) );
  OR2X2 OR2X2_1839 ( .A(u2__abc_44228_n9758), .B(u2__abc_44228_n9744), .Y(u2__abc_44228_n9759_1) );
  OR2X2 OR2X2_184 ( .A(_abc_64468_n753_bF_buf0), .B(\a[91] ), .Y(_abc_64468_n1104) );
  OR2X2 OR2X2_1840 ( .A(u2__abc_44228_n9763), .B(u2__abc_44228_n5259), .Y(u2__abc_44228_n9764_1) );
  OR2X2 OR2X2_1841 ( .A(u2__abc_44228_n9764_1), .B(u2__abc_44228_n5235), .Y(u2__abc_44228_n9765_1) );
  OR2X2 OR2X2_1842 ( .A(u2__abc_44228_n9769), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n9770_1) );
  OR2X2 OR2X2_1843 ( .A(u2__abc_44228_n9770_1), .B(u2__abc_44228_n9762), .Y(u2__abc_44228_n9771) );
  OR2X2 OR2X2_1844 ( .A(u2__abc_44228_n9775_1), .B(u2__abc_44228_n9761), .Y(u2__abc_44228_n9776_1) );
  OR2X2 OR2X2_1845 ( .A(u2__abc_44228_n9783), .B(u2__abc_44228_n9784), .Y(u2__abc_44228_n9785) );
  OR2X2 OR2X2_1846 ( .A(u2__abc_44228_n9786_1), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n9787_1) );
  OR2X2 OR2X2_1847 ( .A(u2__abc_44228_n9787_1), .B(u2__abc_44228_n9779), .Y(u2__abc_44228_n9788) );
  OR2X2 OR2X2_1848 ( .A(u2__abc_44228_n9792_1), .B(u2__abc_44228_n9778), .Y(u2__abc_44228_n9793) );
  OR2X2 OR2X2_1849 ( .A(u2__abc_44228_n9797_1), .B(u2__abc_44228_n5265), .Y(u2__abc_44228_n9798_1) );
  OR2X2 OR2X2_185 ( .A(aNan_bF_buf5), .B(sqrto_168_), .Y(_abc_64468_n1106) );
  OR2X2 OR2X2_1850 ( .A(u2__abc_44228_n9798_1), .B(u2__abc_44228_n5223), .Y(u2__abc_44228_n9801) );
  OR2X2 OR2X2_1851 ( .A(u2__abc_44228_n9803_1), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n9804) );
  OR2X2 OR2X2_1852 ( .A(u2__abc_44228_n9804), .B(u2__abc_44228_n9796), .Y(u2__abc_44228_n9805) );
  OR2X2 OR2X2_1853 ( .A(u2__abc_44228_n9809_1), .B(u2__abc_44228_n9795), .Y(u2__abc_44228_n9810) );
  OR2X2 OR2X2_1854 ( .A(u2__abc_44228_n9799), .B(u2__abc_44228_n5219), .Y(u2__abc_44228_n9815) );
  OR2X2 OR2X2_1855 ( .A(u2__abc_44228_n9818), .B(u2__abc_44228_n9816), .Y(u2__abc_44228_n9819_1) );
  OR2X2 OR2X2_1856 ( .A(u2__abc_44228_n9820_1), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n9821) );
  OR2X2 OR2X2_1857 ( .A(u2__abc_44228_n9821), .B(u2__abc_44228_n9813), .Y(u2__abc_44228_n9822) );
  OR2X2 OR2X2_1858 ( .A(u2__abc_44228_n9826), .B(u2__abc_44228_n9812), .Y(u2__abc_44228_n9827) );
  OR2X2 OR2X2_1859 ( .A(u2__abc_44228_n9830_1), .B(u2__abc_44228_n5268), .Y(u2__abc_44228_n9831_1) );
  OR2X2 OR2X2_186 ( .A(_abc_64468_n753_bF_buf13), .B(\a[92] ), .Y(_abc_64468_n1107) );
  OR2X2 OR2X2_1860 ( .A(u2__abc_44228_n9831_1), .B(u2__abc_44228_n5209), .Y(u2__abc_44228_n9832) );
  OR2X2 OR2X2_1861 ( .A(u2__abc_44228_n7548_1_bF_buf39), .B(u2__abc_44228_n9835), .Y(u2__abc_44228_n9836_1) );
  OR2X2 OR2X2_1862 ( .A(u2__abc_44228_n7547_bF_buf38), .B(u2_remHi_132_), .Y(u2__abc_44228_n9837) );
  OR2X2 OR2X2_1863 ( .A(u2__abc_44228_n9838), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n9839) );
  OR2X2 OR2X2_1864 ( .A(u2__abc_44228_n9843), .B(u2__abc_44228_n9829), .Y(u2__abc_44228_n9844) );
  OR2X2 OR2X2_1865 ( .A(u2__abc_44228_n9833), .B(u2__abc_44228_n5205), .Y(u2__abc_44228_n9847_1) );
  OR2X2 OR2X2_1866 ( .A(u2__abc_44228_n9847_1), .B(u2__abc_44228_n5203), .Y(u2__abc_44228_n9848) );
  OR2X2 OR2X2_1867 ( .A(u2__abc_44228_n9850), .B(u2__abc_44228_n9849), .Y(u2__abc_44228_n9851) );
  OR2X2 OR2X2_1868 ( .A(u2__abc_44228_n9854), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n9855) );
  OR2X2 OR2X2_1869 ( .A(u2__abc_44228_n9855), .B(u2__abc_44228_n9853_1), .Y(u2__abc_44228_n9856) );
  OR2X2 OR2X2_187 ( .A(aNan_bF_buf4), .B(sqrto_169_), .Y(_abc_64468_n1109) );
  OR2X2 OR2X2_1870 ( .A(u2__abc_44228_n9860), .B(u2__abc_44228_n9846), .Y(u2__abc_44228_n9861) );
  OR2X2 OR2X2_1871 ( .A(u2__abc_44228_n9865), .B(u2__abc_44228_n5273), .Y(u2__abc_44228_n9866) );
  OR2X2 OR2X2_1872 ( .A(u2__abc_44228_n9866), .B(u2__abc_44228_n5179), .Y(u2__abc_44228_n9867) );
  OR2X2 OR2X2_1873 ( .A(u2__abc_44228_n9871), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n9872) );
  OR2X2 OR2X2_1874 ( .A(u2__abc_44228_n9872), .B(u2__abc_44228_n9864_1), .Y(u2__abc_44228_n9873) );
  OR2X2 OR2X2_1875 ( .A(u2__abc_44228_n9877), .B(u2__abc_44228_n9863_1), .Y(u2__abc_44228_n9878) );
  OR2X2 OR2X2_1876 ( .A(u2__abc_44228_n9868), .B(u2__abc_44228_n5175), .Y(u2__abc_44228_n9883) );
  OR2X2 OR2X2_1877 ( .A(u2__abc_44228_n9886_1), .B(u2__abc_44228_n9884), .Y(u2__abc_44228_n9887) );
  OR2X2 OR2X2_1878 ( .A(u2__abc_44228_n9888), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n9889) );
  OR2X2 OR2X2_1879 ( .A(u2__abc_44228_n9889), .B(u2__abc_44228_n9881), .Y(u2__abc_44228_n9890) );
  OR2X2 OR2X2_188 ( .A(_abc_64468_n753_bF_buf12), .B(\a[93] ), .Y(_abc_64468_n1110) );
  OR2X2 OR2X2_1880 ( .A(u2__abc_44228_n9894), .B(u2__abc_44228_n9880_1), .Y(u2__abc_44228_n9895) );
  OR2X2 OR2X2_1881 ( .A(u2__abc_44228_n9898), .B(u2__abc_44228_n5276), .Y(u2__abc_44228_n9899) );
  OR2X2 OR2X2_1882 ( .A(u2__abc_44228_n9899), .B(u2__abc_44228_n5193), .Y(u2__abc_44228_n9900) );
  OR2X2 OR2X2_1883 ( .A(u2__abc_44228_n7548_1_bF_buf35), .B(u2__abc_44228_n9903), .Y(u2__abc_44228_n9904) );
  OR2X2 OR2X2_1884 ( .A(u2__abc_44228_n7547_bF_buf34), .B(u2_remHi_136_), .Y(u2__abc_44228_n9905) );
  OR2X2 OR2X2_1885 ( .A(u2__abc_44228_n9906), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n9907_1) );
  OR2X2 OR2X2_1886 ( .A(u2__abc_44228_n9911), .B(u2__abc_44228_n9897_1), .Y(u2__abc_44228_n9912) );
  OR2X2 OR2X2_1887 ( .A(u2__abc_44228_n9901), .B(u2__abc_44228_n5189), .Y(u2__abc_44228_n9916) );
  OR2X2 OR2X2_1888 ( .A(u2__abc_44228_n9917), .B(u2__abc_44228_n9915), .Y(u2__abc_44228_n9918_1) );
  OR2X2 OR2X2_1889 ( .A(u2__abc_44228_n9916), .B(u2__abc_44228_n5187), .Y(u2__abc_44228_n9919_1) );
  OR2X2 OR2X2_189 ( .A(aNan_bF_buf3), .B(sqrto_170_), .Y(_abc_64468_n1112) );
  OR2X2 OR2X2_1890 ( .A(u2__abc_44228_n9922), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n9923) );
  OR2X2 OR2X2_1891 ( .A(u2__abc_44228_n9923), .B(u2__abc_44228_n9921), .Y(u2__abc_44228_n9924_1) );
  OR2X2 OR2X2_1892 ( .A(u2__abc_44228_n9928), .B(u2__abc_44228_n9914), .Y(u2__abc_44228_n9929_1) );
  OR2X2 OR2X2_1893 ( .A(u2__abc_44228_n9932), .B(u2__abc_44228_n5280), .Y(u2__abc_44228_n9933) );
  OR2X2 OR2X2_1894 ( .A(u2__abc_44228_n9933), .B(u2__abc_44228_n5164_1), .Y(u2__abc_44228_n9936) );
  OR2X2 OR2X2_1895 ( .A(u2__abc_44228_n7548_1_bF_buf33), .B(u2__abc_44228_n9937), .Y(u2__abc_44228_n9938) );
  OR2X2 OR2X2_1896 ( .A(u2__abc_44228_n7547_bF_buf32), .B(u2_remHi_138_), .Y(u2__abc_44228_n9939) );
  OR2X2 OR2X2_1897 ( .A(u2__abc_44228_n9940_1), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n9941_1) );
  OR2X2 OR2X2_1898 ( .A(u2__abc_44228_n9945), .B(u2__abc_44228_n9931), .Y(u2__abc_44228_n9946_1) );
  OR2X2 OR2X2_1899 ( .A(u2__abc_44228_n9953), .B(u2__abc_44228_n9950), .Y(u2__abc_44228_n9954) );
  OR2X2 OR2X2_19 ( .A(aNan_bF_buf0), .B(sqrto_85_), .Y(_abc_64468_n857) );
  OR2X2 OR2X2_190 ( .A(_abc_64468_n753_bF_buf11), .B(\a[94] ), .Y(_abc_64468_n1113) );
  OR2X2 OR2X2_1900 ( .A(u2__abc_44228_n9956), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n9957_1) );
  OR2X2 OR2X2_1901 ( .A(u2__abc_44228_n9957_1), .B(u2__abc_44228_n9955), .Y(u2__abc_44228_n9958) );
  OR2X2 OR2X2_1902 ( .A(u2__abc_44228_n9962_1), .B(u2__abc_44228_n9948), .Y(u2__abc_44228_n9963_1) );
  OR2X2 OR2X2_1903 ( .A(u2__abc_44228_n9966), .B(u2__abc_44228_n5156), .Y(u2__abc_44228_n9967) );
  OR2X2 OR2X2_1904 ( .A(u2__abc_44228_n9968_1), .B(u2__abc_44228_n5150), .Y(u2__abc_44228_n9969) );
  OR2X2 OR2X2_1905 ( .A(u2__abc_44228_n9974_1), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n9975) );
  OR2X2 OR2X2_1906 ( .A(u2__abc_44228_n9973_1), .B(u2__abc_44228_n9975), .Y(u2__abc_44228_n9976) );
  OR2X2 OR2X2_1907 ( .A(u2__abc_44228_n9980), .B(u2__abc_44228_n9965), .Y(u2__abc_44228_n9981) );
  OR2X2 OR2X2_1908 ( .A(u2__abc_44228_n9970), .B(u2__abc_44228_n5146_1), .Y(u2__abc_44228_n9985_1) );
  OR2X2 OR2X2_1909 ( .A(u2__abc_44228_n9986), .B(u2__abc_44228_n9984_1), .Y(u2__abc_44228_n9987) );
  OR2X2 OR2X2_191 ( .A(aNan_bF_buf2), .B(sqrto_171_), .Y(_abc_64468_n1115) );
  OR2X2 OR2X2_1910 ( .A(u2__abc_44228_n9985_1), .B(u2__abc_44228_n5144), .Y(u2__abc_44228_n9988) );
  OR2X2 OR2X2_1911 ( .A(u2__abc_44228_n9991), .B(u2__abc_44228_n2983_bF_buf4), .Y(u2__abc_44228_n9992) );
  OR2X2 OR2X2_1912 ( .A(u2__abc_44228_n9990_1), .B(u2__abc_44228_n9992), .Y(u2__abc_44228_n9993) );
  OR2X2 OR2X2_1913 ( .A(u2__abc_44228_n9997), .B(u2__abc_44228_n9983), .Y(u2__abc_44228_n9998) );
  OR2X2 OR2X2_1914 ( .A(u2__abc_44228_n10002), .B(u2__abc_44228_n5291), .Y(u2__abc_44228_n10003) );
  OR2X2 OR2X2_1915 ( .A(u2__abc_44228_n10003), .B(u2__abc_44228_n5133), .Y(u2__abc_44228_n10006_1) );
  OR2X2 OR2X2_1916 ( .A(u2__abc_44228_n10008), .B(u2__abc_44228_n2983_bF_buf2), .Y(u2__abc_44228_n10009) );
  OR2X2 OR2X2_1917 ( .A(u2__abc_44228_n10009), .B(u2__abc_44228_n10001_1), .Y(u2__abc_44228_n10010) );
  OR2X2 OR2X2_1918 ( .A(u2__abc_44228_n10014), .B(u2__abc_44228_n10000), .Y(u2__abc_44228_n10015) );
  OR2X2 OR2X2_1919 ( .A(u2__abc_44228_n10004), .B(u2__abc_44228_n5129), .Y(u2__abc_44228_n10019) );
  OR2X2 OR2X2_192 ( .A(_abc_64468_n753_bF_buf10), .B(\a[95] ), .Y(_abc_64468_n1116) );
  OR2X2 OR2X2_1920 ( .A(u2__abc_44228_n10020), .B(u2__abc_44228_n10018_1), .Y(u2__abc_44228_n10021) );
  OR2X2 OR2X2_1921 ( .A(u2__abc_44228_n10019), .B(u2__abc_44228_n5127_1), .Y(u2__abc_44228_n10022) );
  OR2X2 OR2X2_1922 ( .A(u2__abc_44228_n10025), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n10026) );
  OR2X2 OR2X2_1923 ( .A(u2__abc_44228_n10026), .B(u2__abc_44228_n10024), .Y(u2__abc_44228_n10027) );
  OR2X2 OR2X2_1924 ( .A(u2__abc_44228_n10031), .B(u2__abc_44228_n10017_1), .Y(u2__abc_44228_n10032) );
  OR2X2 OR2X2_1925 ( .A(u2__abc_44228_n10035), .B(u2__abc_44228_n5294), .Y(u2__abc_44228_n10036) );
  OR2X2 OR2X2_1926 ( .A(u2__abc_44228_n10036), .B(u2__abc_44228_n5119), .Y(u2__abc_44228_n10037) );
  OR2X2 OR2X2_1927 ( .A(u2__abc_44228_n7548_1_bF_buf27), .B(u2__abc_44228_n10040_1), .Y(u2__abc_44228_n10041) );
  OR2X2 OR2X2_1928 ( .A(u2__abc_44228_n7547_bF_buf26), .B(u2_remHi_144_), .Y(u2__abc_44228_n10042) );
  OR2X2 OR2X2_1929 ( .A(u2__abc_44228_n10043), .B(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n10044) );
  OR2X2 OR2X2_193 ( .A(aNan_bF_buf1), .B(sqrto_172_), .Y(_abc_64468_n1118) );
  OR2X2 OR2X2_1930 ( .A(u2__abc_44228_n10048), .B(u2__abc_44228_n10034_1), .Y(u2__abc_44228_n10049) );
  OR2X2 OR2X2_1931 ( .A(u2__abc_44228_n10056_1), .B(u2__abc_44228_n10053), .Y(u2__abc_44228_n10057) );
  OR2X2 OR2X2_1932 ( .A(u2__abc_44228_n10059), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n10060) );
  OR2X2 OR2X2_1933 ( .A(u2__abc_44228_n10060), .B(u2__abc_44228_n10058), .Y(u2__abc_44228_n10061_1) );
  OR2X2 OR2X2_1934 ( .A(u2__abc_44228_n10065), .B(u2__abc_44228_n10051_1), .Y(u2__abc_44228_n10066) );
  OR2X2 OR2X2_1935 ( .A(u2__abc_44228_n10069), .B(u2__abc_44228_n5111), .Y(u2__abc_44228_n10070) );
  OR2X2 OR2X2_1936 ( .A(u2__abc_44228_n10071), .B(u2__abc_44228_n5097), .Y(u2__abc_44228_n10074) );
  OR2X2 OR2X2_1937 ( .A(u2__abc_44228_n10075), .B(u2__abc_44228_n7548_1_bF_buf25), .Y(u2__abc_44228_n10076) );
  OR2X2 OR2X2_1938 ( .A(u2__abc_44228_n7547_bF_buf24), .B(u2_remHi_146_), .Y(u2__abc_44228_n10077) );
  OR2X2 OR2X2_1939 ( .A(u2__abc_44228_n10078_1), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n10079) );
  OR2X2 OR2X2_194 ( .A(_abc_64468_n753_bF_buf9), .B(\a[96] ), .Y(_abc_64468_n1119) );
  OR2X2 OR2X2_1940 ( .A(u2__abc_44228_n10083_1), .B(u2__abc_44228_n10068), .Y(u2__abc_44228_n10084_1) );
  OR2X2 OR2X2_1941 ( .A(u2__abc_44228_n10088), .B(u2__abc_44228_n5104), .Y(u2__abc_44228_n10089_1) );
  OR2X2 OR2X2_1942 ( .A(u2__abc_44228_n10087), .B(u2__abc_44228_n10090), .Y(u2__abc_44228_n10091) );
  OR2X2 OR2X2_1943 ( .A(u2__abc_44228_n10094_1), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n10095_1) );
  OR2X2 OR2X2_1944 ( .A(u2__abc_44228_n10093), .B(u2__abc_44228_n10095_1), .Y(u2__abc_44228_n10096) );
  OR2X2 OR2X2_1945 ( .A(u2__abc_44228_n10100_1), .B(u2__abc_44228_n10086), .Y(u2__abc_44228_n10101) );
  OR2X2 OR2X2_1946 ( .A(u2__abc_44228_n10104), .B(u2__abc_44228_n5102), .Y(u2__abc_44228_n10105_1) );
  OR2X2 OR2X2_1947 ( .A(u2__abc_44228_n10106_1), .B(u2__abc_44228_n5090), .Y(u2__abc_44228_n10107) );
  OR2X2 OR2X2_1948 ( .A(u2__abc_44228_n10112), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n10113) );
  OR2X2 OR2X2_1949 ( .A(u2__abc_44228_n10111_1), .B(u2__abc_44228_n10113), .Y(u2__abc_44228_n10114) );
  OR2X2 OR2X2_195 ( .A(aNan_bF_buf0), .B(sqrto_173_), .Y(_abc_64468_n1121) );
  OR2X2 OR2X2_1950 ( .A(u2__abc_44228_n10118), .B(u2__abc_44228_n10103), .Y(u2__abc_44228_n10119) );
  OR2X2 OR2X2_1951 ( .A(u2__abc_44228_n10108), .B(u2__abc_44228_n5086), .Y(u2__abc_44228_n10123) );
  OR2X2 OR2X2_1952 ( .A(u2__abc_44228_n10124), .B(u2__abc_44228_n10122_1), .Y(u2__abc_44228_n10125) );
  OR2X2 OR2X2_1953 ( .A(u2__abc_44228_n10123), .B(u2__abc_44228_n5084), .Y(u2__abc_44228_n10126) );
  OR2X2 OR2X2_1954 ( .A(u2__abc_44228_n10129), .B(u2__abc_44228_n2983_bF_buf132), .Y(u2__abc_44228_n10130) );
  OR2X2 OR2X2_1955 ( .A(u2__abc_44228_n10128_1), .B(u2__abc_44228_n10130), .Y(u2__abc_44228_n10131) );
  OR2X2 OR2X2_1956 ( .A(u2__abc_44228_n10135), .B(u2__abc_44228_n10121), .Y(u2__abc_44228_n10136) );
  OR2X2 OR2X2_1957 ( .A(u2__abc_44228_n10139_1), .B(u2__abc_44228_n5310), .Y(u2__abc_44228_n10140) );
  OR2X2 OR2X2_1958 ( .A(u2__abc_44228_n10140), .B(u2__abc_44228_n5067), .Y(u2__abc_44228_n10141) );
  OR2X2 OR2X2_1959 ( .A(u2__abc_44228_n7548_1_bF_buf21), .B(u2__abc_44228_n10144_1), .Y(u2__abc_44228_n10145) );
  OR2X2 OR2X2_196 ( .A(_abc_64468_n753_bF_buf8), .B(\a[97] ), .Y(_abc_64468_n1122) );
  OR2X2 OR2X2_1960 ( .A(u2__abc_44228_n7547_bF_buf20), .B(u2_remHi_150_), .Y(u2__abc_44228_n10146) );
  OR2X2 OR2X2_1961 ( .A(u2__abc_44228_n10147), .B(u2__abc_44228_n2983_bF_buf130), .Y(u2__abc_44228_n10148) );
  OR2X2 OR2X2_1962 ( .A(u2__abc_44228_n10152), .B(u2__abc_44228_n10138_1), .Y(u2__abc_44228_n10153) );
  OR2X2 OR2X2_1963 ( .A(u2__abc_44228_n10160_1), .B(u2__abc_44228_n10157), .Y(u2__abc_44228_n10161_1) );
  OR2X2 OR2X2_1964 ( .A(u2__abc_44228_n10163), .B(u2__abc_44228_n2983_bF_buf128), .Y(u2__abc_44228_n10164) );
  OR2X2 OR2X2_1965 ( .A(u2__abc_44228_n10164), .B(u2__abc_44228_n10162), .Y(u2__abc_44228_n10165) );
  OR2X2 OR2X2_1966 ( .A(u2__abc_44228_n10169), .B(u2__abc_44228_n10155_1), .Y(u2__abc_44228_n10170) );
  OR2X2 OR2X2_1967 ( .A(u2__abc_44228_n10173), .B(u2__abc_44228_n5072), .Y(u2__abc_44228_n10174) );
  OR2X2 OR2X2_1968 ( .A(u2__abc_44228_n10175), .B(u2__abc_44228_n5060), .Y(u2__abc_44228_n10176) );
  OR2X2 OR2X2_1969 ( .A(u2__abc_44228_n10181), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n10182_1) );
  OR2X2 OR2X2_197 ( .A(aNan_bF_buf10), .B(sqrto_174_), .Y(_abc_64468_n1124) );
  OR2X2 OR2X2_1970 ( .A(u2__abc_44228_n10180), .B(u2__abc_44228_n10182_1), .Y(u2__abc_44228_n10183_1) );
  OR2X2 OR2X2_1971 ( .A(u2__abc_44228_n10187), .B(u2__abc_44228_n10172_1), .Y(u2__abc_44228_n10188_1) );
  OR2X2 OR2X2_1972 ( .A(u2__abc_44228_n10177_1), .B(u2__abc_44228_n5056), .Y(u2__abc_44228_n10192) );
  OR2X2 OR2X2_1973 ( .A(u2__abc_44228_n10193_1), .B(u2__abc_44228_n10191), .Y(u2__abc_44228_n10194_1) );
  OR2X2 OR2X2_1974 ( .A(u2__abc_44228_n10192), .B(u2__abc_44228_n5054), .Y(u2__abc_44228_n10195) );
  OR2X2 OR2X2_1975 ( .A(u2__abc_44228_n10198), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n10199_1) );
  OR2X2 OR2X2_1976 ( .A(u2__abc_44228_n10197), .B(u2__abc_44228_n10199_1), .Y(u2__abc_44228_n10200) );
  OR2X2 OR2X2_1977 ( .A(u2__abc_44228_n10204_1), .B(u2__abc_44228_n10190), .Y(u2__abc_44228_n10205_1) );
  OR2X2 OR2X2_1978 ( .A(u2__abc_44228_n10208), .B(u2__abc_44228_n5319), .Y(u2__abc_44228_n10209) );
  OR2X2 OR2X2_1979 ( .A(u2__abc_44228_n10209), .B(u2__abc_44228_n5045), .Y(u2__abc_44228_n10212) );
  OR2X2 OR2X2_198 ( .A(_abc_64468_n753_bF_buf7), .B(\a[98] ), .Y(_abc_64468_n1125) );
  OR2X2 OR2X2_1980 ( .A(u2__abc_44228_n7548_1_bF_buf17), .B(u2__abc_44228_n10213), .Y(u2__abc_44228_n10214) );
  OR2X2 OR2X2_1981 ( .A(u2__abc_44228_n7547_bF_buf16), .B(u2_remHi_154_), .Y(u2__abc_44228_n10215_1) );
  OR2X2 OR2X2_1982 ( .A(u2__abc_44228_n10216_1), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n10217) );
  OR2X2 OR2X2_1983 ( .A(u2__abc_44228_n10221_1), .B(u2__abc_44228_n10207), .Y(u2__abc_44228_n10222) );
  OR2X2 OR2X2_1984 ( .A(u2__abc_44228_n10226_1), .B(u2__abc_44228_n10225), .Y(u2__abc_44228_n10227_1) );
  OR2X2 OR2X2_1985 ( .A(u2__abc_44228_n10228), .B(u2__abc_44228_n5039), .Y(u2__abc_44228_n10229) );
  OR2X2 OR2X2_1986 ( .A(u2__abc_44228_n10232_1), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n10233) );
  OR2X2 OR2X2_1987 ( .A(u2__abc_44228_n10231), .B(u2__abc_44228_n10233), .Y(u2__abc_44228_n10234) );
  OR2X2 OR2X2_1988 ( .A(u2__abc_44228_n10238_1), .B(u2__abc_44228_n10224), .Y(u2__abc_44228_n10239) );
  OR2X2 OR2X2_1989 ( .A(u2__abc_44228_n10242), .B(u2__abc_44228_n5326), .Y(u2__abc_44228_n10243_1) );
  OR2X2 OR2X2_199 ( .A(aNan_bF_buf9), .B(sqrto_175_), .Y(_abc_64468_n1127) );
  OR2X2 OR2X2_1990 ( .A(u2__abc_44228_n10243_1), .B(u2__abc_44228_n5031), .Y(u2__abc_44228_n10244) );
  OR2X2 OR2X2_1991 ( .A(u2__abc_44228_n10249_1), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n10250) );
  OR2X2 OR2X2_1992 ( .A(u2__abc_44228_n10248_1), .B(u2__abc_44228_n10250), .Y(u2__abc_44228_n10251) );
  OR2X2 OR2X2_1993 ( .A(u2__abc_44228_n10255), .B(u2__abc_44228_n10241), .Y(u2__abc_44228_n10256) );
  OR2X2 OR2X2_1994 ( .A(u2__abc_44228_n10245), .B(u2__abc_44228_n5027), .Y(u2__abc_44228_n10260_1) );
  OR2X2 OR2X2_1995 ( .A(u2__abc_44228_n10261), .B(u2__abc_44228_n10259_1), .Y(u2__abc_44228_n10262) );
  OR2X2 OR2X2_1996 ( .A(u2__abc_44228_n10260_1), .B(u2__abc_44228_n5025), .Y(u2__abc_44228_n10263) );
  OR2X2 OR2X2_1997 ( .A(u2__abc_44228_n10266), .B(u2__abc_44228_n2983_bF_buf118), .Y(u2__abc_44228_n10267) );
  OR2X2 OR2X2_1998 ( .A(u2__abc_44228_n10265_1), .B(u2__abc_44228_n10267), .Y(u2__abc_44228_n10268) );
  OR2X2 OR2X2_1999 ( .A(u2__abc_44228_n10272), .B(u2__abc_44228_n10258), .Y(u2__abc_44228_n10273) );
  OR2X2 OR2X2_2 ( .A(_abc_64468_n753_bF_buf7), .B(\a[0] ), .Y(_abc_64468_n831_1) );
  OR2X2 OR2X2_20 ( .A(_abc_64468_n753_bF_buf12), .B(\a[9] ), .Y(_abc_64468_n858) );
  OR2X2 OR2X2_200 ( .A(_abc_64468_n753_bF_buf6), .B(\a[99] ), .Y(_abc_64468_n1128) );
  OR2X2 OR2X2_2000 ( .A(u2__abc_44228_n10277), .B(u2__abc_44228_n5331), .Y(u2__abc_44228_n10278) );
  OR2X2 OR2X2_2001 ( .A(u2__abc_44228_n10278), .B(u2__abc_44228_n5006), .Y(u2__abc_44228_n10279) );
  OR2X2 OR2X2_2002 ( .A(u2__abc_44228_n10283), .B(u2__abc_44228_n2983_bF_buf116), .Y(u2__abc_44228_n10284) );
  OR2X2 OR2X2_2003 ( .A(u2__abc_44228_n10284), .B(u2__abc_44228_n10276_1), .Y(u2__abc_44228_n10285) );
  OR2X2 OR2X2_2004 ( .A(u2__abc_44228_n10289), .B(u2__abc_44228_n10275), .Y(u2__abc_44228_n10290) );
  OR2X2 OR2X2_2005 ( .A(u2__abc_44228_n10280), .B(u2__abc_44228_n5002), .Y(u2__abc_44228_n10294) );
  OR2X2 OR2X2_2006 ( .A(u2__abc_44228_n10295), .B(u2__abc_44228_n10293_1), .Y(u2__abc_44228_n10296) );
  OR2X2 OR2X2_2007 ( .A(u2__abc_44228_n10294), .B(u2__abc_44228_n5013), .Y(u2__abc_44228_n10297) );
  OR2X2 OR2X2_2008 ( .A(u2__abc_44228_n10300), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n10301) );
  OR2X2 OR2X2_2009 ( .A(u2__abc_44228_n10301), .B(u2__abc_44228_n10299), .Y(u2__abc_44228_n10302) );
  OR2X2 OR2X2_201 ( .A(aNan_bF_buf8), .B(sqrto_176_), .Y(_abc_64468_n1130) );
  OR2X2 OR2X2_2010 ( .A(u2__abc_44228_n10306), .B(u2__abc_44228_n10292_1), .Y(u2__abc_44228_n10307) );
  OR2X2 OR2X2_2011 ( .A(u2__abc_44228_n10310), .B(u2__abc_44228_n5334), .Y(u2__abc_44228_n10311) );
  OR2X2 OR2X2_2012 ( .A(u2__abc_44228_n10311), .B(u2__abc_44228_n4999), .Y(u2__abc_44228_n10312) );
  OR2X2 OR2X2_2013 ( .A(u2__abc_44228_n7548_1_bF_buf11), .B(u2__abc_44228_n10315_1), .Y(u2__abc_44228_n10316) );
  OR2X2 OR2X2_2014 ( .A(u2__abc_44228_n7547_bF_buf10), .B(u2_remHi_160_), .Y(u2__abc_44228_n10317) );
  OR2X2 OR2X2_2015 ( .A(u2__abc_44228_n10318), .B(u2__abc_44228_n2983_bF_buf113), .Y(u2__abc_44228_n10319) );
  OR2X2 OR2X2_2016 ( .A(u2__abc_44228_n10323), .B(u2__abc_44228_n10309_1), .Y(u2__abc_44228_n10324) );
  OR2X2 OR2X2_2017 ( .A(u2__abc_44228_n10313), .B(u2__abc_44228_n4995), .Y(u2__abc_44228_n10327) );
  OR2X2 OR2X2_2018 ( .A(u2__abc_44228_n10327), .B(u2__abc_44228_n4993), .Y(u2__abc_44228_n10328) );
  OR2X2 OR2X2_2019 ( .A(u2__abc_44228_n10330), .B(u2__abc_44228_n10329), .Y(u2__abc_44228_n10331) );
  OR2X2 OR2X2_202 ( .A(_abc_64468_n753_bF_buf5), .B(\a[100] ), .Y(_abc_64468_n1131) );
  OR2X2 OR2X2_2020 ( .A(u2__abc_44228_n10334), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n10335) );
  OR2X2 OR2X2_2021 ( .A(u2__abc_44228_n10335), .B(u2__abc_44228_n10333_1), .Y(u2__abc_44228_n10336) );
  OR2X2 OR2X2_2022 ( .A(u2__abc_44228_n10340_1), .B(u2__abc_44228_n10326_1), .Y(u2__abc_44228_n10341) );
  OR2X2 OR2X2_2023 ( .A(u2__abc_44228_n10344), .B(u2__abc_44228_n5338), .Y(u2__abc_44228_n10345) );
  OR2X2 OR2X2_2024 ( .A(u2__abc_44228_n10345), .B(u2__abc_44228_n4977), .Y(u2__abc_44228_n10348) );
  OR2X2 OR2X2_2025 ( .A(u2__abc_44228_n7548_1_bF_buf9), .B(u2__abc_44228_n10349), .Y(u2__abc_44228_n10350) );
  OR2X2 OR2X2_2026 ( .A(u2__abc_44228_n7547_bF_buf8), .B(u2_remHi_162_), .Y(u2__abc_44228_n10351) );
  OR2X2 OR2X2_2027 ( .A(u2__abc_44228_n10352), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n10353_1) );
  OR2X2 OR2X2_2028 ( .A(u2__abc_44228_n10357), .B(u2__abc_44228_n10343), .Y(u2__abc_44228_n10358) );
  OR2X2 OR2X2_2029 ( .A(u2__abc_44228_n10365), .B(u2__abc_44228_n10362), .Y(u2__abc_44228_n10366) );
  OR2X2 OR2X2_203 ( .A(aNan_bF_buf7), .B(sqrto_177_), .Y(_abc_64468_n1133) );
  OR2X2 OR2X2_2030 ( .A(u2__abc_44228_n10368_1), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n10369) );
  OR2X2 OR2X2_2031 ( .A(u2__abc_44228_n10369), .B(u2__abc_44228_n10367_1), .Y(u2__abc_44228_n10370) );
  OR2X2 OR2X2_2032 ( .A(u2__abc_44228_n10374_1), .B(u2__abc_44228_n10360_1), .Y(u2__abc_44228_n10375_1) );
  OR2X2 OR2X2_2033 ( .A(u2__abc_44228_n10378), .B(u2__abc_44228_n4982), .Y(u2__abc_44228_n10379) );
  OR2X2 OR2X2_2034 ( .A(u2__abc_44228_n10380), .B(u2__abc_44228_n4970), .Y(u2__abc_44228_n10381_1) );
  OR2X2 OR2X2_2035 ( .A(u2__abc_44228_n10386), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n10387) );
  OR2X2 OR2X2_2036 ( .A(u2__abc_44228_n10385), .B(u2__abc_44228_n10387), .Y(u2__abc_44228_n10388_1) );
  OR2X2 OR2X2_2037 ( .A(u2__abc_44228_n10392), .B(u2__abc_44228_n10377), .Y(u2__abc_44228_n10393) );
  OR2X2 OR2X2_2038 ( .A(u2__abc_44228_n10382_1), .B(u2__abc_44228_n4966), .Y(u2__abc_44228_n10397) );
  OR2X2 OR2X2_2039 ( .A(u2__abc_44228_n10398), .B(u2__abc_44228_n10396_1), .Y(u2__abc_44228_n10399) );
  OR2X2 OR2X2_204 ( .A(_abc_64468_n753_bF_buf4), .B(\a[101] ), .Y(_abc_64468_n1134) );
  OR2X2 OR2X2_2040 ( .A(u2__abc_44228_n10397), .B(u2__abc_44228_n4964), .Y(u2__abc_44228_n10400) );
  OR2X2 OR2X2_2041 ( .A(u2__abc_44228_n10403_1), .B(u2__abc_44228_n2983_bF_buf104), .Y(u2__abc_44228_n10404) );
  OR2X2 OR2X2_2042 ( .A(u2__abc_44228_n10402_1), .B(u2__abc_44228_n10404), .Y(u2__abc_44228_n10405) );
  OR2X2 OR2X2_2043 ( .A(u2__abc_44228_n10409_1), .B(u2__abc_44228_n10395_1), .Y(u2__abc_44228_n10410_1) );
  OR2X2 OR2X2_2044 ( .A(u2__abc_44228_n10413), .B(u2__abc_44228_n5348), .Y(u2__abc_44228_n10414) );
  OR2X2 OR2X2_2045 ( .A(u2__abc_44228_n10414), .B(u2__abc_44228_n4947), .Y(u2__abc_44228_n10415) );
  OR2X2 OR2X2_2046 ( .A(u2__abc_44228_n7548_1_bF_buf5), .B(u2__abc_44228_n10418), .Y(u2__abc_44228_n10419) );
  OR2X2 OR2X2_2047 ( .A(u2__abc_44228_n7547_bF_buf4), .B(u2_remHi_166_), .Y(u2__abc_44228_n10420) );
  OR2X2 OR2X2_2048 ( .A(u2__abc_44228_n10421), .B(u2__abc_44228_n2983_bF_buf102), .Y(u2__abc_44228_n10422) );
  OR2X2 OR2X2_2049 ( .A(u2__abc_44228_n10426), .B(u2__abc_44228_n10412), .Y(u2__abc_44228_n10427) );
  OR2X2 OR2X2_205 ( .A(aNan_bF_buf6), .B(sqrto_178_), .Y(_abc_64468_n1136) );
  OR2X2 OR2X2_2050 ( .A(u2__abc_44228_n10434), .B(u2__abc_44228_n10431_1), .Y(u2__abc_44228_n10435) );
  OR2X2 OR2X2_2051 ( .A(u2__abc_44228_n10437_1), .B(u2__abc_44228_n2983_bF_buf100), .Y(u2__abc_44228_n10438_1) );
  OR2X2 OR2X2_2052 ( .A(u2__abc_44228_n10438_1), .B(u2__abc_44228_n10436), .Y(u2__abc_44228_n10439) );
  OR2X2 OR2X2_2053 ( .A(u2__abc_44228_n10443), .B(u2__abc_44228_n10429), .Y(u2__abc_44228_n10444_1) );
  OR2X2 OR2X2_2054 ( .A(u2__abc_44228_n10447), .B(u2__abc_44228_n4952), .Y(u2__abc_44228_n10448) );
  OR2X2 OR2X2_2055 ( .A(u2__abc_44228_n10449), .B(u2__abc_44228_n4940), .Y(u2__abc_44228_n10450) );
  OR2X2 OR2X2_2056 ( .A(u2__abc_44228_n10455), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n10456) );
  OR2X2 OR2X2_2057 ( .A(u2__abc_44228_n10454), .B(u2__abc_44228_n10456), .Y(u2__abc_44228_n10457) );
  OR2X2 OR2X2_2058 ( .A(u2__abc_44228_n10461), .B(u2__abc_44228_n10446), .Y(u2__abc_44228_n10462) );
  OR2X2 OR2X2_2059 ( .A(u2__abc_44228_n10451_1), .B(u2__abc_44228_n4936), .Y(u2__abc_44228_n10466_1) );
  OR2X2 OR2X2_206 ( .A(_abc_64468_n753_bF_buf3), .B(\a[102] ), .Y(_abc_64468_n1137) );
  OR2X2 OR2X2_2060 ( .A(u2__abc_44228_n10467), .B(u2__abc_44228_n10465_1), .Y(u2__abc_44228_n10468) );
  OR2X2 OR2X2_2061 ( .A(u2__abc_44228_n10466_1), .B(u2__abc_44228_n4934), .Y(u2__abc_44228_n10469) );
  OR2X2 OR2X2_2062 ( .A(u2__abc_44228_n10472_1), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n10473_1) );
  OR2X2 OR2X2_2063 ( .A(u2__abc_44228_n10471), .B(u2__abc_44228_n10473_1), .Y(u2__abc_44228_n10474) );
  OR2X2 OR2X2_2064 ( .A(u2__abc_44228_n10478), .B(u2__abc_44228_n10464), .Y(u2__abc_44228_n10479_1) );
  OR2X2 OR2X2_2065 ( .A(u2__abc_44228_n10482), .B(u2__abc_44228_n5357), .Y(u2__abc_44228_n10483) );
  OR2X2 OR2X2_2066 ( .A(u2__abc_44228_n10483), .B(u2__abc_44228_n4918), .Y(u2__abc_44228_n10486_1) );
  OR2X2 OR2X2_2067 ( .A(u2__abc_44228_n7548_1_bF_buf1), .B(u2__abc_44228_n10487_1), .Y(u2__abc_44228_n10488) );
  OR2X2 OR2X2_2068 ( .A(u2__abc_44228_n7547_bF_buf0), .B(u2_remHi_170_), .Y(u2__abc_44228_n10489) );
  OR2X2 OR2X2_2069 ( .A(u2__abc_44228_n10490), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n10491) );
  OR2X2 OR2X2_207 ( .A(aNan_bF_buf5), .B(sqrto_179_), .Y(_abc_64468_n1139) );
  OR2X2 OR2X2_2070 ( .A(u2__abc_44228_n10495), .B(u2__abc_44228_n10481), .Y(u2__abc_44228_n10496) );
  OR2X2 OR2X2_2071 ( .A(u2__abc_44228_n10500_1), .B(u2__abc_44228_n4925), .Y(u2__abc_44228_n10501_1) );
  OR2X2 OR2X2_2072 ( .A(u2__abc_44228_n10499), .B(u2__abc_44228_n10502), .Y(u2__abc_44228_n10503) );
  OR2X2 OR2X2_2073 ( .A(u2__abc_44228_n10506), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n10507_1) );
  OR2X2 OR2X2_2074 ( .A(u2__abc_44228_n10505), .B(u2__abc_44228_n10507_1), .Y(u2__abc_44228_n10508_1) );
  OR2X2 OR2X2_2075 ( .A(u2__abc_44228_n10512), .B(u2__abc_44228_n10498), .Y(u2__abc_44228_n10513) );
  OR2X2 OR2X2_2076 ( .A(u2__abc_44228_n10516), .B(u2__abc_44228_n4923), .Y(u2__abc_44228_n10517) );
  OR2X2 OR2X2_2077 ( .A(u2__abc_44228_n10518), .B(u2__abc_44228_n4911_1), .Y(u2__abc_44228_n10519) );
  OR2X2 OR2X2_2078 ( .A(u2__abc_44228_n10524), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n10525) );
  OR2X2 OR2X2_2079 ( .A(u2__abc_44228_n10523), .B(u2__abc_44228_n10525), .Y(u2__abc_44228_n10526) );
  OR2X2 OR2X2_208 ( .A(_abc_64468_n753_bF_buf2), .B(\a[103] ), .Y(_abc_64468_n1140) );
  OR2X2 OR2X2_2080 ( .A(u2__abc_44228_n10530), .B(u2__abc_44228_n10515_1), .Y(u2__abc_44228_n10531) );
  OR2X2 OR2X2_2081 ( .A(u2__abc_44228_n10520), .B(u2__abc_44228_n4907), .Y(u2__abc_44228_n10535_1) );
  OR2X2 OR2X2_2082 ( .A(u2__abc_44228_n10536_1), .B(u2__abc_44228_n10534), .Y(u2__abc_44228_n10537) );
  OR2X2 OR2X2_2083 ( .A(u2__abc_44228_n10535_1), .B(u2__abc_44228_n4905), .Y(u2__abc_44228_n10538) );
  OR2X2 OR2X2_2084 ( .A(u2__abc_44228_n10541), .B(u2__abc_44228_n2983_bF_buf90), .Y(u2__abc_44228_n10542_1) );
  OR2X2 OR2X2_2085 ( .A(u2__abc_44228_n10540), .B(u2__abc_44228_n10542_1), .Y(u2__abc_44228_n10543_1) );
  OR2X2 OR2X2_2086 ( .A(u2__abc_44228_n10547), .B(u2__abc_44228_n10533), .Y(u2__abc_44228_n10548) );
  OR2X2 OR2X2_2087 ( .A(u2__abc_44228_n10551), .B(u2__abc_44228_n5368), .Y(u2__abc_44228_n10552) );
  OR2X2 OR2X2_2088 ( .A(u2__abc_44228_n10552), .B(u2__abc_44228_n4894), .Y(u2__abc_44228_n10555) );
  OR2X2 OR2X2_2089 ( .A(u2__abc_44228_n7548_1_bF_buf55), .B(u2__abc_44228_n10556_1), .Y(u2__abc_44228_n10557_1) );
  OR2X2 OR2X2_209 ( .A(aNan_bF_buf4), .B(sqrto_180_), .Y(_abc_64468_n1142) );
  OR2X2 OR2X2_2090 ( .A(u2__abc_44228_n7547_bF_buf54), .B(u2_remHi_174_), .Y(u2__abc_44228_n10558) );
  OR2X2 OR2X2_2091 ( .A(u2__abc_44228_n10559), .B(u2__abc_44228_n2983_bF_buf88), .Y(u2__abc_44228_n10560) );
  OR2X2 OR2X2_2092 ( .A(u2__abc_44228_n10564_1), .B(u2__abc_44228_n10550_1), .Y(u2__abc_44228_n10565) );
  OR2X2 OR2X2_2093 ( .A(u2__abc_44228_n10569), .B(u2__abc_44228_n4888), .Y(u2__abc_44228_n10570_1) );
  OR2X2 OR2X2_2094 ( .A(u2__abc_44228_n10568), .B(u2__abc_44228_n10571_1), .Y(u2__abc_44228_n10572) );
  OR2X2 OR2X2_2095 ( .A(u2__abc_44228_n10575), .B(u2__abc_44228_n2983_bF_buf86), .Y(u2__abc_44228_n10576) );
  OR2X2 OR2X2_2096 ( .A(u2__abc_44228_n10576), .B(u2__abc_44228_n10574), .Y(u2__abc_44228_n10577_1) );
  OR2X2 OR2X2_2097 ( .A(u2__abc_44228_n10581), .B(u2__abc_44228_n10567), .Y(u2__abc_44228_n10582) );
  OR2X2 OR2X2_2098 ( .A(u2__abc_44228_n10585_1), .B(u2__abc_44228_n5373), .Y(u2__abc_44228_n10586) );
  OR2X2 OR2X2_2099 ( .A(u2__abc_44228_n10586), .B(u2__abc_44228_n4880), .Y(u2__abc_44228_n10587) );
  OR2X2 OR2X2_21 ( .A(aNan_bF_buf10), .B(sqrto_86_), .Y(_abc_64468_n860) );
  OR2X2 OR2X2_210 ( .A(_abc_64468_n753_bF_buf1), .B(\a[104] ), .Y(_abc_64468_n1143) );
  OR2X2 OR2X2_2100 ( .A(u2__abc_44228_n7548_1_bF_buf53), .B(u2__abc_44228_n10590), .Y(u2__abc_44228_n10591_1) );
  OR2X2 OR2X2_2101 ( .A(u2__abc_44228_n7547_bF_buf52), .B(u2_remHi_176_), .Y(u2__abc_44228_n10592_1) );
  OR2X2 OR2X2_2102 ( .A(u2__abc_44228_n10593), .B(u2__abc_44228_n2983_bF_buf84), .Y(u2__abc_44228_n10594) );
  OR2X2 OR2X2_2103 ( .A(u2__abc_44228_n10598_1), .B(u2__abc_44228_n10584_1), .Y(u2__abc_44228_n10599_1) );
  OR2X2 OR2X2_2104 ( .A(u2__abc_44228_n10588), .B(u2__abc_44228_n4876), .Y(u2__abc_44228_n10603) );
  OR2X2 OR2X2_2105 ( .A(u2__abc_44228_n10604), .B(u2__abc_44228_n10602), .Y(u2__abc_44228_n10605_1) );
  OR2X2 OR2X2_2106 ( .A(u2__abc_44228_n10603), .B(u2__abc_44228_n4874), .Y(u2__abc_44228_n10606_1) );
  OR2X2 OR2X2_2107 ( .A(u2__abc_44228_n10609), .B(u2__abc_44228_n2983_bF_buf82), .Y(u2__abc_44228_n10610) );
  OR2X2 OR2X2_2108 ( .A(u2__abc_44228_n10608), .B(u2__abc_44228_n10610), .Y(u2__abc_44228_n10611) );
  OR2X2 OR2X2_2109 ( .A(u2__abc_44228_n10615), .B(u2__abc_44228_n10601), .Y(u2__abc_44228_n10616) );
  OR2X2 OR2X2_211 ( .A(aNan_bF_buf3), .B(sqrto_181_), .Y(_abc_64468_n1145) );
  OR2X2 OR2X2_2110 ( .A(u2__abc_44228_n10619_1), .B(u2__abc_44228_n5377), .Y(u2__abc_44228_n10620_1) );
  OR2X2 OR2X2_2111 ( .A(u2__abc_44228_n10620_1), .B(u2__abc_44228_n4865), .Y(u2__abc_44228_n10623) );
  OR2X2 OR2X2_2112 ( .A(u2__abc_44228_n7548_1_bF_buf51), .B(u2__abc_44228_n10624), .Y(u2__abc_44228_n10625) );
  OR2X2 OR2X2_2113 ( .A(u2__abc_44228_n7547_bF_buf50), .B(u2_remHi_178_), .Y(u2__abc_44228_n10626_1) );
  OR2X2 OR2X2_2114 ( .A(u2__abc_44228_n10627_1), .B(u2__abc_44228_n2983_bF_buf80), .Y(u2__abc_44228_n10628) );
  OR2X2 OR2X2_2115 ( .A(u2__abc_44228_n10632), .B(u2__abc_44228_n10618), .Y(u2__abc_44228_n10633_1) );
  OR2X2 OR2X2_2116 ( .A(u2__abc_44228_n10637), .B(u2__abc_44228_n10636), .Y(u2__abc_44228_n10638) );
  OR2X2 OR2X2_2117 ( .A(u2__abc_44228_n10639), .B(u2__abc_44228_n4859), .Y(u2__abc_44228_n10640_1) );
  OR2X2 OR2X2_2118 ( .A(u2__abc_44228_n10643), .B(u2__abc_44228_n2983_bF_buf78), .Y(u2__abc_44228_n10644) );
  OR2X2 OR2X2_2119 ( .A(u2__abc_44228_n10642), .B(u2__abc_44228_n10644), .Y(u2__abc_44228_n10645) );
  OR2X2 OR2X2_212 ( .A(_abc_64468_n753_bF_buf0), .B(\a[105] ), .Y(_abc_64468_n1146) );
  OR2X2 OR2X2_2120 ( .A(u2__abc_44228_n10649), .B(u2__abc_44228_n10635), .Y(u2__abc_44228_n10650) );
  OR2X2 OR2X2_2121 ( .A(u2__abc_44228_n10653), .B(u2__abc_44228_n5382), .Y(u2__abc_44228_n10654_1) );
  OR2X2 OR2X2_2122 ( .A(u2__abc_44228_n10654_1), .B(u2__abc_44228_n4851), .Y(u2__abc_44228_n10655_1) );
  OR2X2 OR2X2_2123 ( .A(u2__abc_44228_n10660), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n10661_1) );
  OR2X2 OR2X2_2124 ( .A(u2__abc_44228_n10659), .B(u2__abc_44228_n10661_1), .Y(u2__abc_44228_n10662_1) );
  OR2X2 OR2X2_2125 ( .A(u2__abc_44228_n10666), .B(u2__abc_44228_n10652), .Y(u2__abc_44228_n10667) );
  OR2X2 OR2X2_2126 ( .A(u2__abc_44228_n10656), .B(u2__abc_44228_n4847), .Y(u2__abc_44228_n10671) );
  OR2X2 OR2X2_2127 ( .A(u2__abc_44228_n10672), .B(u2__abc_44228_n10670), .Y(u2__abc_44228_n10673) );
  OR2X2 OR2X2_2128 ( .A(u2__abc_44228_n10671), .B(u2__abc_44228_n4845), .Y(u2__abc_44228_n10674) );
  OR2X2 OR2X2_2129 ( .A(u2__abc_44228_n10677), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n10678) );
  OR2X2 OR2X2_213 ( .A(aNan_bF_buf2), .B(sqrto_182_), .Y(_abc_64468_n1148) );
  OR2X2 OR2X2_2130 ( .A(u2__abc_44228_n10676_1), .B(u2__abc_44228_n10678), .Y(u2__abc_44228_n10679) );
  OR2X2 OR2X2_2131 ( .A(u2__abc_44228_n10683_1), .B(u2__abc_44228_n10669_1), .Y(u2__abc_44228_n10684) );
  OR2X2 OR2X2_2132 ( .A(u2__abc_44228_n10687), .B(u2__abc_44228_n5387), .Y(u2__abc_44228_n10688) );
  OR2X2 OR2X2_2133 ( .A(u2__abc_44228_n10688), .B(u2__abc_44228_n4821), .Y(u2__abc_44228_n10689_1) );
  OR2X2 OR2X2_2134 ( .A(u2__abc_44228_n7548_1_bF_buf47), .B(u2__abc_44228_n10692), .Y(u2__abc_44228_n10693) );
  OR2X2 OR2X2_2135 ( .A(u2__abc_44228_n7547_bF_buf46), .B(u2_remHi_182_), .Y(u2__abc_44228_n10694) );
  OR2X2 OR2X2_2136 ( .A(u2__abc_44228_n10695), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n10696_1) );
  OR2X2 OR2X2_2137 ( .A(u2__abc_44228_n10700), .B(u2__abc_44228_n10686), .Y(u2__abc_44228_n10701) );
  OR2X2 OR2X2_2138 ( .A(u2__abc_44228_n10705), .B(u2__abc_44228_n10704_1), .Y(u2__abc_44228_n10706) );
  OR2X2 OR2X2_2139 ( .A(u2__abc_44228_n10707), .B(u2__abc_44228_n4815), .Y(u2__abc_44228_n10708) );
  OR2X2 OR2X2_214 ( .A(_abc_64468_n753_bF_buf13), .B(\a[106] ), .Y(_abc_64468_n1149) );
  OR2X2 OR2X2_2140 ( .A(u2__abc_44228_n10711_1), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n10712) );
  OR2X2 OR2X2_2141 ( .A(u2__abc_44228_n10710_1), .B(u2__abc_44228_n10712), .Y(u2__abc_44228_n10713) );
  OR2X2 OR2X2_2142 ( .A(u2__abc_44228_n10717_1), .B(u2__abc_44228_n10703_1), .Y(u2__abc_44228_n10718_1) );
  OR2X2 OR2X2_2143 ( .A(u2__abc_44228_n10721), .B(u2__abc_44228_n5400_1), .Y(u2__abc_44228_n10722) );
  OR2X2 OR2X2_2144 ( .A(u2__abc_44228_n10722), .B(u2__abc_44228_n4835), .Y(u2__abc_44228_n10723) );
  OR2X2 OR2X2_2145 ( .A(u2__abc_44228_n10728), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n10729) );
  OR2X2 OR2X2_2146 ( .A(u2__abc_44228_n10727), .B(u2__abc_44228_n10729), .Y(u2__abc_44228_n10730) );
  OR2X2 OR2X2_2147 ( .A(u2__abc_44228_n10734), .B(u2__abc_44228_n10720), .Y(u2__abc_44228_n10735) );
  OR2X2 OR2X2_2148 ( .A(u2__abc_44228_n10739_1), .B(u2__abc_44228_n10738_1), .Y(u2__abc_44228_n10740) );
  OR2X2 OR2X2_2149 ( .A(u2__abc_44228_n10741), .B(u2__abc_44228_n4829), .Y(u2__abc_44228_n10742) );
  OR2X2 OR2X2_215 ( .A(aNan_bF_buf1), .B(sqrto_183_), .Y(_abc_64468_n1151) );
  OR2X2 OR2X2_2150 ( .A(u2__abc_44228_n10745_1), .B(u2__abc_44228_n2983_bF_buf68), .Y(u2__abc_44228_n10746_1) );
  OR2X2 OR2X2_2151 ( .A(u2__abc_44228_n10744), .B(u2__abc_44228_n10746_1), .Y(u2__abc_44228_n10747) );
  OR2X2 OR2X2_2152 ( .A(u2__abc_44228_n10751), .B(u2__abc_44228_n10737), .Y(u2__abc_44228_n10752_1) );
  OR2X2 OR2X2_2153 ( .A(u2__abc_44228_n10755), .B(u2__abc_44228_n4827_1), .Y(u2__abc_44228_n10756) );
  OR2X2 OR2X2_2154 ( .A(u2__abc_44228_n10757), .B(u2__abc_44228_n4806), .Y(u2__abc_44228_n10760_1) );
  OR2X2 OR2X2_2155 ( .A(u2__abc_44228_n10763), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n10764) );
  OR2X2 OR2X2_2156 ( .A(u2__abc_44228_n10762), .B(u2__abc_44228_n10764), .Y(u2__abc_44228_n10765) );
  OR2X2 OR2X2_2157 ( .A(u2__abc_44228_n10769), .B(u2__abc_44228_n10754), .Y(u2__abc_44228_n10770) );
  OR2X2 OR2X2_2158 ( .A(u2__abc_44228_n10774_1), .B(u2__abc_44228_n10773_1), .Y(u2__abc_44228_n10775) );
  OR2X2 OR2X2_2159 ( .A(u2__abc_44228_n10776), .B(u2__abc_44228_n4800), .Y(u2__abc_44228_n10777) );
  OR2X2 OR2X2_216 ( .A(_abc_64468_n753_bF_buf12), .B(\a[107] ), .Y(_abc_64468_n1152) );
  OR2X2 OR2X2_2160 ( .A(u2__abc_44228_n10780_1), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n10781_1) );
  OR2X2 OR2X2_2161 ( .A(u2__abc_44228_n10779), .B(u2__abc_44228_n10781_1), .Y(u2__abc_44228_n10782) );
  OR2X2 OR2X2_2162 ( .A(u2__abc_44228_n10786), .B(u2__abc_44228_n10772), .Y(u2__abc_44228_n10787_1) );
  OR2X2 OR2X2_2163 ( .A(u2__abc_44228_n10790), .B(u2__abc_44228_n5392), .Y(u2__abc_44228_n10791) );
  OR2X2 OR2X2_2164 ( .A(u2__abc_44228_n10791), .B(u2__abc_44228_n4792), .Y(u2__abc_44228_n10792) );
  OR2X2 OR2X2_2165 ( .A(u2__abc_44228_n10797), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n10798) );
  OR2X2 OR2X2_2166 ( .A(u2__abc_44228_n10796), .B(u2__abc_44228_n10798), .Y(u2__abc_44228_n10799) );
  OR2X2 OR2X2_2167 ( .A(u2__abc_44228_n10803), .B(u2__abc_44228_n10789), .Y(u2__abc_44228_n10804) );
  OR2X2 OR2X2_2168 ( .A(u2__abc_44228_n10793), .B(u2__abc_44228_n4788_1), .Y(u2__abc_44228_n10808_1) );
  OR2X2 OR2X2_2169 ( .A(u2__abc_44228_n10809_1), .B(u2__abc_44228_n10807), .Y(u2__abc_44228_n10810) );
  OR2X2 OR2X2_217 ( .A(aNan_bF_buf0), .B(sqrto_184_), .Y(_abc_64468_n1154) );
  OR2X2 OR2X2_2170 ( .A(u2__abc_44228_n10808_1), .B(u2__abc_44228_n4786), .Y(u2__abc_44228_n10811) );
  OR2X2 OR2X2_2171 ( .A(u2__abc_44228_n10814), .B(u2__abc_44228_n2983_bF_buf62), .Y(u2__abc_44228_n10815_1) );
  OR2X2 OR2X2_2172 ( .A(u2__abc_44228_n10813), .B(u2__abc_44228_n10815_1), .Y(u2__abc_44228_n10816_1) );
  OR2X2 OR2X2_2173 ( .A(u2__abc_44228_n10820), .B(u2__abc_44228_n10806), .Y(u2__abc_44228_n10821) );
  OR2X2 OR2X2_2174 ( .A(u2__abc_44228_n10825), .B(u2__abc_44228_n5411), .Y(u2__abc_44228_n10826) );
  OR2X2 OR2X2_2175 ( .A(u2__abc_44228_n10826), .B(u2__abc_44228_n4766), .Y(u2__abc_44228_n10829_1) );
  OR2X2 OR2X2_2176 ( .A(u2__abc_44228_n10831), .B(u2__abc_44228_n2983_bF_buf60), .Y(u2__abc_44228_n10832) );
  OR2X2 OR2X2_2177 ( .A(u2__abc_44228_n10832), .B(u2__abc_44228_n10824), .Y(u2__abc_44228_n10833) );
  OR2X2 OR2X2_2178 ( .A(u2__abc_44228_n10837_1), .B(u2__abc_44228_n10823_1), .Y(u2__abc_44228_n10838) );
  OR2X2 OR2X2_2179 ( .A(u2__abc_44228_n10827), .B(u2__abc_44228_n4762), .Y(u2__abc_44228_n10842) );
  OR2X2 OR2X2_218 ( .A(_abc_64468_n753_bF_buf11), .B(\a[108] ), .Y(_abc_64468_n1155) );
  OR2X2 OR2X2_2180 ( .A(u2__abc_44228_n10843_1), .B(u2__abc_44228_n10841), .Y(u2__abc_44228_n10844_1) );
  OR2X2 OR2X2_2181 ( .A(u2__abc_44228_n10842), .B(u2__abc_44228_n4773), .Y(u2__abc_44228_n10845) );
  OR2X2 OR2X2_2182 ( .A(u2__abc_44228_n10848), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n10849) );
  OR2X2 OR2X2_2183 ( .A(u2__abc_44228_n10849), .B(u2__abc_44228_n10847), .Y(u2__abc_44228_n10850_1) );
  OR2X2 OR2X2_2184 ( .A(u2__abc_44228_n10854), .B(u2__abc_44228_n10840), .Y(u2__abc_44228_n10855) );
  OR2X2 OR2X2_2185 ( .A(u2__abc_44228_n10858_1), .B(u2__abc_44228_n5414), .Y(u2__abc_44228_n10859) );
  OR2X2 OR2X2_2186 ( .A(u2__abc_44228_n10859), .B(u2__abc_44228_n4759), .Y(u2__abc_44228_n10860) );
  OR2X2 OR2X2_2187 ( .A(u2__abc_44228_n7548_1_bF_buf37), .B(u2__abc_44228_n10863), .Y(u2__abc_44228_n10864_1) );
  OR2X2 OR2X2_2188 ( .A(u2__abc_44228_n7547_bF_buf36), .B(u2_remHi_192_), .Y(u2__abc_44228_n10865_1) );
  OR2X2 OR2X2_2189 ( .A(u2__abc_44228_n10866), .B(u2__abc_44228_n2983_bF_buf57), .Y(u2__abc_44228_n10867) );
  OR2X2 OR2X2_219 ( .A(aNan_bF_buf10), .B(sqrto_185_), .Y(_abc_64468_n1157) );
  OR2X2 OR2X2_2190 ( .A(u2__abc_44228_n10871_1), .B(u2__abc_44228_n10857_1), .Y(u2__abc_44228_n10872_1) );
  OR2X2 OR2X2_2191 ( .A(u2__abc_44228_n10861), .B(u2__abc_44228_n4755), .Y(u2__abc_44228_n10875) );
  OR2X2 OR2X2_2192 ( .A(u2__abc_44228_n10877), .B(u2__abc_44228_n10879_1), .Y(u2__abc_44228_n10880) );
  OR2X2 OR2X2_2193 ( .A(u2__abc_44228_n10882), .B(u2__abc_44228_n2983_bF_buf55), .Y(u2__abc_44228_n10883) );
  OR2X2 OR2X2_2194 ( .A(u2__abc_44228_n10883), .B(u2__abc_44228_n10881), .Y(u2__abc_44228_n10884) );
  OR2X2 OR2X2_2195 ( .A(u2__abc_44228_n10888), .B(u2__abc_44228_n10874), .Y(u2__abc_44228_n10889) );
  OR2X2 OR2X2_2196 ( .A(u2__abc_44228_n10892_1), .B(u2__abc_44228_n5418), .Y(u2__abc_44228_n10893_1) );
  OR2X2 OR2X2_2197 ( .A(u2__abc_44228_n10893_1), .B(u2__abc_44228_n4744), .Y(u2__abc_44228_n10896) );
  OR2X2 OR2X2_2198 ( .A(u2__abc_44228_n7548_1_bF_buf35), .B(u2__abc_44228_n10897), .Y(u2__abc_44228_n10898) );
  OR2X2 OR2X2_2199 ( .A(u2__abc_44228_n7547_bF_buf34), .B(u2_remHi_194_), .Y(u2__abc_44228_n10899_1) );
  OR2X2 OR2X2_22 ( .A(_abc_64468_n753_bF_buf11), .B(\a[10] ), .Y(_abc_64468_n861) );
  OR2X2 OR2X2_220 ( .A(_abc_64468_n753_bF_buf10), .B(\a[109] ), .Y(_abc_64468_n1158) );
  OR2X2 OR2X2_2200 ( .A(u2__abc_44228_n10900_1), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n10901) );
  OR2X2 OR2X2_2201 ( .A(u2__abc_44228_n10905), .B(u2__abc_44228_n10891), .Y(u2__abc_44228_n10906_1) );
  OR2X2 OR2X2_2202 ( .A(u2__abc_44228_n10910), .B(u2__abc_44228_n10909), .Y(u2__abc_44228_n10911) );
  OR2X2 OR2X2_2203 ( .A(u2__abc_44228_n10912), .B(u2__abc_44228_n4738), .Y(u2__abc_44228_n10913_1) );
  OR2X2 OR2X2_2204 ( .A(u2__abc_44228_n10916), .B(u2__abc_44228_n2983_bF_buf51), .Y(u2__abc_44228_n10917) );
  OR2X2 OR2X2_2205 ( .A(u2__abc_44228_n10917), .B(u2__abc_44228_n10915), .Y(u2__abc_44228_n10918) );
  OR2X2 OR2X2_2206 ( .A(u2__abc_44228_n10922), .B(u2__abc_44228_n10908), .Y(u2__abc_44228_n10923) );
  OR2X2 OR2X2_2207 ( .A(u2__abc_44228_n10926), .B(u2__abc_44228_n5423), .Y(u2__abc_44228_n10927_1) );
  OR2X2 OR2X2_2208 ( .A(u2__abc_44228_n10927_1), .B(u2__abc_44228_n4730), .Y(u2__abc_44228_n10928_1) );
  OR2X2 OR2X2_2209 ( .A(u2__abc_44228_n7548_1_bF_buf33), .B(u2__abc_44228_n10931), .Y(u2__abc_44228_n10932) );
  OR2X2 OR2X2_221 ( .A(aNan_bF_buf9), .B(sqrto_186_), .Y(_abc_64468_n1160) );
  OR2X2 OR2X2_2210 ( .A(u2__abc_44228_n7547_bF_buf32), .B(u2_remHi_196_), .Y(u2__abc_44228_n10933) );
  OR2X2 OR2X2_2211 ( .A(u2__abc_44228_n10934_1), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n10935_1) );
  OR2X2 OR2X2_2212 ( .A(u2__abc_44228_n10939), .B(u2__abc_44228_n10925), .Y(u2__abc_44228_n10940) );
  OR2X2 OR2X2_2213 ( .A(u2__abc_44228_n10929), .B(u2__abc_44228_n4726), .Y(u2__abc_44228_n10944) );
  OR2X2 OR2X2_2214 ( .A(u2__abc_44228_n10945), .B(u2__abc_44228_n10943), .Y(u2__abc_44228_n10946) );
  OR2X2 OR2X2_2215 ( .A(u2__abc_44228_n10944), .B(u2__abc_44228_n4724), .Y(u2__abc_44228_n10947) );
  OR2X2 OR2X2_2216 ( .A(u2__abc_44228_n10950), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n10951) );
  OR2X2 OR2X2_2217 ( .A(u2__abc_44228_n10949_1), .B(u2__abc_44228_n10951), .Y(u2__abc_44228_n10952) );
  OR2X2 OR2X2_2218 ( .A(u2__abc_44228_n10956_1), .B(u2__abc_44228_n10942_1), .Y(u2__abc_44228_n10957) );
  OR2X2 OR2X2_2219 ( .A(u2__abc_44228_n10960), .B(u2__abc_44228_n5428_1), .Y(u2__abc_44228_n10961) );
  OR2X2 OR2X2_222 ( .A(_abc_64468_n753_bF_buf9), .B(\a[110] ), .Y(_abc_64468_n1161) );
  OR2X2 OR2X2_2220 ( .A(u2__abc_44228_n10961), .B(u2__abc_44228_n4707), .Y(u2__abc_44228_n10962_1) );
  OR2X2 OR2X2_2221 ( .A(u2__abc_44228_n7548_1_bF_buf31), .B(u2__abc_44228_n10965), .Y(u2__abc_44228_n10966) );
  OR2X2 OR2X2_2222 ( .A(u2__abc_44228_n7547_bF_buf30), .B(u2_remHi_198_), .Y(u2__abc_44228_n10967) );
  OR2X2 OR2X2_2223 ( .A(u2__abc_44228_n10968), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n10969_1) );
  OR2X2 OR2X2_2224 ( .A(u2__abc_44228_n10973), .B(u2__abc_44228_n10959), .Y(u2__abc_44228_n10974) );
  OR2X2 OR2X2_2225 ( .A(u2__abc_44228_n10978), .B(u2__abc_44228_n4714), .Y(u2__abc_44228_n10979) );
  OR2X2 OR2X2_2226 ( .A(u2__abc_44228_n10977_1), .B(u2__abc_44228_n10980), .Y(u2__abc_44228_n10981) );
  OR2X2 OR2X2_2227 ( .A(u2__abc_44228_n10984_1), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n10985) );
  OR2X2 OR2X2_2228 ( .A(u2__abc_44228_n10985), .B(u2__abc_44228_n10983_1), .Y(u2__abc_44228_n10986) );
  OR2X2 OR2X2_2229 ( .A(u2__abc_44228_n10990_1), .B(u2__abc_44228_n10976_1), .Y(u2__abc_44228_n10991_1) );
  OR2X2 OR2X2_223 ( .A(aNan_bF_buf8), .B(sqrto_187_), .Y(_abc_64468_n1163) );
  OR2X2 OR2X2_2230 ( .A(u2__abc_44228_n10994), .B(u2__abc_44228_n4712), .Y(u2__abc_44228_n10995) );
  OR2X2 OR2X2_2231 ( .A(u2__abc_44228_n10996), .B(u2__abc_44228_n4700), .Y(u2__abc_44228_n10997_1) );
  OR2X2 OR2X2_2232 ( .A(u2__abc_44228_n11002), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n11003) );
  OR2X2 OR2X2_2233 ( .A(u2__abc_44228_n11001), .B(u2__abc_44228_n11003), .Y(u2__abc_44228_n11004_1) );
  OR2X2 OR2X2_2234 ( .A(u2__abc_44228_n11008), .B(u2__abc_44228_n10993), .Y(u2__abc_44228_n11009) );
  OR2X2 OR2X2_2235 ( .A(u2__abc_44228_n10998_1), .B(u2__abc_44228_n4696), .Y(u2__abc_44228_n11013) );
  OR2X2 OR2X2_2236 ( .A(u2__abc_44228_n11014), .B(u2__abc_44228_n11012_1), .Y(u2__abc_44228_n11015) );
  OR2X2 OR2X2_2237 ( .A(u2__abc_44228_n11013), .B(u2__abc_44228_n4694), .Y(u2__abc_44228_n11016) );
  OR2X2 OR2X2_2238 ( .A(u2__abc_44228_n11019_1), .B(u2__abc_44228_n2983_bF_buf40), .Y(u2__abc_44228_n11020) );
  OR2X2 OR2X2_2239 ( .A(u2__abc_44228_n11018_1), .B(u2__abc_44228_n11020), .Y(u2__abc_44228_n11021) );
  OR2X2 OR2X2_224 ( .A(_abc_64468_n753_bF_buf8), .B(\a[111] ), .Y(_abc_64468_n1164) );
  OR2X2 OR2X2_2240 ( .A(u2__abc_44228_n11025_1), .B(u2__abc_44228_n11011_1), .Y(u2__abc_44228_n11026_1) );
  OR2X2 OR2X2_2241 ( .A(u2__abc_44228_n11029), .B(u2__abc_44228_n5437_1), .Y(u2__abc_44228_n11030) );
  OR2X2 OR2X2_2242 ( .A(u2__abc_44228_n11030), .B(u2__abc_44228_n4685_1), .Y(u2__abc_44228_n11033_1) );
  OR2X2 OR2X2_2243 ( .A(u2__abc_44228_n7548_1_bF_buf27), .B(u2__abc_44228_n11034), .Y(u2__abc_44228_n11035) );
  OR2X2 OR2X2_2244 ( .A(u2__abc_44228_n7547_bF_buf26), .B(u2_remHi_202_), .Y(u2__abc_44228_n11036) );
  OR2X2 OR2X2_2245 ( .A(u2__abc_44228_n11037), .B(u2__abc_44228_n2983_bF_buf38), .Y(u2__abc_44228_n11038) );
  OR2X2 OR2X2_2246 ( .A(u2__abc_44228_n11042), .B(u2__abc_44228_n11028), .Y(u2__abc_44228_n11043) );
  OR2X2 OR2X2_2247 ( .A(u2__abc_44228_n11047_1), .B(u2__abc_44228_n11046_1), .Y(u2__abc_44228_n11048) );
  OR2X2 OR2X2_2248 ( .A(u2__abc_44228_n11049), .B(u2__abc_44228_n4679), .Y(u2__abc_44228_n11050) );
  OR2X2 OR2X2_2249 ( .A(u2__abc_44228_n11053_1), .B(u2__abc_44228_n2983_bF_buf36), .Y(u2__abc_44228_n11054_1) );
  OR2X2 OR2X2_225 ( .A(aNan_bF_buf7), .B(sqrto_188_), .Y(_auto_iopadmap_cc_313_execute_65414_224_) );
  OR2X2 OR2X2_2250 ( .A(u2__abc_44228_n11052), .B(u2__abc_44228_n11054_1), .Y(u2__abc_44228_n11055) );
  OR2X2 OR2X2_2251 ( .A(u2__abc_44228_n11059), .B(u2__abc_44228_n11045), .Y(u2__abc_44228_n11060_1) );
  OR2X2 OR2X2_2252 ( .A(u2__abc_44228_n11063), .B(u2__abc_44228_n5442), .Y(u2__abc_44228_n11064) );
  OR2X2 OR2X2_2253 ( .A(u2__abc_44228_n11064), .B(u2__abc_44228_n4671), .Y(u2__abc_44228_n11065) );
  OR2X2 OR2X2_2254 ( .A(u2__abc_44228_n11070), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n11071) );
  OR2X2 OR2X2_2255 ( .A(u2__abc_44228_n11069), .B(u2__abc_44228_n11071), .Y(u2__abc_44228_n11072) );
  OR2X2 OR2X2_2256 ( .A(u2__abc_44228_n11076), .B(u2__abc_44228_n11062), .Y(u2__abc_44228_n11077) );
  OR2X2 OR2X2_2257 ( .A(u2__abc_44228_n11066), .B(u2__abc_44228_n4667), .Y(u2__abc_44228_n11081_1) );
  OR2X2 OR2X2_2258 ( .A(u2__abc_44228_n11082_1), .B(u2__abc_44228_n11080), .Y(u2__abc_44228_n11083) );
  OR2X2 OR2X2_2259 ( .A(u2__abc_44228_n11081_1), .B(u2__abc_44228_n4665_1), .Y(u2__abc_44228_n11084) );
  OR2X2 OR2X2_226 ( .A(a_112_bF_buf8), .B(\a[0] ), .Y(_abc_64468_n1169) );
  OR2X2 OR2X2_2260 ( .A(u2__abc_44228_n11087), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n11088_1) );
  OR2X2 OR2X2_2261 ( .A(u2__abc_44228_n11086), .B(u2__abc_44228_n11088_1), .Y(u2__abc_44228_n11089_1) );
  OR2X2 OR2X2_2262 ( .A(u2__abc_44228_n11093), .B(u2__abc_44228_n11079), .Y(u2__abc_44228_n11094) );
  OR2X2 OR2X2_2263 ( .A(u2__abc_44228_n11097), .B(u2__abc_44228_n5448), .Y(u2__abc_44228_n11098) );
  OR2X2 OR2X2_2264 ( .A(u2__abc_44228_n11098), .B(u2__abc_44228_n4654), .Y(u2__abc_44228_n11101) );
  OR2X2 OR2X2_2265 ( .A(u2__abc_44228_n7548_1_bF_buf23), .B(u2__abc_44228_n11102_1), .Y(u2__abc_44228_n11103_1) );
  OR2X2 OR2X2_2266 ( .A(u2__abc_44228_n7547_bF_buf22), .B(u2_remHi_206_), .Y(u2__abc_44228_n11104) );
  OR2X2 OR2X2_2267 ( .A(u2__abc_44228_n11105), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n11106) );
  OR2X2 OR2X2_2268 ( .A(u2__abc_44228_n11110_1), .B(u2__abc_44228_n11096_1), .Y(u2__abc_44228_n11111) );
  OR2X2 OR2X2_2269 ( .A(u2__abc_44228_n11115), .B(u2__abc_44228_n4648), .Y(u2__abc_44228_n11116_1) );
  OR2X2 OR2X2_227 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[1] ), .Y(_abc_64468_n1171) );
  OR2X2 OR2X2_2270 ( .A(u2__abc_44228_n11114), .B(u2__abc_44228_n11117_1), .Y(u2__abc_44228_n11118) );
  OR2X2 OR2X2_2271 ( .A(u2__abc_44228_n11121), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n11122) );
  OR2X2 OR2X2_2272 ( .A(u2__abc_44228_n11122), .B(u2__abc_44228_n11120), .Y(u2__abc_44228_n11123_1) );
  OR2X2 OR2X2_2273 ( .A(u2__abc_44228_n11127), .B(u2__abc_44228_n11113), .Y(u2__abc_44228_n11128) );
  OR2X2 OR2X2_2274 ( .A(u2__abc_44228_n11131_1), .B(u2__abc_44228_n5453), .Y(u2__abc_44228_n11132) );
  OR2X2 OR2X2_2275 ( .A(u2__abc_44228_n11132), .B(u2__abc_44228_n4640), .Y(u2__abc_44228_n11133) );
  OR2X2 OR2X2_2276 ( .A(u2__abc_44228_n7548_1_bF_buf21), .B(u2__abc_44228_n11136), .Y(u2__abc_44228_n11137_1) );
  OR2X2 OR2X2_2277 ( .A(u2__abc_44228_n7547_bF_buf20), .B(u2_remHi_208_), .Y(u2__abc_44228_n11138_1) );
  OR2X2 OR2X2_2278 ( .A(u2__abc_44228_n11139), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n11140) );
  OR2X2 OR2X2_2279 ( .A(u2__abc_44228_n11144_1), .B(u2__abc_44228_n11130_1), .Y(u2__abc_44228_n11145_1) );
  OR2X2 OR2X2_228 ( .A(a_112_bF_buf6), .B(\a[1] ), .Y(_abc_64468_n1173) );
  OR2X2 OR2X2_2280 ( .A(u2__abc_44228_n11134), .B(u2__abc_44228_n4636), .Y(u2__abc_44228_n11149) );
  OR2X2 OR2X2_2281 ( .A(u2__abc_44228_n11150), .B(u2__abc_44228_n11148), .Y(u2__abc_44228_n11151_1) );
  OR2X2 OR2X2_2282 ( .A(u2__abc_44228_n11149), .B(u2__abc_44228_n4634), .Y(u2__abc_44228_n11152_1) );
  OR2X2 OR2X2_2283 ( .A(u2__abc_44228_n11155), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n11156) );
  OR2X2 OR2X2_2284 ( .A(u2__abc_44228_n11154), .B(u2__abc_44228_n11156), .Y(u2__abc_44228_n11157) );
  OR2X2 OR2X2_2285 ( .A(u2__abc_44228_n11161), .B(u2__abc_44228_n11147), .Y(u2__abc_44228_n11162) );
  OR2X2 OR2X2_2286 ( .A(u2__abc_44228_n11165_1), .B(u2__abc_44228_n5457), .Y(u2__abc_44228_n11166_1) );
  OR2X2 OR2X2_2287 ( .A(u2__abc_44228_n11166_1), .B(u2__abc_44228_n4618), .Y(u2__abc_44228_n11169) );
  OR2X2 OR2X2_2288 ( .A(u2__abc_44228_n7548_1_bF_buf19), .B(u2__abc_44228_n11170), .Y(u2__abc_44228_n11171) );
  OR2X2 OR2X2_2289 ( .A(u2__abc_44228_n7547_bF_buf18), .B(u2_remHi_210_), .Y(u2__abc_44228_n11172_1) );
  OR2X2 OR2X2_229 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[2] ), .Y(_abc_64468_n1174) );
  OR2X2 OR2X2_2290 ( .A(u2__abc_44228_n11173_1), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n11174) );
  OR2X2 OR2X2_2291 ( .A(u2__abc_44228_n11178), .B(u2__abc_44228_n11164), .Y(u2__abc_44228_n11179_1) );
  OR2X2 OR2X2_2292 ( .A(u2__abc_44228_n11186_1), .B(u2__abc_44228_n11183), .Y(u2__abc_44228_n11187_1) );
  OR2X2 OR2X2_2293 ( .A(u2__abc_44228_n11189), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n11190) );
  OR2X2 OR2X2_2294 ( .A(u2__abc_44228_n11188), .B(u2__abc_44228_n11190), .Y(u2__abc_44228_n11191) );
  OR2X2 OR2X2_2295 ( .A(u2__abc_44228_n11195), .B(u2__abc_44228_n11181), .Y(u2__abc_44228_n11196) );
  OR2X2 OR2X2_2296 ( .A(u2__abc_44228_n11199), .B(u2__abc_44228_n4623), .Y(u2__abc_44228_n11200_1) );
  OR2X2 OR2X2_2297 ( .A(u2__abc_44228_n11201_1), .B(u2__abc_44228_n4611), .Y(u2__abc_44228_n11202) );
  OR2X2 OR2X2_2298 ( .A(u2__abc_44228_n11207_1), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n11208_1) );
  OR2X2 OR2X2_2299 ( .A(u2__abc_44228_n11206), .B(u2__abc_44228_n11208_1), .Y(u2__abc_44228_n11209) );
  OR2X2 OR2X2_23 ( .A(aNan_bF_buf9), .B(sqrto_87_), .Y(_abc_64468_n863) );
  OR2X2 OR2X2_230 ( .A(a_112_bF_buf5), .B(\a[2] ), .Y(_abc_64468_n1176) );
  OR2X2 OR2X2_2300 ( .A(u2__abc_44228_n11213), .B(u2__abc_44228_n11198), .Y(u2__abc_44228_n11214_1) );
  OR2X2 OR2X2_2301 ( .A(u2__abc_44228_n11203), .B(u2__abc_44228_n4607), .Y(u2__abc_44228_n11218) );
  OR2X2 OR2X2_2302 ( .A(u2__abc_44228_n11219), .B(u2__abc_44228_n11217), .Y(u2__abc_44228_n11220) );
  OR2X2 OR2X2_2303 ( .A(u2__abc_44228_n11218), .B(u2__abc_44228_n4605), .Y(u2__abc_44228_n11221_1) );
  OR2X2 OR2X2_2304 ( .A(u2__abc_44228_n11224), .B(u2__abc_44228_n2983_bF_buf18), .Y(u2__abc_44228_n11225) );
  OR2X2 OR2X2_2305 ( .A(u2__abc_44228_n11223), .B(u2__abc_44228_n11225), .Y(u2__abc_44228_n11226) );
  OR2X2 OR2X2_2306 ( .A(u2__abc_44228_n11230), .B(u2__abc_44228_n11216), .Y(u2__abc_44228_n11231) );
  OR2X2 OR2X2_2307 ( .A(u2__abc_44228_n11234), .B(u2__abc_44228_n5467), .Y(u2__abc_44228_n11235_1) );
  OR2X2 OR2X2_2308 ( .A(u2__abc_44228_n11235_1), .B(u2__abc_44228_n4588), .Y(u2__abc_44228_n11236_1) );
  OR2X2 OR2X2_2309 ( .A(u2__abc_44228_n7548_1_bF_buf15), .B(u2__abc_44228_n11239), .Y(u2__abc_44228_n11240) );
  OR2X2 OR2X2_231 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[3] ), .Y(_abc_64468_n1177) );
  OR2X2 OR2X2_2310 ( .A(u2__abc_44228_n7547_bF_buf14), .B(u2_remHi_214_), .Y(u2__abc_44228_n11241) );
  OR2X2 OR2X2_2311 ( .A(u2__abc_44228_n11242_1), .B(u2__abc_44228_n2983_bF_buf16), .Y(u2__abc_44228_n11243_1) );
  OR2X2 OR2X2_2312 ( .A(u2__abc_44228_n11247), .B(u2__abc_44228_n11233), .Y(u2__abc_44228_n11248) );
  OR2X2 OR2X2_2313 ( .A(u2__abc_44228_n11255), .B(u2__abc_44228_n11252), .Y(u2__abc_44228_n11256_1) );
  OR2X2 OR2X2_2314 ( .A(u2__abc_44228_n11258), .B(u2__abc_44228_n2983_bF_buf14), .Y(u2__abc_44228_n11259) );
  OR2X2 OR2X2_2315 ( .A(u2__abc_44228_n11257_1), .B(u2__abc_44228_n11259), .Y(u2__abc_44228_n11260) );
  OR2X2 OR2X2_2316 ( .A(u2__abc_44228_n11264_1), .B(u2__abc_44228_n11250_1), .Y(u2__abc_44228_n11265) );
  OR2X2 OR2X2_2317 ( .A(u2__abc_44228_n11268), .B(u2__abc_44228_n4593), .Y(u2__abc_44228_n11269) );
  OR2X2 OR2X2_2318 ( .A(u2__abc_44228_n11270_1), .B(u2__abc_44228_n4581_1), .Y(u2__abc_44228_n11271_1) );
  OR2X2 OR2X2_2319 ( .A(u2__abc_44228_n11276), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n11277_1) );
  OR2X2 OR2X2_232 ( .A(a_112_bF_buf4), .B(\a[3] ), .Y(_abc_64468_n1179) );
  OR2X2 OR2X2_2320 ( .A(u2__abc_44228_n11275), .B(u2__abc_44228_n11277_1), .Y(u2__abc_44228_n11278_1) );
  OR2X2 OR2X2_2321 ( .A(u2__abc_44228_n11282), .B(u2__abc_44228_n11267), .Y(u2__abc_44228_n11283) );
  OR2X2 OR2X2_2322 ( .A(u2__abc_44228_n11272), .B(u2__abc_44228_n4577), .Y(u2__abc_44228_n11287) );
  OR2X2 OR2X2_2323 ( .A(u2__abc_44228_n11288), .B(u2__abc_44228_n11286), .Y(u2__abc_44228_n11289) );
  OR2X2 OR2X2_2324 ( .A(u2__abc_44228_n11287), .B(u2__abc_44228_n4575), .Y(u2__abc_44228_n11290) );
  OR2X2 OR2X2_2325 ( .A(u2__abc_44228_n11293), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n11294) );
  OR2X2 OR2X2_2326 ( .A(u2__abc_44228_n11292_1), .B(u2__abc_44228_n11294), .Y(u2__abc_44228_n11295) );
  OR2X2 OR2X2_2327 ( .A(u2__abc_44228_n11299_1), .B(u2__abc_44228_n11285_1), .Y(u2__abc_44228_n11300) );
  OR2X2 OR2X2_2328 ( .A(u2__abc_44228_n11303), .B(u2__abc_44228_n5476), .Y(u2__abc_44228_n11304) );
  OR2X2 OR2X2_2329 ( .A(u2__abc_44228_n11304), .B(u2__abc_44228_n4559), .Y(u2__abc_44228_n11307) );
  OR2X2 OR2X2_233 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[4] ), .Y(_abc_64468_n1180) );
  OR2X2 OR2X2_2330 ( .A(u2__abc_44228_n11310), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n11311) );
  OR2X2 OR2X2_2331 ( .A(u2__abc_44228_n11309), .B(u2__abc_44228_n11311), .Y(u2__abc_44228_n11312_1) );
  OR2X2 OR2X2_2332 ( .A(u2__abc_44228_n11316), .B(u2__abc_44228_n11302), .Y(u2__abc_44228_n11317) );
  OR2X2 OR2X2_2333 ( .A(u2__abc_44228_n11321), .B(u2__abc_44228_n4566), .Y(u2__abc_44228_n11322) );
  OR2X2 OR2X2_2334 ( .A(u2__abc_44228_n11320_1), .B(u2__abc_44228_n11323), .Y(u2__abc_44228_n11324) );
  OR2X2 OR2X2_2335 ( .A(u2__abc_44228_n11327_1), .B(u2__abc_44228_n2983_bF_buf8), .Y(u2__abc_44228_n11328) );
  OR2X2 OR2X2_2336 ( .A(u2__abc_44228_n11326_1), .B(u2__abc_44228_n11328), .Y(u2__abc_44228_n11329) );
  OR2X2 OR2X2_2337 ( .A(u2__abc_44228_n11333_1), .B(u2__abc_44228_n11319_1), .Y(u2__abc_44228_n11334_1) );
  OR2X2 OR2X2_2338 ( .A(u2__abc_44228_n11337), .B(u2__abc_44228_n4564), .Y(u2__abc_44228_n11338) );
  OR2X2 OR2X2_2339 ( .A(u2__abc_44228_n11339), .B(u2__abc_44228_n4552), .Y(u2__abc_44228_n11340_1) );
  OR2X2 OR2X2_234 ( .A(a_112_bF_buf3), .B(\a[4] ), .Y(_abc_64468_n1182) );
  OR2X2 OR2X2_2340 ( .A(u2__abc_44228_n11345), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n11346) );
  OR2X2 OR2X2_2341 ( .A(u2__abc_44228_n11344), .B(u2__abc_44228_n11346), .Y(u2__abc_44228_n11347_1) );
  OR2X2 OR2X2_2342 ( .A(u2__abc_44228_n11351), .B(u2__abc_44228_n11336), .Y(u2__abc_44228_n11352) );
  OR2X2 OR2X2_2343 ( .A(u2__abc_44228_n11341_1), .B(u2__abc_44228_n4548), .Y(u2__abc_44228_n11356) );
  OR2X2 OR2X2_2344 ( .A(u2__abc_44228_n11357), .B(u2__abc_44228_n11355_1), .Y(u2__abc_44228_n11358) );
  OR2X2 OR2X2_2345 ( .A(u2__abc_44228_n11356), .B(u2__abc_44228_n4546), .Y(u2__abc_44228_n11359) );
  OR2X2 OR2X2_2346 ( .A(u2__abc_44228_n11362_1), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n11363) );
  OR2X2 OR2X2_2347 ( .A(u2__abc_44228_n11361_1), .B(u2__abc_44228_n11363), .Y(u2__abc_44228_n11364) );
  OR2X2 OR2X2_2348 ( .A(u2__abc_44228_n11368_1), .B(u2__abc_44228_n11354_1), .Y(u2__abc_44228_n11369_1) );
  OR2X2 OR2X2_2349 ( .A(u2__abc_44228_n11372), .B(u2__abc_44228_n5488), .Y(u2__abc_44228_n11373) );
  OR2X2 OR2X2_235 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[5] ), .Y(_abc_64468_n1183) );
  OR2X2 OR2X2_2350 ( .A(u2__abc_44228_n11373), .B(u2__abc_44228_n4527), .Y(u2__abc_44228_n11374) );
  OR2X2 OR2X2_2351 ( .A(u2__abc_44228_n7548_1_bF_buf7), .B(u2__abc_44228_n11377), .Y(u2__abc_44228_n11378) );
  OR2X2 OR2X2_2352 ( .A(u2__abc_44228_n7547_bF_buf6), .B(u2_remHi_222_), .Y(u2__abc_44228_n11379) );
  OR2X2 OR2X2_2353 ( .A(u2__abc_44228_n11380), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n11381) );
  OR2X2 OR2X2_2354 ( .A(u2__abc_44228_n11385), .B(u2__abc_44228_n11371), .Y(u2__abc_44228_n11386) );
  OR2X2 OR2X2_2355 ( .A(u2__abc_44228_n11390_1), .B(u2__abc_44228_n11389_1), .Y(u2__abc_44228_n11391) );
  OR2X2 OR2X2_2356 ( .A(u2__abc_44228_n11392), .B(u2__abc_44228_n4534), .Y(u2__abc_44228_n11393) );
  OR2X2 OR2X2_2357 ( .A(u2__abc_44228_n11396_1), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n11397_1) );
  OR2X2 OR2X2_2358 ( .A(u2__abc_44228_n11397_1), .B(u2__abc_44228_n11395), .Y(u2__abc_44228_n11398) );
  OR2X2 OR2X2_2359 ( .A(u2__abc_44228_n11402), .B(u2__abc_44228_n11388), .Y(u2__abc_44228_n11403_1) );
  OR2X2 OR2X2_236 ( .A(a_112_bF_buf2), .B(\a[5] ), .Y(_abc_64468_n1185) );
  OR2X2 OR2X2_2360 ( .A(u2__abc_44228_n11406), .B(u2__abc_44228_n5493_1), .Y(u2__abc_44228_n11407) );
  OR2X2 OR2X2_2361 ( .A(u2__abc_44228_n11407), .B(u2__abc_44228_n4520), .Y(u2__abc_44228_n11408) );
  OR2X2 OR2X2_2362 ( .A(u2__abc_44228_n7548_1_bF_buf5), .B(u2__abc_44228_n11411_1), .Y(u2__abc_44228_n11412) );
  OR2X2 OR2X2_2363 ( .A(u2__abc_44228_n7547_bF_buf4), .B(u2_remHi_224_), .Y(u2__abc_44228_n11413) );
  OR2X2 OR2X2_2364 ( .A(u2__abc_44228_n11414), .B(u2__abc_44228_n2983_bF_buf0), .Y(u2__abc_44228_n11415) );
  OR2X2 OR2X2_2365 ( .A(u2__abc_44228_n11419), .B(u2__abc_44228_n11405), .Y(u2__abc_44228_n11420) );
  OR2X2 OR2X2_2366 ( .A(u2__abc_44228_n11409), .B(u2__abc_44228_n4516), .Y(u2__abc_44228_n11424_1) );
  OR2X2 OR2X2_2367 ( .A(u2__abc_44228_n11425_1), .B(u2__abc_44228_n11423), .Y(u2__abc_44228_n11426) );
  OR2X2 OR2X2_2368 ( .A(u2__abc_44228_n11424_1), .B(u2__abc_44228_n4514), .Y(u2__abc_44228_n11427) );
  OR2X2 OR2X2_2369 ( .A(u2__abc_44228_n11430), .B(u2__abc_44228_n2983_bF_buf140), .Y(u2__abc_44228_n11431_1) );
  OR2X2 OR2X2_237 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[6] ), .Y(_abc_64468_n1186) );
  OR2X2 OR2X2_2370 ( .A(u2__abc_44228_n11429), .B(u2__abc_44228_n11431_1), .Y(u2__abc_44228_n11432_1) );
  OR2X2 OR2X2_2371 ( .A(u2__abc_44228_n11436), .B(u2__abc_44228_n11422), .Y(u2__abc_44228_n11437) );
  OR2X2 OR2X2_2372 ( .A(u2__abc_44228_n11440), .B(u2__abc_44228_n5497), .Y(u2__abc_44228_n11441) );
  OR2X2 OR2X2_2373 ( .A(u2__abc_44228_n11441), .B(u2__abc_44228_n4498_1), .Y(u2__abc_44228_n11444) );
  OR2X2 OR2X2_2374 ( .A(u2__abc_44228_n7548_1_bF_buf3), .B(u2__abc_44228_n11445_1), .Y(u2__abc_44228_n11446_1) );
  OR2X2 OR2X2_2375 ( .A(u2__abc_44228_n7547_bF_buf2), .B(u2_remHi_226_), .Y(u2__abc_44228_n11447) );
  OR2X2 OR2X2_2376 ( .A(u2__abc_44228_n11448), .B(u2__abc_44228_n2983_bF_buf138), .Y(u2__abc_44228_n11449) );
  OR2X2 OR2X2_2377 ( .A(u2__abc_44228_n11453_1), .B(u2__abc_44228_n11439_1), .Y(u2__abc_44228_n11454) );
  OR2X2 OR2X2_2378 ( .A(u2__abc_44228_n11458), .B(u2__abc_44228_n4505), .Y(u2__abc_44228_n11459_1) );
  OR2X2 OR2X2_2379 ( .A(u2__abc_44228_n11457), .B(u2__abc_44228_n11460_1), .Y(u2__abc_44228_n11461) );
  OR2X2 OR2X2_238 ( .A(a_112_bF_buf1), .B(\a[6] ), .Y(_abc_64468_n1188) );
  OR2X2 OR2X2_2380 ( .A(u2__abc_44228_n11464), .B(u2__abc_44228_n2983_bF_buf136), .Y(u2__abc_44228_n11465) );
  OR2X2 OR2X2_2381 ( .A(u2__abc_44228_n11463), .B(u2__abc_44228_n11465), .Y(u2__abc_44228_n11466_1) );
  OR2X2 OR2X2_2382 ( .A(u2__abc_44228_n11470), .B(u2__abc_44228_n11456), .Y(u2__abc_44228_n11471) );
  OR2X2 OR2X2_2383 ( .A(u2__abc_44228_n11474_1), .B(u2__abc_44228_n4503), .Y(u2__abc_44228_n11475) );
  OR2X2 OR2X2_2384 ( .A(u2__abc_44228_n11476), .B(u2__abc_44228_n4491), .Y(u2__abc_44228_n11477) );
  OR2X2 OR2X2_2385 ( .A(u2__abc_44228_n11482), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n11483) );
  OR2X2 OR2X2_2386 ( .A(u2__abc_44228_n11481_1), .B(u2__abc_44228_n11483), .Y(u2__abc_44228_n11484) );
  OR2X2 OR2X2_2387 ( .A(u2__abc_44228_n11488_1), .B(u2__abc_44228_n11473_1), .Y(u2__abc_44228_n11489) );
  OR2X2 OR2X2_2388 ( .A(u2__abc_44228_n11478), .B(u2__abc_44228_n4487), .Y(u2__abc_44228_n11493) );
  OR2X2 OR2X2_2389 ( .A(u2__abc_44228_n11494_1), .B(u2__abc_44228_n11492), .Y(u2__abc_44228_n11495_1) );
  OR2X2 OR2X2_239 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[7] ), .Y(_abc_64468_n1189) );
  OR2X2 OR2X2_2390 ( .A(u2__abc_44228_n11493), .B(u2__abc_44228_n4485), .Y(u2__abc_44228_n11496) );
  OR2X2 OR2X2_2391 ( .A(u2__abc_44228_n11499), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n11500) );
  OR2X2 OR2X2_2392 ( .A(u2__abc_44228_n11498), .B(u2__abc_44228_n11500), .Y(u2__abc_44228_n11501_1) );
  OR2X2 OR2X2_2393 ( .A(u2__abc_44228_n11505), .B(u2__abc_44228_n11491), .Y(u2__abc_44228_n11506) );
  OR2X2 OR2X2_2394 ( .A(u2__abc_44228_n11509_1), .B(u2__abc_44228_n5507), .Y(u2__abc_44228_n11510) );
  OR2X2 OR2X2_2395 ( .A(u2__abc_44228_n11510), .B(u2__abc_44228_n4461_1), .Y(u2__abc_44228_n11511) );
  OR2X2 OR2X2_2396 ( .A(u2__abc_44228_n7548_1_bF_buf57), .B(u2__abc_44228_n11514), .Y(u2__abc_44228_n11515_1) );
  OR2X2 OR2X2_2397 ( .A(u2__abc_44228_n7547_bF_buf56), .B(u2_remHi_230_), .Y(u2__abc_44228_n11516_1) );
  OR2X2 OR2X2_2398 ( .A(u2__abc_44228_n11517), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n11518) );
  OR2X2 OR2X2_2399 ( .A(u2__abc_44228_n11522_1), .B(u2__abc_44228_n11508_1), .Y(u2__abc_44228_n11523_1) );
  OR2X2 OR2X2_24 ( .A(_abc_64468_n753_bF_buf10), .B(\a[11] ), .Y(_abc_64468_n864) );
  OR2X2 OR2X2_240 ( .A(a_112_bF_buf0), .B(\a[7] ), .Y(_abc_64468_n1191) );
  OR2X2 OR2X2_2400 ( .A(u2__abc_44228_n11527), .B(u2__abc_44228_n11526), .Y(u2__abc_44228_n11528) );
  OR2X2 OR2X2_2401 ( .A(u2__abc_44228_n11529_1), .B(u2__abc_44228_n4455), .Y(u2__abc_44228_n11530_1) );
  OR2X2 OR2X2_2402 ( .A(u2__abc_44228_n11533), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n11534) );
  OR2X2 OR2X2_2403 ( .A(u2__abc_44228_n11532), .B(u2__abc_44228_n11534), .Y(u2__abc_44228_n11535) );
  OR2X2 OR2X2_2404 ( .A(u2__abc_44228_n11539), .B(u2__abc_44228_n11525), .Y(u2__abc_44228_n11540) );
  OR2X2 OR2X2_2405 ( .A(u2__abc_44228_n11543_1), .B(u2__abc_44228_n5512_1), .Y(u2__abc_44228_n11544_1) );
  OR2X2 OR2X2_2406 ( .A(u2__abc_44228_n11544_1), .B(u2__abc_44228_n4475), .Y(u2__abc_44228_n11545) );
  OR2X2 OR2X2_2407 ( .A(u2__abc_44228_n11550_1), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n11551_1) );
  OR2X2 OR2X2_2408 ( .A(u2__abc_44228_n11549), .B(u2__abc_44228_n11551_1), .Y(u2__abc_44228_n11552) );
  OR2X2 OR2X2_2409 ( .A(u2__abc_44228_n11556), .B(u2__abc_44228_n11542), .Y(u2__abc_44228_n11557_1) );
  OR2X2 OR2X2_241 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[8] ), .Y(_abc_64468_n1192) );
  OR2X2 OR2X2_2410 ( .A(u2__abc_44228_n11561), .B(u2__abc_44228_n11560), .Y(u2__abc_44228_n11562) );
  OR2X2 OR2X2_2411 ( .A(u2__abc_44228_n11563), .B(u2__abc_44228_n4469), .Y(u2__abc_44228_n11564_1) );
  OR2X2 OR2X2_2412 ( .A(u2__abc_44228_n11567), .B(u2__abc_44228_n2983_bF_buf126), .Y(u2__abc_44228_n11568) );
  OR2X2 OR2X2_2413 ( .A(u2__abc_44228_n11566), .B(u2__abc_44228_n11568), .Y(u2__abc_44228_n11569) );
  OR2X2 OR2X2_2414 ( .A(u2__abc_44228_n11573), .B(u2__abc_44228_n11559), .Y(u2__abc_44228_n11574) );
  OR2X2 OR2X2_2415 ( .A(u2__abc_44228_n11577), .B(u2__abc_44228_n4467), .Y(u2__abc_44228_n11578_1) );
  OR2X2 OR2X2_2416 ( .A(u2__abc_44228_n11579_1), .B(u2__abc_44228_n4439), .Y(u2__abc_44228_n11582) );
  OR2X2 OR2X2_2417 ( .A(u2__abc_44228_n11585_1), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n11586_1) );
  OR2X2 OR2X2_2418 ( .A(u2__abc_44228_n11584), .B(u2__abc_44228_n11586_1), .Y(u2__abc_44228_n11587) );
  OR2X2 OR2X2_2419 ( .A(u2__abc_44228_n11591), .B(u2__abc_44228_n11576), .Y(u2__abc_44228_n11592_1) );
  OR2X2 OR2X2_242 ( .A(a_112_bF_buf9), .B(\a[8] ), .Y(_abc_64468_n1194) );
  OR2X2 OR2X2_2420 ( .A(u2__abc_44228_n11596), .B(u2__abc_44228_n4446), .Y(u2__abc_44228_n11597) );
  OR2X2 OR2X2_2421 ( .A(u2__abc_44228_n11595), .B(u2__abc_44228_n11598), .Y(u2__abc_44228_n11599_1) );
  OR2X2 OR2X2_2422 ( .A(u2__abc_44228_n11602), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n11603) );
  OR2X2 OR2X2_2423 ( .A(u2__abc_44228_n11601), .B(u2__abc_44228_n11603), .Y(u2__abc_44228_n11604) );
  OR2X2 OR2X2_2424 ( .A(u2__abc_44228_n11608), .B(u2__abc_44228_n11594), .Y(u2__abc_44228_n11609) );
  OR2X2 OR2X2_2425 ( .A(u2__abc_44228_n11612), .B(u2__abc_44228_n4444), .Y(u2__abc_44228_n11613_1) );
  OR2X2 OR2X2_2426 ( .A(u2__abc_44228_n11614_1), .B(u2__abc_44228_n4432_1), .Y(u2__abc_44228_n11617) );
  OR2X2 OR2X2_2427 ( .A(u2__abc_44228_n11620_1), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n11621_1) );
  OR2X2 OR2X2_2428 ( .A(u2__abc_44228_n11619), .B(u2__abc_44228_n11621_1), .Y(u2__abc_44228_n11622) );
  OR2X2 OR2X2_2429 ( .A(u2__abc_44228_n11626), .B(u2__abc_44228_n11611), .Y(u2__abc_44228_n11627_1) );
  OR2X2 OR2X2_243 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[9] ), .Y(_abc_64468_n1195) );
  OR2X2 OR2X2_2430 ( .A(u2__abc_44228_n11615), .B(u2__abc_44228_n4428), .Y(u2__abc_44228_n11631) );
  OR2X2 OR2X2_2431 ( .A(u2__abc_44228_n11632), .B(u2__abc_44228_n11630), .Y(u2__abc_44228_n11633) );
  OR2X2 OR2X2_2432 ( .A(u2__abc_44228_n11631), .B(u2__abc_44228_n4426), .Y(u2__abc_44228_n11634_1) );
  OR2X2 OR2X2_2433 ( .A(u2__abc_44228_n11637), .B(u2__abc_44228_n2983_bF_buf119), .Y(u2__abc_44228_n11638) );
  OR2X2 OR2X2_2434 ( .A(u2__abc_44228_n11636), .B(u2__abc_44228_n11638), .Y(u2__abc_44228_n11639) );
  OR2X2 OR2X2_2435 ( .A(u2__abc_44228_n11643), .B(u2__abc_44228_n11629), .Y(u2__abc_44228_n11644) );
  OR2X2 OR2X2_2436 ( .A(u2__abc_44228_n11647), .B(u2__abc_44228_n5529), .Y(u2__abc_44228_n11648_1) );
  OR2X2 OR2X2_2437 ( .A(u2__abc_44228_n11648_1), .B(u2__abc_44228_n4408), .Y(u2__abc_44228_n11651) );
  OR2X2 OR2X2_2438 ( .A(u2__abc_44228_n7548_1_bF_buf49), .B(u2__abc_44228_n11652), .Y(u2__abc_44228_n11653) );
  OR2X2 OR2X2_2439 ( .A(u2__abc_44228_n7547_bF_buf48), .B(u2_remHi_238_), .Y(u2__abc_44228_n11654) );
  OR2X2 OR2X2_244 ( .A(a_112_bF_buf8), .B(\a[9] ), .Y(_abc_64468_n1197) );
  OR2X2 OR2X2_2440 ( .A(u2__abc_44228_n11655_1), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n11656_1) );
  OR2X2 OR2X2_2441 ( .A(u2__abc_44228_n11660), .B(u2__abc_44228_n11646), .Y(u2__abc_44228_n11661) );
  OR2X2 OR2X2_2442 ( .A(u2__abc_44228_n11665), .B(u2__abc_44228_n11664), .Y(u2__abc_44228_n11666) );
  OR2X2 OR2X2_2443 ( .A(u2__abc_44228_n11667), .B(u2__abc_44228_n4415), .Y(u2__abc_44228_n11668) );
  OR2X2 OR2X2_2444 ( .A(u2__abc_44228_n11671), .B(u2__abc_44228_n2983_bF_buf115), .Y(u2__abc_44228_n11672) );
  OR2X2 OR2X2_2445 ( .A(u2__abc_44228_n11670), .B(u2__abc_44228_n11672), .Y(u2__abc_44228_n11673) );
  OR2X2 OR2X2_2446 ( .A(u2__abc_44228_n11677), .B(u2__abc_44228_n11663_1), .Y(u2__abc_44228_n11678) );
  OR2X2 OR2X2_2447 ( .A(u2__abc_44228_n11681), .B(u2__abc_44228_n4413), .Y(u2__abc_44228_n11682) );
  OR2X2 OR2X2_2448 ( .A(u2__abc_44228_n11683), .B(u2__abc_44228_n4401), .Y(u2__abc_44228_n11684_1) );
  OR2X2 OR2X2_2449 ( .A(u2__abc_44228_n11689), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n11690_1) );
  OR2X2 OR2X2_245 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[10] ), .Y(_abc_64468_n1198) );
  OR2X2 OR2X2_2450 ( .A(u2__abc_44228_n11688), .B(u2__abc_44228_n11690_1), .Y(u2__abc_44228_n11691) );
  OR2X2 OR2X2_2451 ( .A(u2__abc_44228_n11695), .B(u2__abc_44228_n11680), .Y(u2__abc_44228_n11696) );
  OR2X2 OR2X2_2452 ( .A(u2__abc_44228_n11685), .B(u2__abc_44228_n4397), .Y(u2__abc_44228_n11700) );
  OR2X2 OR2X2_2453 ( .A(u2__abc_44228_n11701), .B(u2__abc_44228_n11699), .Y(u2__abc_44228_n11702) );
  OR2X2 OR2X2_2454 ( .A(u2__abc_44228_n11700), .B(u2__abc_44228_n4395), .Y(u2__abc_44228_n11703) );
  OR2X2 OR2X2_2455 ( .A(u2__abc_44228_n11706), .B(u2__abc_44228_n2983_bF_buf112), .Y(u2__abc_44228_n11707) );
  OR2X2 OR2X2_2456 ( .A(u2__abc_44228_n11705), .B(u2__abc_44228_n11707), .Y(u2__abc_44228_n11708) );
  OR2X2 OR2X2_2457 ( .A(u2__abc_44228_n11712), .B(u2__abc_44228_n11698), .Y(u2__abc_44228_n11713) );
  OR2X2 OR2X2_2458 ( .A(u2__abc_44228_n11716), .B(u2__abc_44228_n5556), .Y(u2__abc_44228_n11717) );
  OR2X2 OR2X2_2459 ( .A(u2__abc_44228_n11717), .B(u2__abc_44228_n4379), .Y(u2__abc_44228_n11720) );
  OR2X2 OR2X2_246 ( .A(a_112_bF_buf7), .B(\a[10] ), .Y(_abc_64468_n1200) );
  OR2X2 OR2X2_2460 ( .A(u2__abc_44228_n11723), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n11724) );
  OR2X2 OR2X2_2461 ( .A(u2__abc_44228_n11722), .B(u2__abc_44228_n11724), .Y(u2__abc_44228_n11725) );
  OR2X2 OR2X2_2462 ( .A(u2__abc_44228_n11729), .B(u2__abc_44228_n11715), .Y(u2__abc_44228_n11730) );
  OR2X2 OR2X2_2463 ( .A(u2__abc_44228_n11734_1), .B(u2__abc_44228_n4386_1), .Y(u2__abc_44228_n11735) );
  OR2X2 OR2X2_2464 ( .A(u2__abc_44228_n11733), .B(u2__abc_44228_n11736), .Y(u2__abc_44228_n11737) );
  OR2X2 OR2X2_2465 ( .A(u2__abc_44228_n11740), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n11741_1) );
  OR2X2 OR2X2_2466 ( .A(u2__abc_44228_n11739), .B(u2__abc_44228_n11741_1), .Y(u2__abc_44228_n11742) );
  OR2X2 OR2X2_2467 ( .A(u2__abc_44228_n11746), .B(u2__abc_44228_n11732), .Y(u2__abc_44228_n11747) );
  OR2X2 OR2X2_2468 ( .A(u2__abc_44228_n11750_1), .B(u2__abc_44228_n4384), .Y(u2__abc_44228_n11751) );
  OR2X2 OR2X2_2469 ( .A(u2__abc_44228_n11752), .B(u2__abc_44228_n4372), .Y(u2__abc_44228_n11753) );
  OR2X2 OR2X2_247 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[11] ), .Y(_abc_64468_n1201) );
  OR2X2 OR2X2_2470 ( .A(u2__abc_44228_n11758), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n11759) );
  OR2X2 OR2X2_2471 ( .A(u2__abc_44228_n11757_1), .B(u2__abc_44228_n11759), .Y(u2__abc_44228_n11760) );
  OR2X2 OR2X2_2472 ( .A(u2__abc_44228_n11764), .B(u2__abc_44228_n11749), .Y(u2__abc_44228_n11765_1) );
  OR2X2 OR2X2_2473 ( .A(u2__abc_44228_n11754), .B(u2__abc_44228_n4368_1), .Y(u2__abc_44228_n11769) );
  OR2X2 OR2X2_2474 ( .A(u2__abc_44228_n11770), .B(u2__abc_44228_n11768), .Y(u2__abc_44228_n11771) );
  OR2X2 OR2X2_2475 ( .A(u2__abc_44228_n11769), .B(u2__abc_44228_n4366), .Y(u2__abc_44228_n11772_1) );
  OR2X2 OR2X2_2476 ( .A(u2__abc_44228_n11775), .B(u2__abc_44228_n2983_bF_buf106), .Y(u2__abc_44228_n11776) );
  OR2X2 OR2X2_2477 ( .A(u2__abc_44228_n11774), .B(u2__abc_44228_n11776), .Y(u2__abc_44228_n11777) );
  OR2X2 OR2X2_2478 ( .A(u2__abc_44228_n11781_1), .B(u2__abc_44228_n11767), .Y(u2__abc_44228_n11782) );
  OR2X2 OR2X2_2479 ( .A(u2__abc_44228_n11785), .B(u2__abc_44228_n5566), .Y(u2__abc_44228_n11786) );
  OR2X2 OR2X2_248 ( .A(a_112_bF_buf6), .B(\a[11] ), .Y(_abc_64468_n1203) );
  OR2X2 OR2X2_2480 ( .A(u2__abc_44228_n11786), .B(u2__abc_44228_n4349_1), .Y(u2__abc_44228_n11787) );
  OR2X2 OR2X2_2481 ( .A(u2__abc_44228_n11792), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n11793) );
  OR2X2 OR2X2_2482 ( .A(u2__abc_44228_n11791), .B(u2__abc_44228_n11793), .Y(u2__abc_44228_n11794) );
  OR2X2 OR2X2_2483 ( .A(u2__abc_44228_n11798), .B(u2__abc_44228_n11784), .Y(u2__abc_44228_n11799) );
  OR2X2 OR2X2_2484 ( .A(u2__abc_44228_n11806), .B(u2__abc_44228_n11803_1), .Y(u2__abc_44228_n11807) );
  OR2X2 OR2X2_2485 ( .A(u2__abc_44228_n11809), .B(u2__abc_44228_n2983_bF_buf103), .Y(u2__abc_44228_n11810) );
  OR2X2 OR2X2_2486 ( .A(u2__abc_44228_n11808), .B(u2__abc_44228_n11810), .Y(u2__abc_44228_n11811) );
  OR2X2 OR2X2_2487 ( .A(u2__abc_44228_n11815), .B(u2__abc_44228_n11801), .Y(u2__abc_44228_n11816) );
  OR2X2 OR2X2_2488 ( .A(u2__abc_44228_n11819), .B(u2__abc_44228_n4354), .Y(u2__abc_44228_n11820_1) );
  OR2X2 OR2X2_2489 ( .A(u2__abc_44228_n11821), .B(u2__abc_44228_n4342), .Y(u2__abc_44228_n11822) );
  OR2X2 OR2X2_249 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[12] ), .Y(_abc_64468_n1204) );
  OR2X2 OR2X2_2490 ( .A(u2__abc_44228_n11827), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n11828_1) );
  OR2X2 OR2X2_2491 ( .A(u2__abc_44228_n11826), .B(u2__abc_44228_n11828_1), .Y(u2__abc_44228_n11829) );
  OR2X2 OR2X2_2492 ( .A(u2__abc_44228_n11833), .B(u2__abc_44228_n11818), .Y(u2__abc_44228_n11834) );
  OR2X2 OR2X2_2493 ( .A(u2__abc_44228_n11823), .B(u2__abc_44228_n4338_1), .Y(u2__abc_44228_n11838) );
  OR2X2 OR2X2_2494 ( .A(u2__abc_44228_n11839), .B(u2__abc_44228_n11837), .Y(u2__abc_44228_n11840) );
  OR2X2 OR2X2_2495 ( .A(u2__abc_44228_n11838), .B(u2__abc_44228_n4336), .Y(u2__abc_44228_n11841) );
  OR2X2 OR2X2_2496 ( .A(u2__abc_44228_n11844_1), .B(u2__abc_44228_n2983_bF_buf100), .Y(u2__abc_44228_n11845) );
  OR2X2 OR2X2_2497 ( .A(u2__abc_44228_n11843), .B(u2__abc_44228_n11845), .Y(u2__abc_44228_n11846) );
  OR2X2 OR2X2_2498 ( .A(u2__abc_44228_n11850), .B(u2__abc_44228_n11836), .Y(u2__abc_44228_n11851_1) );
  OR2X2 OR2X2_2499 ( .A(u2__abc_44228_n11854), .B(u2__abc_44228_n5538), .Y(u2__abc_44228_n11855) );
  OR2X2 OR2X2_25 ( .A(aNan_bF_buf8), .B(sqrto_88_), .Y(_abc_64468_n866) );
  OR2X2 OR2X2_250 ( .A(a_112_bF_buf5), .B(\a[12] ), .Y(_abc_64468_n1206) );
  OR2X2 OR2X2_2500 ( .A(u2__abc_44228_n11855), .B(u2__abc_44228_n4320_1), .Y(u2__abc_44228_n11858) );
  OR2X2 OR2X2_2501 ( .A(u2__abc_44228_n11861), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n11862) );
  OR2X2 OR2X2_2502 ( .A(u2__abc_44228_n11860), .B(u2__abc_44228_n11862), .Y(u2__abc_44228_n11863) );
  OR2X2 OR2X2_2503 ( .A(u2__abc_44228_n11867), .B(u2__abc_44228_n11853), .Y(u2__abc_44228_n11868) );
  OR2X2 OR2X2_2504 ( .A(u2__abc_44228_n11875), .B(u2__abc_44228_n11872), .Y(u2__abc_44228_n11876_1) );
  OR2X2 OR2X2_2505 ( .A(u2__abc_44228_n11878), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n11879) );
  OR2X2 OR2X2_2506 ( .A(u2__abc_44228_n11877), .B(u2__abc_44228_n11879), .Y(u2__abc_44228_n11880) );
  OR2X2 OR2X2_2507 ( .A(u2__abc_44228_n11884), .B(u2__abc_44228_n11870), .Y(u2__abc_44228_n11885) );
  OR2X2 OR2X2_2508 ( .A(u2__abc_44228_n11888), .B(u2__abc_44228_n4325), .Y(u2__abc_44228_n11889) );
  OR2X2 OR2X2_2509 ( .A(u2__abc_44228_n11890), .B(u2__abc_44228_n4313), .Y(u2__abc_44228_n11891_1) );
  OR2X2 OR2X2_251 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[13] ), .Y(_abc_64468_n1207) );
  OR2X2 OR2X2_2510 ( .A(u2__abc_44228_n11896), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n11897) );
  OR2X2 OR2X2_2511 ( .A(u2__abc_44228_n11895), .B(u2__abc_44228_n11897), .Y(u2__abc_44228_n11898_1) );
  OR2X2 OR2X2_2512 ( .A(u2__abc_44228_n11902), .B(u2__abc_44228_n11887), .Y(u2__abc_44228_n11903) );
  OR2X2 OR2X2_2513 ( .A(u2__abc_44228_n11892), .B(u2__abc_44228_n4309), .Y(u2__abc_44228_n11907_1) );
  OR2X2 OR2X2_2514 ( .A(u2__abc_44228_n11908), .B(u2__abc_44228_n11906), .Y(u2__abc_44228_n11909) );
  OR2X2 OR2X2_2515 ( .A(u2__abc_44228_n11907_1), .B(u2__abc_44228_n4307), .Y(u2__abc_44228_n11910) );
  OR2X2 OR2X2_2516 ( .A(u2__abc_44228_n11913), .B(u2__abc_44228_n2983_bF_buf94), .Y(u2__abc_44228_n11914_1) );
  OR2X2 OR2X2_2517 ( .A(u2__abc_44228_n11912), .B(u2__abc_44228_n11914_1), .Y(u2__abc_44228_n11915) );
  OR2X2 OR2X2_2518 ( .A(u2__abc_44228_n11919), .B(u2__abc_44228_n11905), .Y(u2__abc_44228_n11920) );
  OR2X2 OR2X2_2519 ( .A(u2__abc_44228_n5572), .B(u2__abc_44228_n6524), .Y(u2__abc_44228_n11924) );
  OR2X2 OR2X2_252 ( .A(a_112_bF_buf4), .B(\a[13] ), .Y(_abc_64468_n1209) );
  OR2X2 OR2X2_2520 ( .A(u2__abc_44228_n11928), .B(u2__abc_44228_n2983_bF_buf92), .Y(u2__abc_44228_n11929_1) );
  OR2X2 OR2X2_2521 ( .A(u2__abc_44228_n11929_1), .B(u2__abc_44228_n11923), .Y(u2__abc_44228_n11930) );
  OR2X2 OR2X2_2522 ( .A(u2__abc_44228_n11934), .B(u2__abc_44228_n11922_1), .Y(u2__abc_44228_n11935) );
  OR2X2 OR2X2_2523 ( .A(u2__abc_44228_n11942), .B(u2__abc_44228_n11943), .Y(u2__abc_44228_n11944) );
  OR2X2 OR2X2_2524 ( .A(u2__abc_44228_n11945), .B(u2__abc_44228_n2983_bF_buf90), .Y(u2__abc_44228_n11946) );
  OR2X2 OR2X2_2525 ( .A(u2__abc_44228_n11946), .B(u2__abc_44228_n11938), .Y(u2__abc_44228_n11947_1) );
  OR2X2 OR2X2_2526 ( .A(u2__abc_44228_n11951), .B(u2__abc_44228_n11937), .Y(u2__abc_44228_n11952) );
  OR2X2 OR2X2_2527 ( .A(u2__abc_44228_n11955_1), .B(u2__abc_44228_n6536), .Y(u2__abc_44228_n11956) );
  OR2X2 OR2X2_2528 ( .A(u2__abc_44228_n11956), .B(u2__abc_44228_n6510), .Y(u2__abc_44228_n11959) );
  OR2X2 OR2X2_2529 ( .A(u2__abc_44228_n7548_1_bF_buf31), .B(u2__abc_44228_n11960), .Y(u2__abc_44228_n11961) );
  OR2X2 OR2X2_253 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[14] ), .Y(_abc_64468_n1210) );
  OR2X2 OR2X2_2530 ( .A(u2__abc_44228_n7547_bF_buf30), .B(u2_remHi_256_), .Y(u2__abc_44228_n11962_1) );
  OR2X2 OR2X2_2531 ( .A(u2__abc_44228_n11963), .B(u2__abc_44228_n2983_bF_buf88), .Y(u2__abc_44228_n11964) );
  OR2X2 OR2X2_2532 ( .A(u2__abc_44228_n11968), .B(u2__abc_44228_n11954), .Y(u2__abc_44228_n11969) );
  OR2X2 OR2X2_2533 ( .A(u2__abc_44228_n11957), .B(u2__abc_44228_n6506), .Y(u2__abc_44228_n11972) );
  OR2X2 OR2X2_2534 ( .A(u2__abc_44228_n11972), .B(u2__abc_44228_n6504), .Y(u2__abc_44228_n11973) );
  OR2X2 OR2X2_2535 ( .A(u2__abc_44228_n11975), .B(u2__abc_44228_n11974), .Y(u2__abc_44228_n11976) );
  OR2X2 OR2X2_2536 ( .A(u2__abc_44228_n11979), .B(u2__abc_44228_n2983_bF_buf86), .Y(u2__abc_44228_n11980) );
  OR2X2 OR2X2_2537 ( .A(u2__abc_44228_n11980), .B(u2__abc_44228_n11978_1), .Y(u2__abc_44228_n11981) );
  OR2X2 OR2X2_2538 ( .A(u2__abc_44228_n11985), .B(u2__abc_44228_n11971_1), .Y(u2__abc_44228_n11986_1) );
  OR2X2 OR2X2_2539 ( .A(u2__abc_44228_n11989), .B(u2__abc_44228_n6540), .Y(u2__abc_44228_n11990) );
  OR2X2 OR2X2_254 ( .A(a_112_bF_buf3), .B(\a[14] ), .Y(_abc_64468_n1212) );
  OR2X2 OR2X2_2540 ( .A(u2__abc_44228_n11990), .B(u2__abc_44228_n6495), .Y(u2__abc_44228_n11991) );
  OR2X2 OR2X2_2541 ( .A(u2__abc_44228_n7548_1_bF_buf29), .B(u2__abc_44228_n11994), .Y(u2__abc_44228_n11995) );
  OR2X2 OR2X2_2542 ( .A(u2__abc_44228_n7547_bF_buf28), .B(u2_remHi_258_), .Y(u2__abc_44228_n11996) );
  OR2X2 OR2X2_2543 ( .A(u2__abc_44228_n11997), .B(u2__abc_44228_n2983_bF_buf84), .Y(u2__abc_44228_n11998) );
  OR2X2 OR2X2_2544 ( .A(u2__abc_44228_n12002), .B(u2__abc_44228_n11988), .Y(u2__abc_44228_n12003_1) );
  OR2X2 OR2X2_2545 ( .A(u2__abc_44228_n12007), .B(u2__abc_44228_n12006), .Y(u2__abc_44228_n12008) );
  OR2X2 OR2X2_2546 ( .A(u2__abc_44228_n12009), .B(u2__abc_44228_n6489_1), .Y(u2__abc_44228_n12010_1) );
  OR2X2 OR2X2_2547 ( .A(u2__abc_44228_n12013), .B(u2__abc_44228_n2983_bF_buf82), .Y(u2__abc_44228_n12014) );
  OR2X2 OR2X2_2548 ( .A(u2__abc_44228_n12014), .B(u2__abc_44228_n12012), .Y(u2__abc_44228_n12015) );
  OR2X2 OR2X2_2549 ( .A(u2__abc_44228_n12019), .B(u2__abc_44228_n12005), .Y(u2__abc_44228_n12020) );
  OR2X2 OR2X2_255 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[15] ), .Y(_abc_64468_n1213) );
  OR2X2 OR2X2_2550 ( .A(u2__abc_44228_n12023), .B(u2__abc_44228_n6545), .Y(u2__abc_44228_n12024) );
  OR2X2 OR2X2_2551 ( .A(u2__abc_44228_n12024), .B(u2__abc_44228_n6481), .Y(u2__abc_44228_n12027) );
  OR2X2 OR2X2_2552 ( .A(u2__abc_44228_n7548_1_bF_buf27), .B(u2__abc_44228_n12028), .Y(u2__abc_44228_n12029) );
  OR2X2 OR2X2_2553 ( .A(u2__abc_44228_n7547_bF_buf26), .B(u2_remHi_260_), .Y(u2__abc_44228_n12030) );
  OR2X2 OR2X2_2554 ( .A(u2__abc_44228_n12031), .B(u2__abc_44228_n2983_bF_buf80), .Y(u2__abc_44228_n12032) );
  OR2X2 OR2X2_2555 ( .A(u2__abc_44228_n12036), .B(u2__abc_44228_n12022), .Y(u2__abc_44228_n12037) );
  OR2X2 OR2X2_2556 ( .A(u2__abc_44228_n12025_1), .B(u2__abc_44228_n6477), .Y(u2__abc_44228_n12041_1) );
  OR2X2 OR2X2_2557 ( .A(u2__abc_44228_n12042), .B(u2__abc_44228_n12040), .Y(u2__abc_44228_n12043) );
  OR2X2 OR2X2_2558 ( .A(u2__abc_44228_n12041_1), .B(u2__abc_44228_n6475), .Y(u2__abc_44228_n12044) );
  OR2X2 OR2X2_2559 ( .A(u2__abc_44228_n12047), .B(u2__abc_44228_n2983_bF_buf78), .Y(u2__abc_44228_n12048) );
  OR2X2 OR2X2_256 ( .A(a_112_bF_buf2), .B(\a[15] ), .Y(_abc_64468_n1215) );
  OR2X2 OR2X2_2560 ( .A(u2__abc_44228_n12046), .B(u2__abc_44228_n12048), .Y(u2__abc_44228_n12049_1) );
  OR2X2 OR2X2_2561 ( .A(u2__abc_44228_n12053), .B(u2__abc_44228_n12039), .Y(u2__abc_44228_n12054) );
  OR2X2 OR2X2_2562 ( .A(u2__abc_44228_n12057), .B(u2__abc_44228_n6550), .Y(u2__abc_44228_n12058) );
  OR2X2 OR2X2_2563 ( .A(u2__abc_44228_n12058), .B(u2__abc_44228_n6465), .Y(u2__abc_44228_n12061) );
  OR2X2 OR2X2_2564 ( .A(u2__abc_44228_n7548_1_bF_buf25), .B(u2__abc_44228_n12062), .Y(u2__abc_44228_n12063) );
  OR2X2 OR2X2_2565 ( .A(u2__abc_44228_n7547_bF_buf24), .B(u2_remHi_262_), .Y(u2__abc_44228_n12064) );
  OR2X2 OR2X2_2566 ( .A(u2__abc_44228_n12065), .B(u2__abc_44228_n2983_bF_buf76), .Y(u2__abc_44228_n12066) );
  OR2X2 OR2X2_2567 ( .A(u2__abc_44228_n12070), .B(u2__abc_44228_n12056_1), .Y(u2__abc_44228_n12071) );
  OR2X2 OR2X2_2568 ( .A(u2__abc_44228_n12075), .B(u2__abc_44228_n12074_1), .Y(u2__abc_44228_n12076) );
  OR2X2 OR2X2_2569 ( .A(u2__abc_44228_n12077), .B(u2__abc_44228_n6459), .Y(u2__abc_44228_n12078) );
  OR2X2 OR2X2_257 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[16] ), .Y(_abc_64468_n1216) );
  OR2X2 OR2X2_2570 ( .A(u2__abc_44228_n12081), .B(u2__abc_44228_n2983_bF_buf74), .Y(u2__abc_44228_n12082_1) );
  OR2X2 OR2X2_2571 ( .A(u2__abc_44228_n12082_1), .B(u2__abc_44228_n12080), .Y(u2__abc_44228_n12083) );
  OR2X2 OR2X2_2572 ( .A(u2__abc_44228_n12087), .B(u2__abc_44228_n12073), .Y(u2__abc_44228_n12088) );
  OR2X2 OR2X2_2573 ( .A(u2__abc_44228_n12091), .B(u2__abc_44228_n6457), .Y(u2__abc_44228_n12092) );
  OR2X2 OR2X2_2574 ( .A(u2__abc_44228_n12093), .B(u2__abc_44228_n6451), .Y(u2__abc_44228_n12096) );
  OR2X2 OR2X2_2575 ( .A(u2__abc_44228_n12099), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n12100) );
  OR2X2 OR2X2_2576 ( .A(u2__abc_44228_n12098_1), .B(u2__abc_44228_n12100), .Y(u2__abc_44228_n12101) );
  OR2X2 OR2X2_2577 ( .A(u2__abc_44228_n12105_1), .B(u2__abc_44228_n12090), .Y(u2__abc_44228_n12106) );
  OR2X2 OR2X2_2578 ( .A(u2__abc_44228_n12094), .B(u2__abc_44228_n6447), .Y(u2__abc_44228_n12110) );
  OR2X2 OR2X2_2579 ( .A(u2__abc_44228_n12111), .B(u2__abc_44228_n12109), .Y(u2__abc_44228_n12112) );
  OR2X2 OR2X2_258 ( .A(a_112_bF_buf1), .B(\a[16] ), .Y(_abc_64468_n1218) );
  OR2X2 OR2X2_2580 ( .A(u2__abc_44228_n12110), .B(u2__abc_44228_n6445_1), .Y(u2__abc_44228_n12113_1) );
  OR2X2 OR2X2_2581 ( .A(u2__abc_44228_n12116), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n12117) );
  OR2X2 OR2X2_2582 ( .A(u2__abc_44228_n12115), .B(u2__abc_44228_n12117), .Y(u2__abc_44228_n12118) );
  OR2X2 OR2X2_2583 ( .A(u2__abc_44228_n12122), .B(u2__abc_44228_n12108), .Y(u2__abc_44228_n12123) );
  OR2X2 OR2X2_2584 ( .A(u2__abc_44228_n12126), .B(u2__abc_44228_n6559), .Y(u2__abc_44228_n12127) );
  OR2X2 OR2X2_2585 ( .A(u2__abc_44228_n12127), .B(u2__abc_44228_n6436), .Y(u2__abc_44228_n12128) );
  OR2X2 OR2X2_2586 ( .A(u2__abc_44228_n7548_1_bF_buf21), .B(u2__abc_44228_n12131), .Y(u2__abc_44228_n12132) );
  OR2X2 OR2X2_2587 ( .A(u2__abc_44228_n7547_bF_buf20), .B(u2_remHi_266_), .Y(u2__abc_44228_n12133) );
  OR2X2 OR2X2_2588 ( .A(u2__abc_44228_n12134), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n12135) );
  OR2X2 OR2X2_2589 ( .A(u2__abc_44228_n12139), .B(u2__abc_44228_n12125), .Y(u2__abc_44228_n12140) );
  OR2X2 OR2X2_259 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[17] ), .Y(_abc_64468_n1219) );
  OR2X2 OR2X2_2590 ( .A(u2__abc_44228_n12144), .B(u2__abc_44228_n12143), .Y(u2__abc_44228_n12145_1) );
  OR2X2 OR2X2_2591 ( .A(u2__abc_44228_n12146), .B(u2__abc_44228_n6430), .Y(u2__abc_44228_n12147) );
  OR2X2 OR2X2_2592 ( .A(u2__abc_44228_n12150), .B(u2__abc_44228_n2983_bF_buf67), .Y(u2__abc_44228_n12151) );
  OR2X2 OR2X2_2593 ( .A(u2__abc_44228_n12149), .B(u2__abc_44228_n12151), .Y(u2__abc_44228_n12152_1) );
  OR2X2 OR2X2_2594 ( .A(u2__abc_44228_n12156), .B(u2__abc_44228_n12142), .Y(u2__abc_44228_n12157) );
  OR2X2 OR2X2_2595 ( .A(u2__abc_44228_n12160), .B(u2__abc_44228_n6564), .Y(u2__abc_44228_n12161_1) );
  OR2X2 OR2X2_2596 ( .A(u2__abc_44228_n12161_1), .B(u2__abc_44228_n6422), .Y(u2__abc_44228_n12164) );
  OR2X2 OR2X2_2597 ( .A(u2__abc_44228_n12167), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n12168_1) );
  OR2X2 OR2X2_2598 ( .A(u2__abc_44228_n12166), .B(u2__abc_44228_n12168_1), .Y(u2__abc_44228_n12169) );
  OR2X2 OR2X2_2599 ( .A(u2__abc_44228_n12173), .B(u2__abc_44228_n12159), .Y(u2__abc_44228_n12174) );
  OR2X2 OR2X2_26 ( .A(_abc_64468_n753_bF_buf9), .B(\a[12] ), .Y(_abc_64468_n867) );
  OR2X2 OR2X2_260 ( .A(a_112_bF_buf0), .B(\a[17] ), .Y(_abc_64468_n1221) );
  OR2X2 OR2X2_2600 ( .A(u2__abc_44228_n12162), .B(u2__abc_44228_n6418), .Y(u2__abc_44228_n12178) );
  OR2X2 OR2X2_2601 ( .A(u2__abc_44228_n12179), .B(u2__abc_44228_n12177), .Y(u2__abc_44228_n12180) );
  OR2X2 OR2X2_2602 ( .A(u2__abc_44228_n12178), .B(u2__abc_44228_n6416), .Y(u2__abc_44228_n12181) );
  OR2X2 OR2X2_2603 ( .A(u2__abc_44228_n12184), .B(u2__abc_44228_n2983_bF_buf64), .Y(u2__abc_44228_n12185) );
  OR2X2 OR2X2_2604 ( .A(u2__abc_44228_n12183_1), .B(u2__abc_44228_n12185), .Y(u2__abc_44228_n12186) );
  OR2X2 OR2X2_2605 ( .A(u2__abc_44228_n12190), .B(u2__abc_44228_n12176_1), .Y(u2__abc_44228_n12191) );
  OR2X2 OR2X2_2606 ( .A(u2__abc_44228_n12194), .B(u2__abc_44228_n6570), .Y(u2__abc_44228_n12195_1) );
  OR2X2 OR2X2_2607 ( .A(u2__abc_44228_n12195_1), .B(u2__abc_44228_n6398), .Y(u2__abc_44228_n12196) );
  OR2X2 OR2X2_2608 ( .A(u2__abc_44228_n7548_1_bF_buf17), .B(u2__abc_44228_n12199), .Y(u2__abc_44228_n12200) );
  OR2X2 OR2X2_2609 ( .A(u2__abc_44228_n7547_bF_buf16), .B(u2_remHi_270_), .Y(u2__abc_44228_n12201) );
  OR2X2 OR2X2_261 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[18] ), .Y(_abc_64468_n1222) );
  OR2X2 OR2X2_2610 ( .A(u2__abc_44228_n12202_1), .B(u2__abc_44228_n2983_bF_buf62), .Y(u2__abc_44228_n12203) );
  OR2X2 OR2X2_2611 ( .A(u2__abc_44228_n12207), .B(u2__abc_44228_n12193), .Y(u2__abc_44228_n12208) );
  OR2X2 OR2X2_2612 ( .A(u2__abc_44228_n12212), .B(u2__abc_44228_n12211), .Y(u2__abc_44228_n12213) );
  OR2X2 OR2X2_2613 ( .A(u2__abc_44228_n12214), .B(u2__abc_44228_n6405), .Y(u2__abc_44228_n12215) );
  OR2X2 OR2X2_2614 ( .A(u2__abc_44228_n12218), .B(u2__abc_44228_n2983_bF_buf60), .Y(u2__abc_44228_n12219) );
  OR2X2 OR2X2_2615 ( .A(u2__abc_44228_n12219), .B(u2__abc_44228_n12217_1), .Y(u2__abc_44228_n12220) );
  OR2X2 OR2X2_2616 ( .A(u2__abc_44228_n12224), .B(u2__abc_44228_n12210_1), .Y(u2__abc_44228_n12225) );
  OR2X2 OR2X2_2617 ( .A(u2__abc_44228_n12228), .B(u2__abc_44228_n6403), .Y(u2__abc_44228_n12229) );
  OR2X2 OR2X2_2618 ( .A(u2__abc_44228_n12230), .B(u2__abc_44228_n6391), .Y(u2__abc_44228_n12233_1) );
  OR2X2 OR2X2_2619 ( .A(u2__abc_44228_n12236), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n12237) );
  OR2X2 OR2X2_262 ( .A(a_112_bF_buf9), .B(\a[18] ), .Y(_abc_64468_n1224) );
  OR2X2 OR2X2_2620 ( .A(u2__abc_44228_n12235), .B(u2__abc_44228_n12237), .Y(u2__abc_44228_n12238) );
  OR2X2 OR2X2_2621 ( .A(u2__abc_44228_n12242), .B(u2__abc_44228_n12227), .Y(u2__abc_44228_n12243) );
  OR2X2 OR2X2_2622 ( .A(u2__abc_44228_n12231), .B(u2__abc_44228_n6387), .Y(u2__abc_44228_n12247) );
  OR2X2 OR2X2_2623 ( .A(u2__abc_44228_n12248_1), .B(u2__abc_44228_n12246), .Y(u2__abc_44228_n12249) );
  OR2X2 OR2X2_2624 ( .A(u2__abc_44228_n12247), .B(u2__abc_44228_n6385), .Y(u2__abc_44228_n12250) );
  OR2X2 OR2X2_2625 ( .A(u2__abc_44228_n12253), .B(u2__abc_44228_n2983_bF_buf57), .Y(u2__abc_44228_n12254) );
  OR2X2 OR2X2_2626 ( .A(u2__abc_44228_n12252), .B(u2__abc_44228_n12254), .Y(u2__abc_44228_n12255) );
  OR2X2 OR2X2_2627 ( .A(u2__abc_44228_n12259), .B(u2__abc_44228_n12245), .Y(u2__abc_44228_n12260) );
  OR2X2 OR2X2_2628 ( .A(u2__abc_44228_n12263), .B(u2__abc_44228_n6579_1), .Y(u2__abc_44228_n12264) );
  OR2X2 OR2X2_2629 ( .A(u2__abc_44228_n12264), .B(u2__abc_44228_n6376), .Y(u2__abc_44228_n12265_1) );
  OR2X2 OR2X2_263 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[19] ), .Y(_abc_64468_n1225) );
  OR2X2 OR2X2_2630 ( .A(u2__abc_44228_n7548_1_bF_buf13), .B(u2__abc_44228_n12268), .Y(u2__abc_44228_n12269) );
  OR2X2 OR2X2_2631 ( .A(u2__abc_44228_n7547_bF_buf12), .B(u2_remHi_274_), .Y(u2__abc_44228_n12270) );
  OR2X2 OR2X2_2632 ( .A(u2__abc_44228_n12271), .B(u2__abc_44228_n2983_bF_buf55), .Y(u2__abc_44228_n12272) );
  OR2X2 OR2X2_2633 ( .A(u2__abc_44228_n12276), .B(u2__abc_44228_n12262), .Y(u2__abc_44228_n12277) );
  OR2X2 OR2X2_2634 ( .A(u2__abc_44228_n12281), .B(u2__abc_44228_n12280_1), .Y(u2__abc_44228_n12282) );
  OR2X2 OR2X2_2635 ( .A(u2__abc_44228_n12283), .B(u2__abc_44228_n6370), .Y(u2__abc_44228_n12284) );
  OR2X2 OR2X2_2636 ( .A(u2__abc_44228_n12287), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n12288) );
  OR2X2 OR2X2_2637 ( .A(u2__abc_44228_n12286), .B(u2__abc_44228_n12288), .Y(u2__abc_44228_n12289_1) );
  OR2X2 OR2X2_2638 ( .A(u2__abc_44228_n12293), .B(u2__abc_44228_n12279), .Y(u2__abc_44228_n12294) );
  OR2X2 OR2X2_2639 ( .A(u2__abc_44228_n12297), .B(u2__abc_44228_n6584), .Y(u2__abc_44228_n12298) );
  OR2X2 OR2X2_264 ( .A(a_112_bF_buf8), .B(\a[19] ), .Y(_abc_64468_n1227) );
  OR2X2 OR2X2_2640 ( .A(u2__abc_44228_n12298), .B(u2__abc_44228_n6362), .Y(u2__abc_44228_n12301) );
  OR2X2 OR2X2_2641 ( .A(u2__abc_44228_n12304_1), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n12305) );
  OR2X2 OR2X2_2642 ( .A(u2__abc_44228_n12303), .B(u2__abc_44228_n12305), .Y(u2__abc_44228_n12306) );
  OR2X2 OR2X2_2643 ( .A(u2__abc_44228_n12310), .B(u2__abc_44228_n12296_1), .Y(u2__abc_44228_n12311_1) );
  OR2X2 OR2X2_2644 ( .A(u2__abc_44228_n12299), .B(u2__abc_44228_n6358), .Y(u2__abc_44228_n12315) );
  OR2X2 OR2X2_2645 ( .A(u2__abc_44228_n12316), .B(u2__abc_44228_n12314), .Y(u2__abc_44228_n12317) );
  OR2X2 OR2X2_2646 ( .A(u2__abc_44228_n12315), .B(u2__abc_44228_n6356), .Y(u2__abc_44228_n12318) );
  OR2X2 OR2X2_2647 ( .A(u2__abc_44228_n12321), .B(u2__abc_44228_n2983_bF_buf50), .Y(u2__abc_44228_n12322_1) );
  OR2X2 OR2X2_2648 ( .A(u2__abc_44228_n12320), .B(u2__abc_44228_n12322_1), .Y(u2__abc_44228_n12323) );
  OR2X2 OR2X2_2649 ( .A(u2__abc_44228_n12327), .B(u2__abc_44228_n12313), .Y(u2__abc_44228_n12328) );
  OR2X2 OR2X2_265 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[20] ), .Y(_abc_64468_n1228) );
  OR2X2 OR2X2_2650 ( .A(u2__abc_44228_n12331), .B(u2__abc_44228_n6589), .Y(u2__abc_44228_n12332) );
  OR2X2 OR2X2_2651 ( .A(u2__abc_44228_n12332), .B(u2__abc_44228_n6332), .Y(u2__abc_44228_n12335) );
  OR2X2 OR2X2_2652 ( .A(u2__abc_44228_n7548_1_bF_buf9), .B(u2__abc_44228_n12336), .Y(u2__abc_44228_n12337_1) );
  OR2X2 OR2X2_2653 ( .A(u2__abc_44228_n7547_bF_buf8), .B(u2_remHi_278_), .Y(u2__abc_44228_n12338) );
  OR2X2 OR2X2_2654 ( .A(u2__abc_44228_n12339), .B(u2__abc_44228_n2983_bF_buf48), .Y(u2__abc_44228_n12340) );
  OR2X2 OR2X2_2655 ( .A(u2__abc_44228_n12344_1), .B(u2__abc_44228_n12330), .Y(u2__abc_44228_n12345) );
  OR2X2 OR2X2_2656 ( .A(u2__abc_44228_n12349), .B(u2__abc_44228_n12348), .Y(u2__abc_44228_n12350) );
  OR2X2 OR2X2_2657 ( .A(u2__abc_44228_n12351), .B(u2__abc_44228_n6326), .Y(u2__abc_44228_n12352) );
  OR2X2 OR2X2_2658 ( .A(u2__abc_44228_n12355), .B(u2__abc_44228_n2983_bF_buf46), .Y(u2__abc_44228_n12356) );
  OR2X2 OR2X2_2659 ( .A(u2__abc_44228_n12354), .B(u2__abc_44228_n12356), .Y(u2__abc_44228_n12357) );
  OR2X2 OR2X2_266 ( .A(a_112_bF_buf7), .B(\a[20] ), .Y(_abc_64468_n1230) );
  OR2X2 OR2X2_2660 ( .A(u2__abc_44228_n12361), .B(u2__abc_44228_n12347), .Y(u2__abc_44228_n12362) );
  OR2X2 OR2X2_2661 ( .A(u2__abc_44228_n12365), .B(u2__abc_44228_n6594), .Y(u2__abc_44228_n12366) );
  OR2X2 OR2X2_2662 ( .A(u2__abc_44228_n12366), .B(u2__abc_44228_n6346), .Y(u2__abc_44228_n12369) );
  OR2X2 OR2X2_2663 ( .A(u2__abc_44228_n12372), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n12373) );
  OR2X2 OR2X2_2664 ( .A(u2__abc_44228_n12371), .B(u2__abc_44228_n12373), .Y(u2__abc_44228_n12374) );
  OR2X2 OR2X2_2665 ( .A(u2__abc_44228_n12378), .B(u2__abc_44228_n12364), .Y(u2__abc_44228_n12379) );
  OR2X2 OR2X2_2666 ( .A(u2__abc_44228_n12383), .B(u2__abc_44228_n12382), .Y(u2__abc_44228_n12384) );
  OR2X2 OR2X2_2667 ( .A(u2__abc_44228_n12385_1), .B(u2__abc_44228_n6340), .Y(u2__abc_44228_n12386) );
  OR2X2 OR2X2_2668 ( .A(u2__abc_44228_n12389), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n12390) );
  OR2X2 OR2X2_2669 ( .A(u2__abc_44228_n12388), .B(u2__abc_44228_n12390), .Y(u2__abc_44228_n12391) );
  OR2X2 OR2X2_267 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[21] ), .Y(_abc_64468_n1231) );
  OR2X2 OR2X2_2670 ( .A(u2__abc_44228_n12395), .B(u2__abc_44228_n12381), .Y(u2__abc_44228_n12396) );
  OR2X2 OR2X2_2671 ( .A(u2__abc_44228_n12399), .B(u2__abc_44228_n6338), .Y(u2__abc_44228_n12400_1) );
  OR2X2 OR2X2_2672 ( .A(u2__abc_44228_n12401), .B(u2__abc_44228_n6317), .Y(u2__abc_44228_n12402) );
  OR2X2 OR2X2_2673 ( .A(u2__abc_44228_n12407_1), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n12408) );
  OR2X2 OR2X2_2674 ( .A(u2__abc_44228_n12406), .B(u2__abc_44228_n12408), .Y(u2__abc_44228_n12409) );
  OR2X2 OR2X2_2675 ( .A(u2__abc_44228_n12413), .B(u2__abc_44228_n12398), .Y(u2__abc_44228_n12414) );
  OR2X2 OR2X2_2676 ( .A(u2__abc_44228_n12421), .B(u2__abc_44228_n12418), .Y(u2__abc_44228_n12422) );
  OR2X2 OR2X2_2677 ( .A(u2__abc_44228_n12424), .B(u2__abc_44228_n2983_bF_buf40), .Y(u2__abc_44228_n12425) );
  OR2X2 OR2X2_2678 ( .A(u2__abc_44228_n12423_1), .B(u2__abc_44228_n12425), .Y(u2__abc_44228_n12426) );
  OR2X2 OR2X2_2679 ( .A(u2__abc_44228_n12430), .B(u2__abc_44228_n12416_1), .Y(u2__abc_44228_n12431_1) );
  OR2X2 OR2X2_268 ( .A(a_112_bF_buf6), .B(\a[21] ), .Y(_abc_64468_n1233) );
  OR2X2 OR2X2_2680 ( .A(u2__abc_44228_n12434), .B(u2__abc_44228_n6309), .Y(u2__abc_44228_n12435) );
  OR2X2 OR2X2_2681 ( .A(u2__abc_44228_n12436), .B(u2__abc_44228_n6303), .Y(u2__abc_44228_n12439) );
  OR2X2 OR2X2_2682 ( .A(u2__abc_44228_n12442), .B(u2__abc_44228_n2983_bF_buf38), .Y(u2__abc_44228_n12443) );
  OR2X2 OR2X2_2683 ( .A(u2__abc_44228_n12441), .B(u2__abc_44228_n12443), .Y(u2__abc_44228_n12444) );
  OR2X2 OR2X2_2684 ( .A(u2__abc_44228_n12448), .B(u2__abc_44228_n12433), .Y(u2__abc_44228_n12449) );
  OR2X2 OR2X2_2685 ( .A(u2__abc_44228_n12437), .B(u2__abc_44228_n6299), .Y(u2__abc_44228_n12453) );
  OR2X2 OR2X2_2686 ( .A(u2__abc_44228_n12454), .B(u2__abc_44228_n12452), .Y(u2__abc_44228_n12455) );
  OR2X2 OR2X2_2687 ( .A(u2__abc_44228_n12453), .B(u2__abc_44228_n6297), .Y(u2__abc_44228_n12456) );
  OR2X2 OR2X2_2688 ( .A(u2__abc_44228_n12459), .B(u2__abc_44228_n2983_bF_buf36), .Y(u2__abc_44228_n12460) );
  OR2X2 OR2X2_2689 ( .A(u2__abc_44228_n12458), .B(u2__abc_44228_n12460), .Y(u2__abc_44228_n12461) );
  OR2X2 OR2X2_269 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[22] ), .Y(_abc_64468_n1234) );
  OR2X2 OR2X2_2690 ( .A(u2__abc_44228_n12465_1), .B(u2__abc_44228_n12451), .Y(u2__abc_44228_n12466) );
  OR2X2 OR2X2_2691 ( .A(u2__abc_44228_n12469), .B(u2__abc_44228_n6612), .Y(u2__abc_44228_n12470) );
  OR2X2 OR2X2_2692 ( .A(u2__abc_44228_n12470), .B(u2__abc_44228_n6285), .Y(u2__abc_44228_n12473) );
  OR2X2 OR2X2_2693 ( .A(u2__abc_44228_n7548_1_bF_buf1), .B(u2__abc_44228_n12474), .Y(u2__abc_44228_n12475) );
  OR2X2 OR2X2_2694 ( .A(u2__abc_44228_n7547_bF_buf0), .B(u2_remHi_286_), .Y(u2__abc_44228_n12476) );
  OR2X2 OR2X2_2695 ( .A(u2__abc_44228_n12477), .B(u2__abc_44228_n2983_bF_buf34), .Y(u2__abc_44228_n12478) );
  OR2X2 OR2X2_2696 ( .A(u2__abc_44228_n12482), .B(u2__abc_44228_n12468), .Y(u2__abc_44228_n12483) );
  OR2X2 OR2X2_2697 ( .A(u2__abc_44228_n12487), .B(u2__abc_44228_n12486), .Y(u2__abc_44228_n12488_1) );
  OR2X2 OR2X2_2698 ( .A(u2__abc_44228_n12489), .B(u2__abc_44228_n6279_1), .Y(u2__abc_44228_n12490) );
  OR2X2 OR2X2_2699 ( .A(u2__abc_44228_n12493), .B(u2__abc_44228_n2983_bF_buf32), .Y(u2__abc_44228_n12494) );
  OR2X2 OR2X2_27 ( .A(aNan_bF_buf7), .B(sqrto_89_), .Y(_abc_64468_n869) );
  OR2X2 OR2X2_270 ( .A(a_112_bF_buf5), .B(\a[22] ), .Y(_abc_64468_n1236) );
  OR2X2 OR2X2_2700 ( .A(u2__abc_44228_n12494), .B(u2__abc_44228_n12492), .Y(u2__abc_44228_n12495) );
  OR2X2 OR2X2_2701 ( .A(u2__abc_44228_n12499), .B(u2__abc_44228_n12485), .Y(u2__abc_44228_n12500) );
  OR2X2 OR2X2_2702 ( .A(u2__abc_44228_n12503_1), .B(u2__abc_44228_n6617), .Y(u2__abc_44228_n12504) );
  OR2X2 OR2X2_2703 ( .A(u2__abc_44228_n12504), .B(u2__abc_44228_n6271), .Y(u2__abc_44228_n12507) );
  OR2X2 OR2X2_2704 ( .A(u2__abc_44228_n7548_1_bF_buf57), .B(u2__abc_44228_n12508), .Y(u2__abc_44228_n12509) );
  OR2X2 OR2X2_2705 ( .A(u2__abc_44228_n7547_bF_buf56), .B(u2_remHi_288_), .Y(u2__abc_44228_n12510) );
  OR2X2 OR2X2_2706 ( .A(u2__abc_44228_n12511), .B(u2__abc_44228_n2983_bF_buf30), .Y(u2__abc_44228_n12512) );
  OR2X2 OR2X2_2707 ( .A(u2__abc_44228_n12516), .B(u2__abc_44228_n12502), .Y(u2__abc_44228_n12517) );
  OR2X2 OR2X2_2708 ( .A(u2__abc_44228_n12505), .B(u2__abc_44228_n6267), .Y(u2__abc_44228_n12521) );
  OR2X2 OR2X2_2709 ( .A(u2__abc_44228_n12522), .B(u2__abc_44228_n12520_1), .Y(u2__abc_44228_n12523) );
  OR2X2 OR2X2_271 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[23] ), .Y(_abc_64468_n1237) );
  OR2X2 OR2X2_2710 ( .A(u2__abc_44228_n12521), .B(u2__abc_44228_n6265), .Y(u2__abc_44228_n12524) );
  OR2X2 OR2X2_2711 ( .A(u2__abc_44228_n12527), .B(u2__abc_44228_n2983_bF_buf28), .Y(u2__abc_44228_n12528_1) );
  OR2X2 OR2X2_2712 ( .A(u2__abc_44228_n12526), .B(u2__abc_44228_n12528_1), .Y(u2__abc_44228_n12529) );
  OR2X2 OR2X2_2713 ( .A(u2__abc_44228_n12533), .B(u2__abc_44228_n12519), .Y(u2__abc_44228_n12534) );
  OR2X2 OR2X2_2714 ( .A(u2__abc_44228_n12537), .B(u2__abc_44228_n6621), .Y(u2__abc_44228_n12538) );
  OR2X2 OR2X2_2715 ( .A(u2__abc_44228_n12538), .B(u2__abc_44228_n6256), .Y(u2__abc_44228_n12539) );
  OR2X2 OR2X2_2716 ( .A(u2__abc_44228_n7548_1_bF_buf55), .B(u2__abc_44228_n12542), .Y(u2__abc_44228_n12543) );
  OR2X2 OR2X2_2717 ( .A(u2__abc_44228_n7547_bF_buf54), .B(u2_remHi_290_), .Y(u2__abc_44228_n12544_1) );
  OR2X2 OR2X2_2718 ( .A(u2__abc_44228_n12545), .B(u2__abc_44228_n2983_bF_buf26), .Y(u2__abc_44228_n12546) );
  OR2X2 OR2X2_2719 ( .A(u2__abc_44228_n12550), .B(u2__abc_44228_n12536), .Y(u2__abc_44228_n12551_1) );
  OR2X2 OR2X2_272 ( .A(a_112_bF_buf4), .B(\a[23] ), .Y(_abc_64468_n1239) );
  OR2X2 OR2X2_2720 ( .A(u2__abc_44228_n12555), .B(u2__abc_44228_n12554), .Y(u2__abc_44228_n12556) );
  OR2X2 OR2X2_2721 ( .A(u2__abc_44228_n12557), .B(u2__abc_44228_n6250), .Y(u2__abc_44228_n12558) );
  OR2X2 OR2X2_2722 ( .A(u2__abc_44228_n12561), .B(u2__abc_44228_n2983_bF_buf24), .Y(u2__abc_44228_n12562) );
  OR2X2 OR2X2_2723 ( .A(u2__abc_44228_n12560), .B(u2__abc_44228_n12562), .Y(u2__abc_44228_n12563) );
  OR2X2 OR2X2_2724 ( .A(u2__abc_44228_n12567), .B(u2__abc_44228_n12553), .Y(u2__abc_44228_n12568) );
  OR2X2 OR2X2_2725 ( .A(u2__abc_44228_n12571), .B(u2__abc_44228_n6626), .Y(u2__abc_44228_n12572) );
  OR2X2 OR2X2_2726 ( .A(u2__abc_44228_n12572), .B(u2__abc_44228_n6242_1), .Y(u2__abc_44228_n12575) );
  OR2X2 OR2X2_2727 ( .A(u2__abc_44228_n12578), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n12579) );
  OR2X2 OR2X2_2728 ( .A(u2__abc_44228_n12577_1), .B(u2__abc_44228_n12579), .Y(u2__abc_44228_n12580) );
  OR2X2 OR2X2_2729 ( .A(u2__abc_44228_n12584_1), .B(u2__abc_44228_n12570), .Y(u2__abc_44228_n12585) );
  OR2X2 OR2X2_273 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[24] ), .Y(_abc_64468_n1240) );
  OR2X2 OR2X2_2730 ( .A(u2__abc_44228_n12573), .B(u2__abc_44228_n6238), .Y(u2__abc_44228_n12589) );
  OR2X2 OR2X2_2731 ( .A(u2__abc_44228_n12590), .B(u2__abc_44228_n12588), .Y(u2__abc_44228_n12591) );
  OR2X2 OR2X2_2732 ( .A(u2__abc_44228_n12589), .B(u2__abc_44228_n6236), .Y(u2__abc_44228_n12592_1) );
  OR2X2 OR2X2_2733 ( .A(u2__abc_44228_n12595), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n12596) );
  OR2X2 OR2X2_2734 ( .A(u2__abc_44228_n12594), .B(u2__abc_44228_n12596), .Y(u2__abc_44228_n12597) );
  OR2X2 OR2X2_2735 ( .A(u2__abc_44228_n12601), .B(u2__abc_44228_n12587), .Y(u2__abc_44228_n12602) );
  OR2X2 OR2X2_2736 ( .A(u2__abc_44228_n12605), .B(u2__abc_44228_n6631), .Y(u2__abc_44228_n12606) );
  OR2X2 OR2X2_2737 ( .A(u2__abc_44228_n12606), .B(u2__abc_44228_n6212), .Y(u2__abc_44228_n12609) );
  OR2X2 OR2X2_2738 ( .A(u2__abc_44228_n7548_1_bF_buf51), .B(u2__abc_44228_n12610), .Y(u2__abc_44228_n12611) );
  OR2X2 OR2X2_2739 ( .A(u2__abc_44228_n7547_bF_buf50), .B(u2_remHi_294_), .Y(u2__abc_44228_n12612) );
  OR2X2 OR2X2_274 ( .A(a_112_bF_buf3), .B(\a[24] ), .Y(_abc_64468_n1242) );
  OR2X2 OR2X2_2740 ( .A(u2__abc_44228_n12613), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n12614) );
  OR2X2 OR2X2_2741 ( .A(u2__abc_44228_n12618), .B(u2__abc_44228_n12604), .Y(u2__abc_44228_n12619) );
  OR2X2 OR2X2_2742 ( .A(u2__abc_44228_n12623_1), .B(u2__abc_44228_n12622), .Y(u2__abc_44228_n12624) );
  OR2X2 OR2X2_2743 ( .A(u2__abc_44228_n12625), .B(u2__abc_44228_n6206_1), .Y(u2__abc_44228_n12626) );
  OR2X2 OR2X2_2744 ( .A(u2__abc_44228_n12629), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n12630_1) );
  OR2X2 OR2X2_2745 ( .A(u2__abc_44228_n12628), .B(u2__abc_44228_n12630_1), .Y(u2__abc_44228_n12631) );
  OR2X2 OR2X2_2746 ( .A(u2__abc_44228_n12635), .B(u2__abc_44228_n12621), .Y(u2__abc_44228_n12636) );
  OR2X2 OR2X2_2747 ( .A(u2__abc_44228_n12639), .B(u2__abc_44228_n6636), .Y(u2__abc_44228_n12640_1) );
  OR2X2 OR2X2_2748 ( .A(u2__abc_44228_n12640_1), .B(u2__abc_44228_n6226), .Y(u2__abc_44228_n12643) );
  OR2X2 OR2X2_2749 ( .A(u2__abc_44228_n12646), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n12647_1) );
  OR2X2 OR2X2_275 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[25] ), .Y(_abc_64468_n1243) );
  OR2X2 OR2X2_2750 ( .A(u2__abc_44228_n12645), .B(u2__abc_44228_n12647_1), .Y(u2__abc_44228_n12648) );
  OR2X2 OR2X2_2751 ( .A(u2__abc_44228_n12652), .B(u2__abc_44228_n12638), .Y(u2__abc_44228_n12653) );
  OR2X2 OR2X2_2752 ( .A(u2__abc_44228_n12657), .B(u2__abc_44228_n12656), .Y(u2__abc_44228_n12658) );
  OR2X2 OR2X2_2753 ( .A(u2__abc_44228_n12659), .B(u2__abc_44228_n6220), .Y(u2__abc_44228_n12660) );
  OR2X2 OR2X2_2754 ( .A(u2__abc_44228_n12663), .B(u2__abc_44228_n2983_bF_buf14), .Y(u2__abc_44228_n12664) );
  OR2X2 OR2X2_2755 ( .A(u2__abc_44228_n12662_1), .B(u2__abc_44228_n12664), .Y(u2__abc_44228_n12665) );
  OR2X2 OR2X2_2756 ( .A(u2__abc_44228_n12669), .B(u2__abc_44228_n12655_1), .Y(u2__abc_44228_n12670) );
  OR2X2 OR2X2_2757 ( .A(u2__abc_44228_n12673), .B(u2__abc_44228_n6218), .Y(u2__abc_44228_n12674) );
  OR2X2 OR2X2_2758 ( .A(u2__abc_44228_n12675), .B(u2__abc_44228_n6197), .Y(u2__abc_44228_n12676) );
  OR2X2 OR2X2_2759 ( .A(u2__abc_44228_n12681), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n12682) );
  OR2X2 OR2X2_276 ( .A(a_112_bF_buf2), .B(\a[25] ), .Y(_abc_64468_n1245) );
  OR2X2 OR2X2_2760 ( .A(u2__abc_44228_n12680), .B(u2__abc_44228_n12682), .Y(u2__abc_44228_n12683) );
  OR2X2 OR2X2_2761 ( .A(u2__abc_44228_n12687), .B(u2__abc_44228_n12672), .Y(u2__abc_44228_n12688) );
  OR2X2 OR2X2_2762 ( .A(u2__abc_44228_n12692), .B(u2__abc_44228_n6191), .Y(u2__abc_44228_n12693_1) );
  OR2X2 OR2X2_2763 ( .A(u2__abc_44228_n12691), .B(u2__abc_44228_n12694), .Y(u2__abc_44228_n12695) );
  OR2X2 OR2X2_2764 ( .A(u2__abc_44228_n12698), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n12699) );
  OR2X2 OR2X2_2765 ( .A(u2__abc_44228_n12697), .B(u2__abc_44228_n12699), .Y(u2__abc_44228_n12700) );
  OR2X2 OR2X2_2766 ( .A(u2__abc_44228_n12704), .B(u2__abc_44228_n12690), .Y(u2__abc_44228_n12705) );
  OR2X2 OR2X2_2767 ( .A(u2__abc_44228_n12708), .B(u2__abc_44228_n6189), .Y(u2__abc_44228_n12709) );
  OR2X2 OR2X2_2768 ( .A(u2__abc_44228_n12710), .B(u2__abc_44228_n6183), .Y(u2__abc_44228_n12713_1) );
  OR2X2 OR2X2_2769 ( .A(u2__abc_44228_n12716), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n12717) );
  OR2X2 OR2X2_277 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[26] ), .Y(_abc_64468_n1246) );
  OR2X2 OR2X2_2770 ( .A(u2__abc_44228_n12715), .B(u2__abc_44228_n12717), .Y(u2__abc_44228_n12718) );
  OR2X2 OR2X2_2771 ( .A(u2__abc_44228_n12722), .B(u2__abc_44228_n12707), .Y(u2__abc_44228_n12723) );
  OR2X2 OR2X2_2772 ( .A(u2__abc_44228_n12711), .B(u2__abc_44228_n6179), .Y(u2__abc_44228_n12727) );
  OR2X2 OR2X2_2773 ( .A(u2__abc_44228_n12728_1), .B(u2__abc_44228_n12726), .Y(u2__abc_44228_n12729) );
  OR2X2 OR2X2_2774 ( .A(u2__abc_44228_n12727), .B(u2__abc_44228_n6177), .Y(u2__abc_44228_n12730) );
  OR2X2 OR2X2_2775 ( .A(u2__abc_44228_n12733), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n12734) );
  OR2X2 OR2X2_2776 ( .A(u2__abc_44228_n12732), .B(u2__abc_44228_n12734), .Y(u2__abc_44228_n12735) );
  OR2X2 OR2X2_2777 ( .A(u2__abc_44228_n12739), .B(u2__abc_44228_n12725), .Y(u2__abc_44228_n12740) );
  OR2X2 OR2X2_2778 ( .A(u2__abc_44228_n12743), .B(u2__abc_44228_n6653_1), .Y(u2__abc_44228_n12744_1) );
  OR2X2 OR2X2_2779 ( .A(u2__abc_44228_n12744_1), .B(u2__abc_44228_n6159_1), .Y(u2__abc_44228_n12745) );
  OR2X2 OR2X2_278 ( .A(a_112_bF_buf1), .B(\a[26] ), .Y(_abc_64468_n1248) );
  OR2X2 OR2X2_2780 ( .A(u2__abc_44228_n7548_1_bF_buf43), .B(u2__abc_44228_n12748), .Y(u2__abc_44228_n12749) );
  OR2X2 OR2X2_2781 ( .A(u2__abc_44228_n7547_bF_buf42), .B(u2_remHi_302_), .Y(u2__abc_44228_n12750) );
  OR2X2 OR2X2_2782 ( .A(u2__abc_44228_n12751), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n12752_1) );
  OR2X2 OR2X2_2783 ( .A(u2__abc_44228_n12756), .B(u2__abc_44228_n12742), .Y(u2__abc_44228_n12757) );
  OR2X2 OR2X2_2784 ( .A(u2__abc_44228_n12760), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n12761) );
  OR2X2 OR2X2_2785 ( .A(u2__abc_44228_n12763), .B(u2__abc_44228_n12762), .Y(u2__abc_44228_n12764) );
  OR2X2 OR2X2_2786 ( .A(u2__abc_44228_n12765), .B(u2__abc_44228_n6166), .Y(u2__abc_44228_n12766) );
  OR2X2 OR2X2_2787 ( .A(u2__abc_44228_n12768), .B(u2__abc_44228_n12761), .Y(u2__abc_44228_n12769_1) );
  OR2X2 OR2X2_2788 ( .A(u2__abc_44228_n12773), .B(u2__abc_44228_n12759_1), .Y(u2__abc_44228_n12774) );
  OR2X2 OR2X2_2789 ( .A(u2__abc_44228_n12777), .B(u2__abc_44228_n6658), .Y(u2__abc_44228_n12778) );
  OR2X2 OR2X2_279 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[27] ), .Y(_abc_64468_n1249) );
  OR2X2 OR2X2_2790 ( .A(u2__abc_44228_n12778), .B(u2__abc_44228_n6152), .Y(u2__abc_44228_n12781) );
  OR2X2 OR2X2_2791 ( .A(u2__abc_44228_n12784_1), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n12785) );
  OR2X2 OR2X2_2792 ( .A(u2__abc_44228_n12783), .B(u2__abc_44228_n12785), .Y(u2__abc_44228_n12786) );
  OR2X2 OR2X2_2793 ( .A(u2__abc_44228_n12790), .B(u2__abc_44228_n12776_1), .Y(u2__abc_44228_n12791_1) );
  OR2X2 OR2X2_2794 ( .A(u2__abc_44228_n12779), .B(u2__abc_44228_n6148), .Y(u2__abc_44228_n12795) );
  OR2X2 OR2X2_2795 ( .A(u2__abc_44228_n12796), .B(u2__abc_44228_n12794), .Y(u2__abc_44228_n12797) );
  OR2X2 OR2X2_2796 ( .A(u2__abc_44228_n12795), .B(u2__abc_44228_n6146), .Y(u2__abc_44228_n12798) );
  OR2X2 OR2X2_2797 ( .A(u2__abc_44228_n12801), .B(u2__abc_44228_n2983_bF_buf1), .Y(u2__abc_44228_n12802) );
  OR2X2 OR2X2_2798 ( .A(u2__abc_44228_n12800_1), .B(u2__abc_44228_n12802), .Y(u2__abc_44228_n12803) );
  OR2X2 OR2X2_2799 ( .A(u2__abc_44228_n12807_1), .B(u2__abc_44228_n12793), .Y(u2__abc_44228_n12808) );
  OR2X2 OR2X2_28 ( .A(_abc_64468_n753_bF_buf8), .B(\a[13] ), .Y(_abc_64468_n870) );
  OR2X2 OR2X2_280 ( .A(a_112_bF_buf0), .B(\a[27] ), .Y(_abc_64468_n1251) );
  OR2X2 OR2X2_2800 ( .A(u2__abc_44228_n12811), .B(u2__abc_44228_n6662), .Y(u2__abc_44228_n12812) );
  OR2X2 OR2X2_2801 ( .A(u2__abc_44228_n12812), .B(u2__abc_44228_n6130), .Y(u2__abc_44228_n12813) );
  OR2X2 OR2X2_2802 ( .A(u2__abc_44228_n12818), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n12819) );
  OR2X2 OR2X2_2803 ( .A(u2__abc_44228_n12817), .B(u2__abc_44228_n12819), .Y(u2__abc_44228_n12820) );
  OR2X2 OR2X2_2804 ( .A(u2__abc_44228_n12824), .B(u2__abc_44228_n12810), .Y(u2__abc_44228_n12825) );
  OR2X2 OR2X2_2805 ( .A(u2__abc_44228_n12828), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n12829) );
  OR2X2 OR2X2_2806 ( .A(u2__abc_44228_n12831), .B(u2__abc_44228_n12830), .Y(u2__abc_44228_n12832) );
  OR2X2 OR2X2_2807 ( .A(u2__abc_44228_n12833_1), .B(u2__abc_44228_n6137), .Y(u2__abc_44228_n12834) );
  OR2X2 OR2X2_2808 ( .A(u2__abc_44228_n12836), .B(u2__abc_44228_n12829), .Y(u2__abc_44228_n12837) );
  OR2X2 OR2X2_2809 ( .A(u2__abc_44228_n12841), .B(u2__abc_44228_n12827), .Y(u2__abc_44228_n12842) );
  OR2X2 OR2X2_281 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[28] ), .Y(_abc_64468_n1252) );
  OR2X2 OR2X2_2810 ( .A(u2__abc_44228_n12845), .B(u2__abc_44228_n6667), .Y(u2__abc_44228_n12846) );
  OR2X2 OR2X2_2811 ( .A(u2__abc_44228_n12846), .B(u2__abc_44228_n6123), .Y(u2__abc_44228_n12849) );
  OR2X2 OR2X2_2812 ( .A(u2__abc_44228_n12852), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n12853) );
  OR2X2 OR2X2_2813 ( .A(u2__abc_44228_n12851), .B(u2__abc_44228_n12853), .Y(u2__abc_44228_n12854) );
  OR2X2 OR2X2_2814 ( .A(u2__abc_44228_n12858), .B(u2__abc_44228_n12844), .Y(u2__abc_44228_n12859) );
  OR2X2 OR2X2_2815 ( .A(u2__abc_44228_n12847), .B(u2__abc_44228_n6119), .Y(u2__abc_44228_n12863) );
  OR2X2 OR2X2_2816 ( .A(u2__abc_44228_n12864_1), .B(u2__abc_44228_n12862), .Y(u2__abc_44228_n12865) );
  OR2X2 OR2X2_2817 ( .A(u2__abc_44228_n12863), .B(u2__abc_44228_n6117), .Y(u2__abc_44228_n12866) );
  OR2X2 OR2X2_2818 ( .A(u2__abc_44228_n12869), .B(u2__abc_44228_n2983_bF_buf138), .Y(u2__abc_44228_n12870) );
  OR2X2 OR2X2_2819 ( .A(u2__abc_44228_n12868), .B(u2__abc_44228_n12870), .Y(u2__abc_44228_n12871_1) );
  OR2X2 OR2X2_282 ( .A(a_112_bF_buf9), .B(\a[28] ), .Y(_abc_64468_n1254) );
  OR2X2 OR2X2_2820 ( .A(u2__abc_44228_n12875), .B(u2__abc_44228_n12861), .Y(u2__abc_44228_n12876) );
  OR2X2 OR2X2_2821 ( .A(u2__abc_44228_n12879_1), .B(u2__abc_44228_n6672), .Y(u2__abc_44228_n12880) );
  OR2X2 OR2X2_2822 ( .A(u2__abc_44228_n12880), .B(u2__abc_44228_n6107), .Y(u2__abc_44228_n12883) );
  OR2X2 OR2X2_2823 ( .A(u2__abc_44228_n12886_1), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n12887) );
  OR2X2 OR2X2_2824 ( .A(u2__abc_44228_n12885), .B(u2__abc_44228_n12887), .Y(u2__abc_44228_n12888) );
  OR2X2 OR2X2_2825 ( .A(u2__abc_44228_n12892), .B(u2__abc_44228_n12878), .Y(u2__abc_44228_n12893) );
  OR2X2 OR2X2_2826 ( .A(u2__abc_44228_n12896_1), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n12897) );
  OR2X2 OR2X2_2827 ( .A(u2__abc_44228_n12899), .B(u2__abc_44228_n12898), .Y(u2__abc_44228_n12900) );
  OR2X2 OR2X2_2828 ( .A(u2__abc_44228_n12901), .B(u2__abc_44228_n6101), .Y(u2__abc_44228_n12902) );
  OR2X2 OR2X2_2829 ( .A(u2__abc_44228_n12904), .B(u2__abc_44228_n12897), .Y(u2__abc_44228_n12905) );
  OR2X2 OR2X2_283 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[29] ), .Y(_abc_64468_n1255) );
  OR2X2 OR2X2_2830 ( .A(u2__abc_44228_n12909), .B(u2__abc_44228_n12895), .Y(u2__abc_44228_n12910) );
  OR2X2 OR2X2_2831 ( .A(u2__abc_44228_n12913), .B(u2__abc_44228_n6677), .Y(u2__abc_44228_n12914) );
  OR2X2 OR2X2_2832 ( .A(u2__abc_44228_n12914), .B(u2__abc_44228_n6093), .Y(u2__abc_44228_n12917) );
  OR2X2 OR2X2_2833 ( .A(u2__abc_44228_n12920), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n12921) );
  OR2X2 OR2X2_2834 ( .A(u2__abc_44228_n12919), .B(u2__abc_44228_n12921), .Y(u2__abc_44228_n12922) );
  OR2X2 OR2X2_2835 ( .A(u2__abc_44228_n12926), .B(u2__abc_44228_n12912), .Y(u2__abc_44228_n12927_1) );
  OR2X2 OR2X2_2836 ( .A(u2__abc_44228_n12931), .B(u2__abc_44228_n12930), .Y(u2__abc_44228_n12932) );
  OR2X2 OR2X2_2837 ( .A(u2__abc_44228_n12933), .B(u2__abc_44228_n6087), .Y(u2__abc_44228_n12934_1) );
  OR2X2 OR2X2_2838 ( .A(u2__abc_44228_n12937), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n12938) );
  OR2X2 OR2X2_2839 ( .A(u2__abc_44228_n12936), .B(u2__abc_44228_n12938), .Y(u2__abc_44228_n12939) );
  OR2X2 OR2X2_284 ( .A(a_112_bF_buf8), .B(\a[29] ), .Y(_abc_64468_n1257) );
  OR2X2 OR2X2_2840 ( .A(u2__abc_44228_n12943), .B(u2__abc_44228_n12929), .Y(u2__abc_44228_n12944) );
  OR2X2 OR2X2_2841 ( .A(u2__abc_44228_n12947), .B(u2__abc_44228_n6085), .Y(u2__abc_44228_n12948) );
  OR2X2 OR2X2_2842 ( .A(u2__abc_44228_n12949_1), .B(u2__abc_44228_n6078_1), .Y(u2__abc_44228_n12952) );
  OR2X2 OR2X2_2843 ( .A(u2__abc_44228_n12955), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n12956) );
  OR2X2 OR2X2_2844 ( .A(u2__abc_44228_n12954), .B(u2__abc_44228_n12956), .Y(u2__abc_44228_n12957) );
  OR2X2 OR2X2_2845 ( .A(u2__abc_44228_n12961_1), .B(u2__abc_44228_n12946), .Y(u2__abc_44228_n12962) );
  OR2X2 OR2X2_2846 ( .A(u2__abc_44228_n12966), .B(u2__abc_44228_n12965), .Y(u2__abc_44228_n12967) );
  OR2X2 OR2X2_2847 ( .A(u2__abc_44228_n12968_1), .B(u2__abc_44228_n6072), .Y(u2__abc_44228_n12969) );
  OR2X2 OR2X2_2848 ( .A(u2__abc_44228_n12972), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n12973) );
  OR2X2 OR2X2_2849 ( .A(u2__abc_44228_n12971), .B(u2__abc_44228_n12973), .Y(u2__abc_44228_n12974) );
  OR2X2 OR2X2_285 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[30] ), .Y(_abc_64468_n1258) );
  OR2X2 OR2X2_2850 ( .A(u2__abc_44228_n12978), .B(u2__abc_44228_n12964), .Y(u2__abc_44228_n12979) );
  OR2X2 OR2X2_2851 ( .A(u2__abc_44228_n12982), .B(u2__abc_44228_n6690), .Y(u2__abc_44228_n12983_1) );
  OR2X2 OR2X2_2852 ( .A(u2__abc_44228_n12983_1), .B(u2__abc_44228_n6064), .Y(u2__abc_44228_n12986) );
  OR2X2 OR2X2_2853 ( .A(u2__abc_44228_n12989), .B(u2__abc_44228_n2983_bF_buf127), .Y(u2__abc_44228_n12990) );
  OR2X2 OR2X2_2854 ( .A(u2__abc_44228_n12988), .B(u2__abc_44228_n12990), .Y(u2__abc_44228_n12991) );
  OR2X2 OR2X2_2855 ( .A(u2__abc_44228_n12995), .B(u2__abc_44228_n12981), .Y(u2__abc_44228_n12996) );
  OR2X2 OR2X2_2856 ( .A(u2__abc_44228_n12984), .B(u2__abc_44228_n6060), .Y(u2__abc_44228_n13000) );
  OR2X2 OR2X2_2857 ( .A(u2__abc_44228_n13001), .B(u2__abc_44228_n12999_1), .Y(u2__abc_44228_n13002) );
  OR2X2 OR2X2_2858 ( .A(u2__abc_44228_n13000), .B(u2__abc_44228_n6058), .Y(u2__abc_44228_n13003) );
  OR2X2 OR2X2_2859 ( .A(u2__abc_44228_n13006), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n13007_1) );
  OR2X2 OR2X2_286 ( .A(a_112_bF_buf7), .B(\a[30] ), .Y(_abc_64468_n1260) );
  OR2X2 OR2X2_2860 ( .A(u2__abc_44228_n13005), .B(u2__abc_44228_n13007_1), .Y(u2__abc_44228_n13008) );
  OR2X2 OR2X2_2861 ( .A(u2__abc_44228_n13012), .B(u2__abc_44228_n12998), .Y(u2__abc_44228_n13013) );
  OR2X2 OR2X2_2862 ( .A(u2__abc_44228_n13016), .B(u2__abc_44228_n6696), .Y(u2__abc_44228_n13017) );
  OR2X2 OR2X2_2863 ( .A(u2__abc_44228_n13017), .B(u2__abc_44228_n6038), .Y(u2__abc_44228_n13020) );
  OR2X2 OR2X2_2864 ( .A(u2__abc_44228_n7548_1_bF_buf27), .B(u2__abc_44228_n13021), .Y(u2__abc_44228_n13022) );
  OR2X2 OR2X2_2865 ( .A(u2__abc_44228_n7547_bF_buf26), .B(u2_remHi_318_), .Y(u2__abc_44228_n13023) );
  OR2X2 OR2X2_2866 ( .A(u2__abc_44228_n13024_1), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n13025) );
  OR2X2 OR2X2_2867 ( .A(u2__abc_44228_n13029), .B(u2__abc_44228_n13015), .Y(u2__abc_44228_n13030) );
  OR2X2 OR2X2_2868 ( .A(u2__abc_44228_n13037), .B(u2__abc_44228_n13034), .Y(u2__abc_44228_n13038) );
  OR2X2 OR2X2_2869 ( .A(u2__abc_44228_n13040), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n13041) );
  OR2X2 OR2X2_287 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[31] ), .Y(_abc_64468_n1261) );
  OR2X2 OR2X2_2870 ( .A(u2__abc_44228_n13041), .B(u2__abc_44228_n13039_1), .Y(u2__abc_44228_n13042) );
  OR2X2 OR2X2_2871 ( .A(u2__abc_44228_n13046_1), .B(u2__abc_44228_n13032), .Y(u2__abc_44228_n13047) );
  OR2X2 OR2X2_2872 ( .A(u2__abc_44228_n13050), .B(u2__abc_44228_n6043), .Y(u2__abc_44228_n13051) );
  OR2X2 OR2X2_2873 ( .A(u2__abc_44228_n13052), .B(u2__abc_44228_n6031_1), .Y(u2__abc_44228_n13055_1) );
  OR2X2 OR2X2_2874 ( .A(u2__abc_44228_n13058), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n13059) );
  OR2X2 OR2X2_2875 ( .A(u2__abc_44228_n13057), .B(u2__abc_44228_n13059), .Y(u2__abc_44228_n13060) );
  OR2X2 OR2X2_2876 ( .A(u2__abc_44228_n13064), .B(u2__abc_44228_n13049), .Y(u2__abc_44228_n13065) );
  OR2X2 OR2X2_2877 ( .A(u2__abc_44228_n13053), .B(u2__abc_44228_n6027), .Y(u2__abc_44228_n13069) );
  OR2X2 OR2X2_2878 ( .A(u2__abc_44228_n13070_1), .B(u2__abc_44228_n13068), .Y(u2__abc_44228_n13071) );
  OR2X2 OR2X2_2879 ( .A(u2__abc_44228_n13069), .B(u2__abc_44228_n6025), .Y(u2__abc_44228_n13072) );
  OR2X2 OR2X2_288 ( .A(a_112_bF_buf6), .B(\a[31] ), .Y(_abc_64468_n1263) );
  OR2X2 OR2X2_2880 ( .A(u2__abc_44228_n13075), .B(u2__abc_44228_n2983_bF_buf118), .Y(u2__abc_44228_n13076) );
  OR2X2 OR2X2_2881 ( .A(u2__abc_44228_n13074), .B(u2__abc_44228_n13076), .Y(u2__abc_44228_n13077_1) );
  OR2X2 OR2X2_2882 ( .A(u2__abc_44228_n13081), .B(u2__abc_44228_n13067), .Y(u2__abc_44228_n13082) );
  OR2X2 OR2X2_2883 ( .A(u2__abc_44228_n13085), .B(u2__abc_44228_n6705), .Y(u2__abc_44228_n13086) );
  OR2X2 OR2X2_2884 ( .A(u2__abc_44228_n13086), .B(u2__abc_44228_n6009), .Y(u2__abc_44228_n13087) );
  OR2X2 OR2X2_2885 ( .A(u2__abc_44228_n7548_1_bF_buf23), .B(u2__abc_44228_n13090), .Y(u2__abc_44228_n13091) );
  OR2X2 OR2X2_2886 ( .A(u2__abc_44228_n7547_bF_buf22), .B(u2_remHi_322_), .Y(u2__abc_44228_n13092) );
  OR2X2 OR2X2_2887 ( .A(u2__abc_44228_n13093), .B(u2__abc_44228_n2983_bF_buf116), .Y(u2__abc_44228_n13094) );
  OR2X2 OR2X2_2888 ( .A(u2__abc_44228_n13098), .B(u2__abc_44228_n13084), .Y(u2__abc_44228_n13099) );
  OR2X2 OR2X2_2889 ( .A(u2__abc_44228_n13103_1), .B(u2__abc_44228_n6016), .Y(u2__abc_44228_n13104) );
  OR2X2 OR2X2_289 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[32] ), .Y(_abc_64468_n1264) );
  OR2X2 OR2X2_2890 ( .A(u2__abc_44228_n13102), .B(u2__abc_44228_n13105), .Y(u2__abc_44228_n13106) );
  OR2X2 OR2X2_2891 ( .A(u2__abc_44228_n13109), .B(u2__abc_44228_n2983_bF_buf114), .Y(u2__abc_44228_n13110_1) );
  OR2X2 OR2X2_2892 ( .A(u2__abc_44228_n13108), .B(u2__abc_44228_n13110_1), .Y(u2__abc_44228_n13111) );
  OR2X2 OR2X2_2893 ( .A(u2__abc_44228_n13115), .B(u2__abc_44228_n13101), .Y(u2__abc_44228_n13116) );
  OR2X2 OR2X2_2894 ( .A(u2__abc_44228_n13119_1), .B(u2__abc_44228_n6014), .Y(u2__abc_44228_n13120) );
  OR2X2 OR2X2_2895 ( .A(u2__abc_44228_n13121), .B(u2__abc_44228_n6002), .Y(u2__abc_44228_n13124) );
  OR2X2 OR2X2_2896 ( .A(u2__abc_44228_n13127), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n13128) );
  OR2X2 OR2X2_2897 ( .A(u2__abc_44228_n13126_1), .B(u2__abc_44228_n13128), .Y(u2__abc_44228_n13129) );
  OR2X2 OR2X2_2898 ( .A(u2__abc_44228_n13133), .B(u2__abc_44228_n13118), .Y(u2__abc_44228_n13134_1) );
  OR2X2 OR2X2_2899 ( .A(u2__abc_44228_n13122), .B(u2__abc_44228_n5998), .Y(u2__abc_44228_n13138) );
  OR2X2 OR2X2_29 ( .A(aNan_bF_buf6), .B(sqrto_90_), .Y(_abc_64468_n872) );
  OR2X2 OR2X2_290 ( .A(a_112_bF_buf5), .B(\a[32] ), .Y(_abc_64468_n1266) );
  OR2X2 OR2X2_2900 ( .A(u2__abc_44228_n13139), .B(u2__abc_44228_n13137), .Y(u2__abc_44228_n13140) );
  OR2X2 OR2X2_2901 ( .A(u2__abc_44228_n13138), .B(u2__abc_44228_n5996), .Y(u2__abc_44228_n13141_1) );
  OR2X2 OR2X2_2902 ( .A(u2__abc_44228_n13144), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n13145) );
  OR2X2 OR2X2_2903 ( .A(u2__abc_44228_n13143), .B(u2__abc_44228_n13145), .Y(u2__abc_44228_n13146) );
  OR2X2 OR2X2_2904 ( .A(u2__abc_44228_n13150), .B(u2__abc_44228_n13136), .Y(u2__abc_44228_n13151_1) );
  OR2X2 OR2X2_2905 ( .A(u2__abc_44228_n13154), .B(u2__abc_44228_n6715), .Y(u2__abc_44228_n13155) );
  OR2X2 OR2X2_2906 ( .A(u2__abc_44228_n13155), .B(u2__abc_44228_n5986), .Y(u2__abc_44228_n13158_1) );
  OR2X2 OR2X2_2907 ( .A(u2__abc_44228_n7548_1_bF_buf19), .B(u2__abc_44228_n13159), .Y(u2__abc_44228_n13160) );
  OR2X2 OR2X2_2908 ( .A(u2__abc_44228_n7547_bF_buf18), .B(u2_remHi_326_), .Y(u2__abc_44228_n13161) );
  OR2X2 OR2X2_2909 ( .A(u2__abc_44228_n13162), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n13163) );
  OR2X2 OR2X2_291 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[33] ), .Y(_abc_64468_n1267) );
  OR2X2 OR2X2_2910 ( .A(u2__abc_44228_n13167), .B(u2__abc_44228_n13153), .Y(u2__abc_44228_n13168) );
  OR2X2 OR2X2_2911 ( .A(u2__abc_44228_n13175), .B(u2__abc_44228_n13172), .Y(u2__abc_44228_n13176) );
  OR2X2 OR2X2_2912 ( .A(u2__abc_44228_n13178), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n13179) );
  OR2X2 OR2X2_2913 ( .A(u2__abc_44228_n13177), .B(u2__abc_44228_n13179), .Y(u2__abc_44228_n13180) );
  OR2X2 OR2X2_2914 ( .A(u2__abc_44228_n13184), .B(u2__abc_44228_n13170), .Y(u2__abc_44228_n13185) );
  OR2X2 OR2X2_2915 ( .A(u2__abc_44228_n13188), .B(u2__abc_44228_n5978), .Y(u2__abc_44228_n13189_1) );
  OR2X2 OR2X2_2916 ( .A(u2__abc_44228_n13190), .B(u2__abc_44228_n5972), .Y(u2__abc_44228_n13193) );
  OR2X2 OR2X2_2917 ( .A(u2__abc_44228_n13196), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n13197_1) );
  OR2X2 OR2X2_2918 ( .A(u2__abc_44228_n13195), .B(u2__abc_44228_n13197_1), .Y(u2__abc_44228_n13198) );
  OR2X2 OR2X2_2919 ( .A(u2__abc_44228_n13202), .B(u2__abc_44228_n13187), .Y(u2__abc_44228_n13203) );
  OR2X2 OR2X2_292 ( .A(a_112_bF_buf4), .B(\a[33] ), .Y(_abc_64468_n1269) );
  OR2X2 OR2X2_2920 ( .A(u2__abc_44228_n13191), .B(u2__abc_44228_n5968), .Y(u2__abc_44228_n13207) );
  OR2X2 OR2X2_2921 ( .A(u2__abc_44228_n13208), .B(u2__abc_44228_n13206), .Y(u2__abc_44228_n13209) );
  OR2X2 OR2X2_2922 ( .A(u2__abc_44228_n13207), .B(u2__abc_44228_n5966_1), .Y(u2__abc_44228_n13210) );
  OR2X2 OR2X2_2923 ( .A(u2__abc_44228_n13213), .B(u2__abc_44228_n2983_bF_buf104), .Y(u2__abc_44228_n13214) );
  OR2X2 OR2X2_2924 ( .A(u2__abc_44228_n13212), .B(u2__abc_44228_n13214), .Y(u2__abc_44228_n13215) );
  OR2X2 OR2X2_2925 ( .A(u2__abc_44228_n13219), .B(u2__abc_44228_n13205), .Y(u2__abc_44228_n13220) );
  OR2X2 OR2X2_2926 ( .A(u2__abc_44228_n13223), .B(u2__abc_44228_n6724), .Y(u2__abc_44228_n13224_1) );
  OR2X2 OR2X2_2927 ( .A(u2__abc_44228_n13224_1), .B(u2__abc_44228_n5957_1), .Y(u2__abc_44228_n13225) );
  OR2X2 OR2X2_2928 ( .A(u2__abc_44228_n13230), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n13231) );
  OR2X2 OR2X2_2929 ( .A(u2__abc_44228_n13229), .B(u2__abc_44228_n13231), .Y(u2__abc_44228_n13232_1) );
  OR2X2 OR2X2_293 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[34] ), .Y(_abc_64468_n1270) );
  OR2X2 OR2X2_2930 ( .A(u2__abc_44228_n13236), .B(u2__abc_44228_n13222), .Y(u2__abc_44228_n13237) );
  OR2X2 OR2X2_2931 ( .A(u2__abc_44228_n13244), .B(u2__abc_44228_n13241), .Y(u2__abc_44228_n13245) );
  OR2X2 OR2X2_2932 ( .A(u2__abc_44228_n13247), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n13248_1) );
  OR2X2 OR2X2_2933 ( .A(u2__abc_44228_n13246), .B(u2__abc_44228_n13248_1), .Y(u2__abc_44228_n13249) );
  OR2X2 OR2X2_2934 ( .A(u2__abc_44228_n13253), .B(u2__abc_44228_n13239_1), .Y(u2__abc_44228_n13254) );
  OR2X2 OR2X2_2935 ( .A(u2__abc_44228_n13257), .B(u2__abc_44228_n5949), .Y(u2__abc_44228_n13258) );
  OR2X2 OR2X2_2936 ( .A(u2__abc_44228_n13259), .B(u2__abc_44228_n5943), .Y(u2__abc_44228_n13262) );
  OR2X2 OR2X2_2937 ( .A(u2__abc_44228_n13265), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n13266) );
  OR2X2 OR2X2_2938 ( .A(u2__abc_44228_n13264), .B(u2__abc_44228_n13266), .Y(u2__abc_44228_n13267) );
  OR2X2 OR2X2_2939 ( .A(u2__abc_44228_n13271), .B(u2__abc_44228_n13256), .Y(u2__abc_44228_n13272) );
  OR2X2 OR2X2_294 ( .A(a_112_bF_buf3), .B(\a[34] ), .Y(_abc_64468_n1272) );
  OR2X2 OR2X2_2940 ( .A(u2__abc_44228_n13260), .B(u2__abc_44228_n5939), .Y(u2__abc_44228_n13276) );
  OR2X2 OR2X2_2941 ( .A(u2__abc_44228_n13277), .B(u2__abc_44228_n13275), .Y(u2__abc_44228_n13278) );
  OR2X2 OR2X2_2942 ( .A(u2__abc_44228_n13276), .B(u2__abc_44228_n5937), .Y(u2__abc_44228_n13279) );
  OR2X2 OR2X2_2943 ( .A(u2__abc_44228_n13282), .B(u2__abc_44228_n2983_bF_buf98), .Y(u2__abc_44228_n13283) );
  OR2X2 OR2X2_2944 ( .A(u2__abc_44228_n13281), .B(u2__abc_44228_n13283), .Y(u2__abc_44228_n13284) );
  OR2X2 OR2X2_2945 ( .A(u2__abc_44228_n13288), .B(u2__abc_44228_n13274), .Y(u2__abc_44228_n13289) );
  OR2X2 OR2X2_2946 ( .A(u2__abc_44228_n13292), .B(u2__abc_44228_n6735_1), .Y(u2__abc_44228_n13293) );
  OR2X2 OR2X2_2947 ( .A(u2__abc_44228_n13293), .B(u2__abc_44228_n5926), .Y(u2__abc_44228_n13294) );
  OR2X2 OR2X2_2948 ( .A(u2__abc_44228_n7548_1_bF_buf11), .B(u2__abc_44228_n13297), .Y(u2__abc_44228_n13298) );
  OR2X2 OR2X2_2949 ( .A(u2__abc_44228_n7547_bF_buf10), .B(u2_remHi_334_), .Y(u2__abc_44228_n13299) );
  OR2X2 OR2X2_295 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[35] ), .Y(_abc_64468_n1273) );
  OR2X2 OR2X2_2950 ( .A(u2__abc_44228_n13300), .B(u2__abc_44228_n2983_bF_buf96), .Y(u2__abc_44228_n13301) );
  OR2X2 OR2X2_2951 ( .A(u2__abc_44228_n13305), .B(u2__abc_44228_n13291), .Y(u2__abc_44228_n13306) );
  OR2X2 OR2X2_2952 ( .A(u2__abc_44228_n13310), .B(u2__abc_44228_n13309), .Y(u2__abc_44228_n13311_1) );
  OR2X2 OR2X2_2953 ( .A(u2__abc_44228_n13312), .B(u2__abc_44228_n5920_1), .Y(u2__abc_44228_n13313) );
  OR2X2 OR2X2_2954 ( .A(u2__abc_44228_n13316), .B(u2__abc_44228_n2983_bF_buf94), .Y(u2__abc_44228_n13317) );
  OR2X2 OR2X2_2955 ( .A(u2__abc_44228_n13315), .B(u2__abc_44228_n13317), .Y(u2__abc_44228_n13318_1) );
  OR2X2 OR2X2_2956 ( .A(u2__abc_44228_n13322), .B(u2__abc_44228_n13308), .Y(u2__abc_44228_n13323) );
  OR2X2 OR2X2_2957 ( .A(u2__abc_44228_n13326_1), .B(u2__abc_44228_n6740), .Y(u2__abc_44228_n13327) );
  OR2X2 OR2X2_2958 ( .A(u2__abc_44228_n13327), .B(u2__abc_44228_n5912), .Y(u2__abc_44228_n13330) );
  OR2X2 OR2X2_2959 ( .A(u2__abc_44228_n13333_1), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n13334) );
  OR2X2 OR2X2_296 ( .A(a_112_bF_buf2), .B(\a[35] ), .Y(_abc_64468_n1275) );
  OR2X2 OR2X2_2960 ( .A(u2__abc_44228_n13332), .B(u2__abc_44228_n13334), .Y(u2__abc_44228_n13335) );
  OR2X2 OR2X2_2961 ( .A(u2__abc_44228_n13339), .B(u2__abc_44228_n13325), .Y(u2__abc_44228_n13340) );
  OR2X2 OR2X2_2962 ( .A(u2__abc_44228_n13328), .B(u2__abc_44228_n5908), .Y(u2__abc_44228_n13344_1) );
  OR2X2 OR2X2_2963 ( .A(u2__abc_44228_n13345), .B(u2__abc_44228_n13343), .Y(u2__abc_44228_n13346) );
  OR2X2 OR2X2_2964 ( .A(u2__abc_44228_n13344_1), .B(u2__abc_44228_n5906), .Y(u2__abc_44228_n13347) );
  OR2X2 OR2X2_2965 ( .A(u2__abc_44228_n13350), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n13351_1) );
  OR2X2 OR2X2_2966 ( .A(u2__abc_44228_n13349), .B(u2__abc_44228_n13351_1), .Y(u2__abc_44228_n13352) );
  OR2X2 OR2X2_2967 ( .A(u2__abc_44228_n13356), .B(u2__abc_44228_n13342), .Y(u2__abc_44228_n13357) );
  OR2X2 OR2X2_2968 ( .A(u2__abc_44228_n13360), .B(u2__abc_44228_n6744), .Y(u2__abc_44228_n13361) );
  OR2X2 OR2X2_2969 ( .A(u2__abc_44228_n13361), .B(u2__abc_44228_n5890), .Y(u2__abc_44228_n13362) );
  OR2X2 OR2X2_297 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[36] ), .Y(_abc_64468_n1276) );
  OR2X2 OR2X2_2970 ( .A(u2__abc_44228_n13367), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n13368) );
  OR2X2 OR2X2_2971 ( .A(u2__abc_44228_n13366_1), .B(u2__abc_44228_n13368), .Y(u2__abc_44228_n13369) );
  OR2X2 OR2X2_2972 ( .A(u2__abc_44228_n13373), .B(u2__abc_44228_n13359_1), .Y(u2__abc_44228_n13374) );
  OR2X2 OR2X2_2973 ( .A(u2__abc_44228_n13381), .B(u2__abc_44228_n13378), .Y(u2__abc_44228_n13382_1) );
  OR2X2 OR2X2_2974 ( .A(u2__abc_44228_n13384), .B(u2__abc_44228_n2983_bF_buf88), .Y(u2__abc_44228_n13385) );
  OR2X2 OR2X2_2975 ( .A(u2__abc_44228_n13383), .B(u2__abc_44228_n13385), .Y(u2__abc_44228_n13386) );
  OR2X2 OR2X2_2976 ( .A(u2__abc_44228_n13390_1), .B(u2__abc_44228_n13376), .Y(u2__abc_44228_n13391) );
  OR2X2 OR2X2_2977 ( .A(u2__abc_44228_n13394), .B(u2__abc_44228_n5895), .Y(u2__abc_44228_n13395) );
  OR2X2 OR2X2_2978 ( .A(u2__abc_44228_n13396), .B(u2__abc_44228_n5883_1), .Y(u2__abc_44228_n13399) );
  OR2X2 OR2X2_2979 ( .A(u2__abc_44228_n13402), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n13403) );
  OR2X2 OR2X2_298 ( .A(a_112_bF_buf1), .B(\a[36] ), .Y(_abc_64468_n1278) );
  OR2X2 OR2X2_2980 ( .A(u2__abc_44228_n13401), .B(u2__abc_44228_n13403), .Y(u2__abc_44228_n13404) );
  OR2X2 OR2X2_2981 ( .A(u2__abc_44228_n13408), .B(u2__abc_44228_n13393), .Y(u2__abc_44228_n13409) );
  OR2X2 OR2X2_2982 ( .A(u2__abc_44228_n13397_1), .B(u2__abc_44228_n5879), .Y(u2__abc_44228_n13413) );
  OR2X2 OR2X2_2983 ( .A(u2__abc_44228_n13414_1), .B(u2__abc_44228_n13412), .Y(u2__abc_44228_n13415) );
  OR2X2 OR2X2_2984 ( .A(u2__abc_44228_n13413), .B(u2__abc_44228_n5877), .Y(u2__abc_44228_n13416) );
  OR2X2 OR2X2_2985 ( .A(u2__abc_44228_n13419), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n13420) );
  OR2X2 OR2X2_2986 ( .A(u2__abc_44228_n13418), .B(u2__abc_44228_n13420), .Y(u2__abc_44228_n13421) );
  OR2X2 OR2X2_2987 ( .A(u2__abc_44228_n13425), .B(u2__abc_44228_n13411), .Y(u2__abc_44228_n13426) );
  OR2X2 OR2X2_2988 ( .A(u2__abc_44228_n13429_1), .B(u2__abc_44228_n6754), .Y(u2__abc_44228_n13430) );
  OR2X2 OR2X2_2989 ( .A(u2__abc_44228_n13430), .B(u2__abc_44228_n5853), .Y(u2__abc_44228_n13433) );
  OR2X2 OR2X2_299 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[37] ), .Y(_abc_64468_n1279) );
  OR2X2 OR2X2_2990 ( .A(u2__abc_44228_n13436), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n13437) );
  OR2X2 OR2X2_2991 ( .A(u2__abc_44228_n13435), .B(u2__abc_44228_n13437), .Y(u2__abc_44228_n13438_1) );
  OR2X2 OR2X2_2992 ( .A(u2__abc_44228_n13442), .B(u2__abc_44228_n13428), .Y(u2__abc_44228_n13443) );
  OR2X2 OR2X2_2993 ( .A(u2__abc_44228_n13447), .B(u2__abc_44228_n13446), .Y(u2__abc_44228_n13448) );
  OR2X2 OR2X2_2994 ( .A(u2__abc_44228_n13449), .B(u2__abc_44228_n5847), .Y(u2__abc_44228_n13450) );
  OR2X2 OR2X2_2995 ( .A(u2__abc_44228_n13453_1), .B(u2__abc_44228_n2983_bF_buf82), .Y(u2__abc_44228_n13454) );
  OR2X2 OR2X2_2996 ( .A(u2__abc_44228_n13452), .B(u2__abc_44228_n13454), .Y(u2__abc_44228_n13455) );
  OR2X2 OR2X2_2997 ( .A(u2__abc_44228_n13459), .B(u2__abc_44228_n13445_1), .Y(u2__abc_44228_n13460_1) );
  OR2X2 OR2X2_2998 ( .A(u2__abc_44228_n13463), .B(u2__abc_44228_n6759), .Y(u2__abc_44228_n13464) );
  OR2X2 OR2X2_2999 ( .A(u2__abc_44228_n13464), .B(u2__abc_44228_n5867), .Y(u2__abc_44228_n13467) );
  OR2X2 OR2X2_3 ( .A(aNan_bF_buf8), .B(sqrto_77_), .Y(_abc_64468_n833) );
  OR2X2 OR2X2_30 ( .A(_abc_64468_n753_bF_buf7), .B(\a[14] ), .Y(_abc_64468_n873) );
  OR2X2 OR2X2_300 ( .A(a_112_bF_buf0), .B(\a[37] ), .Y(_abc_64468_n1281) );
  OR2X2 OR2X2_3000 ( .A(u2__abc_44228_n13470), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n13471) );
  OR2X2 OR2X2_3001 ( .A(u2__abc_44228_n13469), .B(u2__abc_44228_n13471), .Y(u2__abc_44228_n13472_1) );
  OR2X2 OR2X2_3002 ( .A(u2__abc_44228_n13476), .B(u2__abc_44228_n13462), .Y(u2__abc_44228_n13477) );
  OR2X2 OR2X2_3003 ( .A(u2__abc_44228_n13481), .B(u2__abc_44228_n13480), .Y(u2__abc_44228_n13482) );
  OR2X2 OR2X2_3004 ( .A(u2__abc_44228_n13483), .B(u2__abc_44228_n5861), .Y(u2__abc_44228_n13484) );
  OR2X2 OR2X2_3005 ( .A(u2__abc_44228_n13487_1), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n13488) );
  OR2X2 OR2X2_3006 ( .A(u2__abc_44228_n13486), .B(u2__abc_44228_n13488), .Y(u2__abc_44228_n13489) );
  OR2X2 OR2X2_3007 ( .A(u2__abc_44228_n13493), .B(u2__abc_44228_n13479_1), .Y(u2__abc_44228_n13494_1) );
  OR2X2 OR2X2_3008 ( .A(u2__abc_44228_n13497), .B(u2__abc_44228_n5859), .Y(u2__abc_44228_n13498) );
  OR2X2 OR2X2_3009 ( .A(u2__abc_44228_n13499), .B(u2__abc_44228_n5831), .Y(u2__abc_44228_n13500) );
  OR2X2 OR2X2_301 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[38] ), .Y(_abc_64468_n1282) );
  OR2X2 OR2X2_3010 ( .A(u2__abc_44228_n13505), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n13506) );
  OR2X2 OR2X2_3011 ( .A(u2__abc_44228_n13504), .B(u2__abc_44228_n13506), .Y(u2__abc_44228_n13507) );
  OR2X2 OR2X2_3012 ( .A(u2__abc_44228_n13511), .B(u2__abc_44228_n13496), .Y(u2__abc_44228_n13512) );
  OR2X2 OR2X2_3013 ( .A(u2__abc_44228_n13516), .B(u2__abc_44228_n5838_1), .Y(u2__abc_44228_n13517) );
  OR2X2 OR2X2_3014 ( .A(u2__abc_44228_n13515), .B(u2__abc_44228_n13518_1), .Y(u2__abc_44228_n13519) );
  OR2X2 OR2X2_3015 ( .A(u2__abc_44228_n13522), .B(u2__abc_44228_n2983_bF_buf76), .Y(u2__abc_44228_n13523) );
  OR2X2 OR2X2_3016 ( .A(u2__abc_44228_n13521), .B(u2__abc_44228_n13523), .Y(u2__abc_44228_n13524) );
  OR2X2 OR2X2_3017 ( .A(u2__abc_44228_n13528), .B(u2__abc_44228_n13514), .Y(u2__abc_44228_n13529) );
  OR2X2 OR2X2_3018 ( .A(u2__abc_44228_n13532), .B(u2__abc_44228_n5836), .Y(u2__abc_44228_n13533) );
  OR2X2 OR2X2_3019 ( .A(u2__abc_44228_n13534), .B(u2__abc_44228_n5824), .Y(u2__abc_44228_n13537) );
  OR2X2 OR2X2_302 ( .A(a_112_bF_buf9), .B(\a[38] ), .Y(_abc_64468_n1284) );
  OR2X2 OR2X2_3020 ( .A(u2__abc_44228_n13540), .B(u2__abc_44228_n2983_bF_buf74), .Y(u2__abc_44228_n13541) );
  OR2X2 OR2X2_3021 ( .A(u2__abc_44228_n13539), .B(u2__abc_44228_n13541), .Y(u2__abc_44228_n13542_1) );
  OR2X2 OR2X2_3022 ( .A(u2__abc_44228_n13546), .B(u2__abc_44228_n13531), .Y(u2__abc_44228_n13547) );
  OR2X2 OR2X2_3023 ( .A(u2__abc_44228_n13535_1), .B(u2__abc_44228_n5820), .Y(u2__abc_44228_n13551) );
  OR2X2 OR2X2_3024 ( .A(u2__abc_44228_n13552), .B(u2__abc_44228_n13550_1), .Y(u2__abc_44228_n13553) );
  OR2X2 OR2X2_3025 ( .A(u2__abc_44228_n13551), .B(u2__abc_44228_n5818), .Y(u2__abc_44228_n13554) );
  OR2X2 OR2X2_3026 ( .A(u2__abc_44228_n13557_1), .B(u2__abc_44228_n2983_bF_buf72), .Y(u2__abc_44228_n13558) );
  OR2X2 OR2X2_3027 ( .A(u2__abc_44228_n13556), .B(u2__abc_44228_n13558), .Y(u2__abc_44228_n13559) );
  OR2X2 OR2X2_3028 ( .A(u2__abc_44228_n13563), .B(u2__abc_44228_n13549), .Y(u2__abc_44228_n13564) );
  OR2X2 OR2X2_3029 ( .A(u2__abc_44228_n13567), .B(u2__abc_44228_n6777), .Y(u2__abc_44228_n13568) );
  OR2X2 OR2X2_303 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[39] ), .Y(_abc_64468_n1285) );
  OR2X2 OR2X2_3030 ( .A(u2__abc_44228_n13568), .B(u2__abc_44228_n5806), .Y(u2__abc_44228_n13571) );
  OR2X2 OR2X2_3031 ( .A(u2__abc_44228_n7548_1_bF_buf53), .B(u2__abc_44228_n13572), .Y(u2__abc_44228_n13573_1) );
  OR2X2 OR2X2_3032 ( .A(u2__abc_44228_n7547_bF_buf52), .B(u2_remHi_350_), .Y(u2__abc_44228_n13574) );
  OR2X2 OR2X2_3033 ( .A(u2__abc_44228_n13575), .B(u2__abc_44228_n2983_bF_buf70), .Y(u2__abc_44228_n13576) );
  OR2X2 OR2X2_3034 ( .A(u2__abc_44228_n13580), .B(u2__abc_44228_n13566_1), .Y(u2__abc_44228_n13581_1) );
  OR2X2 OR2X2_3035 ( .A(u2__abc_44228_n13585), .B(u2__abc_44228_n13584), .Y(u2__abc_44228_n13586) );
  OR2X2 OR2X2_3036 ( .A(u2__abc_44228_n13587), .B(u2__abc_44228_n5800), .Y(u2__abc_44228_n13588_1) );
  OR2X2 OR2X2_3037 ( .A(u2__abc_44228_n13591), .B(u2__abc_44228_n2983_bF_buf68), .Y(u2__abc_44228_n13592) );
  OR2X2 OR2X2_3038 ( .A(u2__abc_44228_n13590), .B(u2__abc_44228_n13592), .Y(u2__abc_44228_n13593) );
  OR2X2 OR2X2_3039 ( .A(u2__abc_44228_n13597), .B(u2__abc_44228_n13583), .Y(u2__abc_44228_n13598) );
  OR2X2 OR2X2_304 ( .A(a_112_bF_buf8), .B(\a[39] ), .Y(_abc_64468_n1287) );
  OR2X2 OR2X2_3040 ( .A(u2__abc_44228_n13601), .B(u2__abc_44228_n6782), .Y(u2__abc_44228_n13602) );
  OR2X2 OR2X2_3041 ( .A(u2__abc_44228_n13602), .B(u2__abc_44228_n5792), .Y(u2__abc_44228_n13605) );
  OR2X2 OR2X2_3042 ( .A(u2__abc_44228_n13608), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n13609) );
  OR2X2 OR2X2_3043 ( .A(u2__abc_44228_n13607), .B(u2__abc_44228_n13609), .Y(u2__abc_44228_n13610) );
  OR2X2 OR2X2_3044 ( .A(u2__abc_44228_n13614_1), .B(u2__abc_44228_n13600), .Y(u2__abc_44228_n13615) );
  OR2X2 OR2X2_3045 ( .A(u2__abc_44228_n13603), .B(u2__abc_44228_n5788), .Y(u2__abc_44228_n13619) );
  OR2X2 OR2X2_3046 ( .A(u2__abc_44228_n13620), .B(u2__abc_44228_n13618), .Y(u2__abc_44228_n13621_1) );
  OR2X2 OR2X2_3047 ( .A(u2__abc_44228_n13619), .B(u2__abc_44228_n5786), .Y(u2__abc_44228_n13622) );
  OR2X2 OR2X2_3048 ( .A(u2__abc_44228_n13625), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n13626) );
  OR2X2 OR2X2_3049 ( .A(u2__abc_44228_n13624), .B(u2__abc_44228_n13626), .Y(u2__abc_44228_n13627) );
  OR2X2 OR2X2_305 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[40] ), .Y(_abc_64468_n1288) );
  OR2X2 OR2X2_3050 ( .A(u2__abc_44228_n13631), .B(u2__abc_44228_n13617), .Y(u2__abc_44228_n13632) );
  OR2X2 OR2X2_3051 ( .A(u2__abc_44228_n13635), .B(u2__abc_44228_n6786), .Y(u2__abc_44228_n13636) );
  OR2X2 OR2X2_3052 ( .A(u2__abc_44228_n13636), .B(u2__abc_44228_n5770), .Y(u2__abc_44228_n13637_1) );
  OR2X2 OR2X2_3053 ( .A(u2__abc_44228_n13642), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n13643) );
  OR2X2 OR2X2_3054 ( .A(u2__abc_44228_n13641), .B(u2__abc_44228_n13643), .Y(u2__abc_44228_n13644) );
  OR2X2 OR2X2_3055 ( .A(u2__abc_44228_n13648), .B(u2__abc_44228_n13634), .Y(u2__abc_44228_n13649) );
  OR2X2 OR2X2_3056 ( .A(u2__abc_44228_n13656), .B(u2__abc_44228_n13653), .Y(u2__abc_44228_n13657) );
  OR2X2 OR2X2_3057 ( .A(u2__abc_44228_n13659), .B(u2__abc_44228_n2983_bF_buf62), .Y(u2__abc_44228_n13660) );
  OR2X2 OR2X2_3058 ( .A(u2__abc_44228_n13658), .B(u2__abc_44228_n13660), .Y(u2__abc_44228_n13661) );
  OR2X2 OR2X2_3059 ( .A(u2__abc_44228_n13665), .B(u2__abc_44228_n13651), .Y(u2__abc_44228_n13666) );
  OR2X2 OR2X2_306 ( .A(a_112_bF_buf7), .B(\a[40] ), .Y(_abc_64468_n1290) );
  OR2X2 OR2X2_3060 ( .A(u2__abc_44228_n13669_1), .B(u2__abc_44228_n5775), .Y(u2__abc_44228_n13670) );
  OR2X2 OR2X2_3061 ( .A(u2__abc_44228_n13671), .B(u2__abc_44228_n5763), .Y(u2__abc_44228_n13674) );
  OR2X2 OR2X2_3062 ( .A(u2__abc_44228_n13677_1), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n13678) );
  OR2X2 OR2X2_3063 ( .A(u2__abc_44228_n13676), .B(u2__abc_44228_n13678), .Y(u2__abc_44228_n13679) );
  OR2X2 OR2X2_3064 ( .A(u2__abc_44228_n13683), .B(u2__abc_44228_n13668), .Y(u2__abc_44228_n13684_1) );
  OR2X2 OR2X2_3065 ( .A(u2__abc_44228_n13672), .B(u2__abc_44228_n5759), .Y(u2__abc_44228_n13688) );
  OR2X2 OR2X2_3066 ( .A(u2__abc_44228_n13689), .B(u2__abc_44228_n13687), .Y(u2__abc_44228_n13690) );
  OR2X2 OR2X2_3067 ( .A(u2__abc_44228_n13688), .B(u2__abc_44228_n5757), .Y(u2__abc_44228_n13691) );
  OR2X2 OR2X2_3068 ( .A(u2__abc_44228_n13694), .B(u2__abc_44228_n2983_bF_buf59), .Y(u2__abc_44228_n13695) );
  OR2X2 OR2X2_3069 ( .A(u2__abc_44228_n13693_1), .B(u2__abc_44228_n13695), .Y(u2__abc_44228_n13696) );
  OR2X2 OR2X2_307 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[41] ), .Y(_abc_64468_n1291) );
  OR2X2 OR2X2_3070 ( .A(u2__abc_44228_n13700_1), .B(u2__abc_44228_n13686), .Y(u2__abc_44228_n13701) );
  OR2X2 OR2X2_3071 ( .A(u2__abc_44228_n13704), .B(u2__abc_44228_n6796), .Y(u2__abc_44228_n13705) );
  OR2X2 OR2X2_3072 ( .A(u2__abc_44228_n13705), .B(u2__abc_44228_n5733), .Y(u2__abc_44228_n13708) );
  OR2X2 OR2X2_3073 ( .A(u2__abc_44228_n13711), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n13712) );
  OR2X2 OR2X2_3074 ( .A(u2__abc_44228_n13710), .B(u2__abc_44228_n13712), .Y(u2__abc_44228_n13713) );
  OR2X2 OR2X2_3075 ( .A(u2__abc_44228_n13717_1), .B(u2__abc_44228_n13703), .Y(u2__abc_44228_n13718) );
  OR2X2 OR2X2_3076 ( .A(u2__abc_44228_n13722), .B(u2__abc_44228_n13721), .Y(u2__abc_44228_n13723) );
  OR2X2 OR2X2_3077 ( .A(u2__abc_44228_n13724), .B(u2__abc_44228_n5727), .Y(u2__abc_44228_n13725) );
  OR2X2 OR2X2_3078 ( .A(u2__abc_44228_n13728), .B(u2__abc_44228_n2983_bF_buf56), .Y(u2__abc_44228_n13729) );
  OR2X2 OR2X2_3079 ( .A(u2__abc_44228_n13727), .B(u2__abc_44228_n13729), .Y(u2__abc_44228_n13730) );
  OR2X2 OR2X2_308 ( .A(a_112_bF_buf6), .B(\a[41] ), .Y(_abc_64468_n1293) );
  OR2X2 OR2X2_3080 ( .A(u2__abc_44228_n13734), .B(u2__abc_44228_n13720), .Y(u2__abc_44228_n13735) );
  OR2X2 OR2X2_3081 ( .A(u2__abc_44228_n13738), .B(u2__abc_44228_n6801), .Y(u2__abc_44228_n13739) );
  OR2X2 OR2X2_3082 ( .A(u2__abc_44228_n13739), .B(u2__abc_44228_n5747_1), .Y(u2__abc_44228_n13742) );
  OR2X2 OR2X2_3083 ( .A(u2__abc_44228_n13745), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n13746) );
  OR2X2 OR2X2_3084 ( .A(u2__abc_44228_n13744), .B(u2__abc_44228_n13746), .Y(u2__abc_44228_n13747) );
  OR2X2 OR2X2_3085 ( .A(u2__abc_44228_n13751), .B(u2__abc_44228_n13737), .Y(u2__abc_44228_n13752) );
  OR2X2 OR2X2_3086 ( .A(u2__abc_44228_n13756), .B(u2__abc_44228_n13755), .Y(u2__abc_44228_n13757_1) );
  OR2X2 OR2X2_3087 ( .A(u2__abc_44228_n13758), .B(u2__abc_44228_n5741), .Y(u2__abc_44228_n13759) );
  OR2X2 OR2X2_3088 ( .A(u2__abc_44228_n13762), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n13763) );
  OR2X2 OR2X2_3089 ( .A(u2__abc_44228_n13761), .B(u2__abc_44228_n13763), .Y(u2__abc_44228_n13764) );
  OR2X2 OR2X2_309 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[42] ), .Y(_abc_64468_n1294) );
  OR2X2 OR2X2_3090 ( .A(u2__abc_44228_n13768), .B(u2__abc_44228_n13754), .Y(u2__abc_44228_n13769) );
  OR2X2 OR2X2_3091 ( .A(u2__abc_44228_n13772), .B(u2__abc_44228_n5739), .Y(u2__abc_44228_n13773) );
  OR2X2 OR2X2_3092 ( .A(u2__abc_44228_n13774), .B(u2__abc_44228_n5718), .Y(u2__abc_44228_n13775_1) );
  OR2X2 OR2X2_3093 ( .A(u2__abc_44228_n13780), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n13781) );
  OR2X2 OR2X2_3094 ( .A(u2__abc_44228_n13779), .B(u2__abc_44228_n13781), .Y(u2__abc_44228_n13782) );
  OR2X2 OR2X2_3095 ( .A(u2__abc_44228_n13786), .B(u2__abc_44228_n13771), .Y(u2__abc_44228_n13787) );
  OR2X2 OR2X2_3096 ( .A(u2__abc_44228_n13791), .B(u2__abc_44228_n13790), .Y(u2__abc_44228_n13792_1) );
  OR2X2 OR2X2_3097 ( .A(u2__abc_44228_n13793), .B(u2__abc_44228_n5712), .Y(u2__abc_44228_n13794) );
  OR2X2 OR2X2_3098 ( .A(u2__abc_44228_n13797), .B(u2__abc_44228_n2983_bF_buf50), .Y(u2__abc_44228_n13798) );
  OR2X2 OR2X2_3099 ( .A(u2__abc_44228_n13796), .B(u2__abc_44228_n13798), .Y(u2__abc_44228_n13799) );
  OR2X2 OR2X2_31 ( .A(aNan_bF_buf5), .B(sqrto_91_), .Y(_abc_64468_n875) );
  OR2X2 OR2X2_310 ( .A(a_112_bF_buf5), .B(\a[42] ), .Y(_abc_64468_n1296) );
  OR2X2 OR2X2_3100 ( .A(u2__abc_44228_n13803_1), .B(u2__abc_44228_n13789), .Y(u2__abc_44228_n13804) );
  OR2X2 OR2X2_3101 ( .A(u2__abc_44228_n13807), .B(u2__abc_44228_n6814), .Y(u2__abc_44228_n13808) );
  OR2X2 OR2X2_3102 ( .A(u2__abc_44228_n13808), .B(u2__abc_44228_n5704), .Y(u2__abc_44228_n13811_1) );
  OR2X2 OR2X2_3103 ( .A(u2__abc_44228_n13814), .B(u2__abc_44228_n2983_bF_buf48), .Y(u2__abc_44228_n13815) );
  OR2X2 OR2X2_3104 ( .A(u2__abc_44228_n13813), .B(u2__abc_44228_n13815), .Y(u2__abc_44228_n13816) );
  OR2X2 OR2X2_3105 ( .A(u2__abc_44228_n13820_1), .B(u2__abc_44228_n13806), .Y(u2__abc_44228_n13821) );
  OR2X2 OR2X2_3106 ( .A(u2__abc_44228_n13809), .B(u2__abc_44228_n5700_1), .Y(u2__abc_44228_n13825) );
  OR2X2 OR2X2_3107 ( .A(u2__abc_44228_n13826), .B(u2__abc_44228_n13824), .Y(u2__abc_44228_n13827) );
  OR2X2 OR2X2_3108 ( .A(u2__abc_44228_n13825), .B(u2__abc_44228_n5698), .Y(u2__abc_44228_n13828_1) );
  OR2X2 OR2X2_3109 ( .A(u2__abc_44228_n13831), .B(u2__abc_44228_n2983_bF_buf46), .Y(u2__abc_44228_n13832) );
  OR2X2 OR2X2_311 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[43] ), .Y(_abc_64468_n1297) );
  OR2X2 OR2X2_3110 ( .A(u2__abc_44228_n13830), .B(u2__abc_44228_n13832), .Y(u2__abc_44228_n13833) );
  OR2X2 OR2X2_3111 ( .A(u2__abc_44228_n13837), .B(u2__abc_44228_n13823), .Y(u2__abc_44228_n13838_1) );
  OR2X2 OR2X2_3112 ( .A(u2__abc_44228_n13841), .B(u2__abc_44228_n6818), .Y(u2__abc_44228_n13842) );
  OR2X2 OR2X2_3113 ( .A(u2__abc_44228_n13842), .B(u2__abc_44228_n5673), .Y(u2__abc_44228_n13843) );
  OR2X2 OR2X2_3114 ( .A(u2__abc_44228_n13848), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n13849) );
  OR2X2 OR2X2_3115 ( .A(u2__abc_44228_n13847), .B(u2__abc_44228_n13849), .Y(u2__abc_44228_n13850) );
  OR2X2 OR2X2_3116 ( .A(u2__abc_44228_n13854), .B(u2__abc_44228_n13840), .Y(u2__abc_44228_n13855_1) );
  OR2X2 OR2X2_3117 ( .A(u2__abc_44228_n13858), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n13859) );
  OR2X2 OR2X2_3118 ( .A(u2__abc_44228_n13861), .B(u2__abc_44228_n13860), .Y(u2__abc_44228_n13862) );
  OR2X2 OR2X2_3119 ( .A(u2__abc_44228_n13863_1), .B(u2__abc_44228_n5667), .Y(u2__abc_44228_n13864) );
  OR2X2 OR2X2_312 ( .A(a_112_bF_buf4), .B(\a[43] ), .Y(_abc_64468_n1299) );
  OR2X2 OR2X2_3120 ( .A(u2__abc_44228_n13866), .B(u2__abc_44228_n13859), .Y(u2__abc_44228_n13867) );
  OR2X2 OR2X2_3121 ( .A(u2__abc_44228_n13871), .B(u2__abc_44228_n13857), .Y(u2__abc_44228_n13872) );
  OR2X2 OR2X2_3122 ( .A(u2__abc_44228_n13875_1), .B(u2__abc_44228_n6823), .Y(u2__abc_44228_n13876) );
  OR2X2 OR2X2_3123 ( .A(u2__abc_44228_n13876), .B(u2__abc_44228_n5687), .Y(u2__abc_44228_n13879) );
  OR2X2 OR2X2_3124 ( .A(u2__abc_44228_n13882), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n13883_1) );
  OR2X2 OR2X2_3125 ( .A(u2__abc_44228_n13881), .B(u2__abc_44228_n13883_1), .Y(u2__abc_44228_n13884) );
  OR2X2 OR2X2_3126 ( .A(u2__abc_44228_n13888), .B(u2__abc_44228_n13874), .Y(u2__abc_44228_n13889) );
  OR2X2 OR2X2_3127 ( .A(u2__abc_44228_n13893), .B(u2__abc_44228_n13892_1), .Y(u2__abc_44228_n13894) );
  OR2X2 OR2X2_3128 ( .A(u2__abc_44228_n13895), .B(u2__abc_44228_n5681_1), .Y(u2__abc_44228_n13896) );
  OR2X2 OR2X2_3129 ( .A(u2__abc_44228_n13899), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n13900_1) );
  OR2X2 OR2X2_313 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[44] ), .Y(_abc_64468_n1300) );
  OR2X2 OR2X2_3130 ( .A(u2__abc_44228_n13898), .B(u2__abc_44228_n13900_1), .Y(u2__abc_44228_n13901) );
  OR2X2 OR2X2_3131 ( .A(u2__abc_44228_n13905), .B(u2__abc_44228_n13891), .Y(u2__abc_44228_n13906) );
  OR2X2 OR2X2_3132 ( .A(u2__abc_44228_n13909), .B(u2__abc_44228_n5679), .Y(u2__abc_44228_n13910_1) );
  OR2X2 OR2X2_3133 ( .A(u2__abc_44228_n13911), .B(u2__abc_44228_n5651), .Y(u2__abc_44228_n13914) );
  OR2X2 OR2X2_3134 ( .A(u2__abc_44228_n13917), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n13918_1) );
  OR2X2 OR2X2_3135 ( .A(u2__abc_44228_n13916), .B(u2__abc_44228_n13918_1), .Y(u2__abc_44228_n13919) );
  OR2X2 OR2X2_3136 ( .A(u2__abc_44228_n13923), .B(u2__abc_44228_n13908), .Y(u2__abc_44228_n13924) );
  OR2X2 OR2X2_3137 ( .A(u2__abc_44228_n13931), .B(u2__abc_44228_n13928), .Y(u2__abc_44228_n13932) );
  OR2X2 OR2X2_3138 ( .A(u2__abc_44228_n13934), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n13935_1) );
  OR2X2 OR2X2_3139 ( .A(u2__abc_44228_n13933), .B(u2__abc_44228_n13935_1), .Y(u2__abc_44228_n13936) );
  OR2X2 OR2X2_314 ( .A(a_112_bF_buf3), .B(\a[44] ), .Y(_abc_64468_n1302) );
  OR2X2 OR2X2_3140 ( .A(u2__abc_44228_n13940), .B(u2__abc_44228_n13926), .Y(u2__abc_44228_n13941) );
  OR2X2 OR2X2_3141 ( .A(u2__abc_44228_n13944), .B(u2__abc_44228_n5656), .Y(u2__abc_44228_n13945) );
  OR2X2 OR2X2_3142 ( .A(u2__abc_44228_n13946_1), .B(u2__abc_44228_n5644), .Y(u2__abc_44228_n13949) );
  OR2X2 OR2X2_3143 ( .A(u2__abc_44228_n13952), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n13953) );
  OR2X2 OR2X2_3144 ( .A(u2__abc_44228_n13951), .B(u2__abc_44228_n13953), .Y(u2__abc_44228_n13954_1) );
  OR2X2 OR2X2_3145 ( .A(u2__abc_44228_n13958), .B(u2__abc_44228_n13943), .Y(u2__abc_44228_n13959) );
  OR2X2 OR2X2_3146 ( .A(u2__abc_44228_n13947), .B(u2__abc_44228_n5640), .Y(u2__abc_44228_n13963_1) );
  OR2X2 OR2X2_3147 ( .A(u2__abc_44228_n13964), .B(u2__abc_44228_n13962), .Y(u2__abc_44228_n13965) );
  OR2X2 OR2X2_3148 ( .A(u2__abc_44228_n13963_1), .B(u2__abc_44228_n5638), .Y(u2__abc_44228_n13966) );
  OR2X2 OR2X2_3149 ( .A(u2__abc_44228_n13969), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n13970) );
  OR2X2 OR2X2_315 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[45] ), .Y(_abc_64468_n1303) );
  OR2X2 OR2X2_3150 ( .A(u2__abc_44228_n13968), .B(u2__abc_44228_n13970), .Y(u2__abc_44228_n13971_1) );
  OR2X2 OR2X2_3151 ( .A(u2__abc_44228_n13975), .B(u2__abc_44228_n13961), .Y(u2__abc_44228_n13976) );
  OR2X2 OR2X2_3152 ( .A(u2__abc_44228_n13979), .B(u2__abc_44228_n6839), .Y(u2__abc_44228_n13980) );
  OR2X2 OR2X2_3153 ( .A(u2__abc_44228_n13980), .B(u2__abc_44228_n5614), .Y(u2__abc_44228_n13983) );
  OR2X2 OR2X2_3154 ( .A(u2__abc_44228_n13986), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n13987) );
  OR2X2 OR2X2_3155 ( .A(u2__abc_44228_n13985), .B(u2__abc_44228_n13987), .Y(u2__abc_44228_n13988) );
  OR2X2 OR2X2_3156 ( .A(u2__abc_44228_n13992), .B(u2__abc_44228_n13978), .Y(u2__abc_44228_n13993) );
  OR2X2 OR2X2_3157 ( .A(u2__abc_44228_n13997), .B(u2__abc_44228_n13996), .Y(u2__abc_44228_n13998_1) );
  OR2X2 OR2X2_3158 ( .A(u2__abc_44228_n13999), .B(u2__abc_44228_n5608), .Y(u2__abc_44228_n14000) );
  OR2X2 OR2X2_3159 ( .A(u2__abc_44228_n14003), .B(u2__abc_44228_n2983_bF_buf30), .Y(u2__abc_44228_n14004) );
  OR2X2 OR2X2_316 ( .A(a_112_bF_buf2), .B(\a[45] ), .Y(_abc_64468_n1305) );
  OR2X2 OR2X2_3160 ( .A(u2__abc_44228_n14002), .B(u2__abc_44228_n14004), .Y(u2__abc_44228_n14005) );
  OR2X2 OR2X2_3161 ( .A(u2__abc_44228_n14009), .B(u2__abc_44228_n13995), .Y(u2__abc_44228_n14010) );
  OR2X2 OR2X2_3162 ( .A(u2__abc_44228_n14013), .B(u2__abc_44228_n6844), .Y(u2__abc_44228_n14014) );
  OR2X2 OR2X2_3163 ( .A(u2__abc_44228_n14014), .B(u2__abc_44228_n5628), .Y(u2__abc_44228_n14017) );
  OR2X2 OR2X2_3164 ( .A(u2__abc_44228_n14020), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n14021) );
  OR2X2 OR2X2_3165 ( .A(u2__abc_44228_n14019_1), .B(u2__abc_44228_n14021), .Y(u2__abc_44228_n14022) );
  OR2X2 OR2X2_3166 ( .A(u2__abc_44228_n14026), .B(u2__abc_44228_n14012), .Y(u2__abc_44228_n14027_1) );
  OR2X2 OR2X2_3167 ( .A(u2__abc_44228_n14031), .B(u2__abc_44228_n14030), .Y(u2__abc_44228_n14032) );
  OR2X2 OR2X2_3168 ( .A(u2__abc_44228_n14033), .B(u2__abc_44228_n5622), .Y(u2__abc_44228_n14034) );
  OR2X2 OR2X2_3169 ( .A(u2__abc_44228_n14037), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n14038) );
  OR2X2 OR2X2_317 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[46] ), .Y(_abc_64468_n1306) );
  OR2X2 OR2X2_3170 ( .A(u2__abc_44228_n14036_1), .B(u2__abc_44228_n14038), .Y(u2__abc_44228_n14039) );
  OR2X2 OR2X2_3171 ( .A(u2__abc_44228_n14043), .B(u2__abc_44228_n14029), .Y(u2__abc_44228_n14044_1) );
  OR2X2 OR2X2_3172 ( .A(u2__abc_44228_n14047), .B(u2__abc_44228_n5620), .Y(u2__abc_44228_n14048) );
  OR2X2 OR2X2_3173 ( .A(u2__abc_44228_n14049), .B(u2__abc_44228_n5599), .Y(u2__abc_44228_n14052) );
  OR2X2 OR2X2_3174 ( .A(u2__abc_44228_n14055), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n14056) );
  OR2X2 OR2X2_3175 ( .A(u2__abc_44228_n14054_1), .B(u2__abc_44228_n14056), .Y(u2__abc_44228_n14057) );
  OR2X2 OR2X2_3176 ( .A(u2__abc_44228_n14061), .B(u2__abc_44228_n14046), .Y(u2__abc_44228_n14062_1) );
  OR2X2 OR2X2_3177 ( .A(u2__abc_44228_n14069), .B(u2__abc_44228_n14066), .Y(u2__abc_44228_n14070) );
  OR2X2 OR2X2_3178 ( .A(u2__abc_44228_n14072), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n14073) );
  OR2X2 OR2X2_3179 ( .A(u2__abc_44228_n14071_1), .B(u2__abc_44228_n14073), .Y(u2__abc_44228_n14074) );
  OR2X2 OR2X2_318 ( .A(a_112_bF_buf1), .B(\a[46] ), .Y(_abc_64468_n1308) );
  OR2X2 OR2X2_3180 ( .A(u2__abc_44228_n14078), .B(u2__abc_44228_n14064), .Y(u2__abc_44228_n14079_1) );
  OR2X2 OR2X2_3181 ( .A(u2__abc_44228_n14082), .B(u2__abc_44228_n5591), .Y(u2__abc_44228_n14083) );
  OR2X2 OR2X2_3182 ( .A(u2__abc_44228_n14084), .B(u2__abc_44228_n5585), .Y(u2__abc_44228_n14087) );
  OR2X2 OR2X2_3183 ( .A(u2__abc_44228_n14090_1), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n14091) );
  OR2X2 OR2X2_3184 ( .A(u2__abc_44228_n14089), .B(u2__abc_44228_n14091), .Y(u2__abc_44228_n14092) );
  OR2X2 OR2X2_3185 ( .A(u2__abc_44228_n14096), .B(u2__abc_44228_n14081), .Y(u2__abc_44228_n14097) );
  OR2X2 OR2X2_3186 ( .A(u2__abc_44228_n14085), .B(u2__abc_44228_n5581), .Y(u2__abc_44228_n14101) );
  OR2X2 OR2X2_3187 ( .A(u2__abc_44228_n14102), .B(u2__abc_44228_n14100), .Y(u2__abc_44228_n14103) );
  OR2X2 OR2X2_3188 ( .A(u2__abc_44228_n14101), .B(u2__abc_44228_n5579), .Y(u2__abc_44228_n14104) );
  OR2X2 OR2X2_3189 ( .A(u2__abc_44228_n14107_1), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n14108) );
  OR2X2 OR2X2_319 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[47] ), .Y(_abc_64468_n1309) );
  OR2X2 OR2X2_3190 ( .A(u2__abc_44228_n14106), .B(u2__abc_44228_n14108), .Y(u2__abc_44228_n14109) );
  OR2X2 OR2X2_3191 ( .A(u2__abc_44228_n14113), .B(u2__abc_44228_n14099), .Y(u2__abc_44228_n14114) );
  OR2X2 OR2X2_3192 ( .A(u2__abc_44228_n6865), .B(u2__abc_44228_n7338), .Y(u2__abc_44228_n14119) );
  OR2X2 OR2X2_3193 ( .A(u2__abc_44228_n7548_1_bF_buf21), .B(u2__abc_44228_n14120), .Y(u2__abc_44228_n14121) );
  OR2X2 OR2X2_3194 ( .A(u2__abc_44228_n7547_bF_buf20), .B(u2_remHi_382_), .Y(u2__abc_44228_n14122) );
  OR2X2 OR2X2_3195 ( .A(u2__abc_44228_n14123), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n14124) );
  OR2X2 OR2X2_3196 ( .A(u2__abc_44228_n14128), .B(u2__abc_44228_n14116), .Y(u2__abc_44228_n14129) );
  OR2X2 OR2X2_3197 ( .A(u2__abc_44228_n14133_1), .B(u2__abc_44228_n14132), .Y(u2__abc_44228_n14134) );
  OR2X2 OR2X2_3198 ( .A(u2__abc_44228_n14135), .B(u2__abc_44228_n7332), .Y(u2__abc_44228_n14136) );
  OR2X2 OR2X2_3199 ( .A(u2__abc_44228_n14139), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n14140) );
  OR2X2 OR2X2_32 ( .A(_abc_64468_n753_bF_buf6), .B(\a[15] ), .Y(_abc_64468_n876) );
  OR2X2 OR2X2_320 ( .A(a_112_bF_buf0), .B(\a[47] ), .Y(_abc_64468_n1311) );
  OR2X2 OR2X2_3200 ( .A(u2__abc_44228_n14140), .B(u2__abc_44228_n14138), .Y(u2__abc_44228_n14141) );
  OR2X2 OR2X2_3201 ( .A(u2__abc_44228_n14145), .B(u2__abc_44228_n14131), .Y(u2__abc_44228_n14146) );
  OR2X2 OR2X2_3202 ( .A(u2__abc_44228_n14149), .B(u2__abc_44228_n7349), .Y(u2__abc_44228_n14150_1) );
  OR2X2 OR2X2_3203 ( .A(u2__abc_44228_n14150_1), .B(u2__abc_44228_n7324), .Y(u2__abc_44228_n14153) );
  OR2X2 OR2X2_3204 ( .A(u2__abc_44228_n7548_1_bF_buf19), .B(u2__abc_44228_n14154), .Y(u2__abc_44228_n14155) );
  OR2X2 OR2X2_3205 ( .A(u2__abc_44228_n7547_bF_buf18), .B(u2_remHi_384_), .Y(u2__abc_44228_n14156) );
  OR2X2 OR2X2_3206 ( .A(u2__abc_44228_n14157), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n14158) );
  OR2X2 OR2X2_3207 ( .A(u2__abc_44228_n14162_1), .B(u2__abc_44228_n14148), .Y(u2__abc_44228_n14163) );
  OR2X2 OR2X2_3208 ( .A(u2__abc_44228_n14151), .B(u2__abc_44228_n7320), .Y(u2__abc_44228_n14167) );
  OR2X2 OR2X2_3209 ( .A(u2__abc_44228_n14168), .B(u2__abc_44228_n14166), .Y(u2__abc_44228_n14169) );
  OR2X2 OR2X2_321 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[48] ), .Y(_abc_64468_n1312) );
  OR2X2 OR2X2_3210 ( .A(u2__abc_44228_n14167), .B(u2__abc_44228_n7318), .Y(u2__abc_44228_n14170_1) );
  OR2X2 OR2X2_3211 ( .A(u2__abc_44228_n14173), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n14174) );
  OR2X2 OR2X2_3212 ( .A(u2__abc_44228_n14172), .B(u2__abc_44228_n14174), .Y(u2__abc_44228_n14175) );
  OR2X2 OR2X2_3213 ( .A(u2__abc_44228_n14179_1), .B(u2__abc_44228_n14165), .Y(u2__abc_44228_n14180) );
  OR2X2 OR2X2_3214 ( .A(u2__abc_44228_n14183), .B(u2__abc_44228_n7353), .Y(u2__abc_44228_n14184) );
  OR2X2 OR2X2_3215 ( .A(u2__abc_44228_n14184), .B(u2__abc_44228_n7302), .Y(u2__abc_44228_n14185) );
  OR2X2 OR2X2_3216 ( .A(u2__abc_44228_n7548_1_bF_buf17), .B(u2__abc_44228_n14188), .Y(u2__abc_44228_n14189) );
  OR2X2 OR2X2_3217 ( .A(u2__abc_44228_n7547_bF_buf16), .B(u2_remHi_386_), .Y(u2__abc_44228_n14190) );
  OR2X2 OR2X2_3218 ( .A(u2__abc_44228_n14191), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n14192) );
  OR2X2 OR2X2_3219 ( .A(u2__abc_44228_n14196), .B(u2__abc_44228_n14182), .Y(u2__abc_44228_n14197_1) );
  OR2X2 OR2X2_322 ( .A(a_112_bF_buf9), .B(\a[48] ), .Y(_abc_64468_n1314) );
  OR2X2 OR2X2_3220 ( .A(u2__abc_44228_n14201), .B(u2__abc_44228_n7309_1), .Y(u2__abc_44228_n14202) );
  OR2X2 OR2X2_3221 ( .A(u2__abc_44228_n14200), .B(u2__abc_44228_n14203), .Y(u2__abc_44228_n14204) );
  OR2X2 OR2X2_3222 ( .A(u2__abc_44228_n14207), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n14208) );
  OR2X2 OR2X2_3223 ( .A(u2__abc_44228_n14206), .B(u2__abc_44228_n14208), .Y(u2__abc_44228_n14209) );
  OR2X2 OR2X2_3224 ( .A(u2__abc_44228_n14213), .B(u2__abc_44228_n14199), .Y(u2__abc_44228_n14214_1) );
  OR2X2 OR2X2_3225 ( .A(u2__abc_44228_n14217), .B(u2__abc_44228_n7307), .Y(u2__abc_44228_n14218) );
  OR2X2 OR2X2_3226 ( .A(u2__abc_44228_n14219), .B(u2__abc_44228_n7295), .Y(u2__abc_44228_n14222_1) );
  OR2X2 OR2X2_3227 ( .A(u2__abc_44228_n14225), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n14226) );
  OR2X2 OR2X2_3228 ( .A(u2__abc_44228_n14224), .B(u2__abc_44228_n14226), .Y(u2__abc_44228_n14227) );
  OR2X2 OR2X2_3229 ( .A(u2__abc_44228_n14231), .B(u2__abc_44228_n14216), .Y(u2__abc_44228_n14232) );
  OR2X2 OR2X2_323 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[49] ), .Y(_abc_64468_n1315) );
  OR2X2 OR2X2_3230 ( .A(u2__abc_44228_n14220), .B(u2__abc_44228_n7291), .Y(u2__abc_44228_n14236) );
  OR2X2 OR2X2_3231 ( .A(u2__abc_44228_n14237), .B(u2__abc_44228_n14235), .Y(u2__abc_44228_n14238) );
  OR2X2 OR2X2_3232 ( .A(u2__abc_44228_n14236), .B(u2__abc_44228_n7289_1), .Y(u2__abc_44228_n14239) );
  OR2X2 OR2X2_3233 ( .A(u2__abc_44228_n14242), .B(u2__abc_44228_n2983_bF_buf4), .Y(u2__abc_44228_n14243) );
  OR2X2 OR2X2_3234 ( .A(u2__abc_44228_n14241_1), .B(u2__abc_44228_n14243), .Y(u2__abc_44228_n14244) );
  OR2X2 OR2X2_3235 ( .A(u2__abc_44228_n14248), .B(u2__abc_44228_n14234), .Y(u2__abc_44228_n14249) );
  OR2X2 OR2X2_3236 ( .A(u2__abc_44228_n14252), .B(u2__abc_44228_n7363), .Y(u2__abc_44228_n14253) );
  OR2X2 OR2X2_3237 ( .A(u2__abc_44228_n14253), .B(u2__abc_44228_n7272), .Y(u2__abc_44228_n14256) );
  OR2X2 OR2X2_3238 ( .A(u2__abc_44228_n7548_1_bF_buf13), .B(u2__abc_44228_n14257), .Y(u2__abc_44228_n14258_1) );
  OR2X2 OR2X2_3239 ( .A(u2__abc_44228_n7547_bF_buf12), .B(u2_remHi_390_), .Y(u2__abc_44228_n14259) );
  OR2X2 OR2X2_324 ( .A(a_112_bF_buf8), .B(\a[49] ), .Y(_abc_64468_n1317) );
  OR2X2 OR2X2_3240 ( .A(u2__abc_44228_n14260), .B(u2__abc_44228_n2983_bF_buf2), .Y(u2__abc_44228_n14261) );
  OR2X2 OR2X2_3241 ( .A(u2__abc_44228_n14265), .B(u2__abc_44228_n14251), .Y(u2__abc_44228_n14266) );
  OR2X2 OR2X2_3242 ( .A(u2__abc_44228_n14270), .B(u2__abc_44228_n14269), .Y(u2__abc_44228_n14271) );
  OR2X2 OR2X2_3243 ( .A(u2__abc_44228_n14272), .B(u2__abc_44228_n7279), .Y(u2__abc_44228_n14273) );
  OR2X2 OR2X2_3244 ( .A(u2__abc_44228_n14276_1), .B(u2__abc_44228_n2983_bF_buf0), .Y(u2__abc_44228_n14277) );
  OR2X2 OR2X2_3245 ( .A(u2__abc_44228_n14275), .B(u2__abc_44228_n14277), .Y(u2__abc_44228_n14278) );
  OR2X2 OR2X2_3246 ( .A(u2__abc_44228_n14282), .B(u2__abc_44228_n14268_1), .Y(u2__abc_44228_n14283) );
  OR2X2 OR2X2_3247 ( .A(u2__abc_44228_n14286), .B(u2__abc_44228_n7277), .Y(u2__abc_44228_n14287) );
  OR2X2 OR2X2_3248 ( .A(u2__abc_44228_n14288), .B(u2__abc_44228_n7265), .Y(u2__abc_44228_n14291) );
  OR2X2 OR2X2_3249 ( .A(u2__abc_44228_n14294), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n14295) );
  OR2X2 OR2X2_325 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[50] ), .Y(_abc_64468_n1318) );
  OR2X2 OR2X2_3250 ( .A(u2__abc_44228_n14293_1), .B(u2__abc_44228_n14295), .Y(u2__abc_44228_n14296) );
  OR2X2 OR2X2_3251 ( .A(u2__abc_44228_n14300), .B(u2__abc_44228_n14285_1), .Y(u2__abc_44228_n14301) );
  OR2X2 OR2X2_3252 ( .A(u2__abc_44228_n14289), .B(u2__abc_44228_n7261), .Y(u2__abc_44228_n14305) );
  OR2X2 OR2X2_3253 ( .A(u2__abc_44228_n14306), .B(u2__abc_44228_n14304), .Y(u2__abc_44228_n14307_1) );
  OR2X2 OR2X2_3254 ( .A(u2__abc_44228_n14305), .B(u2__abc_44228_n7259), .Y(u2__abc_44228_n14308) );
  OR2X2 OR2X2_3255 ( .A(u2__abc_44228_n14311), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n14312) );
  OR2X2 OR2X2_3256 ( .A(u2__abc_44228_n14310), .B(u2__abc_44228_n14312), .Y(u2__abc_44228_n14313) );
  OR2X2 OR2X2_3257 ( .A(u2__abc_44228_n14317), .B(u2__abc_44228_n14303), .Y(u2__abc_44228_n14318) );
  OR2X2 OR2X2_3258 ( .A(u2__abc_44228_n14321), .B(u2__abc_44228_n7372), .Y(u2__abc_44228_n14322) );
  OR2X2 OR2X2_3259 ( .A(u2__abc_44228_n14322), .B(u2__abc_44228_n7243), .Y(u2__abc_44228_n14323) );
  OR2X2 OR2X2_326 ( .A(a_112_bF_buf7), .B(\a[50] ), .Y(_abc_64468_n1320) );
  OR2X2 OR2X2_3260 ( .A(u2__abc_44228_n14328), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n14329) );
  OR2X2 OR2X2_3261 ( .A(u2__abc_44228_n14327), .B(u2__abc_44228_n14329), .Y(u2__abc_44228_n14330) );
  OR2X2 OR2X2_3262 ( .A(u2__abc_44228_n14334), .B(u2__abc_44228_n14320), .Y(u2__abc_44228_n14335) );
  OR2X2 OR2X2_3263 ( .A(u2__abc_44228_n14342_1), .B(u2__abc_44228_n14339), .Y(u2__abc_44228_n14343) );
  OR2X2 OR2X2_3264 ( .A(u2__abc_44228_n14345), .B(u2__abc_44228_n2983_bF_buf136), .Y(u2__abc_44228_n14346) );
  OR2X2 OR2X2_3265 ( .A(u2__abc_44228_n14344), .B(u2__abc_44228_n14346), .Y(u2__abc_44228_n14347) );
  OR2X2 OR2X2_3266 ( .A(u2__abc_44228_n14351), .B(u2__abc_44228_n14337), .Y(u2__abc_44228_n14352) );
  OR2X2 OR2X2_3267 ( .A(u2__abc_44228_n14355), .B(u2__abc_44228_n7248), .Y(u2__abc_44228_n14356) );
  OR2X2 OR2X2_3268 ( .A(u2__abc_44228_n14357), .B(u2__abc_44228_n7236), .Y(u2__abc_44228_n14360) );
  OR2X2 OR2X2_3269 ( .A(u2__abc_44228_n14363), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n14364) );
  OR2X2 OR2X2_327 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[51] ), .Y(_abc_64468_n1321) );
  OR2X2 OR2X2_3270 ( .A(u2__abc_44228_n14362), .B(u2__abc_44228_n14364), .Y(u2__abc_44228_n14365) );
  OR2X2 OR2X2_3271 ( .A(u2__abc_44228_n14369), .B(u2__abc_44228_n14354), .Y(u2__abc_44228_n14370) );
  OR2X2 OR2X2_3272 ( .A(u2__abc_44228_n14358), .B(u2__abc_44228_n7232), .Y(u2__abc_44228_n14374) );
  OR2X2 OR2X2_3273 ( .A(u2__abc_44228_n14375), .B(u2__abc_44228_n14373), .Y(u2__abc_44228_n14376) );
  OR2X2 OR2X2_3274 ( .A(u2__abc_44228_n14374), .B(u2__abc_44228_n7230), .Y(u2__abc_44228_n14377) );
  OR2X2 OR2X2_3275 ( .A(u2__abc_44228_n14380), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n14381) );
  OR2X2 OR2X2_3276 ( .A(u2__abc_44228_n14379), .B(u2__abc_44228_n14381), .Y(u2__abc_44228_n14382) );
  OR2X2 OR2X2_3277 ( .A(u2__abc_44228_n14386_1), .B(u2__abc_44228_n14372), .Y(u2__abc_44228_n14387) );
  OR2X2 OR2X2_3278 ( .A(u2__abc_44228_n14390), .B(u2__abc_44228_n7383), .Y(u2__abc_44228_n14391) );
  OR2X2 OR2X2_3279 ( .A(u2__abc_44228_n14391), .B(u2__abc_44228_n7212), .Y(u2__abc_44228_n14392) );
  OR2X2 OR2X2_328 ( .A(a_112_bF_buf6), .B(\a[51] ), .Y(_abc_64468_n1323) );
  OR2X2 OR2X2_3280 ( .A(u2__abc_44228_n7548_1_bF_buf5), .B(u2__abc_44228_n14395_1), .Y(u2__abc_44228_n14396) );
  OR2X2 OR2X2_3281 ( .A(u2__abc_44228_n7547_bF_buf4), .B(u2_remHi_398_), .Y(u2__abc_44228_n14397) );
  OR2X2 OR2X2_3282 ( .A(u2__abc_44228_n14398), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n14399) );
  OR2X2 OR2X2_3283 ( .A(u2__abc_44228_n14403_1), .B(u2__abc_44228_n14389), .Y(u2__abc_44228_n14404) );
  OR2X2 OR2X2_3284 ( .A(u2__abc_44228_n14411), .B(u2__abc_44228_n14408), .Y(u2__abc_44228_n14412) );
  OR2X2 OR2X2_3285 ( .A(u2__abc_44228_n14414), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n14415) );
  OR2X2 OR2X2_3286 ( .A(u2__abc_44228_n14413_1), .B(u2__abc_44228_n14415), .Y(u2__abc_44228_n14416) );
  OR2X2 OR2X2_3287 ( .A(u2__abc_44228_n14420), .B(u2__abc_44228_n14406), .Y(u2__abc_44228_n14421_1) );
  OR2X2 OR2X2_3288 ( .A(u2__abc_44228_n14424), .B(u2__abc_44228_n7217), .Y(u2__abc_44228_n14425) );
  OR2X2 OR2X2_3289 ( .A(u2__abc_44228_n14426), .B(u2__abc_44228_n7205), .Y(u2__abc_44228_n14429) );
  OR2X2 OR2X2_329 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[52] ), .Y(_abc_64468_n1324) );
  OR2X2 OR2X2_3290 ( .A(u2__abc_44228_n14432), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n14433) );
  OR2X2 OR2X2_3291 ( .A(u2__abc_44228_n14431), .B(u2__abc_44228_n14433), .Y(u2__abc_44228_n14434) );
  OR2X2 OR2X2_3292 ( .A(u2__abc_44228_n14438_1), .B(u2__abc_44228_n14423), .Y(u2__abc_44228_n14439) );
  OR2X2 OR2X2_3293 ( .A(u2__abc_44228_n14427), .B(u2__abc_44228_n7201), .Y(u2__abc_44228_n14443) );
  OR2X2 OR2X2_3294 ( .A(u2__abc_44228_n14444), .B(u2__abc_44228_n14442), .Y(u2__abc_44228_n14445) );
  OR2X2 OR2X2_3295 ( .A(u2__abc_44228_n14443), .B(u2__abc_44228_n7199), .Y(u2__abc_44228_n14446) );
  OR2X2 OR2X2_3296 ( .A(u2__abc_44228_n14449), .B(u2__abc_44228_n2983_bF_buf126), .Y(u2__abc_44228_n14450_1) );
  OR2X2 OR2X2_3297 ( .A(u2__abc_44228_n14448), .B(u2__abc_44228_n14450_1), .Y(u2__abc_44228_n14451) );
  OR2X2 OR2X2_3298 ( .A(u2__abc_44228_n14455), .B(u2__abc_44228_n14441), .Y(u2__abc_44228_n14456) );
  OR2X2 OR2X2_3299 ( .A(u2__abc_44228_n14459), .B(u2__abc_44228_n7392_1), .Y(u2__abc_44228_n14460) );
  OR2X2 OR2X2_33 ( .A(aNan_bF_buf4), .B(sqrto_92_), .Y(_abc_64468_n878) );
  OR2X2 OR2X2_330 ( .A(a_112_bF_buf5), .B(\a[52] ), .Y(_abc_64468_n1326) );
  OR2X2 OR2X2_3300 ( .A(u2__abc_44228_n14460), .B(u2__abc_44228_n7190), .Y(u2__abc_44228_n14461) );
  OR2X2 OR2X2_3301 ( .A(u2__abc_44228_n14466), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n14467_1) );
  OR2X2 OR2X2_3302 ( .A(u2__abc_44228_n14465), .B(u2__abc_44228_n14467_1), .Y(u2__abc_44228_n14468) );
  OR2X2 OR2X2_3303 ( .A(u2__abc_44228_n14472), .B(u2__abc_44228_n14458_1), .Y(u2__abc_44228_n14473) );
  OR2X2 OR2X2_3304 ( .A(u2__abc_44228_n14477), .B(u2__abc_44228_n14476), .Y(u2__abc_44228_n14478) );
  OR2X2 OR2X2_3305 ( .A(u2__abc_44228_n14479), .B(u2__abc_44228_n7184), .Y(u2__abc_44228_n14480) );
  OR2X2 OR2X2_3306 ( .A(u2__abc_44228_n14483), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n14484) );
  OR2X2 OR2X2_3307 ( .A(u2__abc_44228_n14482), .B(u2__abc_44228_n14484), .Y(u2__abc_44228_n14485_1) );
  OR2X2 OR2X2_3308 ( .A(u2__abc_44228_n14489), .B(u2__abc_44228_n14475_1), .Y(u2__abc_44228_n14490) );
  OR2X2 OR2X2_3309 ( .A(u2__abc_44228_n14493_1), .B(u2__abc_44228_n7397), .Y(u2__abc_44228_n14494) );
  OR2X2 OR2X2_331 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[53] ), .Y(_abc_64468_n1327) );
  OR2X2 OR2X2_3310 ( .A(u2__abc_44228_n14494), .B(u2__abc_44228_n7176), .Y(u2__abc_44228_n14497) );
  OR2X2 OR2X2_3311 ( .A(u2__abc_44228_n14500), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n14501) );
  OR2X2 OR2X2_3312 ( .A(u2__abc_44228_n14499), .B(u2__abc_44228_n14501), .Y(u2__abc_44228_n14502_1) );
  OR2X2 OR2X2_3313 ( .A(u2__abc_44228_n14506), .B(u2__abc_44228_n14492), .Y(u2__abc_44228_n14507) );
  OR2X2 OR2X2_3314 ( .A(u2__abc_44228_n14495), .B(u2__abc_44228_n7172), .Y(u2__abc_44228_n14511) );
  OR2X2 OR2X2_3315 ( .A(u2__abc_44228_n14512), .B(u2__abc_44228_n14510_1), .Y(u2__abc_44228_n14513) );
  OR2X2 OR2X2_3316 ( .A(u2__abc_44228_n14511), .B(u2__abc_44228_n7170_1), .Y(u2__abc_44228_n14514) );
  OR2X2 OR2X2_3317 ( .A(u2__abc_44228_n14517), .B(u2__abc_44228_n2983_bF_buf120), .Y(u2__abc_44228_n14518) );
  OR2X2 OR2X2_3318 ( .A(u2__abc_44228_n14516), .B(u2__abc_44228_n14518), .Y(u2__abc_44228_n14519) );
  OR2X2 OR2X2_3319 ( .A(u2__abc_44228_n14523), .B(u2__abc_44228_n14509), .Y(u2__abc_44228_n14524) );
  OR2X2 OR2X2_332 ( .A(a_112_bF_buf4), .B(\a[53] ), .Y(_abc_64468_n1329) );
  OR2X2 OR2X2_3320 ( .A(u2__abc_44228_n14527), .B(u2__abc_44228_n7402), .Y(u2__abc_44228_n14528) );
  OR2X2 OR2X2_3321 ( .A(u2__abc_44228_n14528), .B(u2__abc_44228_n7160), .Y(u2__abc_44228_n14531) );
  OR2X2 OR2X2_3322 ( .A(u2__abc_44228_n14534), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n14535) );
  OR2X2 OR2X2_3323 ( .A(u2__abc_44228_n14533), .B(u2__abc_44228_n14535), .Y(u2__abc_44228_n14536) );
  OR2X2 OR2X2_3324 ( .A(u2__abc_44228_n14540), .B(u2__abc_44228_n14526), .Y(u2__abc_44228_n14541) );
  OR2X2 OR2X2_3325 ( .A(u2__abc_44228_n14545), .B(u2__abc_44228_n14544), .Y(u2__abc_44228_n14546_1) );
  OR2X2 OR2X2_3326 ( .A(u2__abc_44228_n14547), .B(u2__abc_44228_n7154), .Y(u2__abc_44228_n14548) );
  OR2X2 OR2X2_3327 ( .A(u2__abc_44228_n14551), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n14552) );
  OR2X2 OR2X2_3328 ( .A(u2__abc_44228_n14550), .B(u2__abc_44228_n14552), .Y(u2__abc_44228_n14553) );
  OR2X2 OR2X2_3329 ( .A(u2__abc_44228_n14557), .B(u2__abc_44228_n14543), .Y(u2__abc_44228_n14558) );
  OR2X2 OR2X2_333 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[54] ), .Y(_abc_64468_n1330) );
  OR2X2 OR2X2_3330 ( .A(u2__abc_44228_n14561), .B(u2__abc_44228_n7152), .Y(u2__abc_44228_n14562) );
  OR2X2 OR2X2_3331 ( .A(u2__abc_44228_n14563), .B(u2__abc_44228_n7146), .Y(u2__abc_44228_n14566) );
  OR2X2 OR2X2_3332 ( .A(u2__abc_44228_n14569), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n14570) );
  OR2X2 OR2X2_3333 ( .A(u2__abc_44228_n14568), .B(u2__abc_44228_n14570), .Y(u2__abc_44228_n14571) );
  OR2X2 OR2X2_3334 ( .A(u2__abc_44228_n14575), .B(u2__abc_44228_n14560), .Y(u2__abc_44228_n14576) );
  OR2X2 OR2X2_3335 ( .A(u2__abc_44228_n14564_1), .B(u2__abc_44228_n7142), .Y(u2__abc_44228_n14580) );
  OR2X2 OR2X2_3336 ( .A(u2__abc_44228_n14581_1), .B(u2__abc_44228_n14579), .Y(u2__abc_44228_n14582) );
  OR2X2 OR2X2_3337 ( .A(u2__abc_44228_n14580), .B(u2__abc_44228_n7140), .Y(u2__abc_44228_n14583) );
  OR2X2 OR2X2_3338 ( .A(u2__abc_44228_n14586), .B(u2__abc_44228_n2983_bF_buf114), .Y(u2__abc_44228_n14587) );
  OR2X2 OR2X2_3339 ( .A(u2__abc_44228_n14585), .B(u2__abc_44228_n14587), .Y(u2__abc_44228_n14588) );
  OR2X2 OR2X2_334 ( .A(a_112_bF_buf3), .B(\a[54] ), .Y(_abc_64468_n1332) );
  OR2X2 OR2X2_3340 ( .A(u2__abc_44228_n14592), .B(u2__abc_44228_n14578), .Y(u2__abc_44228_n14593) );
  OR2X2 OR2X2_3341 ( .A(u2__abc_44228_n14596), .B(u2__abc_44228_n7411), .Y(u2__abc_44228_n14597) );
  OR2X2 OR2X2_3342 ( .A(u2__abc_44228_n14597), .B(u2__abc_44228_n7131), .Y(u2__abc_44228_n14598) );
  OR2X2 OR2X2_3343 ( .A(u2__abc_44228_n14603), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n14604) );
  OR2X2 OR2X2_3344 ( .A(u2__abc_44228_n14602_1), .B(u2__abc_44228_n14604), .Y(u2__abc_44228_n14605) );
  OR2X2 OR2X2_3345 ( .A(u2__abc_44228_n14609), .B(u2__abc_44228_n14595), .Y(u2__abc_44228_n14610) );
  OR2X2 OR2X2_3346 ( .A(u2__abc_44228_n14614), .B(u2__abc_44228_n7125_1), .Y(u2__abc_44228_n14615) );
  OR2X2 OR2X2_3347 ( .A(u2__abc_44228_n14613), .B(u2__abc_44228_n14616), .Y(u2__abc_44228_n14617) );
  OR2X2 OR2X2_3348 ( .A(u2__abc_44228_n14620), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n14621) );
  OR2X2 OR2X2_3349 ( .A(u2__abc_44228_n14619_1), .B(u2__abc_44228_n14621), .Y(u2__abc_44228_n14622) );
  OR2X2 OR2X2_335 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[55] ), .Y(_abc_64468_n1333) );
  OR2X2 OR2X2_3350 ( .A(u2__abc_44228_n14626), .B(u2__abc_44228_n14612), .Y(u2__abc_44228_n14627) );
  OR2X2 OR2X2_3351 ( .A(u2__abc_44228_n14630), .B(u2__abc_44228_n7123), .Y(u2__abc_44228_n14631) );
  OR2X2 OR2X2_3352 ( .A(u2__abc_44228_n14632), .B(u2__abc_44228_n7117), .Y(u2__abc_44228_n14635) );
  OR2X2 OR2X2_3353 ( .A(u2__abc_44228_n14638), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n14639) );
  OR2X2 OR2X2_3354 ( .A(u2__abc_44228_n14637_1), .B(u2__abc_44228_n14639), .Y(u2__abc_44228_n14640) );
  OR2X2 OR2X2_3355 ( .A(u2__abc_44228_n14644), .B(u2__abc_44228_n14629_1), .Y(u2__abc_44228_n14645) );
  OR2X2 OR2X2_3356 ( .A(u2__abc_44228_n14633), .B(u2__abc_44228_n7113), .Y(u2__abc_44228_n14649) );
  OR2X2 OR2X2_3357 ( .A(u2__abc_44228_n14650), .B(u2__abc_44228_n14648), .Y(u2__abc_44228_n14651) );
  OR2X2 OR2X2_3358 ( .A(u2__abc_44228_n14649), .B(u2__abc_44228_n7111), .Y(u2__abc_44228_n14652) );
  OR2X2 OR2X2_3359 ( .A(u2__abc_44228_n14655), .B(u2__abc_44228_n2983_bF_buf108), .Y(u2__abc_44228_n14656) );
  OR2X2 OR2X2_336 ( .A(a_112_bF_buf2), .B(\a[55] ), .Y(_abc_64468_n1335) );
  OR2X2 OR2X2_3360 ( .A(u2__abc_44228_n14654_1), .B(u2__abc_44228_n14656), .Y(u2__abc_44228_n14657) );
  OR2X2 OR2X2_3361 ( .A(u2__abc_44228_n14661), .B(u2__abc_44228_n14647), .Y(u2__abc_44228_n14662) );
  OR2X2 OR2X2_3362 ( .A(u2__abc_44228_n14665_1), .B(u2__abc_44228_n7423), .Y(u2__abc_44228_n14666) );
  OR2X2 OR2X2_3363 ( .A(u2__abc_44228_n14666), .B(u2__abc_44228_n7092), .Y(u2__abc_44228_n14669) );
  OR2X2 OR2X2_3364 ( .A(u2__abc_44228_n7548_1_bF_buf47), .B(u2__abc_44228_n14670), .Y(u2__abc_44228_n14671) );
  OR2X2 OR2X2_3365 ( .A(u2__abc_44228_n7547_bF_buf46), .B(u2_remHi_414_), .Y(u2__abc_44228_n14672) );
  OR2X2 OR2X2_3366 ( .A(u2__abc_44228_n14673_1), .B(u2__abc_44228_n2983_bF_buf106), .Y(u2__abc_44228_n14674) );
  OR2X2 OR2X2_3367 ( .A(u2__abc_44228_n14678), .B(u2__abc_44228_n14664), .Y(u2__abc_44228_n14679) );
  OR2X2 OR2X2_3368 ( .A(u2__abc_44228_n14686), .B(u2__abc_44228_n14683), .Y(u2__abc_44228_n14687) );
  OR2X2 OR2X2_3369 ( .A(u2__abc_44228_n14689), .B(u2__abc_44228_n2983_bF_buf104), .Y(u2__abc_44228_n14690_1) );
  OR2X2 OR2X2_337 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[56] ), .Y(_abc_64468_n1336) );
  OR2X2 OR2X2_3370 ( .A(u2__abc_44228_n14688), .B(u2__abc_44228_n14690_1), .Y(u2__abc_44228_n14691) );
  OR2X2 OR2X2_3371 ( .A(u2__abc_44228_n14695), .B(u2__abc_44228_n14681), .Y(u2__abc_44228_n14696) );
  OR2X2 OR2X2_3372 ( .A(u2__abc_44228_n14699), .B(u2__abc_44228_n7097), .Y(u2__abc_44228_n14700_1) );
  OR2X2 OR2X2_3373 ( .A(u2__abc_44228_n14701), .B(u2__abc_44228_n7085), .Y(u2__abc_44228_n14704) );
  OR2X2 OR2X2_3374 ( .A(u2__abc_44228_n14707), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n14708_1) );
  OR2X2 OR2X2_3375 ( .A(u2__abc_44228_n14706), .B(u2__abc_44228_n14708_1), .Y(u2__abc_44228_n14709) );
  OR2X2 OR2X2_3376 ( .A(u2__abc_44228_n14713), .B(u2__abc_44228_n14698), .Y(u2__abc_44228_n14714) );
  OR2X2 OR2X2_3377 ( .A(u2__abc_44228_n14702), .B(u2__abc_44228_n7081), .Y(u2__abc_44228_n14718) );
  OR2X2 OR2X2_3378 ( .A(u2__abc_44228_n14719), .B(u2__abc_44228_n14717_1), .Y(u2__abc_44228_n14720) );
  OR2X2 OR2X2_3379 ( .A(u2__abc_44228_n14718), .B(u2__abc_44228_n7079), .Y(u2__abc_44228_n14721) );
  OR2X2 OR2X2_338 ( .A(a_112_bF_buf1), .B(\a[56] ), .Y(_abc_64468_n1338) );
  OR2X2 OR2X2_3380 ( .A(u2__abc_44228_n14724), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n14725_1) );
  OR2X2 OR2X2_3381 ( .A(u2__abc_44228_n14723), .B(u2__abc_44228_n14725_1), .Y(u2__abc_44228_n14726) );
  OR2X2 OR2X2_3382 ( .A(u2__abc_44228_n14730), .B(u2__abc_44228_n14716), .Y(u2__abc_44228_n14731) );
  OR2X2 OR2X2_3383 ( .A(u2__abc_44228_n14734), .B(u2__abc_44228_n7432), .Y(u2__abc_44228_n14735) );
  OR2X2 OR2X2_3384 ( .A(u2__abc_44228_n14735), .B(u2__abc_44228_n7070), .Y(u2__abc_44228_n14736) );
  OR2X2 OR2X2_3385 ( .A(u2__abc_44228_n14741), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n14742) );
  OR2X2 OR2X2_3386 ( .A(u2__abc_44228_n14740), .B(u2__abc_44228_n14742), .Y(u2__abc_44228_n14743) );
  OR2X2 OR2X2_3387 ( .A(u2__abc_44228_n14747), .B(u2__abc_44228_n14733), .Y(u2__abc_44228_n14748) );
  OR2X2 OR2X2_3388 ( .A(u2__abc_44228_n14752), .B(u2__abc_44228_n14751), .Y(u2__abc_44228_n14753) );
  OR2X2 OR2X2_3389 ( .A(u2__abc_44228_n14754_1), .B(u2__abc_44228_n7064), .Y(u2__abc_44228_n14755) );
  OR2X2 OR2X2_339 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[57] ), .Y(_abc_64468_n1339) );
  OR2X2 OR2X2_3390 ( .A(u2__abc_44228_n14758), .B(u2__abc_44228_n2983_bF_buf98), .Y(u2__abc_44228_n14759) );
  OR2X2 OR2X2_3391 ( .A(u2__abc_44228_n14757), .B(u2__abc_44228_n14759), .Y(u2__abc_44228_n14760) );
  OR2X2 OR2X2_3392 ( .A(u2__abc_44228_n14764), .B(u2__abc_44228_n14750), .Y(u2__abc_44228_n14765) );
  OR2X2 OR2X2_3393 ( .A(u2__abc_44228_n14768), .B(u2__abc_44228_n7437_1), .Y(u2__abc_44228_n14769) );
  OR2X2 OR2X2_3394 ( .A(u2__abc_44228_n14769), .B(u2__abc_44228_n7056), .Y(u2__abc_44228_n14772_1) );
  OR2X2 OR2X2_3395 ( .A(u2__abc_44228_n14775), .B(u2__abc_44228_n8209_bF_buf8), .Y(u2__abc_44228_n14776) );
  OR2X2 OR2X2_3396 ( .A(u2__abc_44228_n14774), .B(u2__abc_44228_n14776), .Y(u2__abc_44228_n14777) );
  OR2X2 OR2X2_3397 ( .A(u2__abc_44228_n14781), .B(u2__abc_44228_n14767), .Y(u2__abc_44228_n14782) );
  OR2X2 OR2X2_3398 ( .A(u2__abc_44228_n14770), .B(u2__abc_44228_n7052), .Y(u2__abc_44228_n14786) );
  OR2X2 OR2X2_3399 ( .A(u2__abc_44228_n14787), .B(u2__abc_44228_n14785), .Y(u2__abc_44228_n14788) );
  OR2X2 OR2X2_34 ( .A(_abc_64468_n753_bF_buf5), .B(\a[16] ), .Y(_abc_64468_n879) );
  OR2X2 OR2X2_340 ( .A(a_112_bF_buf0), .B(\a[57] ), .Y(_abc_64468_n1341) );
  OR2X2 OR2X2_3400 ( .A(u2__abc_44228_n14786), .B(u2__abc_44228_n7050_1), .Y(u2__abc_44228_n14789_1) );
  OR2X2 OR2X2_3401 ( .A(u2__abc_44228_n14792), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n14793) );
  OR2X2 OR2X2_3402 ( .A(u2__abc_44228_n14791), .B(u2__abc_44228_n14793), .Y(u2__abc_44228_n14794) );
  OR2X2 OR2X2_3403 ( .A(u2__abc_44228_n14798), .B(u2__abc_44228_n14784), .Y(u2__abc_44228_n14799) );
  OR2X2 OR2X2_3404 ( .A(u2__abc_44228_n14802), .B(u2__abc_44228_n7442), .Y(u2__abc_44228_n14803) );
  OR2X2 OR2X2_3405 ( .A(u2__abc_44228_n14803), .B(u2__abc_44228_n7040), .Y(u2__abc_44228_n14806) );
  OR2X2 OR2X2_3406 ( .A(u2__abc_44228_n14809), .B(u2__abc_44228_n8209_bF_buf7), .Y(u2__abc_44228_n14810) );
  OR2X2 OR2X2_3407 ( .A(u2__abc_44228_n14808_1), .B(u2__abc_44228_n14810), .Y(u2__abc_44228_n14811) );
  OR2X2 OR2X2_3408 ( .A(u2__abc_44228_n14815), .B(u2__abc_44228_n14801), .Y(u2__abc_44228_n14816_1) );
  OR2X2 OR2X2_3409 ( .A(u2__abc_44228_n14819), .B(u2__abc_44228_n8209_bF_buf6), .Y(u2__abc_44228_n14820) );
  OR2X2 OR2X2_341 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[58] ), .Y(_abc_64468_n1342) );
  OR2X2 OR2X2_3410 ( .A(u2__abc_44228_n14822), .B(u2__abc_44228_n14821), .Y(u2__abc_44228_n14823) );
  OR2X2 OR2X2_3411 ( .A(u2__abc_44228_n14824), .B(u2__abc_44228_n7034), .Y(u2__abc_44228_n14825_1) );
  OR2X2 OR2X2_3412 ( .A(u2__abc_44228_n14827), .B(u2__abc_44228_n14820), .Y(u2__abc_44228_n14828) );
  OR2X2 OR2X2_3413 ( .A(u2__abc_44228_n14832), .B(u2__abc_44228_n14818), .Y(u2__abc_44228_n14833_1) );
  OR2X2 OR2X2_3414 ( .A(u2__abc_44228_n14836), .B(u2__abc_44228_n7447_1), .Y(u2__abc_44228_n14837) );
  OR2X2 OR2X2_3415 ( .A(u2__abc_44228_n14837), .B(u2__abc_44228_n7026), .Y(u2__abc_44228_n14840) );
  OR2X2 OR2X2_3416 ( .A(u2__abc_44228_n14843_1), .B(u2__abc_44228_n8209_bF_buf5), .Y(u2__abc_44228_n14844) );
  OR2X2 OR2X2_3417 ( .A(u2__abc_44228_n14842), .B(u2__abc_44228_n14844), .Y(u2__abc_44228_n14845) );
  OR2X2 OR2X2_3418 ( .A(u2__abc_44228_n14849), .B(u2__abc_44228_n14835), .Y(u2__abc_44228_n14850) );
  OR2X2 OR2X2_3419 ( .A(u2__abc_44228_n14854), .B(u2__abc_44228_n14853), .Y(u2__abc_44228_n14855) );
  OR2X2 OR2X2_342 ( .A(a_112_bF_buf9), .B(\a[58] ), .Y(_abc_64468_n1344) );
  OR2X2 OR2X2_3420 ( .A(u2__abc_44228_n14856), .B(u2__abc_44228_n7020), .Y(u2__abc_44228_n14857) );
  OR2X2 OR2X2_3421 ( .A(u2__abc_44228_n14860_1), .B(u2__abc_44228_n2983_bF_buf90), .Y(u2__abc_44228_n14861) );
  OR2X2 OR2X2_3422 ( .A(u2__abc_44228_n14859), .B(u2__abc_44228_n14861), .Y(u2__abc_44228_n14862) );
  OR2X2 OR2X2_3423 ( .A(u2__abc_44228_n14866), .B(u2__abc_44228_n14852), .Y(u2__abc_44228_n14867) );
  OR2X2 OR2X2_3424 ( .A(u2__abc_44228_n14870), .B(u2__abc_44228_n7018), .Y(u2__abc_44228_n14871) );
  OR2X2 OR2X2_3425 ( .A(u2__abc_44228_n14872), .B(u2__abc_44228_n7011), .Y(u2__abc_44228_n14875) );
  OR2X2 OR2X2_3426 ( .A(u2__abc_44228_n14878), .B(u2__abc_44228_n2983_bF_buf88), .Y(u2__abc_44228_n14879) );
  OR2X2 OR2X2_3427 ( .A(u2__abc_44228_n14877), .B(u2__abc_44228_n14879), .Y(u2__abc_44228_n14880) );
  OR2X2 OR2X2_3428 ( .A(u2__abc_44228_n14884), .B(u2__abc_44228_n14869), .Y(u2__abc_44228_n14885) );
  OR2X2 OR2X2_3429 ( .A(u2__abc_44228_n14892), .B(u2__abc_44228_n14889), .Y(u2__abc_44228_n14893) );
  OR2X2 OR2X2_343 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[59] ), .Y(_abc_64468_n1345) );
  OR2X2 OR2X2_3430 ( .A(u2__abc_44228_n14895), .B(u2__abc_44228_n2983_bF_buf86), .Y(u2__abc_44228_n14896) );
  OR2X2 OR2X2_3431 ( .A(u2__abc_44228_n14894), .B(u2__abc_44228_n14896), .Y(u2__abc_44228_n14897) );
  OR2X2 OR2X2_3432 ( .A(u2__abc_44228_n14901), .B(u2__abc_44228_n14887), .Y(u2__abc_44228_n14902) );
  OR2X2 OR2X2_3433 ( .A(u2__abc_44228_n14905), .B(u2__abc_44228_n7003), .Y(u2__abc_44228_n14906) );
  OR2X2 OR2X2_3434 ( .A(u2__abc_44228_n14907), .B(u2__abc_44228_n6997_1), .Y(u2__abc_44228_n14910) );
  OR2X2 OR2X2_3435 ( .A(u2__abc_44228_n14913), .B(u2__abc_44228_n2983_bF_buf84), .Y(u2__abc_44228_n14914) );
  OR2X2 OR2X2_3436 ( .A(u2__abc_44228_n14912), .B(u2__abc_44228_n14914), .Y(u2__abc_44228_n14915) );
  OR2X2 OR2X2_3437 ( .A(u2__abc_44228_n14919), .B(u2__abc_44228_n14904), .Y(u2__abc_44228_n14920) );
  OR2X2 OR2X2_3438 ( .A(u2__abc_44228_n14908_1), .B(u2__abc_44228_n6993), .Y(u2__abc_44228_n14924) );
  OR2X2 OR2X2_3439 ( .A(u2__abc_44228_n14925), .B(u2__abc_44228_n14923), .Y(u2__abc_44228_n14926_1) );
  OR2X2 OR2X2_344 ( .A(a_112_bF_buf8), .B(\a[59] ), .Y(_abc_64468_n1347) );
  OR2X2 OR2X2_3440 ( .A(u2__abc_44228_n14924), .B(u2__abc_44228_n6991), .Y(u2__abc_44228_n14927) );
  OR2X2 OR2X2_3441 ( .A(u2__abc_44228_n14930), .B(u2__abc_44228_n2983_bF_buf82), .Y(u2__abc_44228_n14931) );
  OR2X2 OR2X2_3442 ( .A(u2__abc_44228_n14929), .B(u2__abc_44228_n14931), .Y(u2__abc_44228_n14932) );
  OR2X2 OR2X2_3443 ( .A(u2__abc_44228_n14936), .B(u2__abc_44228_n14922), .Y(u2__abc_44228_n14937) );
  OR2X2 OR2X2_3444 ( .A(u2__abc_44228_n14940), .B(u2__abc_44228_n7464_1), .Y(u2__abc_44228_n14941) );
  OR2X2 OR2X2_3445 ( .A(u2__abc_44228_n14941), .B(u2__abc_44228_n6966), .Y(u2__abc_44228_n14942) );
  OR2X2 OR2X2_3446 ( .A(u2__abc_44228_n14947), .B(u2__abc_44228_n8209_bF_buf4), .Y(u2__abc_44228_n14948) );
  OR2X2 OR2X2_3447 ( .A(u2__abc_44228_n14946), .B(u2__abc_44228_n14948), .Y(u2__abc_44228_n14949) );
  OR2X2 OR2X2_3448 ( .A(u2__abc_44228_n14953), .B(u2__abc_44228_n14939), .Y(u2__abc_44228_n14954_1) );
  OR2X2 OR2X2_3449 ( .A(u2__abc_44228_n14958), .B(u2__abc_44228_n14957), .Y(u2__abc_44228_n14959) );
  OR2X2 OR2X2_345 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[60] ), .Y(_abc_64468_n1348) );
  OR2X2 OR2X2_3450 ( .A(u2__abc_44228_n14960), .B(u2__abc_44228_n6960), .Y(u2__abc_44228_n14961) );
  OR2X2 OR2X2_3451 ( .A(u2__abc_44228_n14964), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n14965) );
  OR2X2 OR2X2_3452 ( .A(u2__abc_44228_n14963), .B(u2__abc_44228_n14965), .Y(u2__abc_44228_n14966) );
  OR2X2 OR2X2_3453 ( .A(u2__abc_44228_n14970), .B(u2__abc_44228_n14956), .Y(u2__abc_44228_n14971_1) );
  OR2X2 OR2X2_3454 ( .A(u2__abc_44228_n14974), .B(u2__abc_44228_n7469), .Y(u2__abc_44228_n14975) );
  OR2X2 OR2X2_3455 ( .A(u2__abc_44228_n14975), .B(u2__abc_44228_n6980), .Y(u2__abc_44228_n14978) );
  OR2X2 OR2X2_3456 ( .A(u2__abc_44228_n14981), .B(u2__abc_44228_n8209_bF_buf3), .Y(u2__abc_44228_n14982) );
  OR2X2 OR2X2_3457 ( .A(u2__abc_44228_n14980), .B(u2__abc_44228_n14982), .Y(u2__abc_44228_n14983) );
  OR2X2 OR2X2_3458 ( .A(u2__abc_44228_n14987), .B(u2__abc_44228_n14973), .Y(u2__abc_44228_n14988) );
  OR2X2 OR2X2_3459 ( .A(u2__abc_44228_n14992), .B(u2__abc_44228_n14991), .Y(u2__abc_44228_n14993) );
  OR2X2 OR2X2_346 ( .A(a_112_bF_buf7), .B(\a[60] ), .Y(_abc_64468_n1350) );
  OR2X2 OR2X2_3460 ( .A(u2__abc_44228_n14994), .B(u2__abc_44228_n6974), .Y(u2__abc_44228_n14995) );
  OR2X2 OR2X2_3461 ( .A(u2__abc_44228_n14998), .B(u2__abc_44228_n2983_bF_buf76), .Y(u2__abc_44228_n14999) );
  OR2X2 OR2X2_3462 ( .A(u2__abc_44228_n14997_1), .B(u2__abc_44228_n14999), .Y(u2__abc_44228_n15000) );
  OR2X2 OR2X2_3463 ( .A(u2__abc_44228_n15004), .B(u2__abc_44228_n14990), .Y(u2__abc_44228_n15005) );
  OR2X2 OR2X2_3464 ( .A(u2__abc_44228_n15008), .B(u2__abc_44228_n6972), .Y(u2__abc_44228_n15009) );
  OR2X2 OR2X2_3465 ( .A(u2__abc_44228_n15010), .B(u2__abc_44228_n6944), .Y(u2__abc_44228_n15011) );
  OR2X2 OR2X2_3466 ( .A(u2__abc_44228_n15016), .B(u2__abc_44228_n8209_bF_buf2), .Y(u2__abc_44228_n15017) );
  OR2X2 OR2X2_3467 ( .A(u2__abc_44228_n15015), .B(u2__abc_44228_n15017), .Y(u2__abc_44228_n15018) );
  OR2X2 OR2X2_3468 ( .A(u2__abc_44228_n15022), .B(u2__abc_44228_n15007), .Y(u2__abc_44228_n15023) );
  OR2X2 OR2X2_3469 ( .A(u2__abc_44228_n15027), .B(u2__abc_44228_n6951), .Y(u2__abc_44228_n15028) );
  OR2X2 OR2X2_347 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[61] ), .Y(_abc_64468_n1351) );
  OR2X2 OR2X2_3470 ( .A(u2__abc_44228_n15026_1), .B(u2__abc_44228_n15029), .Y(u2__abc_44228_n15030) );
  OR2X2 OR2X2_3471 ( .A(u2__abc_44228_n15033), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n15034_1) );
  OR2X2 OR2X2_3472 ( .A(u2__abc_44228_n15032), .B(u2__abc_44228_n15034_1), .Y(u2__abc_44228_n15035) );
  OR2X2 OR2X2_3473 ( .A(u2__abc_44228_n15039), .B(u2__abc_44228_n15025), .Y(u2__abc_44228_n15040) );
  OR2X2 OR2X2_3474 ( .A(u2__abc_44228_n15043_1), .B(u2__abc_44228_n6949), .Y(u2__abc_44228_n15044) );
  OR2X2 OR2X2_3475 ( .A(u2__abc_44228_n15045), .B(u2__abc_44228_n6937), .Y(u2__abc_44228_n15048) );
  OR2X2 OR2X2_3476 ( .A(u2__abc_44228_n15051_1), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n15052) );
  OR2X2 OR2X2_3477 ( .A(u2__abc_44228_n15050), .B(u2__abc_44228_n15052), .Y(u2__abc_44228_n15053) );
  OR2X2 OR2X2_3478 ( .A(u2__abc_44228_n15057), .B(u2__abc_44228_n15042), .Y(u2__abc_44228_n15058) );
  OR2X2 OR2X2_3479 ( .A(u2__abc_44228_n15046), .B(u2__abc_44228_n6933), .Y(u2__abc_44228_n15062) );
  OR2X2 OR2X2_348 ( .A(a_112_bF_buf6), .B(\a[61] ), .Y(_abc_64468_n1353) );
  OR2X2 OR2X2_3480 ( .A(u2__abc_44228_n15063), .B(u2__abc_44228_n15061_1), .Y(u2__abc_44228_n15064) );
  OR2X2 OR2X2_3481 ( .A(u2__abc_44228_n15062), .B(u2__abc_44228_n6931), .Y(u2__abc_44228_n15065) );
  OR2X2 OR2X2_3482 ( .A(u2__abc_44228_n15068), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n15069_1) );
  OR2X2 OR2X2_3483 ( .A(u2__abc_44228_n15067), .B(u2__abc_44228_n15069_1), .Y(u2__abc_44228_n15070) );
  OR2X2 OR2X2_3484 ( .A(u2__abc_44228_n15074), .B(u2__abc_44228_n15060), .Y(u2__abc_44228_n15075) );
  OR2X2 OR2X2_3485 ( .A(u2__abc_44228_n15078_1), .B(u2__abc_44228_n7485), .Y(u2__abc_44228_n15079) );
  OR2X2 OR2X2_3486 ( .A(u2__abc_44228_n15079), .B(u2__abc_44228_n6921), .Y(u2__abc_44228_n15082) );
  OR2X2 OR2X2_3487 ( .A(u2__abc_44228_n15085), .B(u2__abc_44228_n8209_bF_buf1), .Y(u2__abc_44228_n15086_1) );
  OR2X2 OR2X2_3488 ( .A(u2__abc_44228_n15084), .B(u2__abc_44228_n15086_1), .Y(u2__abc_44228_n15087) );
  OR2X2 OR2X2_3489 ( .A(u2__abc_44228_n15091), .B(u2__abc_44228_n15077), .Y(u2__abc_44228_n15092) );
  OR2X2 OR2X2_349 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[62] ), .Y(_abc_64468_n1354) );
  OR2X2 OR2X2_3490 ( .A(u2__abc_44228_n15099), .B(u2__abc_44228_n15096), .Y(u2__abc_44228_n15100) );
  OR2X2 OR2X2_3491 ( .A(u2__abc_44228_n15102), .B(u2__abc_44228_n2983_bF_buf66), .Y(u2__abc_44228_n15103) );
  OR2X2 OR2X2_3492 ( .A(u2__abc_44228_n15101), .B(u2__abc_44228_n15103), .Y(u2__abc_44228_n15104) );
  OR2X2 OR2X2_3493 ( .A(u2__abc_44228_n15108), .B(u2__abc_44228_n15094), .Y(u2__abc_44228_n15109) );
  OR2X2 OR2X2_3494 ( .A(u2__abc_44228_n15112), .B(u2__abc_44228_n6913), .Y(u2__abc_44228_n15113) );
  OR2X2 OR2X2_3495 ( .A(u2__abc_44228_n15114_1), .B(u2__abc_44228_n6907), .Y(u2__abc_44228_n15117) );
  OR2X2 OR2X2_3496 ( .A(u2__abc_44228_n15120), .B(u2__abc_44228_n8209_bF_buf0), .Y(u2__abc_44228_n15121) );
  OR2X2 OR2X2_3497 ( .A(u2__abc_44228_n15119), .B(u2__abc_44228_n15121), .Y(u2__abc_44228_n15122_1) );
  OR2X2 OR2X2_3498 ( .A(u2__abc_44228_n15126), .B(u2__abc_44228_n15111), .Y(u2__abc_44228_n15127) );
  OR2X2 OR2X2_3499 ( .A(u2__abc_44228_n15115), .B(u2__abc_44228_n6903), .Y(u2__abc_44228_n15131) );
  OR2X2 OR2X2_35 ( .A(aNan_bF_buf3), .B(sqrto_93_), .Y(_abc_64468_n881) );
  OR2X2 OR2X2_350 ( .A(a_112_bF_buf5), .B(\a[62] ), .Y(_abc_64468_n1356) );
  OR2X2 OR2X2_3500 ( .A(u2__abc_44228_n15132_1), .B(u2__abc_44228_n15130), .Y(u2__abc_44228_n15133) );
  OR2X2 OR2X2_3501 ( .A(u2__abc_44228_n15131), .B(u2__abc_44228_n6901), .Y(u2__abc_44228_n15134) );
  OR2X2 OR2X2_3502 ( .A(u2__abc_44228_n15137), .B(u2__abc_44228_n2983_bF_buf63), .Y(u2__abc_44228_n15138) );
  OR2X2 OR2X2_3503 ( .A(u2__abc_44228_n15136), .B(u2__abc_44228_n15138), .Y(u2__abc_44228_n15139) );
  OR2X2 OR2X2_3504 ( .A(u2__abc_44228_n15143), .B(u2__abc_44228_n15129), .Y(u2__abc_44228_n15144) );
  OR2X2 OR2X2_3505 ( .A(u2__abc_44228_n15147), .B(u2__abc_44228_n7494), .Y(u2__abc_44228_n15148) );
  OR2X2 OR2X2_3506 ( .A(u2__abc_44228_n15148), .B(u2__abc_44228_n6892), .Y(u2__abc_44228_n15149_1) );
  OR2X2 OR2X2_3507 ( .A(u2__abc_44228_n15154), .B(u2__abc_44228_n8209_bF_buf9), .Y(u2__abc_44228_n15155) );
  OR2X2 OR2X2_3508 ( .A(u2__abc_44228_n15153), .B(u2__abc_44228_n15155), .Y(u2__abc_44228_n15156) );
  OR2X2 OR2X2_3509 ( .A(u2__abc_44228_n15160), .B(u2__abc_44228_n15146), .Y(u2__abc_44228_n15161) );
  OR2X2 OR2X2_351 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[63] ), .Y(_abc_64468_n1357) );
  OR2X2 OR2X2_3510 ( .A(u2__abc_44228_n15165), .B(u2__abc_44228_n15164), .Y(u2__abc_44228_n15166) );
  OR2X2 OR2X2_3511 ( .A(u2__abc_44228_n15167), .B(u2__abc_44228_n6886), .Y(u2__abc_44228_n15168) );
  OR2X2 OR2X2_3512 ( .A(u2__abc_44228_n15171), .B(u2__abc_44228_n2983_bF_buf60), .Y(u2__abc_44228_n15172) );
  OR2X2 OR2X2_3513 ( .A(u2__abc_44228_n15170_1), .B(u2__abc_44228_n15172), .Y(u2__abc_44228_n15173) );
  OR2X2 OR2X2_3514 ( .A(u2__abc_44228_n15177), .B(u2__abc_44228_n15163), .Y(u2__abc_44228_n15178_1) );
  OR2X2 OR2X2_3515 ( .A(u2__abc_44228_n15181), .B(u2__abc_44228_n7499), .Y(u2__abc_44228_n15182) );
  OR2X2 OR2X2_3516 ( .A(u2__abc_44228_n15182), .B(u2__abc_44228_n6878_1), .Y(u2__abc_44228_n15185) );
  OR2X2 OR2X2_3517 ( .A(u2__abc_44228_n15188), .B(u2__abc_44228_n2983_bF_buf58), .Y(u2__abc_44228_n15189) );
  OR2X2 OR2X2_3518 ( .A(u2__abc_44228_n15187_1), .B(u2__abc_44228_n15189), .Y(u2__abc_44228_n15190) );
  OR2X2 OR2X2_3519 ( .A(u2__abc_44228_n15194), .B(u2__abc_44228_n15180), .Y(u2__abc_44228_n15195_1) );
  OR2X2 OR2X2_352 ( .A(a_112_bF_buf4), .B(\a[63] ), .Y(_abc_64468_n1359) );
  OR2X2 OR2X2_3520 ( .A(u2__abc_44228_n15183), .B(u2__abc_44228_n6874), .Y(u2__abc_44228_n15199) );
  OR2X2 OR2X2_3521 ( .A(u2__abc_44228_n15200), .B(u2__abc_44228_n15198), .Y(u2__abc_44228_n15201) );
  OR2X2 OR2X2_3522 ( .A(u2__abc_44228_n15199), .B(u2__abc_44228_n6872), .Y(u2__abc_44228_n15202) );
  OR2X2 OR2X2_3523 ( .A(u2__abc_44228_n15205_1), .B(u2__abc_44228_n2983_bF_buf56), .Y(u2__abc_44228_n15206) );
  OR2X2 OR2X2_3524 ( .A(u2__abc_44228_n15204), .B(u2__abc_44228_n15206), .Y(u2__abc_44228_n15207) );
  OR2X2 OR2X2_3525 ( .A(u2__abc_44228_n15211), .B(u2__abc_44228_n15197), .Y(u2__abc_44228_n15212) );
  OR2X2 OR2X2_3526 ( .A(u2__abc_44228_n7508), .B(u2__abc_44228_n7528), .Y(u2__abc_44228_n15215) );
  OR2X2 OR2X2_3527 ( .A(u2__abc_44228_n7548_1_bF_buf15), .B(u2__abc_44228_n15218), .Y(u2__abc_44228_n15219) );
  OR2X2 OR2X2_3528 ( .A(u2__abc_44228_n7547_bF_buf14), .B(u2_remHi_446_), .Y(u2__abc_44228_n15220) );
  OR2X2 OR2X2_3529 ( .A(u2__abc_44228_n15221), .B(u2__abc_44228_n2983_bF_buf54), .Y(u2__abc_44228_n15222_1) );
  OR2X2 OR2X2_353 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[64] ), .Y(_abc_64468_n1360) );
  OR2X2 OR2X2_3530 ( .A(u2__abc_44228_n15226), .B(u2__abc_44228_n15214), .Y(u2__abc_44228_n15227) );
  OR2X2 OR2X2_3531 ( .A(u2__abc_44228_n15231), .B(u2__abc_44228_n15230_1), .Y(u2__abc_44228_n15232) );
  OR2X2 OR2X2_3532 ( .A(u2__abc_44228_n15233), .B(u2__abc_44228_n7535), .Y(u2__abc_44228_n15234) );
  OR2X2 OR2X2_3533 ( .A(u2__abc_44228_n15237), .B(u2__abc_44228_n2983_bF_buf52), .Y(u2__abc_44228_n15238) );
  OR2X2 OR2X2_3534 ( .A(u2__abc_44228_n15236), .B(u2__abc_44228_n15238), .Y(u2__abc_44228_n15239) );
  OR2X2 OR2X2_3535 ( .A(u2__abc_44228_n15243), .B(u2__abc_44228_n15229), .Y(u2__abc_44228_n15244) );
  OR2X2 OR2X2_3536 ( .A(u2__abc_44228_n15246), .B(u2__abc_44228_n3062_bF_buf14), .Y(u2__abc_44228_n15247) );
  OR2X2 OR2X2_3537 ( .A(u2__abc_44228_n15252), .B(u2__abc_44228_n15254), .Y(u2__abc_44228_n15255) );
  OR2X2 OR2X2_3538 ( .A(u2__abc_44228_n15257), .B(u2__abc_44228_n15259), .Y(u2__abc_44228_n15260) );
  OR2X2 OR2X2_3539 ( .A(u2__abc_44228_n15262), .B(u2__abc_44228_n15264), .Y(u2__abc_44228_n15265) );
  OR2X2 OR2X2_354 ( .A(a_112_bF_buf3), .B(\a[64] ), .Y(_abc_64468_n1362) );
  OR2X2 OR2X2_3540 ( .A(u2__abc_44228_n15267), .B(u2__abc_44228_n15269), .Y(u2__abc_44228_n15270) );
  OR2X2 OR2X2_3541 ( .A(u2__abc_44228_n15272), .B(u2__abc_44228_n15274), .Y(u2__abc_44228_n15275) );
  OR2X2 OR2X2_3542 ( .A(u2__abc_44228_n15277), .B(u2__abc_44228_n15279), .Y(u2__abc_44228_n15280) );
  OR2X2 OR2X2_3543 ( .A(u2__abc_44228_n15282), .B(u2__abc_44228_n15284_1), .Y(u2__abc_44228_n15285) );
  OR2X2 OR2X2_3544 ( .A(u2__abc_44228_n15287), .B(u2__abc_44228_n15289), .Y(u2__abc_44228_n15290) );
  OR2X2 OR2X2_3545 ( .A(u2__abc_44228_n15292), .B(u2__abc_44228_n15294), .Y(u2__abc_44228_n15295) );
  OR2X2 OR2X2_3546 ( .A(u2__abc_44228_n15297), .B(u2__abc_44228_n15299), .Y(u2__abc_44228_n15300) );
  OR2X2 OR2X2_3547 ( .A(u2__abc_44228_n15302), .B(u2__abc_44228_n15304), .Y(u2__abc_44228_n15305) );
  OR2X2 OR2X2_3548 ( .A(u2__abc_44228_n15307), .B(u2__abc_44228_n15309), .Y(u2__abc_44228_n15310) );
  OR2X2 OR2X2_3549 ( .A(u2__abc_44228_n15312), .B(u2__abc_44228_n15314), .Y(u2__abc_44228_n15315) );
  OR2X2 OR2X2_355 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[65] ), .Y(_abc_64468_n1363) );
  OR2X2 OR2X2_3550 ( .A(u2__abc_44228_n15317), .B(u2__abc_44228_n15319), .Y(u2__abc_44228_n15320) );
  OR2X2 OR2X2_3551 ( .A(u2__abc_44228_n15322), .B(u2__abc_44228_n15324), .Y(u2__abc_44228_n15325) );
  OR2X2 OR2X2_3552 ( .A(u2__abc_44228_n15327), .B(u2__abc_44228_n15329), .Y(u2__abc_44228_n15330_1) );
  OR2X2 OR2X2_3553 ( .A(u2__abc_44228_n15332), .B(u2__abc_44228_n15334), .Y(u2__abc_44228_n15335) );
  OR2X2 OR2X2_3554 ( .A(u2__abc_44228_n15337), .B(u2__abc_44228_n15339), .Y(u2__abc_44228_n15340) );
  OR2X2 OR2X2_3555 ( .A(u2__abc_44228_n15342), .B(u2__abc_44228_n15344), .Y(u2__abc_44228_n15345) );
  OR2X2 OR2X2_3556 ( .A(u2__abc_44228_n15347), .B(u2__abc_44228_n15349), .Y(u2__abc_44228_n15350) );
  OR2X2 OR2X2_3557 ( .A(u2__abc_44228_n15352), .B(u2__abc_44228_n15354), .Y(u2__abc_44228_n15355) );
  OR2X2 OR2X2_3558 ( .A(u2__abc_44228_n15357), .B(u2__abc_44228_n15359), .Y(u2__abc_44228_n15360) );
  OR2X2 OR2X2_3559 ( .A(u2__abc_44228_n15362), .B(u2__abc_44228_n15364), .Y(u2__abc_44228_n15365_1) );
  OR2X2 OR2X2_356 ( .A(a_112_bF_buf2), .B(\a[65] ), .Y(_abc_64468_n1365) );
  OR2X2 OR2X2_3560 ( .A(u2__abc_44228_n15367), .B(u2__abc_44228_n15369), .Y(u2__abc_44228_n15370) );
  OR2X2 OR2X2_3561 ( .A(u2__abc_44228_n15372), .B(u2__abc_44228_n15374), .Y(u2__abc_44228_n15375) );
  OR2X2 OR2X2_3562 ( .A(u2__abc_44228_n15377), .B(u2__abc_44228_n15379), .Y(u2__abc_44228_n15380) );
  OR2X2 OR2X2_3563 ( .A(u2__abc_44228_n15382), .B(u2__abc_44228_n15384_1), .Y(u2__abc_44228_n15385) );
  OR2X2 OR2X2_3564 ( .A(u2__abc_44228_n15387), .B(u2__abc_44228_n15389), .Y(u2__abc_44228_n15390) );
  OR2X2 OR2X2_3565 ( .A(u2__abc_44228_n15392_1), .B(u2__abc_44228_n15394), .Y(u2__abc_44228_n15395) );
  OR2X2 OR2X2_3566 ( .A(u2__abc_44228_n15397), .B(u2__abc_44228_n15399), .Y(u2__abc_44228_n15400) );
  OR2X2 OR2X2_3567 ( .A(u2__abc_44228_n15246), .B(u2__abc_44228_n2963), .Y(u2__abc_44228_n15403) );
  OR2X2 OR2X2_3568 ( .A(u2__abc_44228_n15404), .B(u2__abc_44228_n15402_bF_buf3), .Y(u2__abc_44228_n15405) );
  OR2X2 OR2X2_3569 ( .A(u2__abc_44228_n15409_1), .B(u2__abc_44228_n15407), .Y(u2__abc_44228_n15410) );
  OR2X2 OR2X2_357 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[66] ), .Y(_abc_64468_n1366) );
  OR2X2 OR2X2_3570 ( .A(u2__abc_44228_n15406), .B(u2__abc_44228_n15411), .Y(u2_remLo_32__FF_INPUT) );
  OR2X2 OR2X2_3571 ( .A(u2__abc_44228_n15415), .B(u2__abc_44228_n15414), .Y(u2__abc_44228_n15416) );
  OR2X2 OR2X2_3572 ( .A(u2__abc_44228_n15413), .B(u2__abc_44228_n15417), .Y(u2_remLo_33__FF_INPUT) );
  OR2X2 OR2X2_3573 ( .A(u2__abc_44228_n15421), .B(u2__abc_44228_n15420), .Y(u2__abc_44228_n15422) );
  OR2X2 OR2X2_3574 ( .A(u2__abc_44228_n15419_1), .B(u2__abc_44228_n15423), .Y(u2_remLo_34__FF_INPUT) );
  OR2X2 OR2X2_3575 ( .A(u2__abc_44228_n15426), .B(u2__abc_44228_n15427_1), .Y(u2__abc_44228_n15428) );
  OR2X2 OR2X2_3576 ( .A(u2__abc_44228_n15425), .B(u2__abc_44228_n15429), .Y(u2_remLo_35__FF_INPUT) );
  OR2X2 OR2X2_3577 ( .A(u2__abc_44228_n15431), .B(u2__abc_44228_n15432), .Y(u2__abc_44228_n15433) );
  OR2X2 OR2X2_3578 ( .A(u2__abc_44228_n15435_1), .B(u2__abc_44228_n15436), .Y(u2__abc_44228_n15437) );
  OR2X2 OR2X2_3579 ( .A(u2__abc_44228_n15434), .B(u2__abc_44228_n15437), .Y(u2_remLo_36__FF_INPUT) );
  OR2X2 OR2X2_358 ( .A(a_112_bF_buf1), .B(\a[66] ), .Y(_abc_64468_n1368) );
  OR2X2 OR2X2_3580 ( .A(u2__abc_44228_n15440), .B(u2__abc_44228_n15441), .Y(u2__abc_44228_n15442_1) );
  OR2X2 OR2X2_3581 ( .A(u2__abc_44228_n15439), .B(u2__abc_44228_n15443), .Y(u2_remLo_37__FF_INPUT) );
  OR2X2 OR2X2_3582 ( .A(u2__abc_44228_n15446), .B(u2__abc_44228_n15447), .Y(u2__abc_44228_n15448) );
  OR2X2 OR2X2_3583 ( .A(u2__abc_44228_n15445), .B(u2__abc_44228_n15449), .Y(u2_remLo_38__FF_INPUT) );
  OR2X2 OR2X2_3584 ( .A(u2__abc_44228_n15452), .B(u2__abc_44228_n15453), .Y(u2__abc_44228_n15454) );
  OR2X2 OR2X2_3585 ( .A(u2__abc_44228_n15451), .B(u2__abc_44228_n15455_1), .Y(u2_remLo_39__FF_INPUT) );
  OR2X2 OR2X2_3586 ( .A(u2__abc_44228_n15459), .B(u2__abc_44228_n15458), .Y(u2__abc_44228_n15460) );
  OR2X2 OR2X2_3587 ( .A(u2__abc_44228_n15457), .B(u2__abc_44228_n15461), .Y(u2_remLo_40__FF_INPUT) );
  OR2X2 OR2X2_3588 ( .A(u2__abc_44228_n15464), .B(u2__abc_44228_n15465), .Y(u2__abc_44228_n15466) );
  OR2X2 OR2X2_3589 ( .A(u2__abc_44228_n15463_1), .B(u2__abc_44228_n15467), .Y(u2_remLo_41__FF_INPUT) );
  OR2X2 OR2X2_359 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[67] ), .Y(_abc_64468_n1369) );
  OR2X2 OR2X2_3590 ( .A(u2__abc_44228_n15471), .B(u2__abc_44228_n15470), .Y(u2__abc_44228_n15472_1) );
  OR2X2 OR2X2_3591 ( .A(u2__abc_44228_n15469), .B(u2__abc_44228_n15473_1), .Y(u2_remLo_42__FF_INPUT) );
  OR2X2 OR2X2_3592 ( .A(u2__abc_44228_n15476), .B(u2__abc_44228_n15477), .Y(u2__abc_44228_n15478) );
  OR2X2 OR2X2_3593 ( .A(u2__abc_44228_n15475), .B(u2__abc_44228_n15479), .Y(u2_remLo_43__FF_INPUT) );
  OR2X2 OR2X2_3594 ( .A(u2__abc_44228_n15482), .B(u2__abc_44228_n15483), .Y(u2__abc_44228_n15484) );
  OR2X2 OR2X2_3595 ( .A(u2__abc_44228_n15481_1), .B(u2__abc_44228_n15485), .Y(u2_remLo_44__FF_INPUT) );
  OR2X2 OR2X2_3596 ( .A(u2__abc_44228_n15488), .B(u2__abc_44228_n15489), .Y(u2__abc_44228_n15490) );
  OR2X2 OR2X2_3597 ( .A(u2__abc_44228_n15487), .B(u2__abc_44228_n15491), .Y(u2_remLo_45__FF_INPUT) );
  OR2X2 OR2X2_3598 ( .A(u2__abc_44228_n15494), .B(u2__abc_44228_n15495), .Y(u2__abc_44228_n15496) );
  OR2X2 OR2X2_3599 ( .A(u2__abc_44228_n15493), .B(u2__abc_44228_n15497), .Y(u2_remLo_46__FF_INPUT) );
  OR2X2 OR2X2_36 ( .A(_abc_64468_n753_bF_buf4), .B(\a[17] ), .Y(_abc_64468_n882) );
  OR2X2 OR2X2_360 ( .A(a_112_bF_buf0), .B(\a[67] ), .Y(_abc_64468_n1371) );
  OR2X2 OR2X2_3600 ( .A(u2__abc_44228_n15501), .B(u2__abc_44228_n15500), .Y(u2__abc_44228_n15502) );
  OR2X2 OR2X2_3601 ( .A(u2__abc_44228_n15499), .B(u2__abc_44228_n15503), .Y(u2_remLo_47__FF_INPUT) );
  OR2X2 OR2X2_3602 ( .A(u2__abc_44228_n15506), .B(u2__abc_44228_n15507), .Y(u2__abc_44228_n15508) );
  OR2X2 OR2X2_3603 ( .A(u2__abc_44228_n15505), .B(u2__abc_44228_n15509), .Y(u2_remLo_48__FF_INPUT) );
  OR2X2 OR2X2_3604 ( .A(u2__abc_44228_n15512), .B(u2__abc_44228_n15513), .Y(u2__abc_44228_n15514) );
  OR2X2 OR2X2_3605 ( .A(u2__abc_44228_n15511), .B(u2__abc_44228_n15515), .Y(u2_remLo_49__FF_INPUT) );
  OR2X2 OR2X2_3606 ( .A(u2__abc_44228_n15519), .B(u2__abc_44228_n15518), .Y(u2__abc_44228_n15520) );
  OR2X2 OR2X2_3607 ( .A(u2__abc_44228_n15517), .B(u2__abc_44228_n15521), .Y(u2_remLo_50__FF_INPUT) );
  OR2X2 OR2X2_3608 ( .A(u2__abc_44228_n15525), .B(u2__abc_44228_n15524), .Y(u2__abc_44228_n15526) );
  OR2X2 OR2X2_3609 ( .A(u2__abc_44228_n15523), .B(u2__abc_44228_n15527), .Y(u2_remLo_51__FF_INPUT) );
  OR2X2 OR2X2_361 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[68] ), .Y(_abc_64468_n1372) );
  OR2X2 OR2X2_3610 ( .A(u2__abc_44228_n15531), .B(u2__abc_44228_n15530), .Y(u2__abc_44228_n15532) );
  OR2X2 OR2X2_3611 ( .A(u2__abc_44228_n15529), .B(u2__abc_44228_n15533), .Y(u2_remLo_52__FF_INPUT) );
  OR2X2 OR2X2_3612 ( .A(u2__abc_44228_n15536), .B(u2__abc_44228_n15537), .Y(u2__abc_44228_n15538) );
  OR2X2 OR2X2_3613 ( .A(u2__abc_44228_n15535), .B(u2__abc_44228_n15539), .Y(u2_remLo_53__FF_INPUT) );
  OR2X2 OR2X2_3614 ( .A(u2__abc_44228_n15542), .B(u2__abc_44228_n15541), .Y(u2__abc_44228_n15543) );
  OR2X2 OR2X2_3615 ( .A(u2__abc_44228_n15545), .B(u2__abc_44228_n15546), .Y(u2__abc_44228_n15547) );
  OR2X2 OR2X2_3616 ( .A(u2__abc_44228_n15544), .B(u2__abc_44228_n15547), .Y(u2_remLo_54__FF_INPUT) );
  OR2X2 OR2X2_3617 ( .A(u2__abc_44228_n15550), .B(u2__abc_44228_n15551), .Y(u2__abc_44228_n15552) );
  OR2X2 OR2X2_3618 ( .A(u2__abc_44228_n15549), .B(u2__abc_44228_n15553), .Y(u2_remLo_55__FF_INPUT) );
  OR2X2 OR2X2_3619 ( .A(u2__abc_44228_n15556), .B(u2__abc_44228_n15557), .Y(u2__abc_44228_n15558) );
  OR2X2 OR2X2_362 ( .A(a_112_bF_buf9), .B(\a[68] ), .Y(_abc_64468_n1374) );
  OR2X2 OR2X2_3620 ( .A(u2__abc_44228_n15555), .B(u2__abc_44228_n15559), .Y(u2_remLo_56__FF_INPUT) );
  OR2X2 OR2X2_3621 ( .A(u2__abc_44228_n15562), .B(u2__abc_44228_n15563), .Y(u2__abc_44228_n15564) );
  OR2X2 OR2X2_3622 ( .A(u2__abc_44228_n15561), .B(u2__abc_44228_n15565), .Y(u2_remLo_57__FF_INPUT) );
  OR2X2 OR2X2_3623 ( .A(u2__abc_44228_n15569), .B(u2__abc_44228_n15568), .Y(u2__abc_44228_n15570) );
  OR2X2 OR2X2_3624 ( .A(u2__abc_44228_n15567), .B(u2__abc_44228_n15571), .Y(u2_remLo_58__FF_INPUT) );
  OR2X2 OR2X2_3625 ( .A(u2__abc_44228_n15575), .B(u2__abc_44228_n15574), .Y(u2__abc_44228_n15576) );
  OR2X2 OR2X2_3626 ( .A(u2__abc_44228_n15573), .B(u2__abc_44228_n15577), .Y(u2_remLo_59__FF_INPUT) );
  OR2X2 OR2X2_3627 ( .A(u2__abc_44228_n15580), .B(u2__abc_44228_n15581), .Y(u2__abc_44228_n15582) );
  OR2X2 OR2X2_3628 ( .A(u2__abc_44228_n15579), .B(u2__abc_44228_n15583), .Y(u2_remLo_60__FF_INPUT) );
  OR2X2 OR2X2_3629 ( .A(u2__abc_44228_n15586), .B(u2__abc_44228_n15587), .Y(u2__abc_44228_n15588) );
  OR2X2 OR2X2_363 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[69] ), .Y(_abc_64468_n1375) );
  OR2X2 OR2X2_3630 ( .A(u2__abc_44228_n15585), .B(u2__abc_44228_n15589), .Y(u2_remLo_61__FF_INPUT) );
  OR2X2 OR2X2_3631 ( .A(u2__abc_44228_n15593), .B(u2__abc_44228_n15592), .Y(u2__abc_44228_n15594) );
  OR2X2 OR2X2_3632 ( .A(u2__abc_44228_n15591), .B(u2__abc_44228_n15595), .Y(u2_remLo_62__FF_INPUT) );
  OR2X2 OR2X2_3633 ( .A(u2__abc_44228_n15599), .B(u2__abc_44228_n15598), .Y(u2__abc_44228_n15600) );
  OR2X2 OR2X2_3634 ( .A(u2__abc_44228_n15597), .B(u2__abc_44228_n15601), .Y(u2_remLo_63__FF_INPUT) );
  OR2X2 OR2X2_3635 ( .A(u2__abc_44228_n15604), .B(u2__abc_44228_n15605), .Y(u2__abc_44228_n15606) );
  OR2X2 OR2X2_3636 ( .A(u2__abc_44228_n15603), .B(u2__abc_44228_n15607), .Y(u2_remLo_64__FF_INPUT) );
  OR2X2 OR2X2_3637 ( .A(u2__abc_44228_n15611), .B(u2__abc_44228_n15610), .Y(u2__abc_44228_n15612) );
  OR2X2 OR2X2_3638 ( .A(u2__abc_44228_n15609), .B(u2__abc_44228_n15613), .Y(u2_remLo_65__FF_INPUT) );
  OR2X2 OR2X2_3639 ( .A(u2__abc_44228_n15616), .B(u2__abc_44228_n15617), .Y(u2__abc_44228_n15618) );
  OR2X2 OR2X2_364 ( .A(a_112_bF_buf8), .B(\a[69] ), .Y(_abc_64468_n1377) );
  OR2X2 OR2X2_3640 ( .A(u2__abc_44228_n15615), .B(u2__abc_44228_n15619), .Y(u2_remLo_66__FF_INPUT) );
  OR2X2 OR2X2_3641 ( .A(u2__abc_44228_n15622), .B(u2__abc_44228_n15623), .Y(u2__abc_44228_n15624) );
  OR2X2 OR2X2_3642 ( .A(u2__abc_44228_n15621), .B(u2__abc_44228_n15625), .Y(u2_remLo_67__FF_INPUT) );
  OR2X2 OR2X2_3643 ( .A(u2__abc_44228_n15629), .B(u2__abc_44228_n15628), .Y(u2__abc_44228_n15630) );
  OR2X2 OR2X2_3644 ( .A(u2__abc_44228_n15627), .B(u2__abc_44228_n15631), .Y(u2_remLo_68__FF_INPUT) );
  OR2X2 OR2X2_3645 ( .A(u2__abc_44228_n15634), .B(u2__abc_44228_n15635), .Y(u2__abc_44228_n15636) );
  OR2X2 OR2X2_3646 ( .A(u2__abc_44228_n15633), .B(u2__abc_44228_n15637), .Y(u2_remLo_69__FF_INPUT) );
  OR2X2 OR2X2_3647 ( .A(u2__abc_44228_n15640), .B(u2__abc_44228_n15641), .Y(u2__abc_44228_n15642) );
  OR2X2 OR2X2_3648 ( .A(u2__abc_44228_n15639), .B(u2__abc_44228_n15643), .Y(u2_remLo_70__FF_INPUT) );
  OR2X2 OR2X2_3649 ( .A(u2__abc_44228_n15646), .B(u2__abc_44228_n15647), .Y(u2__abc_44228_n15648) );
  OR2X2 OR2X2_365 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[70] ), .Y(_abc_64468_n1378) );
  OR2X2 OR2X2_3650 ( .A(u2__abc_44228_n15645), .B(u2__abc_44228_n15649), .Y(u2_remLo_71__FF_INPUT) );
  OR2X2 OR2X2_3651 ( .A(u2__abc_44228_n15652), .B(u2__abc_44228_n15653), .Y(u2__abc_44228_n15654) );
  OR2X2 OR2X2_3652 ( .A(u2__abc_44228_n15651), .B(u2__abc_44228_n15655), .Y(u2_remLo_72__FF_INPUT) );
  OR2X2 OR2X2_3653 ( .A(u2__abc_44228_n15658), .B(u2__abc_44228_n15659), .Y(u2__abc_44228_n15660) );
  OR2X2 OR2X2_3654 ( .A(u2__abc_44228_n15657), .B(u2__abc_44228_n15661), .Y(u2_remLo_73__FF_INPUT) );
  OR2X2 OR2X2_3655 ( .A(u2__abc_44228_n15665), .B(u2__abc_44228_n15664), .Y(u2__abc_44228_n15666) );
  OR2X2 OR2X2_3656 ( .A(u2__abc_44228_n15663), .B(u2__abc_44228_n15667), .Y(u2_remLo_74__FF_INPUT) );
  OR2X2 OR2X2_3657 ( .A(u2__abc_44228_n15670), .B(u2__abc_44228_n15671), .Y(u2__abc_44228_n15672) );
  OR2X2 OR2X2_3658 ( .A(u2__abc_44228_n15669), .B(u2__abc_44228_n15673), .Y(u2_remLo_75__FF_INPUT) );
  OR2X2 OR2X2_3659 ( .A(u2__abc_44228_n15676), .B(u2__abc_44228_n15677), .Y(u2__abc_44228_n15678) );
  OR2X2 OR2X2_366 ( .A(a_112_bF_buf7), .B(\a[70] ), .Y(_abc_64468_n1380) );
  OR2X2 OR2X2_3660 ( .A(u2__abc_44228_n15675), .B(u2__abc_44228_n15679), .Y(u2_remLo_76__FF_INPUT) );
  OR2X2 OR2X2_3661 ( .A(u2__abc_44228_n15682), .B(u2__abc_44228_n15683), .Y(u2__abc_44228_n15684) );
  OR2X2 OR2X2_3662 ( .A(u2__abc_44228_n15681), .B(u2__abc_44228_n15685), .Y(u2_remLo_77__FF_INPUT) );
  OR2X2 OR2X2_3663 ( .A(u2__abc_44228_n15689), .B(u2__abc_44228_n15688), .Y(u2__abc_44228_n15690) );
  OR2X2 OR2X2_3664 ( .A(u2__abc_44228_n15687), .B(u2__abc_44228_n15691), .Y(u2_remLo_78__FF_INPUT) );
  OR2X2 OR2X2_3665 ( .A(u2__abc_44228_n15695), .B(u2__abc_44228_n15694), .Y(u2__abc_44228_n15696) );
  OR2X2 OR2X2_3666 ( .A(u2__abc_44228_n15693), .B(u2__abc_44228_n15697), .Y(u2_remLo_79__FF_INPUT) );
  OR2X2 OR2X2_3667 ( .A(u2__abc_44228_n15700), .B(u2__abc_44228_n15701), .Y(u2__abc_44228_n15702) );
  OR2X2 OR2X2_3668 ( .A(u2__abc_44228_n15699), .B(u2__abc_44228_n15703), .Y(u2_remLo_80__FF_INPUT) );
  OR2X2 OR2X2_3669 ( .A(u2__abc_44228_n15706), .B(u2__abc_44228_n15707), .Y(u2__abc_44228_n15708) );
  OR2X2 OR2X2_367 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[71] ), .Y(_abc_64468_n1381) );
  OR2X2 OR2X2_3670 ( .A(u2__abc_44228_n15705), .B(u2__abc_44228_n15709), .Y(u2_remLo_81__FF_INPUT) );
  OR2X2 OR2X2_3671 ( .A(u2__abc_44228_n15713), .B(u2__abc_44228_n15712), .Y(u2__abc_44228_n15714) );
  OR2X2 OR2X2_3672 ( .A(u2__abc_44228_n15711), .B(u2__abc_44228_n15715), .Y(u2_remLo_82__FF_INPUT) );
  OR2X2 OR2X2_3673 ( .A(u2__abc_44228_n15719), .B(u2__abc_44228_n15718), .Y(u2__abc_44228_n15720) );
  OR2X2 OR2X2_3674 ( .A(u2__abc_44228_n15717), .B(u2__abc_44228_n15721), .Y(u2_remLo_83__FF_INPUT) );
  OR2X2 OR2X2_3675 ( .A(u2__abc_44228_n15725), .B(u2__abc_44228_n15724), .Y(u2__abc_44228_n15726) );
  OR2X2 OR2X2_3676 ( .A(u2__abc_44228_n15723), .B(u2__abc_44228_n15727), .Y(u2_remLo_84__FF_INPUT) );
  OR2X2 OR2X2_3677 ( .A(u2__abc_44228_n15730), .B(u2__abc_44228_n15731), .Y(u2__abc_44228_n15732) );
  OR2X2 OR2X2_3678 ( .A(u2__abc_44228_n15729), .B(u2__abc_44228_n15733), .Y(u2_remLo_85__FF_INPUT) );
  OR2X2 OR2X2_3679 ( .A(u2__abc_44228_n15736), .B(u2__abc_44228_n15735), .Y(u2__abc_44228_n15737) );
  OR2X2 OR2X2_368 ( .A(a_112_bF_buf6), .B(\a[71] ), .Y(_abc_64468_n1383) );
  OR2X2 OR2X2_3680 ( .A(u2__abc_44228_n15739), .B(u2__abc_44228_n15740), .Y(u2__abc_44228_n15741) );
  OR2X2 OR2X2_3681 ( .A(u2__abc_44228_n15738), .B(u2__abc_44228_n15741), .Y(u2_remLo_86__FF_INPUT) );
  OR2X2 OR2X2_3682 ( .A(u2__abc_44228_n15744), .B(u2__abc_44228_n15745), .Y(u2__abc_44228_n15746) );
  OR2X2 OR2X2_3683 ( .A(u2__abc_44228_n15743), .B(u2__abc_44228_n15747), .Y(u2_remLo_87__FF_INPUT) );
  OR2X2 OR2X2_3684 ( .A(u2__abc_44228_n15750), .B(u2__abc_44228_n15751), .Y(u2__abc_44228_n15752) );
  OR2X2 OR2X2_3685 ( .A(u2__abc_44228_n15749), .B(u2__abc_44228_n15753), .Y(u2_remLo_88__FF_INPUT) );
  OR2X2 OR2X2_3686 ( .A(u2__abc_44228_n15757), .B(u2__abc_44228_n15756), .Y(u2__abc_44228_n15758) );
  OR2X2 OR2X2_3687 ( .A(u2__abc_44228_n15755), .B(u2__abc_44228_n15759), .Y(u2_remLo_89__FF_INPUT) );
  OR2X2 OR2X2_3688 ( .A(u2__abc_44228_n15761), .B(u2__abc_44228_n15762), .Y(u2__abc_44228_n15763) );
  OR2X2 OR2X2_3689 ( .A(u2__abc_44228_n15765), .B(u2__abc_44228_n15766), .Y(u2__abc_44228_n15767) );
  OR2X2 OR2X2_369 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[72] ), .Y(_abc_64468_n1384) );
  OR2X2 OR2X2_3690 ( .A(u2__abc_44228_n15764), .B(u2__abc_44228_n15767), .Y(u2_remLo_90__FF_INPUT) );
  OR2X2 OR2X2_3691 ( .A(u2__abc_44228_n15771), .B(u2__abc_44228_n15770), .Y(u2__abc_44228_n15772) );
  OR2X2 OR2X2_3692 ( .A(u2__abc_44228_n15769), .B(u2__abc_44228_n15773), .Y(u2_remLo_91__FF_INPUT) );
  OR2X2 OR2X2_3693 ( .A(u2__abc_44228_n15776), .B(u2__abc_44228_n15777), .Y(u2__abc_44228_n15778) );
  OR2X2 OR2X2_3694 ( .A(u2__abc_44228_n15775), .B(u2__abc_44228_n15779), .Y(u2_remLo_92__FF_INPUT) );
  OR2X2 OR2X2_3695 ( .A(u2__abc_44228_n15782), .B(u2__abc_44228_n15783), .Y(u2__abc_44228_n15784) );
  OR2X2 OR2X2_3696 ( .A(u2__abc_44228_n15781), .B(u2__abc_44228_n15785), .Y(u2_remLo_93__FF_INPUT) );
  OR2X2 OR2X2_3697 ( .A(u2__abc_44228_n15789), .B(u2__abc_44228_n15788), .Y(u2__abc_44228_n15790) );
  OR2X2 OR2X2_3698 ( .A(u2__abc_44228_n15787), .B(u2__abc_44228_n15791), .Y(u2_remLo_94__FF_INPUT) );
  OR2X2 OR2X2_3699 ( .A(u2__abc_44228_n15795), .B(u2__abc_44228_n15794), .Y(u2__abc_44228_n15796) );
  OR2X2 OR2X2_37 ( .A(aNan_bF_buf2), .B(sqrto_94_), .Y(_abc_64468_n884) );
  OR2X2 OR2X2_370 ( .A(a_112_bF_buf5), .B(\a[72] ), .Y(_abc_64468_n1386) );
  OR2X2 OR2X2_3700 ( .A(u2__abc_44228_n15793), .B(u2__abc_44228_n15797), .Y(u2_remLo_95__FF_INPUT) );
  OR2X2 OR2X2_3701 ( .A(u2__abc_44228_n15800), .B(u2__abc_44228_n15801), .Y(u2__abc_44228_n15802) );
  OR2X2 OR2X2_3702 ( .A(u2__abc_44228_n15799), .B(u2__abc_44228_n15803), .Y(u2_remLo_96__FF_INPUT) );
  OR2X2 OR2X2_3703 ( .A(u2__abc_44228_n15806), .B(u2__abc_44228_n15807), .Y(u2__abc_44228_n15808) );
  OR2X2 OR2X2_3704 ( .A(u2__abc_44228_n15805), .B(u2__abc_44228_n15809), .Y(u2_remLo_97__FF_INPUT) );
  OR2X2 OR2X2_3705 ( .A(u2__abc_44228_n15812), .B(u2__abc_44228_n15813), .Y(u2__abc_44228_n15814) );
  OR2X2 OR2X2_3706 ( .A(u2__abc_44228_n15811), .B(u2__abc_44228_n15815), .Y(u2_remLo_98__FF_INPUT) );
  OR2X2 OR2X2_3707 ( .A(u2__abc_44228_n15818), .B(u2__abc_44228_n15819), .Y(u2__abc_44228_n15820) );
  OR2X2 OR2X2_3708 ( .A(u2__abc_44228_n15817), .B(u2__abc_44228_n15821), .Y(u2_remLo_99__FF_INPUT) );
  OR2X2 OR2X2_3709 ( .A(u2__abc_44228_n15825), .B(u2__abc_44228_n15824), .Y(u2__abc_44228_n15826) );
  OR2X2 OR2X2_371 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[73] ), .Y(_abc_64468_n1387) );
  OR2X2 OR2X2_3710 ( .A(u2__abc_44228_n15823), .B(u2__abc_44228_n15827), .Y(u2_remLo_100__FF_INPUT) );
  OR2X2 OR2X2_3711 ( .A(u2__abc_44228_n15830), .B(u2__abc_44228_n15831), .Y(u2__abc_44228_n15832) );
  OR2X2 OR2X2_3712 ( .A(u2__abc_44228_n15829), .B(u2__abc_44228_n15833), .Y(u2_remLo_101__FF_INPUT) );
  OR2X2 OR2X2_3713 ( .A(u2__abc_44228_n15836), .B(u2__abc_44228_n15837), .Y(u2__abc_44228_n15838) );
  OR2X2 OR2X2_3714 ( .A(u2__abc_44228_n15835), .B(u2__abc_44228_n15839), .Y(u2_remLo_102__FF_INPUT) );
  OR2X2 OR2X2_3715 ( .A(u2__abc_44228_n15842), .B(u2__abc_44228_n15843), .Y(u2__abc_44228_n15844) );
  OR2X2 OR2X2_3716 ( .A(u2__abc_44228_n15841), .B(u2__abc_44228_n15845), .Y(u2_remLo_103__FF_INPUT) );
  OR2X2 OR2X2_3717 ( .A(u2__abc_44228_n15849), .B(u2__abc_44228_n15848), .Y(u2__abc_44228_n15850) );
  OR2X2 OR2X2_3718 ( .A(u2__abc_44228_n15847), .B(u2__abc_44228_n15851), .Y(u2_remLo_104__FF_INPUT) );
  OR2X2 OR2X2_3719 ( .A(u2__abc_44228_n15854), .B(u2__abc_44228_n15855), .Y(u2__abc_44228_n15856) );
  OR2X2 OR2X2_372 ( .A(a_112_bF_buf4), .B(\a[73] ), .Y(_abc_64468_n1389) );
  OR2X2 OR2X2_3720 ( .A(u2__abc_44228_n15853), .B(u2__abc_44228_n15857), .Y(u2_remLo_105__FF_INPUT) );
  OR2X2 OR2X2_3721 ( .A(u2__abc_44228_n15860), .B(u2__abc_44228_n15861), .Y(u2__abc_44228_n15862) );
  OR2X2 OR2X2_3722 ( .A(u2__abc_44228_n15859), .B(u2__abc_44228_n15863), .Y(u2_remLo_106__FF_INPUT) );
  OR2X2 OR2X2_3723 ( .A(u2__abc_44228_n15866), .B(u2__abc_44228_n15867), .Y(u2__abc_44228_n15868) );
  OR2X2 OR2X2_3724 ( .A(u2__abc_44228_n15865), .B(u2__abc_44228_n15869), .Y(u2_remLo_107__FF_INPUT) );
  OR2X2 OR2X2_3725 ( .A(u2__abc_44228_n15872), .B(u2__abc_44228_n15873), .Y(u2__abc_44228_n15874) );
  OR2X2 OR2X2_3726 ( .A(u2__abc_44228_n15871), .B(u2__abc_44228_n15875), .Y(u2_remLo_108__FF_INPUT) );
  OR2X2 OR2X2_3727 ( .A(u2__abc_44228_n15878), .B(u2__abc_44228_n15879), .Y(u2__abc_44228_n15880) );
  OR2X2 OR2X2_3728 ( .A(u2__abc_44228_n15877), .B(u2__abc_44228_n15881), .Y(u2_remLo_109__FF_INPUT) );
  OR2X2 OR2X2_3729 ( .A(u2__abc_44228_n15885), .B(u2__abc_44228_n15884), .Y(u2__abc_44228_n15886) );
  OR2X2 OR2X2_373 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[74] ), .Y(_abc_64468_n1390) );
  OR2X2 OR2X2_3730 ( .A(u2__abc_44228_n15883), .B(u2__abc_44228_n15887), .Y(u2_remLo_110__FF_INPUT) );
  OR2X2 OR2X2_3731 ( .A(u2__abc_44228_n15891), .B(u2__abc_44228_n15890), .Y(u2__abc_44228_n15892) );
  OR2X2 OR2X2_3732 ( .A(u2__abc_44228_n15889), .B(u2__abc_44228_n15893), .Y(u2_remLo_111__FF_INPUT) );
  OR2X2 OR2X2_3733 ( .A(u2__abc_44228_n15897), .B(u2__abc_44228_n15896), .Y(u2__abc_44228_n15898) );
  OR2X2 OR2X2_3734 ( .A(u2__abc_44228_n15895), .B(u2__abc_44228_n15899), .Y(u2_remLo_112__FF_INPUT) );
  OR2X2 OR2X2_3735 ( .A(u2__abc_44228_n15902), .B(u2__abc_44228_n15903), .Y(u2__abc_44228_n15904) );
  OR2X2 OR2X2_3736 ( .A(u2__abc_44228_n15901), .B(u2__abc_44228_n15905), .Y(u2_remLo_113__FF_INPUT) );
  OR2X2 OR2X2_3737 ( .A(u2__abc_44228_n15909), .B(u2__abc_44228_n15908), .Y(u2__abc_44228_n15910) );
  OR2X2 OR2X2_3738 ( .A(u2__abc_44228_n15907), .B(u2__abc_44228_n15911), .Y(u2_remLo_114__FF_INPUT) );
  OR2X2 OR2X2_3739 ( .A(u2__abc_44228_n15914), .B(u2__abc_44228_n15915), .Y(u2__abc_44228_n15916) );
  OR2X2 OR2X2_374 ( .A(a_112_bF_buf3), .B(\a[74] ), .Y(_abc_64468_n1392) );
  OR2X2 OR2X2_3740 ( .A(u2__abc_44228_n15913), .B(u2__abc_44228_n15917), .Y(u2_remLo_115__FF_INPUT) );
  OR2X2 OR2X2_3741 ( .A(u2__abc_44228_n15921), .B(u2__abc_44228_n15920), .Y(u2__abc_44228_n15922) );
  OR2X2 OR2X2_3742 ( .A(u2__abc_44228_n15919), .B(u2__abc_44228_n15923), .Y(u2_remLo_116__FF_INPUT) );
  OR2X2 OR2X2_3743 ( .A(u2__abc_44228_n15926), .B(u2__abc_44228_n15927), .Y(u2__abc_44228_n15928) );
  OR2X2 OR2X2_3744 ( .A(u2__abc_44228_n15925), .B(u2__abc_44228_n15929), .Y(u2_remLo_117__FF_INPUT) );
  OR2X2 OR2X2_3745 ( .A(u2__abc_44228_n15932), .B(u2__abc_44228_n15931), .Y(u2__abc_44228_n15933) );
  OR2X2 OR2X2_3746 ( .A(u2__abc_44228_n15935), .B(u2__abc_44228_n15936), .Y(u2__abc_44228_n15937) );
  OR2X2 OR2X2_3747 ( .A(u2__abc_44228_n15934), .B(u2__abc_44228_n15937), .Y(u2_remLo_118__FF_INPUT) );
  OR2X2 OR2X2_3748 ( .A(u2__abc_44228_n15940), .B(u2__abc_44228_n15941), .Y(u2__abc_44228_n15942) );
  OR2X2 OR2X2_3749 ( .A(u2__abc_44228_n15939), .B(u2__abc_44228_n15943), .Y(u2_remLo_119__FF_INPUT) );
  OR2X2 OR2X2_375 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[75] ), .Y(_abc_64468_n1393) );
  OR2X2 OR2X2_3750 ( .A(u2__abc_44228_n15946), .B(u2__abc_44228_n15947), .Y(u2__abc_44228_n15948) );
  OR2X2 OR2X2_3751 ( .A(u2__abc_44228_n15945), .B(u2__abc_44228_n15949), .Y(u2_remLo_120__FF_INPUT) );
  OR2X2 OR2X2_3752 ( .A(u2__abc_44228_n15952), .B(u2__abc_44228_n15953), .Y(u2__abc_44228_n15954) );
  OR2X2 OR2X2_3753 ( .A(u2__abc_44228_n15951), .B(u2__abc_44228_n15955), .Y(u2_remLo_121__FF_INPUT) );
  OR2X2 OR2X2_3754 ( .A(u2__abc_44228_n15959), .B(u2__abc_44228_n15958), .Y(u2__abc_44228_n15960) );
  OR2X2 OR2X2_3755 ( .A(u2__abc_44228_n15957), .B(u2__abc_44228_n15961), .Y(u2_remLo_122__FF_INPUT) );
  OR2X2 OR2X2_3756 ( .A(u2__abc_44228_n15965), .B(u2__abc_44228_n15964), .Y(u2__abc_44228_n15966) );
  OR2X2 OR2X2_3757 ( .A(u2__abc_44228_n15963), .B(u2__abc_44228_n15967), .Y(u2_remLo_123__FF_INPUT) );
  OR2X2 OR2X2_3758 ( .A(u2__abc_44228_n15970), .B(u2__abc_44228_n15971), .Y(u2__abc_44228_n15972) );
  OR2X2 OR2X2_3759 ( .A(u2__abc_44228_n15969), .B(u2__abc_44228_n15973), .Y(u2_remLo_124__FF_INPUT) );
  OR2X2 OR2X2_376 ( .A(a_112_bF_buf2), .B(\a[75] ), .Y(_abc_64468_n1395) );
  OR2X2 OR2X2_3760 ( .A(u2__abc_44228_n15976), .B(u2__abc_44228_n15977), .Y(u2__abc_44228_n15978) );
  OR2X2 OR2X2_3761 ( .A(u2__abc_44228_n15975), .B(u2__abc_44228_n15979), .Y(u2_remLo_125__FF_INPUT) );
  OR2X2 OR2X2_3762 ( .A(u2__abc_44228_n15982), .B(u2__abc_44228_n15983), .Y(u2__abc_44228_n15984) );
  OR2X2 OR2X2_3763 ( .A(u2__abc_44228_n15981), .B(u2__abc_44228_n15985), .Y(u2_remLo_126__FF_INPUT) );
  OR2X2 OR2X2_3764 ( .A(u2__abc_44228_n15987), .B(u2__abc_44228_n15988), .Y(u2__abc_44228_n15989) );
  OR2X2 OR2X2_3765 ( .A(u2__abc_44228_n15991), .B(u2__abc_44228_n15992), .Y(u2__abc_44228_n15993) );
  OR2X2 OR2X2_3766 ( .A(u2__abc_44228_n15990), .B(u2__abc_44228_n15993), .Y(u2_remLo_127__FF_INPUT) );
  OR2X2 OR2X2_3767 ( .A(u2__abc_44228_n15996), .B(u2__abc_44228_n15997), .Y(u2__abc_44228_n15998) );
  OR2X2 OR2X2_3768 ( .A(u2__abc_44228_n15995), .B(u2__abc_44228_n15999), .Y(u2_remLo_128__FF_INPUT) );
  OR2X2 OR2X2_3769 ( .A(u2__abc_44228_n16003), .B(u2__abc_44228_n16002), .Y(u2__abc_44228_n16004) );
  OR2X2 OR2X2_377 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[76] ), .Y(_abc_64468_n1396) );
  OR2X2 OR2X2_3770 ( .A(u2__abc_44228_n16001), .B(u2__abc_44228_n16005), .Y(u2_remLo_129__FF_INPUT) );
  OR2X2 OR2X2_3771 ( .A(u2__abc_44228_n16009), .B(u2__abc_44228_n16008), .Y(u2__abc_44228_n16010) );
  OR2X2 OR2X2_3772 ( .A(u2__abc_44228_n16007), .B(u2__abc_44228_n16011), .Y(u2_remLo_130__FF_INPUT) );
  OR2X2 OR2X2_3773 ( .A(u2__abc_44228_n16014), .B(u2__abc_44228_n16015), .Y(u2__abc_44228_n16016) );
  OR2X2 OR2X2_3774 ( .A(u2__abc_44228_n16013), .B(u2__abc_44228_n16017), .Y(u2_remLo_131__FF_INPUT) );
  OR2X2 OR2X2_3775 ( .A(u2__abc_44228_n16021), .B(u2__abc_44228_n16020), .Y(u2__abc_44228_n16022) );
  OR2X2 OR2X2_3776 ( .A(u2__abc_44228_n16019), .B(u2__abc_44228_n16023), .Y(u2_remLo_132__FF_INPUT) );
  OR2X2 OR2X2_3777 ( .A(u2__abc_44228_n16026), .B(u2__abc_44228_n16027), .Y(u2__abc_44228_n16028) );
  OR2X2 OR2X2_3778 ( .A(u2__abc_44228_n16025), .B(u2__abc_44228_n16029), .Y(u2_remLo_133__FF_INPUT) );
  OR2X2 OR2X2_3779 ( .A(u2__abc_44228_n16032), .B(u2__abc_44228_n16033), .Y(u2__abc_44228_n16034) );
  OR2X2 OR2X2_378 ( .A(a_112_bF_buf1), .B(\a[76] ), .Y(_abc_64468_n1398) );
  OR2X2 OR2X2_3780 ( .A(u2__abc_44228_n16031), .B(u2__abc_44228_n16035), .Y(u2_remLo_134__FF_INPUT) );
  OR2X2 OR2X2_3781 ( .A(u2__abc_44228_n16038), .B(u2__abc_44228_n16039), .Y(u2__abc_44228_n16040) );
  OR2X2 OR2X2_3782 ( .A(u2__abc_44228_n16037), .B(u2__abc_44228_n16041), .Y(u2_remLo_135__FF_INPUT) );
  OR2X2 OR2X2_3783 ( .A(u2__abc_44228_n16045), .B(u2__abc_44228_n16044), .Y(u2__abc_44228_n16046) );
  OR2X2 OR2X2_3784 ( .A(u2__abc_44228_n16043), .B(u2__abc_44228_n16047), .Y(u2_remLo_136__FF_INPUT) );
  OR2X2 OR2X2_3785 ( .A(u2__abc_44228_n16050), .B(u2__abc_44228_n16051), .Y(u2__abc_44228_n16052) );
  OR2X2 OR2X2_3786 ( .A(u2__abc_44228_n16049), .B(u2__abc_44228_n16053), .Y(u2_remLo_137__FF_INPUT) );
  OR2X2 OR2X2_3787 ( .A(u2__abc_44228_n16057), .B(u2__abc_44228_n16056), .Y(u2__abc_44228_n16058) );
  OR2X2 OR2X2_3788 ( .A(u2__abc_44228_n16055), .B(u2__abc_44228_n16059), .Y(u2_remLo_138__FF_INPUT) );
  OR2X2 OR2X2_3789 ( .A(u2__abc_44228_n16062), .B(u2__abc_44228_n16063), .Y(u2__abc_44228_n16064) );
  OR2X2 OR2X2_379 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[77] ), .Y(_abc_64468_n1399) );
  OR2X2 OR2X2_3790 ( .A(u2__abc_44228_n16061), .B(u2__abc_44228_n16065), .Y(u2_remLo_139__FF_INPUT) );
  OR2X2 OR2X2_3791 ( .A(u2__abc_44228_n16068), .B(u2__abc_44228_n16069), .Y(u2__abc_44228_n16070) );
  OR2X2 OR2X2_3792 ( .A(u2__abc_44228_n16067), .B(u2__abc_44228_n16071), .Y(u2_remLo_140__FF_INPUT) );
  OR2X2 OR2X2_3793 ( .A(u2__abc_44228_n16074), .B(u2__abc_44228_n16075), .Y(u2__abc_44228_n16076) );
  OR2X2 OR2X2_3794 ( .A(u2__abc_44228_n16073), .B(u2__abc_44228_n16077), .Y(u2_remLo_141__FF_INPUT) );
  OR2X2 OR2X2_3795 ( .A(u2__abc_44228_n16081), .B(u2__abc_44228_n16080), .Y(u2__abc_44228_n16082) );
  OR2X2 OR2X2_3796 ( .A(u2__abc_44228_n16079), .B(u2__abc_44228_n16083), .Y(u2_remLo_142__FF_INPUT) );
  OR2X2 OR2X2_3797 ( .A(u2__abc_44228_n16087), .B(u2__abc_44228_n16086), .Y(u2__abc_44228_n16088) );
  OR2X2 OR2X2_3798 ( .A(u2__abc_44228_n16085), .B(u2__abc_44228_n16089), .Y(u2_remLo_143__FF_INPUT) );
  OR2X2 OR2X2_3799 ( .A(u2__abc_44228_n16092), .B(u2__abc_44228_n16093), .Y(u2__abc_44228_n16094) );
  OR2X2 OR2X2_38 ( .A(_abc_64468_n753_bF_buf3), .B(\a[18] ), .Y(_abc_64468_n885) );
  OR2X2 OR2X2_380 ( .A(a_112_bF_buf0), .B(\a[77] ), .Y(_abc_64468_n1401) );
  OR2X2 OR2X2_3800 ( .A(u2__abc_44228_n16091), .B(u2__abc_44228_n16095), .Y(u2_remLo_144__FF_INPUT) );
  OR2X2 OR2X2_3801 ( .A(u2__abc_44228_n16098), .B(u2__abc_44228_n16097), .Y(u2__abc_44228_n16099) );
  OR2X2 OR2X2_3802 ( .A(u2__abc_44228_n16101), .B(u2__abc_44228_n16102), .Y(u2__abc_44228_n16103) );
  OR2X2 OR2X2_3803 ( .A(u2__abc_44228_n16100), .B(u2__abc_44228_n16103), .Y(u2_remLo_145__FF_INPUT) );
  OR2X2 OR2X2_3804 ( .A(u2__abc_44228_n16106), .B(u2__abc_44228_n16105), .Y(u2__abc_44228_n16107) );
  OR2X2 OR2X2_3805 ( .A(u2__abc_44228_n16109), .B(u2__abc_44228_n16110), .Y(u2__abc_44228_n16111) );
  OR2X2 OR2X2_3806 ( .A(u2__abc_44228_n16108), .B(u2__abc_44228_n16111), .Y(u2_remLo_146__FF_INPUT) );
  OR2X2 OR2X2_3807 ( .A(u2__abc_44228_n16115), .B(u2__abc_44228_n16114), .Y(u2__abc_44228_n16116) );
  OR2X2 OR2X2_3808 ( .A(u2__abc_44228_n16113), .B(u2__abc_44228_n16117), .Y(u2_remLo_147__FF_INPUT) );
  OR2X2 OR2X2_3809 ( .A(u2__abc_44228_n16121), .B(u2__abc_44228_n16120), .Y(u2__abc_44228_n16122) );
  OR2X2 OR2X2_381 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[78] ), .Y(_abc_64468_n1402) );
  OR2X2 OR2X2_3810 ( .A(u2__abc_44228_n16119), .B(u2__abc_44228_n16123), .Y(u2_remLo_148__FF_INPUT) );
  OR2X2 OR2X2_3811 ( .A(u2__abc_44228_n16126), .B(u2__abc_44228_n16127), .Y(u2__abc_44228_n16128) );
  OR2X2 OR2X2_3812 ( .A(u2__abc_44228_n16125), .B(u2__abc_44228_n16129), .Y(u2_remLo_149__FF_INPUT) );
  OR2X2 OR2X2_3813 ( .A(u2__abc_44228_n16132), .B(u2__abc_44228_n16131), .Y(u2__abc_44228_n16133) );
  OR2X2 OR2X2_3814 ( .A(u2__abc_44228_n16135), .B(u2__abc_44228_n16136), .Y(u2__abc_44228_n16137) );
  OR2X2 OR2X2_3815 ( .A(u2__abc_44228_n16134), .B(u2__abc_44228_n16137), .Y(u2_remLo_150__FF_INPUT) );
  OR2X2 OR2X2_3816 ( .A(u2__abc_44228_n16140), .B(u2__abc_44228_n16141), .Y(u2__abc_44228_n16142) );
  OR2X2 OR2X2_3817 ( .A(u2__abc_44228_n16139), .B(u2__abc_44228_n16143), .Y(u2_remLo_151__FF_INPUT) );
  OR2X2 OR2X2_3818 ( .A(u2__abc_44228_n16146), .B(u2__abc_44228_n16147), .Y(u2__abc_44228_n16148) );
  OR2X2 OR2X2_3819 ( .A(u2__abc_44228_n16145), .B(u2__abc_44228_n16149), .Y(u2_remLo_152__FF_INPUT) );
  OR2X2 OR2X2_382 ( .A(a_112_bF_buf9), .B(\a[78] ), .Y(_abc_64468_n1404) );
  OR2X2 OR2X2_3820 ( .A(u2__abc_44228_n16152), .B(u2__abc_44228_n16153), .Y(u2__abc_44228_n16154) );
  OR2X2 OR2X2_3821 ( .A(u2__abc_44228_n16151), .B(u2__abc_44228_n16155), .Y(u2_remLo_153__FF_INPUT) );
  OR2X2 OR2X2_3822 ( .A(u2__abc_44228_n16159), .B(u2__abc_44228_n16158), .Y(u2__abc_44228_n16160) );
  OR2X2 OR2X2_3823 ( .A(u2__abc_44228_n16157), .B(u2__abc_44228_n16161), .Y(u2_remLo_154__FF_INPUT) );
  OR2X2 OR2X2_3824 ( .A(u2__abc_44228_n16165), .B(u2__abc_44228_n16164), .Y(u2__abc_44228_n16166) );
  OR2X2 OR2X2_3825 ( .A(u2__abc_44228_n16163), .B(u2__abc_44228_n16167), .Y(u2_remLo_155__FF_INPUT) );
  OR2X2 OR2X2_3826 ( .A(u2__abc_44228_n16170), .B(u2__abc_44228_n16171), .Y(u2__abc_44228_n16172) );
  OR2X2 OR2X2_3827 ( .A(u2__abc_44228_n16169), .B(u2__abc_44228_n16173), .Y(u2_remLo_156__FF_INPUT) );
  OR2X2 OR2X2_3828 ( .A(u2__abc_44228_n16176), .B(u2__abc_44228_n16177), .Y(u2__abc_44228_n16178) );
  OR2X2 OR2X2_3829 ( .A(u2__abc_44228_n16175), .B(u2__abc_44228_n16179), .Y(u2_remLo_157__FF_INPUT) );
  OR2X2 OR2X2_383 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[79] ), .Y(_abc_64468_n1405) );
  OR2X2 OR2X2_3830 ( .A(u2__abc_44228_n16183), .B(u2__abc_44228_n16182), .Y(u2__abc_44228_n16184) );
  OR2X2 OR2X2_3831 ( .A(u2__abc_44228_n16181), .B(u2__abc_44228_n16185), .Y(u2_remLo_158__FF_INPUT) );
  OR2X2 OR2X2_3832 ( .A(u2__abc_44228_n16188), .B(u2__abc_44228_n16189), .Y(u2__abc_44228_n16190) );
  OR2X2 OR2X2_3833 ( .A(u2__abc_44228_n16187), .B(u2__abc_44228_n16191), .Y(u2_remLo_159__FF_INPUT) );
  OR2X2 OR2X2_3834 ( .A(u2__abc_44228_n16195), .B(u2__abc_44228_n16194), .Y(u2__abc_44228_n16196) );
  OR2X2 OR2X2_3835 ( .A(u2__abc_44228_n16193), .B(u2__abc_44228_n16197), .Y(u2_remLo_160__FF_INPUT) );
  OR2X2 OR2X2_3836 ( .A(u2__abc_44228_n16201), .B(u2__abc_44228_n16200), .Y(u2__abc_44228_n16202) );
  OR2X2 OR2X2_3837 ( .A(u2__abc_44228_n16199), .B(u2__abc_44228_n16203), .Y(u2_remLo_161__FF_INPUT) );
  OR2X2 OR2X2_3838 ( .A(u2__abc_44228_n16206), .B(u2__abc_44228_n16207), .Y(u2__abc_44228_n16208) );
  OR2X2 OR2X2_3839 ( .A(u2__abc_44228_n16205), .B(u2__abc_44228_n16209), .Y(u2_remLo_162__FF_INPUT) );
  OR2X2 OR2X2_384 ( .A(a_112_bF_buf8), .B(\a[79] ), .Y(_abc_64468_n1407) );
  OR2X2 OR2X2_3840 ( .A(u2__abc_44228_n16212), .B(u2__abc_44228_n16213), .Y(u2__abc_44228_n16214) );
  OR2X2 OR2X2_3841 ( .A(u2__abc_44228_n16211), .B(u2__abc_44228_n16215), .Y(u2_remLo_163__FF_INPUT) );
  OR2X2 OR2X2_3842 ( .A(u2__abc_44228_n16219), .B(u2__abc_44228_n16218), .Y(u2__abc_44228_n16220) );
  OR2X2 OR2X2_3843 ( .A(u2__abc_44228_n16217), .B(u2__abc_44228_n16221), .Y(u2_remLo_164__FF_INPUT) );
  OR2X2 OR2X2_3844 ( .A(u2__abc_44228_n16224), .B(u2__abc_44228_n16225), .Y(u2__abc_44228_n16226) );
  OR2X2 OR2X2_3845 ( .A(u2__abc_44228_n16223), .B(u2__abc_44228_n16227), .Y(u2_remLo_165__FF_INPUT) );
  OR2X2 OR2X2_3846 ( .A(u2__abc_44228_n16230), .B(u2__abc_44228_n16231), .Y(u2__abc_44228_n16232) );
  OR2X2 OR2X2_3847 ( .A(u2__abc_44228_n16229), .B(u2__abc_44228_n16233), .Y(u2_remLo_166__FF_INPUT) );
  OR2X2 OR2X2_3848 ( .A(u2__abc_44228_n16236), .B(u2__abc_44228_n16237), .Y(u2__abc_44228_n16238) );
  OR2X2 OR2X2_3849 ( .A(u2__abc_44228_n16235), .B(u2__abc_44228_n16239), .Y(u2_remLo_167__FF_INPUT) );
  OR2X2 OR2X2_385 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[80] ), .Y(_abc_64468_n1408) );
  OR2X2 OR2X2_3850 ( .A(u2__abc_44228_n16243), .B(u2__abc_44228_n16242), .Y(u2__abc_44228_n16244) );
  OR2X2 OR2X2_3851 ( .A(u2__abc_44228_n16241), .B(u2__abc_44228_n16245), .Y(u2_remLo_168__FF_INPUT) );
  OR2X2 OR2X2_3852 ( .A(u2__abc_44228_n16248), .B(u2__abc_44228_n16249), .Y(u2__abc_44228_n16250) );
  OR2X2 OR2X2_3853 ( .A(u2__abc_44228_n16247), .B(u2__abc_44228_n16251), .Y(u2_remLo_169__FF_INPUT) );
  OR2X2 OR2X2_3854 ( .A(u2__abc_44228_n16254), .B(u2__abc_44228_n16255), .Y(u2__abc_44228_n16256) );
  OR2X2 OR2X2_3855 ( .A(u2__abc_44228_n16253), .B(u2__abc_44228_n16257), .Y(u2_remLo_170__FF_INPUT) );
  OR2X2 OR2X2_3856 ( .A(u2__abc_44228_n16260), .B(u2__abc_44228_n16261), .Y(u2__abc_44228_n16262) );
  OR2X2 OR2X2_3857 ( .A(u2__abc_44228_n16259), .B(u2__abc_44228_n16263), .Y(u2_remLo_171__FF_INPUT) );
  OR2X2 OR2X2_3858 ( .A(u2__abc_44228_n16266), .B(u2__abc_44228_n16267), .Y(u2__abc_44228_n16268) );
  OR2X2 OR2X2_3859 ( .A(u2__abc_44228_n16265), .B(u2__abc_44228_n16269), .Y(u2_remLo_172__FF_INPUT) );
  OR2X2 OR2X2_386 ( .A(a_112_bF_buf7), .B(\a[80] ), .Y(_abc_64468_n1410) );
  OR2X2 OR2X2_3860 ( .A(u2__abc_44228_n16272), .B(u2__abc_44228_n16273), .Y(u2__abc_44228_n16274) );
  OR2X2 OR2X2_3861 ( .A(u2__abc_44228_n16271), .B(u2__abc_44228_n16275), .Y(u2_remLo_173__FF_INPUT) );
  OR2X2 OR2X2_3862 ( .A(u2__abc_44228_n16279), .B(u2__abc_44228_n16278), .Y(u2__abc_44228_n16280) );
  OR2X2 OR2X2_3863 ( .A(u2__abc_44228_n16277), .B(u2__abc_44228_n16281), .Y(u2_remLo_174__FF_INPUT) );
  OR2X2 OR2X2_3864 ( .A(u2__abc_44228_n16284), .B(u2__abc_44228_n16283), .Y(u2__abc_44228_n16285) );
  OR2X2 OR2X2_3865 ( .A(u2__abc_44228_n16287), .B(u2__abc_44228_n16288), .Y(u2__abc_44228_n16289) );
  OR2X2 OR2X2_3866 ( .A(u2__abc_44228_n16286), .B(u2__abc_44228_n16289), .Y(u2_remLo_175__FF_INPUT) );
  OR2X2 OR2X2_3867 ( .A(u2__abc_44228_n16292), .B(u2__abc_44228_n16293), .Y(u2__abc_44228_n16294) );
  OR2X2 OR2X2_3868 ( .A(u2__abc_44228_n16291), .B(u2__abc_44228_n16295), .Y(u2_remLo_176__FF_INPUT) );
  OR2X2 OR2X2_3869 ( .A(u2__abc_44228_n16298), .B(u2__abc_44228_n16297), .Y(u2__abc_44228_n16299) );
  OR2X2 OR2X2_387 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[81] ), .Y(_abc_64468_n1411) );
  OR2X2 OR2X2_3870 ( .A(u2__abc_44228_n16301), .B(u2__abc_44228_n16302), .Y(u2__abc_44228_n16303) );
  OR2X2 OR2X2_3871 ( .A(u2__abc_44228_n16300), .B(u2__abc_44228_n16303), .Y(u2_remLo_177__FF_INPUT) );
  OR2X2 OR2X2_3872 ( .A(u2__abc_44228_n16306), .B(u2__abc_44228_n16305), .Y(u2__abc_44228_n16307) );
  OR2X2 OR2X2_3873 ( .A(u2__abc_44228_n16309), .B(u2__abc_44228_n16310), .Y(u2__abc_44228_n16311) );
  OR2X2 OR2X2_3874 ( .A(u2__abc_44228_n16308), .B(u2__abc_44228_n16311), .Y(u2_remLo_178__FF_INPUT) );
  OR2X2 OR2X2_3875 ( .A(u2__abc_44228_n16314), .B(u2__abc_44228_n16315), .Y(u2__abc_44228_n16316) );
  OR2X2 OR2X2_3876 ( .A(u2__abc_44228_n16313), .B(u2__abc_44228_n16317), .Y(u2_remLo_179__FF_INPUT) );
  OR2X2 OR2X2_3877 ( .A(u2__abc_44228_n16320), .B(u2__abc_44228_n16321), .Y(u2__abc_44228_n16322) );
  OR2X2 OR2X2_3878 ( .A(u2__abc_44228_n16319), .B(u2__abc_44228_n16323), .Y(u2_remLo_180__FF_INPUT) );
  OR2X2 OR2X2_3879 ( .A(u2__abc_44228_n16326), .B(u2__abc_44228_n16327), .Y(u2__abc_44228_n16328) );
  OR2X2 OR2X2_388 ( .A(a_112_bF_buf6), .B(\a[81] ), .Y(_abc_64468_n1413) );
  OR2X2 OR2X2_3880 ( .A(u2__abc_44228_n16325), .B(u2__abc_44228_n16329), .Y(u2_remLo_181__FF_INPUT) );
  OR2X2 OR2X2_3881 ( .A(u2__abc_44228_n16332), .B(u2__abc_44228_n16331), .Y(u2__abc_44228_n16333) );
  OR2X2 OR2X2_3882 ( .A(u2__abc_44228_n16335), .B(u2__abc_44228_n16336), .Y(u2__abc_44228_n16337) );
  OR2X2 OR2X2_3883 ( .A(u2__abc_44228_n16334), .B(u2__abc_44228_n16337), .Y(u2_remLo_182__FF_INPUT) );
  OR2X2 OR2X2_3884 ( .A(u2__abc_44228_n16340), .B(u2__abc_44228_n16341), .Y(u2__abc_44228_n16342) );
  OR2X2 OR2X2_3885 ( .A(u2__abc_44228_n16339), .B(u2__abc_44228_n16343), .Y(u2_remLo_183__FF_INPUT) );
  OR2X2 OR2X2_3886 ( .A(u2__abc_44228_n16346), .B(u2__abc_44228_n16347), .Y(u2__abc_44228_n16348) );
  OR2X2 OR2X2_3887 ( .A(u2__abc_44228_n16345), .B(u2__abc_44228_n16349), .Y(u2_remLo_184__FF_INPUT) );
  OR2X2 OR2X2_3888 ( .A(u2__abc_44228_n16352), .B(u2__abc_44228_n16353), .Y(u2__abc_44228_n16354) );
  OR2X2 OR2X2_3889 ( .A(u2__abc_44228_n16351), .B(u2__abc_44228_n16355), .Y(u2_remLo_185__FF_INPUT) );
  OR2X2 OR2X2_389 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[82] ), .Y(_abc_64468_n1414) );
  OR2X2 OR2X2_3890 ( .A(u2__abc_44228_n16359), .B(u2__abc_44228_n16358), .Y(u2__abc_44228_n16360) );
  OR2X2 OR2X2_3891 ( .A(u2__abc_44228_n16357), .B(u2__abc_44228_n16361), .Y(u2_remLo_186__FF_INPUT) );
  OR2X2 OR2X2_3892 ( .A(u2__abc_44228_n16365), .B(u2__abc_44228_n16364), .Y(u2__abc_44228_n16366) );
  OR2X2 OR2X2_3893 ( .A(u2__abc_44228_n16363), .B(u2__abc_44228_n16367), .Y(u2_remLo_187__FF_INPUT) );
  OR2X2 OR2X2_3894 ( .A(u2__abc_44228_n16370), .B(u2__abc_44228_n16371), .Y(u2__abc_44228_n16372) );
  OR2X2 OR2X2_3895 ( .A(u2__abc_44228_n16369), .B(u2__abc_44228_n16373), .Y(u2_remLo_188__FF_INPUT) );
  OR2X2 OR2X2_3896 ( .A(u2__abc_44228_n16376), .B(u2__abc_44228_n16377), .Y(u2__abc_44228_n16378) );
  OR2X2 OR2X2_3897 ( .A(u2__abc_44228_n16375), .B(u2__abc_44228_n16379), .Y(u2_remLo_189__FF_INPUT) );
  OR2X2 OR2X2_3898 ( .A(u2__abc_44228_n16383), .B(u2__abc_44228_n16382), .Y(u2__abc_44228_n16384) );
  OR2X2 OR2X2_3899 ( .A(u2__abc_44228_n16381), .B(u2__abc_44228_n16385), .Y(u2_remLo_190__FF_INPUT) );
  OR2X2 OR2X2_39 ( .A(aNan_bF_buf1), .B(sqrto_95_), .Y(_abc_64468_n887) );
  OR2X2 OR2X2_390 ( .A(a_112_bF_buf5), .B(\a[82] ), .Y(_abc_64468_n1416) );
  OR2X2 OR2X2_3900 ( .A(u2__abc_44228_n16388), .B(u2__abc_44228_n16389), .Y(u2__abc_44228_n16390) );
  OR2X2 OR2X2_3901 ( .A(u2__abc_44228_n16387), .B(u2__abc_44228_n16391), .Y(u2_remLo_191__FF_INPUT) );
  OR2X2 OR2X2_3902 ( .A(u2__abc_44228_n16394), .B(u2__abc_44228_n16395), .Y(u2__abc_44228_n16396) );
  OR2X2 OR2X2_3903 ( .A(u2__abc_44228_n16393), .B(u2__abc_44228_n16397), .Y(u2_remLo_192__FF_INPUT) );
  OR2X2 OR2X2_3904 ( .A(u2__abc_44228_n16401), .B(u2__abc_44228_n16400), .Y(u2__abc_44228_n16402) );
  OR2X2 OR2X2_3905 ( .A(u2__abc_44228_n16399), .B(u2__abc_44228_n16403), .Y(u2_remLo_193__FF_INPUT) );
  OR2X2 OR2X2_3906 ( .A(u2__abc_44228_n16406), .B(u2__abc_44228_n16407), .Y(u2__abc_44228_n16408) );
  OR2X2 OR2X2_3907 ( .A(u2__abc_44228_n16405), .B(u2__abc_44228_n16409), .Y(u2_remLo_194__FF_INPUT) );
  OR2X2 OR2X2_3908 ( .A(u2__abc_44228_n16412), .B(u2__abc_44228_n16413), .Y(u2__abc_44228_n16414) );
  OR2X2 OR2X2_3909 ( .A(u2__abc_44228_n16411), .B(u2__abc_44228_n16415), .Y(u2_remLo_195__FF_INPUT) );
  OR2X2 OR2X2_391 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[83] ), .Y(_abc_64468_n1417) );
  OR2X2 OR2X2_3910 ( .A(u2__abc_44228_n16419), .B(u2__abc_44228_n16418), .Y(u2__abc_44228_n16420) );
  OR2X2 OR2X2_3911 ( .A(u2__abc_44228_n16417), .B(u2__abc_44228_n16421), .Y(u2_remLo_196__FF_INPUT) );
  OR2X2 OR2X2_3912 ( .A(u2__abc_44228_n16424), .B(u2__abc_44228_n16425), .Y(u2__abc_44228_n16426) );
  OR2X2 OR2X2_3913 ( .A(u2__abc_44228_n16423), .B(u2__abc_44228_n16427), .Y(u2_remLo_197__FF_INPUT) );
  OR2X2 OR2X2_3914 ( .A(u2__abc_44228_n16430), .B(u2__abc_44228_n16431), .Y(u2__abc_44228_n16432) );
  OR2X2 OR2X2_3915 ( .A(u2__abc_44228_n16429), .B(u2__abc_44228_n16433), .Y(u2_remLo_198__FF_INPUT) );
  OR2X2 OR2X2_3916 ( .A(u2__abc_44228_n16436), .B(u2__abc_44228_n16437), .Y(u2__abc_44228_n16438) );
  OR2X2 OR2X2_3917 ( .A(u2__abc_44228_n16435), .B(u2__abc_44228_n16439), .Y(u2_remLo_199__FF_INPUT) );
  OR2X2 OR2X2_3918 ( .A(u2__abc_44228_n16443), .B(u2__abc_44228_n16442), .Y(u2__abc_44228_n16444) );
  OR2X2 OR2X2_3919 ( .A(u2__abc_44228_n16441), .B(u2__abc_44228_n16445), .Y(u2_remLo_200__FF_INPUT) );
  OR2X2 OR2X2_392 ( .A(a_112_bF_buf4), .B(\a[83] ), .Y(_abc_64468_n1419) );
  OR2X2 OR2X2_3920 ( .A(u2__abc_44228_n16448), .B(u2__abc_44228_n16449), .Y(u2__abc_44228_n16450) );
  OR2X2 OR2X2_3921 ( .A(u2__abc_44228_n16447), .B(u2__abc_44228_n16451), .Y(u2_remLo_201__FF_INPUT) );
  OR2X2 OR2X2_3922 ( .A(u2__abc_44228_n16455), .B(u2__abc_44228_n16454), .Y(u2__abc_44228_n16456) );
  OR2X2 OR2X2_3923 ( .A(u2__abc_44228_n16453), .B(u2__abc_44228_n16457), .Y(u2_remLo_202__FF_INPUT) );
  OR2X2 OR2X2_3924 ( .A(u2__abc_44228_n16460), .B(u2__abc_44228_n16461), .Y(u2__abc_44228_n16462) );
  OR2X2 OR2X2_3925 ( .A(u2__abc_44228_n16459), .B(u2__abc_44228_n16463), .Y(u2_remLo_203__FF_INPUT) );
  OR2X2 OR2X2_3926 ( .A(u2__abc_44228_n16466), .B(u2__abc_44228_n16467), .Y(u2__abc_44228_n16468) );
  OR2X2 OR2X2_3927 ( .A(u2__abc_44228_n16465), .B(u2__abc_44228_n16469), .Y(u2_remLo_204__FF_INPUT) );
  OR2X2 OR2X2_3928 ( .A(u2__abc_44228_n16472), .B(u2__abc_44228_n16473), .Y(u2__abc_44228_n16474) );
  OR2X2 OR2X2_3929 ( .A(u2__abc_44228_n16471), .B(u2__abc_44228_n16475), .Y(u2_remLo_205__FF_INPUT) );
  OR2X2 OR2X2_393 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[84] ), .Y(_abc_64468_n1420) );
  OR2X2 OR2X2_3930 ( .A(u2__abc_44228_n16479), .B(u2__abc_44228_n16478), .Y(u2__abc_44228_n16480) );
  OR2X2 OR2X2_3931 ( .A(u2__abc_44228_n16477), .B(u2__abc_44228_n16481), .Y(u2_remLo_206__FF_INPUT) );
  OR2X2 OR2X2_3932 ( .A(u2__abc_44228_n16485), .B(u2__abc_44228_n16484), .Y(u2__abc_44228_n16486) );
  OR2X2 OR2X2_3933 ( .A(u2__abc_44228_n16483), .B(u2__abc_44228_n16487), .Y(u2_remLo_207__FF_INPUT) );
  OR2X2 OR2X2_3934 ( .A(u2__abc_44228_n16490), .B(u2__abc_44228_n16491), .Y(u2__abc_44228_n16492) );
  OR2X2 OR2X2_3935 ( .A(u2__abc_44228_n16489), .B(u2__abc_44228_n16493), .Y(u2_remLo_208__FF_INPUT) );
  OR2X2 OR2X2_3936 ( .A(u2__abc_44228_n16496), .B(u2__abc_44228_n16497), .Y(u2__abc_44228_n16498) );
  OR2X2 OR2X2_3937 ( .A(u2__abc_44228_n16495), .B(u2__abc_44228_n16499), .Y(u2_remLo_209__FF_INPUT) );
  OR2X2 OR2X2_3938 ( .A(u2__abc_44228_n16502), .B(u2__abc_44228_n16501), .Y(u2__abc_44228_n16503) );
  OR2X2 OR2X2_3939 ( .A(u2__abc_44228_n16505), .B(u2__abc_44228_n16506), .Y(u2__abc_44228_n16507) );
  OR2X2 OR2X2_394 ( .A(a_112_bF_buf3), .B(\a[84] ), .Y(_abc_64468_n1422) );
  OR2X2 OR2X2_3940 ( .A(u2__abc_44228_n16504), .B(u2__abc_44228_n16507), .Y(u2_remLo_210__FF_INPUT) );
  OR2X2 OR2X2_3941 ( .A(u2__abc_44228_n16511), .B(u2__abc_44228_n16510), .Y(u2__abc_44228_n16512) );
  OR2X2 OR2X2_3942 ( .A(u2__abc_44228_n16509), .B(u2__abc_44228_n16513), .Y(u2_remLo_211__FF_INPUT) );
  OR2X2 OR2X2_3943 ( .A(u2__abc_44228_n16517), .B(u2__abc_44228_n16516), .Y(u2__abc_44228_n16518) );
  OR2X2 OR2X2_3944 ( .A(u2__abc_44228_n16515), .B(u2__abc_44228_n16519), .Y(u2_remLo_212__FF_INPUT) );
  OR2X2 OR2X2_3945 ( .A(u2__abc_44228_n16522), .B(u2__abc_44228_n16523), .Y(u2__abc_44228_n16524) );
  OR2X2 OR2X2_3946 ( .A(u2__abc_44228_n16521), .B(u2__abc_44228_n16525), .Y(u2_remLo_213__FF_INPUT) );
  OR2X2 OR2X2_3947 ( .A(u2__abc_44228_n16528), .B(u2__abc_44228_n16527), .Y(u2__abc_44228_n16529) );
  OR2X2 OR2X2_3948 ( .A(u2__abc_44228_n16531), .B(u2__abc_44228_n16532), .Y(u2__abc_44228_n16533) );
  OR2X2 OR2X2_3949 ( .A(u2__abc_44228_n16530), .B(u2__abc_44228_n16533), .Y(u2_remLo_214__FF_INPUT) );
  OR2X2 OR2X2_395 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[85] ), .Y(_abc_64468_n1423) );
  OR2X2 OR2X2_3950 ( .A(u2__abc_44228_n16536), .B(u2__abc_44228_n16537), .Y(u2__abc_44228_n16538) );
  OR2X2 OR2X2_3951 ( .A(u2__abc_44228_n16535), .B(u2__abc_44228_n16539), .Y(u2_remLo_215__FF_INPUT) );
  OR2X2 OR2X2_3952 ( .A(u2__abc_44228_n16542), .B(u2__abc_44228_n16543), .Y(u2__abc_44228_n16544) );
  OR2X2 OR2X2_3953 ( .A(u2__abc_44228_n16541), .B(u2__abc_44228_n16545), .Y(u2_remLo_216__FF_INPUT) );
  OR2X2 OR2X2_3954 ( .A(u2__abc_44228_n16548), .B(u2__abc_44228_n16549), .Y(u2__abc_44228_n16550) );
  OR2X2 OR2X2_3955 ( .A(u2__abc_44228_n16547), .B(u2__abc_44228_n16551), .Y(u2_remLo_217__FF_INPUT) );
  OR2X2 OR2X2_3956 ( .A(u2__abc_44228_n16553), .B(u2__abc_44228_n16554), .Y(u2__abc_44228_n16555) );
  OR2X2 OR2X2_3957 ( .A(u2__abc_44228_n16557), .B(u2__abc_44228_n16558), .Y(u2__abc_44228_n16559) );
  OR2X2 OR2X2_3958 ( .A(u2__abc_44228_n16556), .B(u2__abc_44228_n16559), .Y(u2_remLo_218__FF_INPUT) );
  OR2X2 OR2X2_3959 ( .A(u2__abc_44228_n16562), .B(u2__abc_44228_n16563), .Y(u2__abc_44228_n16564) );
  OR2X2 OR2X2_396 ( .A(a_112_bF_buf2), .B(\a[85] ), .Y(_abc_64468_n1425) );
  OR2X2 OR2X2_3960 ( .A(u2__abc_44228_n16561), .B(u2__abc_44228_n16565), .Y(u2_remLo_219__FF_INPUT) );
  OR2X2 OR2X2_3961 ( .A(u2__abc_44228_n16568), .B(u2__abc_44228_n16569), .Y(u2__abc_44228_n16570) );
  OR2X2 OR2X2_3962 ( .A(u2__abc_44228_n16567), .B(u2__abc_44228_n16571), .Y(u2_remLo_220__FF_INPUT) );
  OR2X2 OR2X2_3963 ( .A(u2__abc_44228_n16574), .B(u2__abc_44228_n16575), .Y(u2__abc_44228_n16576) );
  OR2X2 OR2X2_3964 ( .A(u2__abc_44228_n16573), .B(u2__abc_44228_n16577), .Y(u2_remLo_221__FF_INPUT) );
  OR2X2 OR2X2_3965 ( .A(u2__abc_44228_n16579), .B(u2__abc_44228_n16580), .Y(u2__abc_44228_n16581) );
  OR2X2 OR2X2_3966 ( .A(u2__abc_44228_n16583), .B(u2__abc_44228_n16584), .Y(u2__abc_44228_n16585) );
  OR2X2 OR2X2_3967 ( .A(u2__abc_44228_n16582), .B(u2__abc_44228_n16585), .Y(u2_remLo_222__FF_INPUT) );
  OR2X2 OR2X2_3968 ( .A(u2__abc_44228_n16589), .B(u2__abc_44228_n16588), .Y(u2__abc_44228_n16590) );
  OR2X2 OR2X2_3969 ( .A(u2__abc_44228_n16587), .B(u2__abc_44228_n16591), .Y(u2_remLo_223__FF_INPUT) );
  OR2X2 OR2X2_397 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[86] ), .Y(_abc_64468_n1426) );
  OR2X2 OR2X2_3970 ( .A(u2__abc_44228_n16594), .B(u2__abc_44228_n16595), .Y(u2__abc_44228_n16596) );
  OR2X2 OR2X2_3971 ( .A(u2__abc_44228_n16593), .B(u2__abc_44228_n16597), .Y(u2_remLo_224__FF_INPUT) );
  OR2X2 OR2X2_3972 ( .A(u2__abc_44228_n16600), .B(u2__abc_44228_n16601), .Y(u2__abc_44228_n16602) );
  OR2X2 OR2X2_3973 ( .A(u2__abc_44228_n16599), .B(u2__abc_44228_n16603), .Y(u2_remLo_225__FF_INPUT) );
  OR2X2 OR2X2_3974 ( .A(u2__abc_44228_n16607), .B(u2__abc_44228_n16606), .Y(u2__abc_44228_n16608) );
  OR2X2 OR2X2_3975 ( .A(u2__abc_44228_n16605), .B(u2__abc_44228_n16609), .Y(u2_remLo_226__FF_INPUT) );
  OR2X2 OR2X2_3976 ( .A(u2__abc_44228_n16612), .B(u2__abc_44228_n16613), .Y(u2__abc_44228_n16614) );
  OR2X2 OR2X2_3977 ( .A(u2__abc_44228_n16611), .B(u2__abc_44228_n16615), .Y(u2_remLo_227__FF_INPUT) );
  OR2X2 OR2X2_3978 ( .A(u2__abc_44228_n16619), .B(u2__abc_44228_n16618), .Y(u2__abc_44228_n16620) );
  OR2X2 OR2X2_3979 ( .A(u2__abc_44228_n16617), .B(u2__abc_44228_n16621), .Y(u2_remLo_228__FF_INPUT) );
  OR2X2 OR2X2_398 ( .A(a_112_bF_buf1), .B(\a[86] ), .Y(_abc_64468_n1428) );
  OR2X2 OR2X2_3980 ( .A(u2__abc_44228_n16624), .B(u2__abc_44228_n16625), .Y(u2__abc_44228_n16626) );
  OR2X2 OR2X2_3981 ( .A(u2__abc_44228_n16623), .B(u2__abc_44228_n16627), .Y(u2_remLo_229__FF_INPUT) );
  OR2X2 OR2X2_3982 ( .A(u2__abc_44228_n16630), .B(u2__abc_44228_n16631), .Y(u2__abc_44228_n16632) );
  OR2X2 OR2X2_3983 ( .A(u2__abc_44228_n16629), .B(u2__abc_44228_n16633), .Y(u2_remLo_230__FF_INPUT) );
  OR2X2 OR2X2_3984 ( .A(u2__abc_44228_n16636), .B(u2__abc_44228_n16637), .Y(u2__abc_44228_n16638) );
  OR2X2 OR2X2_3985 ( .A(u2__abc_44228_n16635), .B(u2__abc_44228_n16639), .Y(u2_remLo_231__FF_INPUT) );
  OR2X2 OR2X2_3986 ( .A(u2__abc_44228_n16643), .B(u2__abc_44228_n16642), .Y(u2__abc_44228_n16644) );
  OR2X2 OR2X2_3987 ( .A(u2__abc_44228_n16641), .B(u2__abc_44228_n16645), .Y(u2_remLo_232__FF_INPUT) );
  OR2X2 OR2X2_3988 ( .A(u2__abc_44228_n16648), .B(u2__abc_44228_n16649), .Y(u2__abc_44228_n16650) );
  OR2X2 OR2X2_3989 ( .A(u2__abc_44228_n16647), .B(u2__abc_44228_n16651), .Y(u2_remLo_233__FF_INPUT) );
  OR2X2 OR2X2_399 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[87] ), .Y(_abc_64468_n1429) );
  OR2X2 OR2X2_3990 ( .A(u2__abc_44228_n16655), .B(u2__abc_44228_n16654), .Y(u2__abc_44228_n16656) );
  OR2X2 OR2X2_3991 ( .A(u2__abc_44228_n16653), .B(u2__abc_44228_n16657), .Y(u2_remLo_234__FF_INPUT) );
  OR2X2 OR2X2_3992 ( .A(u2__abc_44228_n16660), .B(u2__abc_44228_n16661), .Y(u2__abc_44228_n16662) );
  OR2X2 OR2X2_3993 ( .A(u2__abc_44228_n16659), .B(u2__abc_44228_n16663), .Y(u2_remLo_235__FF_INPUT) );
  OR2X2 OR2X2_3994 ( .A(u2__abc_44228_n16666), .B(u2__abc_44228_n16667), .Y(u2__abc_44228_n16668) );
  OR2X2 OR2X2_3995 ( .A(u2__abc_44228_n16665), .B(u2__abc_44228_n16669), .Y(u2_remLo_236__FF_INPUT) );
  OR2X2 OR2X2_3996 ( .A(u2__abc_44228_n16672), .B(u2__abc_44228_n16673), .Y(u2__abc_44228_n16674) );
  OR2X2 OR2X2_3997 ( .A(u2__abc_44228_n16671), .B(u2__abc_44228_n16675), .Y(u2_remLo_237__FF_INPUT) );
  OR2X2 OR2X2_3998 ( .A(u2__abc_44228_n16678), .B(u2__abc_44228_n16679), .Y(u2__abc_44228_n16680) );
  OR2X2 OR2X2_3999 ( .A(u2__abc_44228_n16677), .B(u2__abc_44228_n16681), .Y(u2_remLo_238__FF_INPUT) );
  OR2X2 OR2X2_4 ( .A(_abc_64468_n753_bF_buf6), .B(\a[1] ), .Y(_abc_64468_n834) );
  OR2X2 OR2X2_40 ( .A(_abc_64468_n753_bF_buf2), .B(\a[19] ), .Y(_abc_64468_n888) );
  OR2X2 OR2X2_400 ( .A(a_112_bF_buf0), .B(\a[87] ), .Y(_abc_64468_n1431) );
  OR2X2 OR2X2_4000 ( .A(u2__abc_44228_n16685), .B(u2__abc_44228_n16684), .Y(u2__abc_44228_n16686) );
  OR2X2 OR2X2_4001 ( .A(u2__abc_44228_n16683), .B(u2__abc_44228_n16687), .Y(u2_remLo_239__FF_INPUT) );
  OR2X2 OR2X2_4002 ( .A(u2__abc_44228_n16690), .B(u2__abc_44228_n16691), .Y(u2__abc_44228_n16692) );
  OR2X2 OR2X2_4003 ( .A(u2__abc_44228_n16689), .B(u2__abc_44228_n16693), .Y(u2_remLo_240__FF_INPUT) );
  OR2X2 OR2X2_4004 ( .A(u2__abc_44228_n16696), .B(u2__abc_44228_n16697), .Y(u2__abc_44228_n16698) );
  OR2X2 OR2X2_4005 ( .A(u2__abc_44228_n16695), .B(u2__abc_44228_n16699), .Y(u2_remLo_241__FF_INPUT) );
  OR2X2 OR2X2_4006 ( .A(u2__abc_44228_n16702), .B(u2__abc_44228_n16701), .Y(u2__abc_44228_n16703) );
  OR2X2 OR2X2_4007 ( .A(u2__abc_44228_n16705), .B(u2__abc_44228_n16706), .Y(u2__abc_44228_n16707) );
  OR2X2 OR2X2_4008 ( .A(u2__abc_44228_n16704), .B(u2__abc_44228_n16707), .Y(u2_remLo_242__FF_INPUT) );
  OR2X2 OR2X2_4009 ( .A(u2__abc_44228_n16711), .B(u2__abc_44228_n16710), .Y(u2__abc_44228_n16712) );
  OR2X2 OR2X2_401 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[88] ), .Y(_abc_64468_n1432) );
  OR2X2 OR2X2_4010 ( .A(u2__abc_44228_n16709), .B(u2__abc_44228_n16713), .Y(u2_remLo_243__FF_INPUT) );
  OR2X2 OR2X2_4011 ( .A(u2__abc_44228_n16717), .B(u2__abc_44228_n16716), .Y(u2__abc_44228_n16718) );
  OR2X2 OR2X2_4012 ( .A(u2__abc_44228_n16715), .B(u2__abc_44228_n16719), .Y(u2_remLo_244__FF_INPUT) );
  OR2X2 OR2X2_4013 ( .A(u2__abc_44228_n16722), .B(u2__abc_44228_n16723), .Y(u2__abc_44228_n16724) );
  OR2X2 OR2X2_4014 ( .A(u2__abc_44228_n16721), .B(u2__abc_44228_n16725), .Y(u2_remLo_245__FF_INPUT) );
  OR2X2 OR2X2_4015 ( .A(u2__abc_44228_n16728), .B(u2__abc_44228_n16727), .Y(u2__abc_44228_n16729) );
  OR2X2 OR2X2_4016 ( .A(u2__abc_44228_n16731), .B(u2__abc_44228_n16732), .Y(u2__abc_44228_n16733) );
  OR2X2 OR2X2_4017 ( .A(u2__abc_44228_n16730), .B(u2__abc_44228_n16733), .Y(u2_remLo_246__FF_INPUT) );
  OR2X2 OR2X2_4018 ( .A(u2__abc_44228_n16736), .B(u2__abc_44228_n16737), .Y(u2__abc_44228_n16738) );
  OR2X2 OR2X2_4019 ( .A(u2__abc_44228_n16735), .B(u2__abc_44228_n16739), .Y(u2_remLo_247__FF_INPUT) );
  OR2X2 OR2X2_402 ( .A(a_112_bF_buf9), .B(\a[88] ), .Y(_abc_64468_n1434) );
  OR2X2 OR2X2_4020 ( .A(u2__abc_44228_n16742), .B(u2__abc_44228_n16743), .Y(u2__abc_44228_n16744) );
  OR2X2 OR2X2_4021 ( .A(u2__abc_44228_n16741), .B(u2__abc_44228_n16745), .Y(u2_remLo_248__FF_INPUT) );
  OR2X2 OR2X2_4022 ( .A(u2__abc_44228_n16748), .B(u2__abc_44228_n16749), .Y(u2__abc_44228_n16750) );
  OR2X2 OR2X2_4023 ( .A(u2__abc_44228_n16747), .B(u2__abc_44228_n16751), .Y(u2_remLo_249__FF_INPUT) );
  OR2X2 OR2X2_4024 ( .A(u2__abc_44228_n16755), .B(u2__abc_44228_n16754), .Y(u2__abc_44228_n16756) );
  OR2X2 OR2X2_4025 ( .A(u2__abc_44228_n16753), .B(u2__abc_44228_n16757), .Y(u2_remLo_250__FF_INPUT) );
  OR2X2 OR2X2_4026 ( .A(u2__abc_44228_n16759), .B(u2__abc_44228_n16760), .Y(u2__abc_44228_n16761) );
  OR2X2 OR2X2_4027 ( .A(u2__abc_44228_n16763), .B(u2__abc_44228_n16764), .Y(u2__abc_44228_n16765) );
  OR2X2 OR2X2_4028 ( .A(u2__abc_44228_n16762), .B(u2__abc_44228_n16765), .Y(u2_remLo_251__FF_INPUT) );
  OR2X2 OR2X2_4029 ( .A(u2__abc_44228_n16768), .B(u2__abc_44228_n16769), .Y(u2__abc_44228_n16770) );
  OR2X2 OR2X2_403 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[89] ), .Y(_abc_64468_n1435) );
  OR2X2 OR2X2_4030 ( .A(u2__abc_44228_n16767), .B(u2__abc_44228_n16771), .Y(u2_remLo_252__FF_INPUT) );
  OR2X2 OR2X2_4031 ( .A(u2__abc_44228_n16774), .B(u2__abc_44228_n16775), .Y(u2__abc_44228_n16776) );
  OR2X2 OR2X2_4032 ( .A(u2__abc_44228_n16773), .B(u2__abc_44228_n16777), .Y(u2_remLo_253__FF_INPUT) );
  OR2X2 OR2X2_4033 ( .A(u2__abc_44228_n16781), .B(u2__abc_44228_n16780), .Y(u2__abc_44228_n16782) );
  OR2X2 OR2X2_4034 ( .A(u2__abc_44228_n16779), .B(u2__abc_44228_n16783), .Y(u2_remLo_254__FF_INPUT) );
  OR2X2 OR2X2_4035 ( .A(u2__abc_44228_n16786), .B(u2__abc_44228_n16787), .Y(u2__abc_44228_n16788) );
  OR2X2 OR2X2_4036 ( .A(u2__abc_44228_n16785), .B(u2__abc_44228_n16789), .Y(u2_remLo_255__FF_INPUT) );
  OR2X2 OR2X2_4037 ( .A(u2__abc_44228_n16793), .B(u2__abc_44228_n16792), .Y(u2__abc_44228_n16794) );
  OR2X2 OR2X2_4038 ( .A(u2__abc_44228_n16791), .B(u2__abc_44228_n16795), .Y(u2_remLo_256__FF_INPUT) );
  OR2X2 OR2X2_4039 ( .A(u2__abc_44228_n16799), .B(u2__abc_44228_n16798), .Y(u2__abc_44228_n16800) );
  OR2X2 OR2X2_404 ( .A(a_112_bF_buf8), .B(\a[89] ), .Y(_abc_64468_n1437) );
  OR2X2 OR2X2_4040 ( .A(u2__abc_44228_n16797), .B(u2__abc_44228_n16801), .Y(u2_remLo_257__FF_INPUT) );
  OR2X2 OR2X2_4041 ( .A(u2__abc_44228_n16803), .B(u2__abc_44228_n16805), .Y(u2__abc_44228_n16806) );
  OR2X2 OR2X2_4042 ( .A(u2__abc_44228_n16808), .B(u2__abc_44228_n16810), .Y(u2__abc_44228_n16811) );
  OR2X2 OR2X2_4043 ( .A(u2__abc_44228_n16813), .B(u2__abc_44228_n16815), .Y(u2__abc_44228_n16816) );
  OR2X2 OR2X2_4044 ( .A(u2__abc_44228_n16818), .B(u2__abc_44228_n16820), .Y(u2__abc_44228_n16821) );
  OR2X2 OR2X2_4045 ( .A(u2__abc_44228_n16823), .B(u2__abc_44228_n16825), .Y(u2__abc_44228_n16826) );
  OR2X2 OR2X2_4046 ( .A(u2__abc_44228_n16828), .B(u2__abc_44228_n16830), .Y(u2__abc_44228_n16831) );
  OR2X2 OR2X2_4047 ( .A(u2__abc_44228_n16833), .B(u2__abc_44228_n16835), .Y(u2__abc_44228_n16836) );
  OR2X2 OR2X2_4048 ( .A(u2__abc_44228_n16838), .B(u2__abc_44228_n16840), .Y(u2__abc_44228_n16841) );
  OR2X2 OR2X2_4049 ( .A(u2__abc_44228_n16843), .B(u2__abc_44228_n16845), .Y(u2__abc_44228_n16846) );
  OR2X2 OR2X2_405 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[90] ), .Y(_abc_64468_n1438) );
  OR2X2 OR2X2_4050 ( .A(u2__abc_44228_n16848), .B(u2__abc_44228_n16850), .Y(u2__abc_44228_n16851) );
  OR2X2 OR2X2_4051 ( .A(u2__abc_44228_n16853), .B(u2__abc_44228_n16855), .Y(u2__abc_44228_n16856) );
  OR2X2 OR2X2_4052 ( .A(u2__abc_44228_n16858), .B(u2__abc_44228_n16860), .Y(u2__abc_44228_n16861) );
  OR2X2 OR2X2_4053 ( .A(u2__abc_44228_n16863), .B(u2__abc_44228_n16865), .Y(u2__abc_44228_n16866) );
  OR2X2 OR2X2_4054 ( .A(u2__abc_44228_n16868), .B(u2__abc_44228_n16870), .Y(u2__abc_44228_n16871) );
  OR2X2 OR2X2_4055 ( .A(u2__abc_44228_n16873), .B(u2__abc_44228_n16875), .Y(u2__abc_44228_n16876) );
  OR2X2 OR2X2_4056 ( .A(u2__abc_44228_n16878), .B(u2__abc_44228_n16880), .Y(u2__abc_44228_n16881) );
  OR2X2 OR2X2_4057 ( .A(u2__abc_44228_n16883), .B(u2__abc_44228_n16885), .Y(u2__abc_44228_n16886) );
  OR2X2 OR2X2_4058 ( .A(u2__abc_44228_n16888), .B(u2__abc_44228_n16890), .Y(u2__abc_44228_n16891) );
  OR2X2 OR2X2_4059 ( .A(u2__abc_44228_n16893), .B(u2__abc_44228_n16895), .Y(u2__abc_44228_n16896) );
  OR2X2 OR2X2_406 ( .A(a_112_bF_buf7), .B(\a[90] ), .Y(_abc_64468_n1440) );
  OR2X2 OR2X2_4060 ( .A(u2__abc_44228_n16898), .B(u2__abc_44228_n16900), .Y(u2__abc_44228_n16901) );
  OR2X2 OR2X2_4061 ( .A(u2__abc_44228_n16903), .B(u2__abc_44228_n16905), .Y(u2__abc_44228_n16906) );
  OR2X2 OR2X2_4062 ( .A(u2__abc_44228_n16908), .B(u2__abc_44228_n16910), .Y(u2__abc_44228_n16911) );
  OR2X2 OR2X2_4063 ( .A(u2__abc_44228_n16913), .B(u2__abc_44228_n16915), .Y(u2__abc_44228_n16916) );
  OR2X2 OR2X2_4064 ( .A(u2__abc_44228_n16918), .B(u2__abc_44228_n16920), .Y(u2__abc_44228_n16921) );
  OR2X2 OR2X2_4065 ( .A(u2__abc_44228_n16923), .B(u2__abc_44228_n16925), .Y(u2__abc_44228_n16926) );
  OR2X2 OR2X2_4066 ( .A(u2__abc_44228_n16928), .B(u2__abc_44228_n16930), .Y(u2__abc_44228_n16931) );
  OR2X2 OR2X2_4067 ( .A(u2__abc_44228_n16933), .B(u2__abc_44228_n16935), .Y(u2__abc_44228_n16936) );
  OR2X2 OR2X2_4068 ( .A(u2__abc_44228_n16938), .B(u2__abc_44228_n16940), .Y(u2__abc_44228_n16941) );
  OR2X2 OR2X2_4069 ( .A(u2__abc_44228_n16943), .B(u2__abc_44228_n16945), .Y(u2__abc_44228_n16946) );
  OR2X2 OR2X2_407 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[91] ), .Y(_abc_64468_n1441) );
  OR2X2 OR2X2_4070 ( .A(u2__abc_44228_n16948), .B(u2__abc_44228_n16950), .Y(u2__abc_44228_n16951) );
  OR2X2 OR2X2_4071 ( .A(u2__abc_44228_n16953), .B(u2__abc_44228_n16955), .Y(u2__abc_44228_n16956) );
  OR2X2 OR2X2_4072 ( .A(u2__abc_44228_n16958), .B(u2__abc_44228_n16960), .Y(u2__abc_44228_n16961) );
  OR2X2 OR2X2_4073 ( .A(u2__abc_44228_n16963), .B(u2__abc_44228_n16965), .Y(u2__abc_44228_n16966) );
  OR2X2 OR2X2_4074 ( .A(u2__abc_44228_n16968), .B(u2__abc_44228_n16970), .Y(u2__abc_44228_n16971) );
  OR2X2 OR2X2_4075 ( .A(u2__abc_44228_n16973), .B(u2__abc_44228_n16975), .Y(u2__abc_44228_n16976) );
  OR2X2 OR2X2_4076 ( .A(u2__abc_44228_n16978), .B(u2__abc_44228_n16980), .Y(u2__abc_44228_n16981) );
  OR2X2 OR2X2_4077 ( .A(u2__abc_44228_n16983), .B(u2__abc_44228_n16985), .Y(u2__abc_44228_n16986) );
  OR2X2 OR2X2_4078 ( .A(u2__abc_44228_n16988), .B(u2__abc_44228_n16990), .Y(u2__abc_44228_n16991) );
  OR2X2 OR2X2_4079 ( .A(u2__abc_44228_n16993), .B(u2__abc_44228_n16995), .Y(u2__abc_44228_n16996) );
  OR2X2 OR2X2_408 ( .A(a_112_bF_buf6), .B(\a[91] ), .Y(_abc_64468_n1443) );
  OR2X2 OR2X2_4080 ( .A(u2__abc_44228_n16998), .B(u2__abc_44228_n17000), .Y(u2__abc_44228_n17001) );
  OR2X2 OR2X2_4081 ( .A(u2__abc_44228_n17003), .B(u2__abc_44228_n17005), .Y(u2__abc_44228_n17006) );
  OR2X2 OR2X2_4082 ( .A(u2__abc_44228_n17008), .B(u2__abc_44228_n17010), .Y(u2__abc_44228_n17011) );
  OR2X2 OR2X2_4083 ( .A(u2__abc_44228_n17013), .B(u2__abc_44228_n17015), .Y(u2__abc_44228_n17016) );
  OR2X2 OR2X2_4084 ( .A(u2__abc_44228_n17018), .B(u2__abc_44228_n17020), .Y(u2__abc_44228_n17021) );
  OR2X2 OR2X2_4085 ( .A(u2__abc_44228_n17023), .B(u2__abc_44228_n17025), .Y(u2__abc_44228_n17026) );
  OR2X2 OR2X2_4086 ( .A(u2__abc_44228_n17028), .B(u2__abc_44228_n17030), .Y(u2__abc_44228_n17031) );
  OR2X2 OR2X2_4087 ( .A(u2__abc_44228_n17033), .B(u2__abc_44228_n17035), .Y(u2__abc_44228_n17036) );
  OR2X2 OR2X2_4088 ( .A(u2__abc_44228_n17038), .B(u2__abc_44228_n17040), .Y(u2__abc_44228_n17041) );
  OR2X2 OR2X2_4089 ( .A(u2__abc_44228_n17043), .B(u2__abc_44228_n17045), .Y(u2__abc_44228_n17046) );
  OR2X2 OR2X2_409 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[92] ), .Y(_abc_64468_n1444) );
  OR2X2 OR2X2_4090 ( .A(u2__abc_44228_n17048), .B(u2__abc_44228_n17050), .Y(u2__abc_44228_n17051) );
  OR2X2 OR2X2_4091 ( .A(u2__abc_44228_n17053), .B(u2__abc_44228_n17055), .Y(u2__abc_44228_n17056) );
  OR2X2 OR2X2_4092 ( .A(u2__abc_44228_n17058), .B(u2__abc_44228_n17060), .Y(u2__abc_44228_n17061) );
  OR2X2 OR2X2_4093 ( .A(u2__abc_44228_n17063), .B(u2__abc_44228_n17065), .Y(u2__abc_44228_n17066) );
  OR2X2 OR2X2_4094 ( .A(u2__abc_44228_n17068), .B(u2__abc_44228_n17070), .Y(u2__abc_44228_n17071) );
  OR2X2 OR2X2_4095 ( .A(u2__abc_44228_n17073), .B(u2__abc_44228_n17075), .Y(u2__abc_44228_n17076) );
  OR2X2 OR2X2_4096 ( .A(u2__abc_44228_n17078), .B(u2__abc_44228_n17080), .Y(u2__abc_44228_n17081) );
  OR2X2 OR2X2_4097 ( .A(u2__abc_44228_n17083), .B(u2__abc_44228_n17085), .Y(u2__abc_44228_n17086) );
  OR2X2 OR2X2_4098 ( .A(u2__abc_44228_n17088), .B(u2__abc_44228_n17090), .Y(u2__abc_44228_n17091) );
  OR2X2 OR2X2_4099 ( .A(u2__abc_44228_n17093), .B(u2__abc_44228_n17095), .Y(u2__abc_44228_n17096) );
  OR2X2 OR2X2_41 ( .A(aNan_bF_buf0), .B(sqrto_96_), .Y(_abc_64468_n890) );
  OR2X2 OR2X2_410 ( .A(a_112_bF_buf5), .B(\a[92] ), .Y(_abc_64468_n1446) );
  OR2X2 OR2X2_4100 ( .A(u2__abc_44228_n17098), .B(u2__abc_44228_n17100), .Y(u2__abc_44228_n17101) );
  OR2X2 OR2X2_4101 ( .A(u2__abc_44228_n17103), .B(u2__abc_44228_n17105), .Y(u2__abc_44228_n17106) );
  OR2X2 OR2X2_4102 ( .A(u2__abc_44228_n17108), .B(u2__abc_44228_n17110), .Y(u2__abc_44228_n17111) );
  OR2X2 OR2X2_4103 ( .A(u2__abc_44228_n17113), .B(u2__abc_44228_n17115), .Y(u2__abc_44228_n17116) );
  OR2X2 OR2X2_4104 ( .A(u2__abc_44228_n17118), .B(u2__abc_44228_n17120), .Y(u2__abc_44228_n17121) );
  OR2X2 OR2X2_4105 ( .A(u2__abc_44228_n17123), .B(u2__abc_44228_n17125), .Y(u2__abc_44228_n17126) );
  OR2X2 OR2X2_4106 ( .A(u2__abc_44228_n17128), .B(u2__abc_44228_n17130), .Y(u2__abc_44228_n17131) );
  OR2X2 OR2X2_4107 ( .A(u2__abc_44228_n17133), .B(u2__abc_44228_n17135), .Y(u2__abc_44228_n17136) );
  OR2X2 OR2X2_4108 ( .A(u2__abc_44228_n17138), .B(u2__abc_44228_n17140), .Y(u2__abc_44228_n17141) );
  OR2X2 OR2X2_4109 ( .A(u2__abc_44228_n17143), .B(u2__abc_44228_n17145), .Y(u2__abc_44228_n17146) );
  OR2X2 OR2X2_411 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[93] ), .Y(_abc_64468_n1447) );
  OR2X2 OR2X2_4110 ( .A(u2__abc_44228_n17148), .B(u2__abc_44228_n17150), .Y(u2__abc_44228_n17151) );
  OR2X2 OR2X2_4111 ( .A(u2__abc_44228_n17153), .B(u2__abc_44228_n17155), .Y(u2__abc_44228_n17156) );
  OR2X2 OR2X2_4112 ( .A(u2__abc_44228_n17158), .B(u2__abc_44228_n17160), .Y(u2__abc_44228_n17161) );
  OR2X2 OR2X2_4113 ( .A(u2__abc_44228_n17163), .B(u2__abc_44228_n17165), .Y(u2__abc_44228_n17166) );
  OR2X2 OR2X2_4114 ( .A(u2__abc_44228_n17168), .B(u2__abc_44228_n17170), .Y(u2__abc_44228_n17171) );
  OR2X2 OR2X2_4115 ( .A(u2__abc_44228_n17173), .B(u2__abc_44228_n17175), .Y(u2__abc_44228_n17176) );
  OR2X2 OR2X2_4116 ( .A(u2__abc_44228_n17178), .B(u2__abc_44228_n17180), .Y(u2__abc_44228_n17181) );
  OR2X2 OR2X2_4117 ( .A(u2__abc_44228_n17183), .B(u2__abc_44228_n17185), .Y(u2__abc_44228_n17186) );
  OR2X2 OR2X2_4118 ( .A(u2__abc_44228_n17188), .B(u2__abc_44228_n17190), .Y(u2__abc_44228_n17191) );
  OR2X2 OR2X2_4119 ( .A(u2__abc_44228_n17193), .B(u2__abc_44228_n17195), .Y(u2__abc_44228_n17196) );
  OR2X2 OR2X2_412 ( .A(a_112_bF_buf4), .B(\a[93] ), .Y(_abc_64468_n1449) );
  OR2X2 OR2X2_4120 ( .A(u2__abc_44228_n17198), .B(u2__abc_44228_n17200), .Y(u2__abc_44228_n17201) );
  OR2X2 OR2X2_4121 ( .A(u2__abc_44228_n17203), .B(u2__abc_44228_n17205), .Y(u2__abc_44228_n17206) );
  OR2X2 OR2X2_4122 ( .A(u2__abc_44228_n17208), .B(u2__abc_44228_n17210), .Y(u2__abc_44228_n17211) );
  OR2X2 OR2X2_4123 ( .A(u2__abc_44228_n17213), .B(u2__abc_44228_n17215), .Y(u2__abc_44228_n17216) );
  OR2X2 OR2X2_4124 ( .A(u2__abc_44228_n17218), .B(u2__abc_44228_n17220), .Y(u2__abc_44228_n17221) );
  OR2X2 OR2X2_4125 ( .A(u2__abc_44228_n17223), .B(u2__abc_44228_n17225), .Y(u2__abc_44228_n17226) );
  OR2X2 OR2X2_4126 ( .A(u2__abc_44228_n17228), .B(u2__abc_44228_n17230), .Y(u2__abc_44228_n17231) );
  OR2X2 OR2X2_4127 ( .A(u2__abc_44228_n17233), .B(u2__abc_44228_n17235), .Y(u2__abc_44228_n17236) );
  OR2X2 OR2X2_4128 ( .A(u2__abc_44228_n17238), .B(u2__abc_44228_n17240), .Y(u2__abc_44228_n17241) );
  OR2X2 OR2X2_4129 ( .A(u2__abc_44228_n17243), .B(u2__abc_44228_n17245), .Y(u2__abc_44228_n17246) );
  OR2X2 OR2X2_413 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[94] ), .Y(_abc_64468_n1450) );
  OR2X2 OR2X2_4130 ( .A(u2__abc_44228_n17248), .B(u2__abc_44228_n17250), .Y(u2__abc_44228_n17251) );
  OR2X2 OR2X2_4131 ( .A(u2__abc_44228_n17253), .B(u2__abc_44228_n17255), .Y(u2__abc_44228_n17256) );
  OR2X2 OR2X2_4132 ( .A(u2__abc_44228_n17258), .B(u2__abc_44228_n17260), .Y(u2__abc_44228_n17261) );
  OR2X2 OR2X2_4133 ( .A(u2__abc_44228_n17263), .B(u2__abc_44228_n17265), .Y(u2__abc_44228_n17266) );
  OR2X2 OR2X2_4134 ( .A(u2__abc_44228_n17268), .B(u2__abc_44228_n17270), .Y(u2__abc_44228_n17271) );
  OR2X2 OR2X2_4135 ( .A(u2__abc_44228_n17273), .B(u2__abc_44228_n17275), .Y(u2__abc_44228_n17276) );
  OR2X2 OR2X2_4136 ( .A(u2__abc_44228_n17278), .B(u2__abc_44228_n17280), .Y(u2__abc_44228_n17281) );
  OR2X2 OR2X2_4137 ( .A(u2__abc_44228_n17283), .B(u2__abc_44228_n17285), .Y(u2__abc_44228_n17286) );
  OR2X2 OR2X2_4138 ( .A(u2__abc_44228_n17288), .B(u2__abc_44228_n17290), .Y(u2__abc_44228_n17291) );
  OR2X2 OR2X2_4139 ( .A(u2__abc_44228_n17293), .B(u2__abc_44228_n17295), .Y(u2__abc_44228_n17296) );
  OR2X2 OR2X2_414 ( .A(a_112_bF_buf3), .B(\a[94] ), .Y(_abc_64468_n1452) );
  OR2X2 OR2X2_4140 ( .A(u2__abc_44228_n17298), .B(u2__abc_44228_n17300), .Y(u2__abc_44228_n17301) );
  OR2X2 OR2X2_4141 ( .A(u2__abc_44228_n17303), .B(u2__abc_44228_n17305), .Y(u2__abc_44228_n17306) );
  OR2X2 OR2X2_4142 ( .A(u2__abc_44228_n17308), .B(u2__abc_44228_n17310), .Y(u2__abc_44228_n17311) );
  OR2X2 OR2X2_4143 ( .A(u2__abc_44228_n17313), .B(u2__abc_44228_n17315), .Y(u2__abc_44228_n17316) );
  OR2X2 OR2X2_4144 ( .A(u2__abc_44228_n17318), .B(u2__abc_44228_n17320), .Y(u2__abc_44228_n17321) );
  OR2X2 OR2X2_4145 ( .A(u2__abc_44228_n17323), .B(u2__abc_44228_n17325), .Y(u2__abc_44228_n17326) );
  OR2X2 OR2X2_4146 ( .A(u2__abc_44228_n17328), .B(u2__abc_44228_n17330), .Y(u2__abc_44228_n17331) );
  OR2X2 OR2X2_4147 ( .A(u2__abc_44228_n17333), .B(u2__abc_44228_n17335), .Y(u2__abc_44228_n17336) );
  OR2X2 OR2X2_4148 ( .A(u2__abc_44228_n17338), .B(u2__abc_44228_n17340), .Y(u2__abc_44228_n17341) );
  OR2X2 OR2X2_4149 ( .A(u2__abc_44228_n17343), .B(u2__abc_44228_n17345), .Y(u2__abc_44228_n17346) );
  OR2X2 OR2X2_415 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[95] ), .Y(_abc_64468_n1453) );
  OR2X2 OR2X2_4150 ( .A(u2__abc_44228_n17348), .B(u2__abc_44228_n17350), .Y(u2__abc_44228_n17351) );
  OR2X2 OR2X2_4151 ( .A(u2__abc_44228_n17353), .B(u2__abc_44228_n17355), .Y(u2__abc_44228_n17356) );
  OR2X2 OR2X2_4152 ( .A(u2__abc_44228_n17358), .B(u2__abc_44228_n17360), .Y(u2__abc_44228_n17361) );
  OR2X2 OR2X2_4153 ( .A(u2__abc_44228_n17363), .B(u2__abc_44228_n17365), .Y(u2__abc_44228_n17366) );
  OR2X2 OR2X2_4154 ( .A(u2__abc_44228_n17368), .B(u2__abc_44228_n17370), .Y(u2__abc_44228_n17371) );
  OR2X2 OR2X2_4155 ( .A(u2__abc_44228_n17373), .B(u2__abc_44228_n17375), .Y(u2__abc_44228_n17376) );
  OR2X2 OR2X2_4156 ( .A(u2__abc_44228_n17378), .B(u2__abc_44228_n17380), .Y(u2__abc_44228_n17381) );
  OR2X2 OR2X2_4157 ( .A(u2__abc_44228_n17383), .B(u2__abc_44228_n17385), .Y(u2__abc_44228_n17386) );
  OR2X2 OR2X2_4158 ( .A(u2__abc_44228_n17388), .B(u2__abc_44228_n17390), .Y(u2__abc_44228_n17391) );
  OR2X2 OR2X2_4159 ( .A(u2__abc_44228_n17393), .B(u2__abc_44228_n17395), .Y(u2__abc_44228_n17396) );
  OR2X2 OR2X2_416 ( .A(a_112_bF_buf2), .B(\a[95] ), .Y(_abc_64468_n1455) );
  OR2X2 OR2X2_4160 ( .A(u2__abc_44228_n17398), .B(u2__abc_44228_n17400), .Y(u2__abc_44228_n17401) );
  OR2X2 OR2X2_4161 ( .A(u2__abc_44228_n17403), .B(u2__abc_44228_n17405), .Y(u2__abc_44228_n17406) );
  OR2X2 OR2X2_4162 ( .A(u2__abc_44228_n17408), .B(u2__abc_44228_n17410), .Y(u2__abc_44228_n17411) );
  OR2X2 OR2X2_4163 ( .A(u2__abc_44228_n17413), .B(u2__abc_44228_n17415), .Y(u2__abc_44228_n17416) );
  OR2X2 OR2X2_4164 ( .A(u2__abc_44228_n17418), .B(u2__abc_44228_n17420), .Y(u2__abc_44228_n17421) );
  OR2X2 OR2X2_4165 ( .A(u2__abc_44228_n17423), .B(u2__abc_44228_n17425), .Y(u2__abc_44228_n17426) );
  OR2X2 OR2X2_4166 ( .A(u2__abc_44228_n17428), .B(u2__abc_44228_n17430), .Y(u2__abc_44228_n17431) );
  OR2X2 OR2X2_4167 ( .A(u2__abc_44228_n17433), .B(u2__abc_44228_n17435), .Y(u2__abc_44228_n17436) );
  OR2X2 OR2X2_4168 ( .A(u2__abc_44228_n17438), .B(u2__abc_44228_n17440), .Y(u2__abc_44228_n17441) );
  OR2X2 OR2X2_4169 ( .A(u2__abc_44228_n17443), .B(u2__abc_44228_n17445), .Y(u2__abc_44228_n17446) );
  OR2X2 OR2X2_417 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[96] ), .Y(_abc_64468_n1456) );
  OR2X2 OR2X2_4170 ( .A(u2__abc_44228_n17448), .B(u2__abc_44228_n17450), .Y(u2__abc_44228_n17451) );
  OR2X2 OR2X2_4171 ( .A(u2__abc_44228_n17453), .B(u2__abc_44228_n17455), .Y(u2__abc_44228_n17456) );
  OR2X2 OR2X2_4172 ( .A(u2__abc_44228_n17458), .B(u2__abc_44228_n17460), .Y(u2__abc_44228_n17461) );
  OR2X2 OR2X2_4173 ( .A(u2__abc_44228_n17463), .B(u2__abc_44228_n17465), .Y(u2__abc_44228_n17466) );
  OR2X2 OR2X2_4174 ( .A(u2__abc_44228_n17468), .B(u2__abc_44228_n17470), .Y(u2__abc_44228_n17471) );
  OR2X2 OR2X2_4175 ( .A(u2__abc_44228_n17473), .B(u2__abc_44228_n17475), .Y(u2__abc_44228_n17476) );
  OR2X2 OR2X2_4176 ( .A(u2__abc_44228_n17478), .B(u2__abc_44228_n17480), .Y(u2__abc_44228_n17481) );
  OR2X2 OR2X2_4177 ( .A(u2__abc_44228_n17483), .B(u2__abc_44228_n17485), .Y(u2__abc_44228_n17486) );
  OR2X2 OR2X2_4178 ( .A(u2__abc_44228_n17488), .B(u2__abc_44228_n17490), .Y(u2__abc_44228_n17491) );
  OR2X2 OR2X2_4179 ( .A(u2__abc_44228_n17493), .B(u2__abc_44228_n17495), .Y(u2__abc_44228_n17496) );
  OR2X2 OR2X2_418 ( .A(a_112_bF_buf1), .B(\a[96] ), .Y(_abc_64468_n1458) );
  OR2X2 OR2X2_4180 ( .A(u2__abc_44228_n17498), .B(u2__abc_44228_n17500), .Y(u2__abc_44228_n17501) );
  OR2X2 OR2X2_4181 ( .A(u2__abc_44228_n17503), .B(u2__abc_44228_n17505), .Y(u2__abc_44228_n17506) );
  OR2X2 OR2X2_4182 ( .A(u2__abc_44228_n17508), .B(u2__abc_44228_n17510), .Y(u2__abc_44228_n17511) );
  OR2X2 OR2X2_4183 ( .A(u2__abc_44228_n17513), .B(u2__abc_44228_n17515), .Y(u2__abc_44228_n17516) );
  OR2X2 OR2X2_4184 ( .A(u2__abc_44228_n17518), .B(u2__abc_44228_n17520), .Y(u2__abc_44228_n17521) );
  OR2X2 OR2X2_4185 ( .A(u2__abc_44228_n17523), .B(u2__abc_44228_n17525), .Y(u2__abc_44228_n17526) );
  OR2X2 OR2X2_4186 ( .A(u2__abc_44228_n17528), .B(u2__abc_44228_n17530), .Y(u2__abc_44228_n17531) );
  OR2X2 OR2X2_4187 ( .A(u2__abc_44228_n17533), .B(u2__abc_44228_n17535), .Y(u2__abc_44228_n17536) );
  OR2X2 OR2X2_4188 ( .A(u2__abc_44228_n17538), .B(u2__abc_44228_n17540), .Y(u2__abc_44228_n17541) );
  OR2X2 OR2X2_4189 ( .A(u2__abc_44228_n17543), .B(u2__abc_44228_n17545), .Y(u2__abc_44228_n17546) );
  OR2X2 OR2X2_419 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[97] ), .Y(_abc_64468_n1459) );
  OR2X2 OR2X2_4190 ( .A(u2__abc_44228_n17548), .B(u2__abc_44228_n17550), .Y(u2__abc_44228_n17551) );
  OR2X2 OR2X2_4191 ( .A(u2__abc_44228_n17553), .B(u2__abc_44228_n17555), .Y(u2__abc_44228_n17556) );
  OR2X2 OR2X2_4192 ( .A(u2__abc_44228_n17558), .B(u2__abc_44228_n17560), .Y(u2__abc_44228_n17561) );
  OR2X2 OR2X2_4193 ( .A(u2__abc_44228_n17563), .B(u2__abc_44228_n17565), .Y(u2__abc_44228_n17566) );
  OR2X2 OR2X2_4194 ( .A(u2__abc_44228_n17568), .B(u2__abc_44228_n17570), .Y(u2__abc_44228_n17571) );
  OR2X2 OR2X2_4195 ( .A(u2__abc_44228_n17573), .B(u2__abc_44228_n17575), .Y(u2__abc_44228_n17576) );
  OR2X2 OR2X2_4196 ( .A(u2__abc_44228_n17578), .B(u2__abc_44228_n17580), .Y(u2__abc_44228_n17581) );
  OR2X2 OR2X2_4197 ( .A(u2__abc_44228_n17583), .B(u2__abc_44228_n17585), .Y(u2__abc_44228_n17586) );
  OR2X2 OR2X2_4198 ( .A(u2__abc_44228_n17588), .B(u2__abc_44228_n17590), .Y(u2__abc_44228_n17591) );
  OR2X2 OR2X2_4199 ( .A(u2__abc_44228_n17593), .B(u2__abc_44228_n17595), .Y(u2__abc_44228_n17596) );
  OR2X2 OR2X2_42 ( .A(_abc_64468_n753_bF_buf1), .B(\a[20] ), .Y(_abc_64468_n891) );
  OR2X2 OR2X2_420 ( .A(a_112_bF_buf0), .B(\a[97] ), .Y(_abc_64468_n1461) );
  OR2X2 OR2X2_4200 ( .A(u2__abc_44228_n17598), .B(u2__abc_44228_n17600), .Y(u2__abc_44228_n17601) );
  OR2X2 OR2X2_4201 ( .A(u2__abc_44228_n17603), .B(u2__abc_44228_n17605), .Y(u2__abc_44228_n17606) );
  OR2X2 OR2X2_4202 ( .A(u2__abc_44228_n17608), .B(u2__abc_44228_n17610), .Y(u2__abc_44228_n17611) );
  OR2X2 OR2X2_4203 ( .A(u2__abc_44228_n17613), .B(u2__abc_44228_n17615), .Y(u2__abc_44228_n17616) );
  OR2X2 OR2X2_4204 ( .A(u2__abc_44228_n17618), .B(u2__abc_44228_n17620), .Y(u2__abc_44228_n17621) );
  OR2X2 OR2X2_4205 ( .A(u2__abc_44228_n17623), .B(u2__abc_44228_n17625), .Y(u2__abc_44228_n17626) );
  OR2X2 OR2X2_4206 ( .A(u2__abc_44228_n17628), .B(u2__abc_44228_n17630), .Y(u2__abc_44228_n17631) );
  OR2X2 OR2X2_4207 ( .A(u2__abc_44228_n17633), .B(u2__abc_44228_n17635), .Y(u2__abc_44228_n17636) );
  OR2X2 OR2X2_4208 ( .A(u2__abc_44228_n17638), .B(u2__abc_44228_n17640), .Y(u2__abc_44228_n17641) );
  OR2X2 OR2X2_4209 ( .A(u2__abc_44228_n17643), .B(u2__abc_44228_n17645), .Y(u2__abc_44228_n17646) );
  OR2X2 OR2X2_421 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[98] ), .Y(_abc_64468_n1462) );
  OR2X2 OR2X2_4210 ( .A(u2__abc_44228_n17648), .B(u2__abc_44228_n17650), .Y(u2__abc_44228_n17651) );
  OR2X2 OR2X2_4211 ( .A(u2__abc_44228_n17653), .B(u2__abc_44228_n17655), .Y(u2__abc_44228_n17656) );
  OR2X2 OR2X2_4212 ( .A(u2__abc_44228_n17658), .B(u2__abc_44228_n17660), .Y(u2__abc_44228_n17661) );
  OR2X2 OR2X2_4213 ( .A(u2__abc_44228_n17663), .B(u2__abc_44228_n17665), .Y(u2__abc_44228_n17666) );
  OR2X2 OR2X2_4214 ( .A(u2__abc_44228_n17668), .B(u2__abc_44228_n17670), .Y(u2__abc_44228_n17671) );
  OR2X2 OR2X2_4215 ( .A(u2__abc_44228_n17673), .B(u2__abc_44228_n17675), .Y(u2__abc_44228_n17676) );
  OR2X2 OR2X2_4216 ( .A(u2__abc_44228_n17678), .B(u2__abc_44228_n17680), .Y(u2__abc_44228_n17681) );
  OR2X2 OR2X2_4217 ( .A(u2__abc_44228_n17683), .B(u2__abc_44228_n17685), .Y(u2__abc_44228_n17686) );
  OR2X2 OR2X2_4218 ( .A(u2__abc_44228_n17688), .B(u2__abc_44228_n17690), .Y(u2__abc_44228_n17691) );
  OR2X2 OR2X2_4219 ( .A(u2__abc_44228_n17693), .B(u2__abc_44228_n17695), .Y(u2__abc_44228_n17696) );
  OR2X2 OR2X2_422 ( .A(a_112_bF_buf9), .B(\a[98] ), .Y(_abc_64468_n1464) );
  OR2X2 OR2X2_4220 ( .A(u2__abc_44228_n17698), .B(u2__abc_44228_n17700), .Y(u2__abc_44228_n17701) );
  OR2X2 OR2X2_4221 ( .A(u2__abc_44228_n17703), .B(u2__abc_44228_n17705), .Y(u2__abc_44228_n17706) );
  OR2X2 OR2X2_4222 ( .A(u2__abc_44228_n17708), .B(u2__abc_44228_n17710), .Y(u2__abc_44228_n17711) );
  OR2X2 OR2X2_4223 ( .A(u2__abc_44228_n17713), .B(u2__abc_44228_n17715), .Y(u2__abc_44228_n17716) );
  OR2X2 OR2X2_4224 ( .A(u2__abc_44228_n17718), .B(u2__abc_44228_n17720), .Y(u2__abc_44228_n17721) );
  OR2X2 OR2X2_4225 ( .A(u2__abc_44228_n17723), .B(u2__abc_44228_n17725), .Y(u2__abc_44228_n17726) );
  OR2X2 OR2X2_4226 ( .A(u2__abc_44228_n17728), .B(u2__abc_44228_n17730), .Y(u2__abc_44228_n17731) );
  OR2X2 OR2X2_4227 ( .A(u2__abc_44228_n17733), .B(u2__abc_44228_n17735), .Y(u2__abc_44228_n17736) );
  OR2X2 OR2X2_4228 ( .A(u2__abc_44228_n17738), .B(u2__abc_44228_n17740), .Y(u2__abc_44228_n17741) );
  OR2X2 OR2X2_4229 ( .A(u2__abc_44228_n17743), .B(u2__abc_44228_n17745), .Y(u2__abc_44228_n17746) );
  OR2X2 OR2X2_423 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[99] ), .Y(_abc_64468_n1465) );
  OR2X2 OR2X2_4230 ( .A(u2__abc_44228_n17748), .B(u2__abc_44228_n17750), .Y(u2__abc_44228_n17751) );
  OR2X2 OR2X2_4231 ( .A(u2__abc_44228_n17753), .B(u2__abc_44228_n17755), .Y(u2__abc_44228_n17756) );
  OR2X2 OR2X2_4232 ( .A(u2__abc_44228_n17758), .B(u2__abc_44228_n17760), .Y(u2__abc_44228_n17761) );
  OR2X2 OR2X2_4233 ( .A(u2__abc_44228_n17763), .B(u2__abc_44228_n17765), .Y(u2__abc_44228_n17766) );
  OR2X2 OR2X2_4234 ( .A(u2__abc_44228_n17768), .B(u2__abc_44228_n17770), .Y(u2__abc_44228_n17771) );
  OR2X2 OR2X2_4235 ( .A(u2__abc_44228_n7547_bF_buf11), .B(u2_root_0_), .Y(u2__abc_44228_n17778) );
  OR2X2 OR2X2_4236 ( .A(u2__abc_44228_n17779), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n17780) );
  OR2X2 OR2X2_4237 ( .A(u2__abc_44228_n17784), .B(u2__abc_44228_n17775), .Y(u2__abc_44228_n17785) );
  OR2X2 OR2X2_4238 ( .A(u2__abc_44228_n17776), .B(sqrto_0_), .Y(u2__abc_44228_n17788) );
  OR2X2 OR2X2_4239 ( .A(u2__abc_44228_n17791), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n17792) );
  OR2X2 OR2X2_424 ( .A(a_112_bF_buf8), .B(\a[99] ), .Y(_abc_64468_n1467) );
  OR2X2 OR2X2_4240 ( .A(u2__abc_44228_n17796), .B(u2__abc_44228_n17787), .Y(u2__abc_44228_n17797) );
  OR2X2 OR2X2_4241 ( .A(u2__abc_44228_n17789), .B(sqrto_1_), .Y(u2__abc_44228_n17800) );
  OR2X2 OR2X2_4242 ( .A(u2__abc_44228_n17803), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n17804) );
  OR2X2 OR2X2_4243 ( .A(u2__abc_44228_n17808), .B(u2__abc_44228_n17799), .Y(u2__abc_44228_n17809) );
  OR2X2 OR2X2_4244 ( .A(u2__abc_44228_n17801), .B(sqrto_2_), .Y(u2__abc_44228_n17812) );
  OR2X2 OR2X2_4245 ( .A(u2__abc_44228_n17815), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n17816) );
  OR2X2 OR2X2_4246 ( .A(u2__abc_44228_n17820), .B(u2__abc_44228_n17811), .Y(u2__abc_44228_n17821) );
  OR2X2 OR2X2_4247 ( .A(u2__abc_44228_n17813), .B(sqrto_3_), .Y(u2__abc_44228_n17824) );
  OR2X2 OR2X2_4248 ( .A(u2__abc_44228_n17827), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n17828) );
  OR2X2 OR2X2_4249 ( .A(u2__abc_44228_n17832), .B(u2__abc_44228_n17823), .Y(u2__abc_44228_n17833) );
  OR2X2 OR2X2_425 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[100] ), .Y(_abc_64468_n1468) );
  OR2X2 OR2X2_4250 ( .A(u2__abc_44228_n17825), .B(sqrto_4_), .Y(u2__abc_44228_n17836) );
  OR2X2 OR2X2_4251 ( .A(u2__abc_44228_n17839), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n17840) );
  OR2X2 OR2X2_4252 ( .A(u2__abc_44228_n17844), .B(u2__abc_44228_n17835), .Y(u2__abc_44228_n17845) );
  OR2X2 OR2X2_4253 ( .A(u2__abc_44228_n17837), .B(sqrto_5_), .Y(u2__abc_44228_n17848) );
  OR2X2 OR2X2_4254 ( .A(u2__abc_44228_n17851), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n17852) );
  OR2X2 OR2X2_4255 ( .A(u2__abc_44228_n17856), .B(u2__abc_44228_n17847), .Y(u2__abc_44228_n17857) );
  OR2X2 OR2X2_4256 ( .A(u2__abc_44228_n17849), .B(sqrto_6_), .Y(u2__abc_44228_n17860) );
  OR2X2 OR2X2_4257 ( .A(u2__abc_44228_n17863), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n17864) );
  OR2X2 OR2X2_4258 ( .A(u2__abc_44228_n17868), .B(u2__abc_44228_n17859), .Y(u2__abc_44228_n17869) );
  OR2X2 OR2X2_4259 ( .A(u2__abc_44228_n17861), .B(sqrto_7_), .Y(u2__abc_44228_n17872) );
  OR2X2 OR2X2_426 ( .A(a_112_bF_buf7), .B(\a[100] ), .Y(_abc_64468_n1470) );
  OR2X2 OR2X2_4260 ( .A(u2__abc_44228_n17875), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n17876) );
  OR2X2 OR2X2_4261 ( .A(u2__abc_44228_n17880), .B(u2__abc_44228_n17871), .Y(u2__abc_44228_n17881) );
  OR2X2 OR2X2_4262 ( .A(u2__abc_44228_n17873), .B(sqrto_8_), .Y(u2__abc_44228_n17884) );
  OR2X2 OR2X2_4263 ( .A(u2__abc_44228_n17887), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n17888) );
  OR2X2 OR2X2_4264 ( .A(u2__abc_44228_n17892), .B(u2__abc_44228_n17883), .Y(u2__abc_44228_n17893) );
  OR2X2 OR2X2_4265 ( .A(u2__abc_44228_n17885), .B(sqrto_9_), .Y(u2__abc_44228_n17896) );
  OR2X2 OR2X2_4266 ( .A(u2__abc_44228_n17899), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n17900) );
  OR2X2 OR2X2_4267 ( .A(u2__abc_44228_n17904), .B(u2__abc_44228_n17895), .Y(u2__abc_44228_n17905) );
  OR2X2 OR2X2_4268 ( .A(u2__abc_44228_n17897), .B(sqrto_10_), .Y(u2__abc_44228_n17908) );
  OR2X2 OR2X2_4269 ( .A(u2__abc_44228_n17911), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n17912) );
  OR2X2 OR2X2_427 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[101] ), .Y(_abc_64468_n1471) );
  OR2X2 OR2X2_4270 ( .A(u2__abc_44228_n17916), .B(u2__abc_44228_n17907), .Y(u2__abc_44228_n17917) );
  OR2X2 OR2X2_4271 ( .A(u2__abc_44228_n17909), .B(sqrto_11_), .Y(u2__abc_44228_n17920) );
  OR2X2 OR2X2_4272 ( .A(u2__abc_44228_n17923), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n17924) );
  OR2X2 OR2X2_4273 ( .A(u2__abc_44228_n17928), .B(u2__abc_44228_n17919), .Y(u2__abc_44228_n17929) );
  OR2X2 OR2X2_4274 ( .A(u2__abc_44228_n17921), .B(sqrto_12_), .Y(u2__abc_44228_n17932) );
  OR2X2 OR2X2_4275 ( .A(u2__abc_44228_n17935), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n17936) );
  OR2X2 OR2X2_4276 ( .A(u2__abc_44228_n17940), .B(u2__abc_44228_n17931), .Y(u2__abc_44228_n17941) );
  OR2X2 OR2X2_4277 ( .A(u2__abc_44228_n17933), .B(sqrto_13_), .Y(u2__abc_44228_n17944) );
  OR2X2 OR2X2_4278 ( .A(u2__abc_44228_n17947), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n17948) );
  OR2X2 OR2X2_4279 ( .A(u2__abc_44228_n17952), .B(u2__abc_44228_n17943), .Y(u2__abc_44228_n17953) );
  OR2X2 OR2X2_428 ( .A(a_112_bF_buf6), .B(\a[101] ), .Y(_abc_64468_n1473) );
  OR2X2 OR2X2_4280 ( .A(u2__abc_44228_n17945), .B(sqrto_14_), .Y(u2__abc_44228_n17956) );
  OR2X2 OR2X2_4281 ( .A(u2__abc_44228_n17959), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n17960) );
  OR2X2 OR2X2_4282 ( .A(u2__abc_44228_n17964), .B(u2__abc_44228_n17955), .Y(u2__abc_44228_n17965) );
  OR2X2 OR2X2_4283 ( .A(u2__abc_44228_n17957), .B(sqrto_15_), .Y(u2__abc_44228_n17968) );
  OR2X2 OR2X2_4284 ( .A(u2__abc_44228_n17971), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n17972) );
  OR2X2 OR2X2_4285 ( .A(u2__abc_44228_n17976), .B(u2__abc_44228_n17967), .Y(u2__abc_44228_n17977) );
  OR2X2 OR2X2_4286 ( .A(u2__abc_44228_n17969), .B(sqrto_16_), .Y(u2__abc_44228_n17980) );
  OR2X2 OR2X2_4287 ( .A(u2__abc_44228_n17983), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n17984) );
  OR2X2 OR2X2_4288 ( .A(u2__abc_44228_n17988), .B(u2__abc_44228_n17979), .Y(u2__abc_44228_n17989) );
  OR2X2 OR2X2_4289 ( .A(u2__abc_44228_n17981), .B(sqrto_17_), .Y(u2__abc_44228_n17992) );
  OR2X2 OR2X2_429 ( .A(_abc_64468_n1170_bF_buf8), .B(\a[102] ), .Y(_abc_64468_n1474) );
  OR2X2 OR2X2_4290 ( .A(u2__abc_44228_n17995), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n17996) );
  OR2X2 OR2X2_4291 ( .A(u2__abc_44228_n18000), .B(u2__abc_44228_n17991), .Y(u2__abc_44228_n18001) );
  OR2X2 OR2X2_4292 ( .A(u2__abc_44228_n17993), .B(sqrto_18_), .Y(u2__abc_44228_n18004) );
  OR2X2 OR2X2_4293 ( .A(u2__abc_44228_n18007), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n18008) );
  OR2X2 OR2X2_4294 ( .A(u2__abc_44228_n18012), .B(u2__abc_44228_n18003), .Y(u2__abc_44228_n18013) );
  OR2X2 OR2X2_4295 ( .A(u2__abc_44228_n18005), .B(sqrto_19_), .Y(u2__abc_44228_n18016) );
  OR2X2 OR2X2_4296 ( .A(u2__abc_44228_n18019), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n18020) );
  OR2X2 OR2X2_4297 ( .A(u2__abc_44228_n18024), .B(u2__abc_44228_n18015), .Y(u2__abc_44228_n18025) );
  OR2X2 OR2X2_4298 ( .A(u2__abc_44228_n18017), .B(sqrto_20_), .Y(u2__abc_44228_n18028) );
  OR2X2 OR2X2_4299 ( .A(u2__abc_44228_n18031), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n18032) );
  OR2X2 OR2X2_43 ( .A(aNan_bF_buf10), .B(sqrto_97_), .Y(_abc_64468_n893) );
  OR2X2 OR2X2_430 ( .A(a_112_bF_buf5), .B(\a[102] ), .Y(_abc_64468_n1476) );
  OR2X2 OR2X2_4300 ( .A(u2__abc_44228_n18036), .B(u2__abc_44228_n18027), .Y(u2__abc_44228_n18037) );
  OR2X2 OR2X2_4301 ( .A(u2__abc_44228_n18029), .B(sqrto_21_), .Y(u2__abc_44228_n18040) );
  OR2X2 OR2X2_4302 ( .A(u2__abc_44228_n18043), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n18044) );
  OR2X2 OR2X2_4303 ( .A(u2__abc_44228_n18048), .B(u2__abc_44228_n18039), .Y(u2__abc_44228_n18049) );
  OR2X2 OR2X2_4304 ( .A(u2__abc_44228_n18041), .B(sqrto_22_), .Y(u2__abc_44228_n18052) );
  OR2X2 OR2X2_4305 ( .A(u2__abc_44228_n18055), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n18056) );
  OR2X2 OR2X2_4306 ( .A(u2__abc_44228_n18060), .B(u2__abc_44228_n18051), .Y(u2__abc_44228_n18061) );
  OR2X2 OR2X2_4307 ( .A(u2__abc_44228_n18053), .B(sqrto_23_), .Y(u2__abc_44228_n18064) );
  OR2X2 OR2X2_4308 ( .A(u2__abc_44228_n18067), .B(u2__abc_44228_n2983_bF_buf1), .Y(u2__abc_44228_n18068) );
  OR2X2 OR2X2_4309 ( .A(u2__abc_44228_n18072), .B(u2__abc_44228_n18063), .Y(u2__abc_44228_n18073) );
  OR2X2 OR2X2_431 ( .A(_abc_64468_n1170_bF_buf7), .B(\a[103] ), .Y(_abc_64468_n1477) );
  OR2X2 OR2X2_4310 ( .A(u2__abc_44228_n18065), .B(sqrto_24_), .Y(u2__abc_44228_n18076) );
  OR2X2 OR2X2_4311 ( .A(u2__abc_44228_n18079), .B(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n18080) );
  OR2X2 OR2X2_4312 ( .A(u2__abc_44228_n18084), .B(u2__abc_44228_n18075), .Y(u2__abc_44228_n18085) );
  OR2X2 OR2X2_4313 ( .A(u2__abc_44228_n18077), .B(sqrto_25_), .Y(u2__abc_44228_n18088) );
  OR2X2 OR2X2_4314 ( .A(u2__abc_44228_n18091), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n18092) );
  OR2X2 OR2X2_4315 ( .A(u2__abc_44228_n18096), .B(u2__abc_44228_n18087), .Y(u2__abc_44228_n18097) );
  OR2X2 OR2X2_4316 ( .A(u2__abc_44228_n18089), .B(sqrto_26_), .Y(u2__abc_44228_n18100) );
  OR2X2 OR2X2_4317 ( .A(u2__abc_44228_n18103), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n18104) );
  OR2X2 OR2X2_4318 ( .A(u2__abc_44228_n18108), .B(u2__abc_44228_n18099), .Y(u2__abc_44228_n18109) );
  OR2X2 OR2X2_4319 ( .A(u2__abc_44228_n18101), .B(sqrto_27_), .Y(u2__abc_44228_n18112) );
  OR2X2 OR2X2_432 ( .A(a_112_bF_buf4), .B(\a[103] ), .Y(_abc_64468_n1479) );
  OR2X2 OR2X2_4320 ( .A(u2__abc_44228_n18115), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n18116) );
  OR2X2 OR2X2_4321 ( .A(u2__abc_44228_n18120), .B(u2__abc_44228_n18111), .Y(u2__abc_44228_n18121) );
  OR2X2 OR2X2_4322 ( .A(u2__abc_44228_n18113), .B(sqrto_28_), .Y(u2__abc_44228_n18124) );
  OR2X2 OR2X2_4323 ( .A(u2__abc_44228_n18127), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n18128) );
  OR2X2 OR2X2_4324 ( .A(u2__abc_44228_n18132), .B(u2__abc_44228_n18123), .Y(u2__abc_44228_n18133) );
  OR2X2 OR2X2_4325 ( .A(u2__abc_44228_n18125), .B(sqrto_29_), .Y(u2__abc_44228_n18136) );
  OR2X2 OR2X2_4326 ( .A(u2__abc_44228_n18139), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n18140) );
  OR2X2 OR2X2_4327 ( .A(u2__abc_44228_n18144), .B(u2__abc_44228_n18135), .Y(u2__abc_44228_n18145) );
  OR2X2 OR2X2_4328 ( .A(u2__abc_44228_n18137), .B(sqrto_30_), .Y(u2__abc_44228_n18148) );
  OR2X2 OR2X2_4329 ( .A(u2__abc_44228_n18151), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n18152) );
  OR2X2 OR2X2_433 ( .A(_abc_64468_n1170_bF_buf6), .B(\a[104] ), .Y(_abc_64468_n1480) );
  OR2X2 OR2X2_4330 ( .A(u2__abc_44228_n18156), .B(u2__abc_44228_n18147), .Y(u2__abc_44228_n18157) );
  OR2X2 OR2X2_4331 ( .A(u2__abc_44228_n18149), .B(sqrto_31_), .Y(u2__abc_44228_n18160) );
  OR2X2 OR2X2_4332 ( .A(u2__abc_44228_n18163), .B(u2__abc_44228_n2983_bF_buf127), .Y(u2__abc_44228_n18164) );
  OR2X2 OR2X2_4333 ( .A(u2__abc_44228_n18168), .B(u2__abc_44228_n18159), .Y(u2__abc_44228_n18169) );
  OR2X2 OR2X2_4334 ( .A(u2__abc_44228_n18161), .B(sqrto_32_), .Y(u2__abc_44228_n18172) );
  OR2X2 OR2X2_4335 ( .A(u2__abc_44228_n18175), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n18176) );
  OR2X2 OR2X2_4336 ( .A(u2__abc_44228_n18180), .B(u2__abc_44228_n18171), .Y(u2__abc_44228_n18181) );
  OR2X2 OR2X2_4337 ( .A(u2__abc_44228_n18173), .B(sqrto_33_), .Y(u2__abc_44228_n18184) );
  OR2X2 OR2X2_4338 ( .A(u2__abc_44228_n18187), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n18188) );
  OR2X2 OR2X2_4339 ( .A(u2__abc_44228_n18192), .B(u2__abc_44228_n18183), .Y(u2__abc_44228_n18193) );
  OR2X2 OR2X2_434 ( .A(a_112_bF_buf3), .B(\a[104] ), .Y(_abc_64468_n1482) );
  OR2X2 OR2X2_4340 ( .A(u2__abc_44228_n18185), .B(sqrto_34_), .Y(u2__abc_44228_n18196) );
  OR2X2 OR2X2_4341 ( .A(u2__abc_44228_n18199), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n18200) );
  OR2X2 OR2X2_4342 ( .A(u2__abc_44228_n18204), .B(u2__abc_44228_n18195), .Y(u2__abc_44228_n18205) );
  OR2X2 OR2X2_4343 ( .A(u2__abc_44228_n18197), .B(sqrto_35_), .Y(u2__abc_44228_n18208) );
  OR2X2 OR2X2_4344 ( .A(u2__abc_44228_n18211), .B(u2__abc_44228_n2983_bF_buf119), .Y(u2__abc_44228_n18212) );
  OR2X2 OR2X2_4345 ( .A(u2__abc_44228_n18216), .B(u2__abc_44228_n18207), .Y(u2__abc_44228_n18217) );
  OR2X2 OR2X2_4346 ( .A(u2__abc_44228_n18209), .B(sqrto_36_), .Y(u2__abc_44228_n18220) );
  OR2X2 OR2X2_4347 ( .A(u2__abc_44228_n18223), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n18224) );
  OR2X2 OR2X2_4348 ( .A(u2__abc_44228_n18228), .B(u2__abc_44228_n18219), .Y(u2__abc_44228_n18229) );
  OR2X2 OR2X2_4349 ( .A(u2__abc_44228_n18221), .B(sqrto_37_), .Y(u2__abc_44228_n18232) );
  OR2X2 OR2X2_435 ( .A(_abc_64468_n1170_bF_buf5), .B(\a[105] ), .Y(_abc_64468_n1483) );
  OR2X2 OR2X2_4350 ( .A(u2__abc_44228_n18235), .B(u2__abc_44228_n2983_bF_buf115), .Y(u2__abc_44228_n18236) );
  OR2X2 OR2X2_4351 ( .A(u2__abc_44228_n18240), .B(u2__abc_44228_n18231), .Y(u2__abc_44228_n18241) );
  OR2X2 OR2X2_4352 ( .A(u2__abc_44228_n18233), .B(sqrto_38_), .Y(u2__abc_44228_n18244) );
  OR2X2 OR2X2_4353 ( .A(u2__abc_44228_n18247), .B(u2__abc_44228_n2983_bF_buf113), .Y(u2__abc_44228_n18248) );
  OR2X2 OR2X2_4354 ( .A(u2__abc_44228_n18252), .B(u2__abc_44228_n18243), .Y(u2__abc_44228_n18253) );
  OR2X2 OR2X2_4355 ( .A(u2__abc_44228_n18245), .B(sqrto_39_), .Y(u2__abc_44228_n18256) );
  OR2X2 OR2X2_4356 ( .A(u2__abc_44228_n18259), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n18260) );
  OR2X2 OR2X2_4357 ( .A(u2__abc_44228_n18264), .B(u2__abc_44228_n18255), .Y(u2__abc_44228_n18265) );
  OR2X2 OR2X2_4358 ( .A(u2__abc_44228_n18257), .B(sqrto_40_), .Y(u2__abc_44228_n18268) );
  OR2X2 OR2X2_4359 ( .A(u2__abc_44228_n18271), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n18272) );
  OR2X2 OR2X2_436 ( .A(a_112_bF_buf2), .B(\a[105] ), .Y(_abc_64468_n1485) );
  OR2X2 OR2X2_4360 ( .A(u2__abc_44228_n18276), .B(u2__abc_44228_n18267), .Y(u2__abc_44228_n18277) );
  OR2X2 OR2X2_4361 ( .A(u2__abc_44228_n18269), .B(sqrto_41_), .Y(u2__abc_44228_n18280) );
  OR2X2 OR2X2_4362 ( .A(u2__abc_44228_n18283), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n18284) );
  OR2X2 OR2X2_4363 ( .A(u2__abc_44228_n18288), .B(u2__abc_44228_n18279), .Y(u2__abc_44228_n18289) );
  OR2X2 OR2X2_4364 ( .A(u2__abc_44228_n18281), .B(sqrto_42_), .Y(u2__abc_44228_n18292) );
  OR2X2 OR2X2_4365 ( .A(u2__abc_44228_n18295), .B(u2__abc_44228_n2983_bF_buf105), .Y(u2__abc_44228_n18296) );
  OR2X2 OR2X2_4366 ( .A(u2__abc_44228_n18300), .B(u2__abc_44228_n18291), .Y(u2__abc_44228_n18301) );
  OR2X2 OR2X2_4367 ( .A(u2__abc_44228_n18293), .B(sqrto_43_), .Y(u2__abc_44228_n18304) );
  OR2X2 OR2X2_4368 ( .A(u2__abc_44228_n18307), .B(u2__abc_44228_n2983_bF_buf103), .Y(u2__abc_44228_n18308) );
  OR2X2 OR2X2_4369 ( .A(u2__abc_44228_n18312), .B(u2__abc_44228_n18303), .Y(u2__abc_44228_n18313) );
  OR2X2 OR2X2_437 ( .A(_abc_64468_n1170_bF_buf4), .B(\a[106] ), .Y(_abc_64468_n1486) );
  OR2X2 OR2X2_4370 ( .A(u2__abc_44228_n18305), .B(sqrto_44_), .Y(u2__abc_44228_n18316) );
  OR2X2 OR2X2_4371 ( .A(u2__abc_44228_n18319), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n18320) );
  OR2X2 OR2X2_4372 ( .A(u2__abc_44228_n18324), .B(u2__abc_44228_n18315), .Y(u2__abc_44228_n18325) );
  OR2X2 OR2X2_4373 ( .A(u2__abc_44228_n18317), .B(sqrto_45_), .Y(u2__abc_44228_n18328) );
  OR2X2 OR2X2_4374 ( .A(u2__abc_44228_n18331), .B(u2__abc_44228_n2983_bF_buf99), .Y(u2__abc_44228_n18332) );
  OR2X2 OR2X2_4375 ( .A(u2__abc_44228_n18336), .B(u2__abc_44228_n18327), .Y(u2__abc_44228_n18337) );
  OR2X2 OR2X2_4376 ( .A(u2__abc_44228_n18329), .B(sqrto_46_), .Y(u2__abc_44228_n18340) );
  OR2X2 OR2X2_4377 ( .A(u2__abc_44228_n18343), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n18344) );
  OR2X2 OR2X2_4378 ( .A(u2__abc_44228_n18348), .B(u2__abc_44228_n18339), .Y(u2__abc_44228_n18349) );
  OR2X2 OR2X2_4379 ( .A(u2__abc_44228_n18341), .B(sqrto_47_), .Y(u2__abc_44228_n18352) );
  OR2X2 OR2X2_438 ( .A(a_112_bF_buf1), .B(\a[106] ), .Y(_abc_64468_n1488) );
  OR2X2 OR2X2_4380 ( .A(u2__abc_44228_n18355), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n18356) );
  OR2X2 OR2X2_4381 ( .A(u2__abc_44228_n18360), .B(u2__abc_44228_n18351), .Y(u2__abc_44228_n18361) );
  OR2X2 OR2X2_4382 ( .A(u2__abc_44228_n18353), .B(sqrto_48_), .Y(u2__abc_44228_n18364) );
  OR2X2 OR2X2_4383 ( .A(u2__abc_44228_n18367), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n18368) );
  OR2X2 OR2X2_4384 ( .A(u2__abc_44228_n18372), .B(u2__abc_44228_n18363), .Y(u2__abc_44228_n18373) );
  OR2X2 OR2X2_4385 ( .A(u2__abc_44228_n18365), .B(sqrto_49_), .Y(u2__abc_44228_n18376) );
  OR2X2 OR2X2_4386 ( .A(u2__abc_44228_n18379), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n18380) );
  OR2X2 OR2X2_4387 ( .A(u2__abc_44228_n18384), .B(u2__abc_44228_n18375), .Y(u2__abc_44228_n18385) );
  OR2X2 OR2X2_4388 ( .A(u2__abc_44228_n18377), .B(sqrto_50_), .Y(u2__abc_44228_n18388) );
  OR2X2 OR2X2_4389 ( .A(u2__abc_44228_n18391), .B(u2__abc_44228_n2983_bF_buf89), .Y(u2__abc_44228_n18392) );
  OR2X2 OR2X2_439 ( .A(_abc_64468_n1170_bF_buf3), .B(\a[107] ), .Y(_abc_64468_n1489) );
  OR2X2 OR2X2_4390 ( .A(u2__abc_44228_n18396), .B(u2__abc_44228_n18387), .Y(u2__abc_44228_n18397) );
  OR2X2 OR2X2_4391 ( .A(u2__abc_44228_n18389), .B(sqrto_51_), .Y(u2__abc_44228_n18400) );
  OR2X2 OR2X2_4392 ( .A(u2__abc_44228_n18403), .B(u2__abc_44228_n2983_bF_buf87), .Y(u2__abc_44228_n18404) );
  OR2X2 OR2X2_4393 ( .A(u2__abc_44228_n18408), .B(u2__abc_44228_n18399), .Y(u2__abc_44228_n18409) );
  OR2X2 OR2X2_4394 ( .A(u2__abc_44228_n18401), .B(sqrto_52_), .Y(u2__abc_44228_n18412) );
  OR2X2 OR2X2_4395 ( .A(u2__abc_44228_n18415), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n18416) );
  OR2X2 OR2X2_4396 ( .A(u2__abc_44228_n18420), .B(u2__abc_44228_n18411), .Y(u2__abc_44228_n18421) );
  OR2X2 OR2X2_4397 ( .A(u2__abc_44228_n18413), .B(sqrto_53_), .Y(u2__abc_44228_n18424) );
  OR2X2 OR2X2_4398 ( .A(u2__abc_44228_n18427), .B(u2__abc_44228_n2983_bF_buf83), .Y(u2__abc_44228_n18428) );
  OR2X2 OR2X2_4399 ( .A(u2__abc_44228_n18432), .B(u2__abc_44228_n18423), .Y(u2__abc_44228_n18433) );
  OR2X2 OR2X2_44 ( .A(_abc_64468_n753_bF_buf0), .B(\a[21] ), .Y(_abc_64468_n894) );
  OR2X2 OR2X2_440 ( .A(a_112_bF_buf0), .B(\a[107] ), .Y(_abc_64468_n1491) );
  OR2X2 OR2X2_4400 ( .A(u2__abc_44228_n18425), .B(sqrto_54_), .Y(u2__abc_44228_n18436) );
  OR2X2 OR2X2_4401 ( .A(u2__abc_44228_n18439), .B(u2__abc_44228_n2983_bF_buf81), .Y(u2__abc_44228_n18440) );
  OR2X2 OR2X2_4402 ( .A(u2__abc_44228_n18444), .B(u2__abc_44228_n18435), .Y(u2__abc_44228_n18445) );
  OR2X2 OR2X2_4403 ( .A(u2__abc_44228_n18437), .B(sqrto_55_), .Y(u2__abc_44228_n18448) );
  OR2X2 OR2X2_4404 ( .A(u2__abc_44228_n18451), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n18452) );
  OR2X2 OR2X2_4405 ( .A(u2__abc_44228_n18456), .B(u2__abc_44228_n18447), .Y(u2__abc_44228_n18457) );
  OR2X2 OR2X2_4406 ( .A(u2__abc_44228_n18449), .B(sqrto_56_), .Y(u2__abc_44228_n18460) );
  OR2X2 OR2X2_4407 ( .A(u2__abc_44228_n18463), .B(u2__abc_44228_n2983_bF_buf77), .Y(u2__abc_44228_n18464) );
  OR2X2 OR2X2_4408 ( .A(u2__abc_44228_n18468), .B(u2__abc_44228_n18459), .Y(u2__abc_44228_n18469) );
  OR2X2 OR2X2_4409 ( .A(u2__abc_44228_n18461), .B(sqrto_57_), .Y(u2__abc_44228_n18472) );
  OR2X2 OR2X2_441 ( .A(_abc_64468_n1170_bF_buf2), .B(\a[108] ), .Y(_abc_64468_n1492) );
  OR2X2 OR2X2_4410 ( .A(u2__abc_44228_n18475), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n18476) );
  OR2X2 OR2X2_4411 ( .A(u2__abc_44228_n18480), .B(u2__abc_44228_n18471), .Y(u2__abc_44228_n18481) );
  OR2X2 OR2X2_4412 ( .A(u2__abc_44228_n18473), .B(sqrto_58_), .Y(u2__abc_44228_n18484) );
  OR2X2 OR2X2_4413 ( .A(u2__abc_44228_n18487), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n18488) );
  OR2X2 OR2X2_4414 ( .A(u2__abc_44228_n18492), .B(u2__abc_44228_n18483), .Y(u2__abc_44228_n18493) );
  OR2X2 OR2X2_4415 ( .A(u2__abc_44228_n18485), .B(sqrto_59_), .Y(u2__abc_44228_n18496) );
  OR2X2 OR2X2_4416 ( .A(u2__abc_44228_n18499), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n18500) );
  OR2X2 OR2X2_4417 ( .A(u2__abc_44228_n18504), .B(u2__abc_44228_n18495), .Y(u2__abc_44228_n18505) );
  OR2X2 OR2X2_4418 ( .A(u2__abc_44228_n18497), .B(sqrto_60_), .Y(u2__abc_44228_n18508) );
  OR2X2 OR2X2_4419 ( .A(u2__abc_44228_n18511), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n18512) );
  OR2X2 OR2X2_442 ( .A(a_112_bF_buf9), .B(\a[108] ), .Y(_abc_64468_n1494) );
  OR2X2 OR2X2_4420 ( .A(u2__abc_44228_n18516), .B(u2__abc_44228_n18507), .Y(u2__abc_44228_n18517) );
  OR2X2 OR2X2_4421 ( .A(u2__abc_44228_n18509), .B(sqrto_61_), .Y(u2__abc_44228_n18520) );
  OR2X2 OR2X2_4422 ( .A(u2__abc_44228_n18523), .B(u2__abc_44228_n2983_bF_buf67), .Y(u2__abc_44228_n18524) );
  OR2X2 OR2X2_4423 ( .A(u2__abc_44228_n18528), .B(u2__abc_44228_n18519), .Y(u2__abc_44228_n18529) );
  OR2X2 OR2X2_4424 ( .A(u2__abc_44228_n18521), .B(sqrto_62_), .Y(u2__abc_44228_n18532) );
  OR2X2 OR2X2_4425 ( .A(u2__abc_44228_n18535), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n18536) );
  OR2X2 OR2X2_4426 ( .A(u2__abc_44228_n18540), .B(u2__abc_44228_n18531), .Y(u2__abc_44228_n18541) );
  OR2X2 OR2X2_4427 ( .A(u2__abc_44228_n18533), .B(sqrto_63_), .Y(u2__abc_44228_n18544) );
  OR2X2 OR2X2_4428 ( .A(u2__abc_44228_n18547), .B(u2__abc_44228_n2983_bF_buf63), .Y(u2__abc_44228_n18548) );
  OR2X2 OR2X2_4429 ( .A(u2__abc_44228_n18552), .B(u2__abc_44228_n18543), .Y(u2__abc_44228_n18553) );
  OR2X2 OR2X2_443 ( .A(_abc_64468_n1170_bF_buf1), .B(\a[109] ), .Y(_abc_64468_n1495) );
  OR2X2 OR2X2_4430 ( .A(u2__abc_44228_n18545), .B(sqrto_64_), .Y(u2__abc_44228_n18556) );
  OR2X2 OR2X2_4431 ( .A(u2__abc_44228_n18559), .B(u2__abc_44228_n2983_bF_buf61), .Y(u2__abc_44228_n18560) );
  OR2X2 OR2X2_4432 ( .A(u2__abc_44228_n18564), .B(u2__abc_44228_n18555), .Y(u2__abc_44228_n18565) );
  OR2X2 OR2X2_4433 ( .A(u2__abc_44228_n18557), .B(sqrto_65_), .Y(u2__abc_44228_n18568) );
  OR2X2 OR2X2_4434 ( .A(u2__abc_44228_n18571), .B(u2__abc_44228_n2983_bF_buf59), .Y(u2__abc_44228_n18572) );
  OR2X2 OR2X2_4435 ( .A(u2__abc_44228_n18576), .B(u2__abc_44228_n18567), .Y(u2__abc_44228_n18577) );
  OR2X2 OR2X2_4436 ( .A(u2__abc_44228_n18569), .B(sqrto_66_), .Y(u2__abc_44228_n18580) );
  OR2X2 OR2X2_4437 ( .A(u2__abc_44228_n18583), .B(u2__abc_44228_n2983_bF_buf57), .Y(u2__abc_44228_n18584) );
  OR2X2 OR2X2_4438 ( .A(u2__abc_44228_n18588), .B(u2__abc_44228_n18579), .Y(u2__abc_44228_n18589) );
  OR2X2 OR2X2_4439 ( .A(u2__abc_44228_n18581), .B(sqrto_67_), .Y(u2__abc_44228_n18592) );
  OR2X2 OR2X2_444 ( .A(a_112_bF_buf8), .B(\a[109] ), .Y(_abc_64468_n1497) );
  OR2X2 OR2X2_4440 ( .A(u2__abc_44228_n18595), .B(u2__abc_44228_n2983_bF_buf55), .Y(u2__abc_44228_n18596) );
  OR2X2 OR2X2_4441 ( .A(u2__abc_44228_n18600), .B(u2__abc_44228_n18591), .Y(u2__abc_44228_n18601) );
  OR2X2 OR2X2_4442 ( .A(u2__abc_44228_n18593), .B(sqrto_68_), .Y(u2__abc_44228_n18604) );
  OR2X2 OR2X2_4443 ( .A(u2__abc_44228_n18607), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n18608) );
  OR2X2 OR2X2_4444 ( .A(u2__abc_44228_n18612), .B(u2__abc_44228_n18603), .Y(u2__abc_44228_n18613) );
  OR2X2 OR2X2_4445 ( .A(u2__abc_44228_n18605), .B(sqrto_69_), .Y(u2__abc_44228_n18616) );
  OR2X2 OR2X2_4446 ( .A(u2__abc_44228_n18619), .B(u2__abc_44228_n2983_bF_buf51), .Y(u2__abc_44228_n18620) );
  OR2X2 OR2X2_4447 ( .A(u2__abc_44228_n18624), .B(u2__abc_44228_n18615), .Y(u2__abc_44228_n18625) );
  OR2X2 OR2X2_4448 ( .A(u2__abc_44228_n18617), .B(sqrto_70_), .Y(u2__abc_44228_n18628) );
  OR2X2 OR2X2_4449 ( .A(u2__abc_44228_n18631), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n18632) );
  OR2X2 OR2X2_445 ( .A(_abc_64468_n1170_bF_buf0), .B(\a[110] ), .Y(_abc_64468_n1498) );
  OR2X2 OR2X2_4450 ( .A(u2__abc_44228_n18636), .B(u2__abc_44228_n18627), .Y(u2__abc_44228_n18637) );
  OR2X2 OR2X2_4451 ( .A(u2__abc_44228_n18629), .B(sqrto_71_), .Y(u2__abc_44228_n18640) );
  OR2X2 OR2X2_4452 ( .A(u2__abc_44228_n18643), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n18644) );
  OR2X2 OR2X2_4453 ( .A(u2__abc_44228_n18648), .B(u2__abc_44228_n18639), .Y(u2__abc_44228_n18649) );
  OR2X2 OR2X2_4454 ( .A(u2__abc_44228_n18641), .B(sqrto_72_), .Y(u2__abc_44228_n18652) );
  OR2X2 OR2X2_4455 ( .A(u2__abc_44228_n18655), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n18656) );
  OR2X2 OR2X2_4456 ( .A(u2__abc_44228_n18660), .B(u2__abc_44228_n18651), .Y(u2__abc_44228_n18661) );
  OR2X2 OR2X2_4457 ( .A(u2__abc_44228_n18653), .B(sqrto_73_), .Y(u2__abc_44228_n18664) );
  OR2X2 OR2X2_4458 ( .A(u2__abc_44228_n18667), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n18668) );
  OR2X2 OR2X2_4459 ( .A(u2__abc_44228_n18672), .B(u2__abc_44228_n18663), .Y(u2__abc_44228_n18673) );
  OR2X2 OR2X2_446 ( .A(a_112_bF_buf7), .B(\a[110] ), .Y(_abc_64468_n1500) );
  OR2X2 OR2X2_4460 ( .A(u2__abc_44228_n18665), .B(sqrto_74_), .Y(u2__abc_44228_n18676) );
  OR2X2 OR2X2_4461 ( .A(u2__abc_44228_n18679), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n18680) );
  OR2X2 OR2X2_4462 ( .A(u2__abc_44228_n18684), .B(u2__abc_44228_n18675), .Y(u2__abc_44228_n18685) );
  OR2X2 OR2X2_4463 ( .A(u2__abc_44228_n18677), .B(sqrto_75_), .Y(u2__abc_44228_n18688) );
  OR2X2 OR2X2_4464 ( .A(u2__abc_44228_n18691), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n18692) );
  OR2X2 OR2X2_4465 ( .A(u2__abc_44228_n18696), .B(u2__abc_44228_n18687), .Y(u2__abc_44228_n18697) );
  OR2X2 OR2X2_4466 ( .A(u2__abc_44228_n18689), .B(sqrto_76_), .Y(u2__abc_44228_n18700) );
  OR2X2 OR2X2_4467 ( .A(u2__abc_44228_n18703), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n18704) );
  OR2X2 OR2X2_4468 ( .A(u2__abc_44228_n18708), .B(u2__abc_44228_n18699), .Y(u2__abc_44228_n18709) );
  OR2X2 OR2X2_4469 ( .A(u2__abc_44228_n18701), .B(sqrto_77_), .Y(u2__abc_44228_n18712) );
  OR2X2 OR2X2_447 ( .A(_abc_64468_n1170_bF_buf9), .B(\a[111] ), .Y(_abc_64468_n1501) );
  OR2X2 OR2X2_4470 ( .A(u2__abc_44228_n18715), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n18716) );
  OR2X2 OR2X2_4471 ( .A(u2__abc_44228_n18720), .B(u2__abc_44228_n18711), .Y(u2__abc_44228_n18721) );
  OR2X2 OR2X2_4472 ( .A(u2__abc_44228_n18713), .B(sqrto_78_), .Y(u2__abc_44228_n18724) );
  OR2X2 OR2X2_4473 ( .A(u2__abc_44228_n18727), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n18728) );
  OR2X2 OR2X2_4474 ( .A(u2__abc_44228_n18732), .B(u2__abc_44228_n18723), .Y(u2__abc_44228_n18733) );
  OR2X2 OR2X2_4475 ( .A(u2__abc_44228_n18725), .B(sqrto_79_), .Y(u2__abc_44228_n18736) );
  OR2X2 OR2X2_4476 ( .A(u2__abc_44228_n18739), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n18740) );
  OR2X2 OR2X2_4477 ( .A(u2__abc_44228_n18744), .B(u2__abc_44228_n18735), .Y(u2__abc_44228_n18745) );
  OR2X2 OR2X2_4478 ( .A(u2__abc_44228_n18737), .B(sqrto_80_), .Y(u2__abc_44228_n18748) );
  OR2X2 OR2X2_4479 ( .A(u2__abc_44228_n18751), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n18752) );
  OR2X2 OR2X2_448 ( .A(a_112_bF_buf6), .B(\a[111] ), .Y(_abc_64468_n1503) );
  OR2X2 OR2X2_4480 ( .A(u2__abc_44228_n18756), .B(u2__abc_44228_n18747), .Y(u2__abc_44228_n18757) );
  OR2X2 OR2X2_4481 ( .A(u2__abc_44228_n18749), .B(sqrto_81_), .Y(u2__abc_44228_n18760) );
  OR2X2 OR2X2_4482 ( .A(u2__abc_44228_n18763), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n18764) );
  OR2X2 OR2X2_4483 ( .A(u2__abc_44228_n18768), .B(u2__abc_44228_n18759), .Y(u2__abc_44228_n18769) );
  OR2X2 OR2X2_4484 ( .A(u2__abc_44228_n18761), .B(sqrto_82_), .Y(u2__abc_44228_n18772) );
  OR2X2 OR2X2_4485 ( .A(u2__abc_44228_n18775), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n18776) );
  OR2X2 OR2X2_4486 ( .A(u2__abc_44228_n18780), .B(u2__abc_44228_n18771), .Y(u2__abc_44228_n18781) );
  OR2X2 OR2X2_4487 ( .A(u2__abc_44228_n18773), .B(sqrto_83_), .Y(u2__abc_44228_n18784) );
  OR2X2 OR2X2_4488 ( .A(u2__abc_44228_n18787), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n18788) );
  OR2X2 OR2X2_4489 ( .A(u2__abc_44228_n18792), .B(u2__abc_44228_n18783), .Y(u2__abc_44228_n18793) );
  OR2X2 OR2X2_449 ( .A(_abc_64468_n1170_bF_buf8), .B(fracta_112_), .Y(_abc_64468_n1504) );
  OR2X2 OR2X2_4490 ( .A(u2__abc_44228_n18785), .B(sqrto_84_), .Y(u2__abc_44228_n18796) );
  OR2X2 OR2X2_4491 ( .A(u2__abc_44228_n18799), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n18800) );
  OR2X2 OR2X2_4492 ( .A(u2__abc_44228_n18804), .B(u2__abc_44228_n18795), .Y(u2__abc_44228_n18805) );
  OR2X2 OR2X2_4493 ( .A(u2__abc_44228_n18797), .B(sqrto_85_), .Y(u2__abc_44228_n18808) );
  OR2X2 OR2X2_4494 ( .A(u2__abc_44228_n18811), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n18812) );
  OR2X2 OR2X2_4495 ( .A(u2__abc_44228_n18816), .B(u2__abc_44228_n18807), .Y(u2__abc_44228_n18817) );
  OR2X2 OR2X2_4496 ( .A(u2__abc_44228_n18809), .B(sqrto_86_), .Y(u2__abc_44228_n18820) );
  OR2X2 OR2X2_4497 ( .A(u2__abc_44228_n18823), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n18824) );
  OR2X2 OR2X2_4498 ( .A(u2__abc_44228_n18828), .B(u2__abc_44228_n18819), .Y(u2__abc_44228_n18829) );
  OR2X2 OR2X2_4499 ( .A(u2__abc_44228_n18821), .B(sqrto_87_), .Y(u2__abc_44228_n18832) );
  OR2X2 OR2X2_45 ( .A(aNan_bF_buf9), .B(sqrto_98_), .Y(_abc_64468_n896) );
  OR2X2 OR2X2_450 ( .A(_abc_64468_n753_bF_buf6), .B(a_112_bF_buf5), .Y(_abc_64468_n1507) );
  OR2X2 OR2X2_4500 ( .A(u2__abc_44228_n18835), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n18836) );
  OR2X2 OR2X2_4501 ( .A(u2__abc_44228_n18840), .B(u2__abc_44228_n18831), .Y(u2__abc_44228_n18841) );
  OR2X2 OR2X2_4502 ( .A(u2__abc_44228_n18833), .B(sqrto_88_), .Y(u2__abc_44228_n18844) );
  OR2X2 OR2X2_4503 ( .A(u2__abc_44228_n18847), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n18848) );
  OR2X2 OR2X2_4504 ( .A(u2__abc_44228_n18852), .B(u2__abc_44228_n18843), .Y(u2__abc_44228_n18853) );
  OR2X2 OR2X2_4505 ( .A(u2__abc_44228_n18845), .B(sqrto_89_), .Y(u2__abc_44228_n18856) );
  OR2X2 OR2X2_4506 ( .A(u2__abc_44228_n18859), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n18860) );
  OR2X2 OR2X2_4507 ( .A(u2__abc_44228_n18864), .B(u2__abc_44228_n18855), .Y(u2__abc_44228_n18865) );
  OR2X2 OR2X2_4508 ( .A(u2__abc_44228_n18857), .B(sqrto_90_), .Y(u2__abc_44228_n18868) );
  OR2X2 OR2X2_4509 ( .A(u2__abc_44228_n18871), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n18872) );
  OR2X2 OR2X2_451 ( .A(_abc_64468_n1510), .B(aNan_bF_buf6), .Y(_abc_64468_n1511) );
  OR2X2 OR2X2_4510 ( .A(u2__abc_44228_n18876), .B(u2__abc_44228_n18867), .Y(u2__abc_44228_n18877) );
  OR2X2 OR2X2_4511 ( .A(u2__abc_44228_n18869), .B(sqrto_91_), .Y(u2__abc_44228_n18880) );
  OR2X2 OR2X2_4512 ( .A(u2__abc_44228_n18883), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n18884) );
  OR2X2 OR2X2_4513 ( .A(u2__abc_44228_n18888), .B(u2__abc_44228_n18879), .Y(u2__abc_44228_n18889) );
  OR2X2 OR2X2_4514 ( .A(u2__abc_44228_n18881), .B(sqrto_92_), .Y(u2__abc_44228_n18892) );
  OR2X2 OR2X2_4515 ( .A(u2__abc_44228_n18895), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n18896) );
  OR2X2 OR2X2_4516 ( .A(u2__abc_44228_n18900), .B(u2__abc_44228_n18891), .Y(u2__abc_44228_n18901) );
  OR2X2 OR2X2_4517 ( .A(u2__abc_44228_n18893), .B(sqrto_93_), .Y(u2__abc_44228_n18904) );
  OR2X2 OR2X2_4518 ( .A(u2__abc_44228_n18907), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n18908) );
  OR2X2 OR2X2_4519 ( .A(u2__abc_44228_n18912), .B(u2__abc_44228_n18903), .Y(u2__abc_44228_n18913) );
  OR2X2 OR2X2_452 ( .A(_abc_64468_n1511), .B(_abc_64468_n1509), .Y(_abc_64468_n1512) );
  OR2X2 OR2X2_4520 ( .A(u2__abc_44228_n18905), .B(sqrto_94_), .Y(u2__abc_44228_n18916) );
  OR2X2 OR2X2_4521 ( .A(u2__abc_44228_n18919), .B(u2__abc_44228_n2983_bF_buf1), .Y(u2__abc_44228_n18920) );
  OR2X2 OR2X2_4522 ( .A(u2__abc_44228_n18924), .B(u2__abc_44228_n18915), .Y(u2__abc_44228_n18925) );
  OR2X2 OR2X2_4523 ( .A(u2__abc_44228_n18917), .B(sqrto_95_), .Y(u2__abc_44228_n18928) );
  OR2X2 OR2X2_4524 ( .A(u2__abc_44228_n18931), .B(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n18932) );
  OR2X2 OR2X2_4525 ( .A(u2__abc_44228_n18936), .B(u2__abc_44228_n18927), .Y(u2__abc_44228_n18937) );
  OR2X2 OR2X2_4526 ( .A(u2__abc_44228_n18929), .B(sqrto_96_), .Y(u2__abc_44228_n18940) );
  OR2X2 OR2X2_4527 ( .A(u2__abc_44228_n18943), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n18944) );
  OR2X2 OR2X2_4528 ( .A(u2__abc_44228_n18948), .B(u2__abc_44228_n18939), .Y(u2__abc_44228_n18949) );
  OR2X2 OR2X2_4529 ( .A(u2__abc_44228_n18941), .B(sqrto_97_), .Y(u2__abc_44228_n18952) );
  OR2X2 OR2X2_453 ( .A(_abc_64468_n1509), .B(\a[114] ), .Y(_abc_64468_n1514) );
  OR2X2 OR2X2_4530 ( .A(u2__abc_44228_n18955), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n18956) );
  OR2X2 OR2X2_4531 ( .A(u2__abc_44228_n18960), .B(u2__abc_44228_n18951), .Y(u2__abc_44228_n18961) );
  OR2X2 OR2X2_4532 ( .A(u2__abc_44228_n18953), .B(sqrto_98_), .Y(u2__abc_44228_n18964) );
  OR2X2 OR2X2_4533 ( .A(u2__abc_44228_n18967), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n18968) );
  OR2X2 OR2X2_4534 ( .A(u2__abc_44228_n18972), .B(u2__abc_44228_n18963), .Y(u2__abc_44228_n18973) );
  OR2X2 OR2X2_4535 ( .A(u2__abc_44228_n18965), .B(sqrto_99_), .Y(u2__abc_44228_n18976) );
  OR2X2 OR2X2_4536 ( .A(u2__abc_44228_n18979), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n18980) );
  OR2X2 OR2X2_4537 ( .A(u2__abc_44228_n18984), .B(u2__abc_44228_n18975), .Y(u2__abc_44228_n18985) );
  OR2X2 OR2X2_4538 ( .A(u2__abc_44228_n18977), .B(sqrto_100_), .Y(u2__abc_44228_n18988) );
  OR2X2 OR2X2_4539 ( .A(u2__abc_44228_n18991), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n18992) );
  OR2X2 OR2X2_454 ( .A(_abc_64468_n1518), .B(a_112_bF_buf3), .Y(_abc_64468_n1519) );
  OR2X2 OR2X2_4540 ( .A(u2__abc_44228_n18996), .B(u2__abc_44228_n18987), .Y(u2__abc_44228_n18997) );
  OR2X2 OR2X2_4541 ( .A(u2__abc_44228_n18989), .B(sqrto_101_), .Y(u2__abc_44228_n19000) );
  OR2X2 OR2X2_4542 ( .A(u2__abc_44228_n19003), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n19004) );
  OR2X2 OR2X2_4543 ( .A(u2__abc_44228_n19008), .B(u2__abc_44228_n18999), .Y(u2__abc_44228_n19009) );
  OR2X2 OR2X2_4544 ( .A(u2__abc_44228_n19001), .B(sqrto_102_), .Y(u2__abc_44228_n19012) );
  OR2X2 OR2X2_4545 ( .A(u2__abc_44228_n19015), .B(u2__abc_44228_n2983_bF_buf127), .Y(u2__abc_44228_n19016) );
  OR2X2 OR2X2_4546 ( .A(u2__abc_44228_n19020), .B(u2__abc_44228_n19011), .Y(u2__abc_44228_n19021) );
  OR2X2 OR2X2_4547 ( .A(u2__abc_44228_n19013), .B(sqrto_103_), .Y(u2__abc_44228_n19024) );
  OR2X2 OR2X2_4548 ( .A(u2__abc_44228_n19027), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n19028) );
  OR2X2 OR2X2_4549 ( .A(u2__abc_44228_n19032), .B(u2__abc_44228_n19023), .Y(u2__abc_44228_n19033) );
  OR2X2 OR2X2_455 ( .A(_abc_64468_n1520), .B(\a[113] ), .Y(_abc_64468_n1521) );
  OR2X2 OR2X2_4550 ( .A(u2__abc_44228_n19025), .B(sqrto_104_), .Y(u2__abc_44228_n19036) );
  OR2X2 OR2X2_4551 ( .A(u2__abc_44228_n19039), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n19040) );
  OR2X2 OR2X2_4552 ( .A(u2__abc_44228_n19044), .B(u2__abc_44228_n19035), .Y(u2__abc_44228_n19045) );
  OR2X2 OR2X2_4553 ( .A(u2__abc_44228_n19037), .B(sqrto_105_), .Y(u2__abc_44228_n19048) );
  OR2X2 OR2X2_4554 ( .A(u2__abc_44228_n19051), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n19052) );
  OR2X2 OR2X2_4555 ( .A(u2__abc_44228_n19056), .B(u2__abc_44228_n19047), .Y(u2__abc_44228_n19057) );
  OR2X2 OR2X2_4556 ( .A(u2__abc_44228_n19049), .B(sqrto_106_), .Y(u2__abc_44228_n19060) );
  OR2X2 OR2X2_4557 ( .A(u2__abc_44228_n19063), .B(u2__abc_44228_n2983_bF_buf119), .Y(u2__abc_44228_n19064) );
  OR2X2 OR2X2_4558 ( .A(u2__abc_44228_n19068), .B(u2__abc_44228_n19059), .Y(u2__abc_44228_n19069) );
  OR2X2 OR2X2_4559 ( .A(u2__abc_44228_n19061), .B(sqrto_107_), .Y(u2__abc_44228_n19072) );
  OR2X2 OR2X2_456 ( .A(_abc_64468_n1510), .B(_abc_64468_n1518), .Y(_abc_64468_n1523) );
  OR2X2 OR2X2_4560 ( .A(u2__abc_44228_n19075), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n19076) );
  OR2X2 OR2X2_4561 ( .A(u2__abc_44228_n19080), .B(u2__abc_44228_n19071), .Y(u2__abc_44228_n19081) );
  OR2X2 OR2X2_4562 ( .A(u2__abc_44228_n19073), .B(sqrto_108_), .Y(u2__abc_44228_n19084) );
  OR2X2 OR2X2_4563 ( .A(u2__abc_44228_n19087), .B(u2__abc_44228_n2983_bF_buf115), .Y(u2__abc_44228_n19088) );
  OR2X2 OR2X2_4564 ( .A(u2__abc_44228_n19092), .B(u2__abc_44228_n19083), .Y(u2__abc_44228_n19093) );
  OR2X2 OR2X2_4565 ( .A(u2__abc_44228_n19085), .B(sqrto_109_), .Y(u2__abc_44228_n19096) );
  OR2X2 OR2X2_4566 ( .A(u2__abc_44228_n19099), .B(u2__abc_44228_n2983_bF_buf113), .Y(u2__abc_44228_n19100) );
  OR2X2 OR2X2_4567 ( .A(u2__abc_44228_n19104), .B(u2__abc_44228_n19095), .Y(u2__abc_44228_n19105) );
  OR2X2 OR2X2_4568 ( .A(u2__abc_44228_n19097), .B(sqrto_110_), .Y(u2__abc_44228_n19108) );
  OR2X2 OR2X2_4569 ( .A(u2__abc_44228_n19111), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n19112) );
  OR2X2 OR2X2_457 ( .A(_abc_64468_n1526), .B(_abc_64468_n1525), .Y(_abc_64468_n1527) );
  OR2X2 OR2X2_4570 ( .A(u2__abc_44228_n19116), .B(u2__abc_44228_n19107), .Y(u2__abc_44228_n19117) );
  OR2X2 OR2X2_4571 ( .A(u2__abc_44228_n19109), .B(sqrto_111_), .Y(u2__abc_44228_n19120) );
  OR2X2 OR2X2_4572 ( .A(u2__abc_44228_n19123), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n19124) );
  OR2X2 OR2X2_4573 ( .A(u2__abc_44228_n19128), .B(u2__abc_44228_n19119), .Y(u2__abc_44228_n19129) );
  OR2X2 OR2X2_4574 ( .A(u2__abc_44228_n19121), .B(sqrto_112_), .Y(u2__abc_44228_n19132) );
  OR2X2 OR2X2_4575 ( .A(u2__abc_44228_n19135), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n19136) );
  OR2X2 OR2X2_4576 ( .A(u2__abc_44228_n19140), .B(u2__abc_44228_n19131), .Y(u2__abc_44228_n19141) );
  OR2X2 OR2X2_4577 ( .A(u2__abc_44228_n19133), .B(sqrto_113_), .Y(u2__abc_44228_n19144) );
  OR2X2 OR2X2_4578 ( .A(u2__abc_44228_n19147), .B(u2__abc_44228_n2983_bF_buf105), .Y(u2__abc_44228_n19148) );
  OR2X2 OR2X2_4579 ( .A(u2__abc_44228_n19152), .B(u2__abc_44228_n19143), .Y(u2__abc_44228_n19153) );
  OR2X2 OR2X2_458 ( .A(_abc_64468_n1531), .B(_abc_64468_n1533), .Y(_abc_64468_n1534) );
  OR2X2 OR2X2_4580 ( .A(u2__abc_44228_n19145), .B(sqrto_114_), .Y(u2__abc_44228_n19156) );
  OR2X2 OR2X2_4581 ( .A(u2__abc_44228_n19159), .B(u2__abc_44228_n2983_bF_buf103), .Y(u2__abc_44228_n19160) );
  OR2X2 OR2X2_4582 ( .A(u2__abc_44228_n19164), .B(u2__abc_44228_n19155), .Y(u2__abc_44228_n19165) );
  OR2X2 OR2X2_4583 ( .A(u2__abc_44228_n19157), .B(sqrto_115_), .Y(u2__abc_44228_n19168) );
  OR2X2 OR2X2_4584 ( .A(u2__abc_44228_n19171), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n19172) );
  OR2X2 OR2X2_4585 ( .A(u2__abc_44228_n19176), .B(u2__abc_44228_n19167), .Y(u2__abc_44228_n19177) );
  OR2X2 OR2X2_4586 ( .A(u2__abc_44228_n19169), .B(sqrto_116_), .Y(u2__abc_44228_n19180) );
  OR2X2 OR2X2_4587 ( .A(u2__abc_44228_n19183), .B(u2__abc_44228_n2983_bF_buf99), .Y(u2__abc_44228_n19184) );
  OR2X2 OR2X2_4588 ( .A(u2__abc_44228_n19188), .B(u2__abc_44228_n19179), .Y(u2__abc_44228_n19189) );
  OR2X2 OR2X2_4589 ( .A(u2__abc_44228_n19181), .B(sqrto_117_), .Y(u2__abc_44228_n19192) );
  OR2X2 OR2X2_459 ( .A(_abc_64468_n1535), .B(_abc_64468_n1536), .Y(_auto_iopadmap_cc_313_execute_65414_228_) );
  OR2X2 OR2X2_4590 ( .A(u2__abc_44228_n19195), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n19196) );
  OR2X2 OR2X2_4591 ( .A(u2__abc_44228_n19200), .B(u2__abc_44228_n19191), .Y(u2__abc_44228_n19201) );
  OR2X2 OR2X2_4592 ( .A(u2__abc_44228_n19193), .B(sqrto_118_), .Y(u2__abc_44228_n19204) );
  OR2X2 OR2X2_4593 ( .A(u2__abc_44228_n19207), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n19208) );
  OR2X2 OR2X2_4594 ( .A(u2__abc_44228_n19212), .B(u2__abc_44228_n19203), .Y(u2__abc_44228_n19213) );
  OR2X2 OR2X2_4595 ( .A(u2__abc_44228_n19205), .B(sqrto_119_), .Y(u2__abc_44228_n19216) );
  OR2X2 OR2X2_4596 ( .A(u2__abc_44228_n19219), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n19220) );
  OR2X2 OR2X2_4597 ( .A(u2__abc_44228_n19224), .B(u2__abc_44228_n19215), .Y(u2__abc_44228_n19225) );
  OR2X2 OR2X2_4598 ( .A(u2__abc_44228_n19217), .B(sqrto_120_), .Y(u2__abc_44228_n19228) );
  OR2X2 OR2X2_4599 ( .A(u2__abc_44228_n19231), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n19232) );
  OR2X2 OR2X2_46 ( .A(_abc_64468_n753_bF_buf13), .B(\a[22] ), .Y(_abc_64468_n897) );
  OR2X2 OR2X2_460 ( .A(_abc_64468_n1539), .B(_abc_64468_n1538), .Y(_abc_64468_n1540) );
  OR2X2 OR2X2_4600 ( .A(u2__abc_44228_n19236), .B(u2__abc_44228_n19227), .Y(u2__abc_44228_n19237) );
  OR2X2 OR2X2_4601 ( .A(u2__abc_44228_n19229), .B(sqrto_121_), .Y(u2__abc_44228_n19240) );
  OR2X2 OR2X2_4602 ( .A(u2__abc_44228_n19243), .B(u2__abc_44228_n2983_bF_buf89), .Y(u2__abc_44228_n19244) );
  OR2X2 OR2X2_4603 ( .A(u2__abc_44228_n19248), .B(u2__abc_44228_n19239), .Y(u2__abc_44228_n19249) );
  OR2X2 OR2X2_4604 ( .A(u2__abc_44228_n19241), .B(sqrto_122_), .Y(u2__abc_44228_n19252) );
  OR2X2 OR2X2_4605 ( .A(u2__abc_44228_n19255), .B(u2__abc_44228_n2983_bF_buf87), .Y(u2__abc_44228_n19256) );
  OR2X2 OR2X2_4606 ( .A(u2__abc_44228_n19260), .B(u2__abc_44228_n19251), .Y(u2__abc_44228_n19261) );
  OR2X2 OR2X2_4607 ( .A(u2__abc_44228_n19253), .B(sqrto_123_), .Y(u2__abc_44228_n19264) );
  OR2X2 OR2X2_4608 ( .A(u2__abc_44228_n19267), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n19268) );
  OR2X2 OR2X2_4609 ( .A(u2__abc_44228_n19272), .B(u2__abc_44228_n19263), .Y(u2__abc_44228_n19273) );
  OR2X2 OR2X2_461 ( .A(_abc_64468_n1547), .B(_abc_64468_n1544), .Y(_abc_64468_n1548) );
  OR2X2 OR2X2_4610 ( .A(u2__abc_44228_n19265), .B(sqrto_124_), .Y(u2__abc_44228_n19276) );
  OR2X2 OR2X2_4611 ( .A(u2__abc_44228_n19279), .B(u2__abc_44228_n2983_bF_buf83), .Y(u2__abc_44228_n19280) );
  OR2X2 OR2X2_4612 ( .A(u2__abc_44228_n19284), .B(u2__abc_44228_n19275), .Y(u2__abc_44228_n19285) );
  OR2X2 OR2X2_4613 ( .A(u2__abc_44228_n19277), .B(sqrto_125_), .Y(u2__abc_44228_n19288) );
  OR2X2 OR2X2_4614 ( .A(u2__abc_44228_n19291), .B(u2__abc_44228_n2983_bF_buf81), .Y(u2__abc_44228_n19292) );
  OR2X2 OR2X2_4615 ( .A(u2__abc_44228_n19296), .B(u2__abc_44228_n19287), .Y(u2__abc_44228_n19297) );
  OR2X2 OR2X2_4616 ( .A(u2__abc_44228_n19289), .B(sqrto_126_), .Y(u2__abc_44228_n19300) );
  OR2X2 OR2X2_4617 ( .A(u2__abc_44228_n19303), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n19304) );
  OR2X2 OR2X2_4618 ( .A(u2__abc_44228_n19308), .B(u2__abc_44228_n19299), .Y(u2__abc_44228_n19309) );
  OR2X2 OR2X2_4619 ( .A(u2__abc_44228_n19301), .B(sqrto_127_), .Y(u2__abc_44228_n19312) );
  OR2X2 OR2X2_462 ( .A(_abc_64468_n1548), .B(aNan_bF_buf4), .Y(_abc_64468_n1549) );
  OR2X2 OR2X2_4620 ( .A(u2__abc_44228_n19315), .B(u2__abc_44228_n2983_bF_buf77), .Y(u2__abc_44228_n19316) );
  OR2X2 OR2X2_4621 ( .A(u2__abc_44228_n19320), .B(u2__abc_44228_n19311), .Y(u2__abc_44228_n19321) );
  OR2X2 OR2X2_4622 ( .A(u2__abc_44228_n19313), .B(sqrto_128_), .Y(u2__abc_44228_n19324) );
  OR2X2 OR2X2_4623 ( .A(u2__abc_44228_n19327), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n19328) );
  OR2X2 OR2X2_4624 ( .A(u2__abc_44228_n19332), .B(u2__abc_44228_n19323), .Y(u2__abc_44228_n19333) );
  OR2X2 OR2X2_4625 ( .A(u2__abc_44228_n19325), .B(sqrto_129_), .Y(u2__abc_44228_n19336) );
  OR2X2 OR2X2_4626 ( .A(u2__abc_44228_n19339), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n19340) );
  OR2X2 OR2X2_4627 ( .A(u2__abc_44228_n19344), .B(u2__abc_44228_n19335), .Y(u2__abc_44228_n19345) );
  OR2X2 OR2X2_4628 ( .A(u2__abc_44228_n19337), .B(sqrto_130_), .Y(u2__abc_44228_n19348) );
  OR2X2 OR2X2_4629 ( .A(u2__abc_44228_n19351), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n19352) );
  OR2X2 OR2X2_463 ( .A(_abc_64468_n753_bF_buf2), .B(\a[115] ), .Y(_abc_64468_n1550) );
  OR2X2 OR2X2_4630 ( .A(u2__abc_44228_n19356), .B(u2__abc_44228_n19347), .Y(u2__abc_44228_n19357) );
  OR2X2 OR2X2_4631 ( .A(u2__abc_44228_n19349), .B(sqrto_131_), .Y(u2__abc_44228_n19360) );
  OR2X2 OR2X2_4632 ( .A(u2__abc_44228_n19363), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n19364) );
  OR2X2 OR2X2_4633 ( .A(u2__abc_44228_n19368), .B(u2__abc_44228_n19359), .Y(u2__abc_44228_n19369) );
  OR2X2 OR2X2_4634 ( .A(u2__abc_44228_n19361), .B(sqrto_132_), .Y(u2__abc_44228_n19372) );
  OR2X2 OR2X2_4635 ( .A(u2__abc_44228_n19375), .B(u2__abc_44228_n2983_bF_buf67), .Y(u2__abc_44228_n19376) );
  OR2X2 OR2X2_4636 ( .A(u2__abc_44228_n19380), .B(u2__abc_44228_n19371), .Y(u2__abc_44228_n19381) );
  OR2X2 OR2X2_4637 ( .A(u2__abc_44228_n19373), .B(sqrto_133_), .Y(u2__abc_44228_n19384) );
  OR2X2 OR2X2_4638 ( .A(u2__abc_44228_n19387), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n19388) );
  OR2X2 OR2X2_4639 ( .A(u2__abc_44228_n19392), .B(u2__abc_44228_n19383), .Y(u2__abc_44228_n19393) );
  OR2X2 OR2X2_464 ( .A(_abc_64468_n1557), .B(_abc_64468_n1554), .Y(_abc_64468_n1558) );
  OR2X2 OR2X2_4640 ( .A(u2__abc_44228_n19385), .B(sqrto_134_), .Y(u2__abc_44228_n19396) );
  OR2X2 OR2X2_4641 ( .A(u2__abc_44228_n19399), .B(u2__abc_44228_n2983_bF_buf63), .Y(u2__abc_44228_n19400) );
  OR2X2 OR2X2_4642 ( .A(u2__abc_44228_n19404), .B(u2__abc_44228_n19395), .Y(u2__abc_44228_n19405) );
  OR2X2 OR2X2_4643 ( .A(u2__abc_44228_n19397), .B(sqrto_135_), .Y(u2__abc_44228_n19408) );
  OR2X2 OR2X2_4644 ( .A(u2__abc_44228_n19411), .B(u2__abc_44228_n2983_bF_buf61), .Y(u2__abc_44228_n19412) );
  OR2X2 OR2X2_4645 ( .A(u2__abc_44228_n19416), .B(u2__abc_44228_n19407), .Y(u2__abc_44228_n19417) );
  OR2X2 OR2X2_4646 ( .A(u2__abc_44228_n19409), .B(sqrto_136_), .Y(u2__abc_44228_n19420) );
  OR2X2 OR2X2_4647 ( .A(u2__abc_44228_n19423), .B(u2__abc_44228_n2983_bF_buf59), .Y(u2__abc_44228_n19424) );
  OR2X2 OR2X2_4648 ( .A(u2__abc_44228_n19428), .B(u2__abc_44228_n19419), .Y(u2__abc_44228_n19429) );
  OR2X2 OR2X2_4649 ( .A(u2__abc_44228_n19421), .B(sqrto_137_), .Y(u2__abc_44228_n19432) );
  OR2X2 OR2X2_465 ( .A(_abc_64468_n1561), .B(aNan_bF_buf3), .Y(_abc_64468_n1562) );
  OR2X2 OR2X2_4650 ( .A(u2__abc_44228_n19435), .B(u2__abc_44228_n2983_bF_buf57), .Y(u2__abc_44228_n19436) );
  OR2X2 OR2X2_4651 ( .A(u2__abc_44228_n19440), .B(u2__abc_44228_n19431), .Y(u2__abc_44228_n19441) );
  OR2X2 OR2X2_4652 ( .A(u2__abc_44228_n19433), .B(sqrto_138_), .Y(u2__abc_44228_n19444) );
  OR2X2 OR2X2_4653 ( .A(u2__abc_44228_n19447), .B(u2__abc_44228_n2983_bF_buf55), .Y(u2__abc_44228_n19448) );
  OR2X2 OR2X2_4654 ( .A(u2__abc_44228_n19452), .B(u2__abc_44228_n19443), .Y(u2__abc_44228_n19453) );
  OR2X2 OR2X2_4655 ( .A(u2__abc_44228_n19445), .B(sqrto_139_), .Y(u2__abc_44228_n19456) );
  OR2X2 OR2X2_4656 ( .A(u2__abc_44228_n19459), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n19460) );
  OR2X2 OR2X2_4657 ( .A(u2__abc_44228_n19464), .B(u2__abc_44228_n19455), .Y(u2__abc_44228_n19465) );
  OR2X2 OR2X2_4658 ( .A(u2__abc_44228_n19457), .B(sqrto_140_), .Y(u2__abc_44228_n19468) );
  OR2X2 OR2X2_4659 ( .A(u2__abc_44228_n19471), .B(u2__abc_44228_n2983_bF_buf51), .Y(u2__abc_44228_n19472) );
  OR2X2 OR2X2_466 ( .A(_abc_64468_n1562), .B(_abc_64468_n1560), .Y(_abc_64468_n1563) );
  OR2X2 OR2X2_4660 ( .A(u2__abc_44228_n19476), .B(u2__abc_44228_n19467), .Y(u2__abc_44228_n19477) );
  OR2X2 OR2X2_4661 ( .A(u2__abc_44228_n19469), .B(sqrto_141_), .Y(u2__abc_44228_n19480) );
  OR2X2 OR2X2_4662 ( .A(u2__abc_44228_n19483), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n19484) );
  OR2X2 OR2X2_4663 ( .A(u2__abc_44228_n19488), .B(u2__abc_44228_n19479), .Y(u2__abc_44228_n19489) );
  OR2X2 OR2X2_4664 ( .A(u2__abc_44228_n19481), .B(sqrto_142_), .Y(u2__abc_44228_n19492) );
  OR2X2 OR2X2_4665 ( .A(u2__abc_44228_n19495), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n19496) );
  OR2X2 OR2X2_4666 ( .A(u2__abc_44228_n19500), .B(u2__abc_44228_n19491), .Y(u2__abc_44228_n19501) );
  OR2X2 OR2X2_4667 ( .A(u2__abc_44228_n19493), .B(sqrto_143_), .Y(u2__abc_44228_n19504) );
  OR2X2 OR2X2_4668 ( .A(u2__abc_44228_n19507), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n19508) );
  OR2X2 OR2X2_4669 ( .A(u2__abc_44228_n19512), .B(u2__abc_44228_n19503), .Y(u2__abc_44228_n19513) );
  OR2X2 OR2X2_467 ( .A(_abc_64468_n753_bF_buf1), .B(\a[116] ), .Y(_abc_64468_n1564) );
  OR2X2 OR2X2_4670 ( .A(u2__abc_44228_n19505), .B(sqrto_144_), .Y(u2__abc_44228_n19516) );
  OR2X2 OR2X2_4671 ( .A(u2__abc_44228_n19519), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n19520) );
  OR2X2 OR2X2_4672 ( .A(u2__abc_44228_n19524), .B(u2__abc_44228_n19515), .Y(u2__abc_44228_n19525) );
  OR2X2 OR2X2_4673 ( .A(u2__abc_44228_n19517), .B(sqrto_145_), .Y(u2__abc_44228_n19528) );
  OR2X2 OR2X2_4674 ( .A(u2__abc_44228_n19531), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n19532) );
  OR2X2 OR2X2_4675 ( .A(u2__abc_44228_n19536), .B(u2__abc_44228_n19527), .Y(u2__abc_44228_n19537) );
  OR2X2 OR2X2_4676 ( .A(u2__abc_44228_n19529), .B(sqrto_146_), .Y(u2__abc_44228_n19540) );
  OR2X2 OR2X2_4677 ( .A(u2__abc_44228_n19543), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n19544) );
  OR2X2 OR2X2_4678 ( .A(u2__abc_44228_n19548), .B(u2__abc_44228_n19539), .Y(u2__abc_44228_n19549) );
  OR2X2 OR2X2_4679 ( .A(u2__abc_44228_n19541), .B(sqrto_147_), .Y(u2__abc_44228_n19552) );
  OR2X2 OR2X2_468 ( .A(_abc_64468_n1554), .B(_abc_64468_n1568), .Y(_abc_64468_n1569) );
  OR2X2 OR2X2_4680 ( .A(u2__abc_44228_n19555), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n19556) );
  OR2X2 OR2X2_4681 ( .A(u2__abc_44228_n19560), .B(u2__abc_44228_n19551), .Y(u2__abc_44228_n19561) );
  OR2X2 OR2X2_4682 ( .A(u2__abc_44228_n19553), .B(sqrto_148_), .Y(u2__abc_44228_n19564) );
  OR2X2 OR2X2_4683 ( .A(u2__abc_44228_n19567), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n19568) );
  OR2X2 OR2X2_4684 ( .A(u2__abc_44228_n19572), .B(u2__abc_44228_n19563), .Y(u2__abc_44228_n19573) );
  OR2X2 OR2X2_4685 ( .A(u2__abc_44228_n19565), .B(sqrto_149_), .Y(u2__abc_44228_n19576) );
  OR2X2 OR2X2_4686 ( .A(u2__abc_44228_n19579), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n19580) );
  OR2X2 OR2X2_4687 ( .A(u2__abc_44228_n19584), .B(u2__abc_44228_n19575), .Y(u2__abc_44228_n19585) );
  OR2X2 OR2X2_4688 ( .A(u2__abc_44228_n19577), .B(sqrto_150_), .Y(u2__abc_44228_n19588) );
  OR2X2 OR2X2_4689 ( .A(u2__abc_44228_n19591), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n19592) );
  OR2X2 OR2X2_469 ( .A(_abc_64468_n1574), .B(_abc_64468_n1575), .Y(_abc_64468_n1576) );
  OR2X2 OR2X2_4690 ( .A(u2__abc_44228_n19596), .B(u2__abc_44228_n19587), .Y(u2__abc_44228_n19597) );
  OR2X2 OR2X2_4691 ( .A(u2__abc_44228_n19589), .B(sqrto_151_), .Y(u2__abc_44228_n19600) );
  OR2X2 OR2X2_4692 ( .A(u2__abc_44228_n19603), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n19604) );
  OR2X2 OR2X2_4693 ( .A(u2__abc_44228_n19608), .B(u2__abc_44228_n19599), .Y(u2__abc_44228_n19609) );
  OR2X2 OR2X2_4694 ( .A(u2__abc_44228_n19601), .B(sqrto_152_), .Y(u2__abc_44228_n19612) );
  OR2X2 OR2X2_4695 ( .A(u2__abc_44228_n19615), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n19616) );
  OR2X2 OR2X2_4696 ( .A(u2__abc_44228_n19620), .B(u2__abc_44228_n19611), .Y(u2__abc_44228_n19621) );
  OR2X2 OR2X2_4697 ( .A(u2__abc_44228_n19613), .B(sqrto_153_), .Y(u2__abc_44228_n19624) );
  OR2X2 OR2X2_4698 ( .A(u2__abc_44228_n19627), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n19628) );
  OR2X2 OR2X2_4699 ( .A(u2__abc_44228_n19632), .B(u2__abc_44228_n19623), .Y(u2__abc_44228_n19633) );
  OR2X2 OR2X2_47 ( .A(aNan_bF_buf8), .B(sqrto_99_), .Y(_abc_64468_n899) );
  OR2X2 OR2X2_470 ( .A(_abc_64468_n1577), .B(_abc_64468_n1566), .Y(_auto_iopadmap_cc_313_execute_65414_231_) );
  OR2X2 OR2X2_4700 ( .A(u2__abc_44228_n19625), .B(sqrto_154_), .Y(u2__abc_44228_n19636) );
  OR2X2 OR2X2_4701 ( .A(u2__abc_44228_n19639), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n19640) );
  OR2X2 OR2X2_4702 ( .A(u2__abc_44228_n19644), .B(u2__abc_44228_n19635), .Y(u2__abc_44228_n19645) );
  OR2X2 OR2X2_4703 ( .A(u2__abc_44228_n19637), .B(sqrto_155_), .Y(u2__abc_44228_n19648) );
  OR2X2 OR2X2_4704 ( .A(u2__abc_44228_n19651), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n19652) );
  OR2X2 OR2X2_4705 ( .A(u2__abc_44228_n19656), .B(u2__abc_44228_n19647), .Y(u2__abc_44228_n19657) );
  OR2X2 OR2X2_4706 ( .A(u2__abc_44228_n19649), .B(sqrto_156_), .Y(u2__abc_44228_n19660) );
  OR2X2 OR2X2_4707 ( .A(u2__abc_44228_n19663), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n19664) );
  OR2X2 OR2X2_4708 ( .A(u2__abc_44228_n19668), .B(u2__abc_44228_n19659), .Y(u2__abc_44228_n19669) );
  OR2X2 OR2X2_4709 ( .A(u2__abc_44228_n19661), .B(sqrto_157_), .Y(u2__abc_44228_n19672) );
  OR2X2 OR2X2_471 ( .A(_abc_64468_n1581), .B(_abc_64468_n1580), .Y(_abc_64468_n1582) );
  OR2X2 OR2X2_4710 ( .A(u2__abc_44228_n19675), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n19676) );
  OR2X2 OR2X2_4711 ( .A(u2__abc_44228_n19680), .B(u2__abc_44228_n19671), .Y(u2__abc_44228_n19681) );
  OR2X2 OR2X2_4712 ( .A(u2__abc_44228_n19673), .B(sqrto_158_), .Y(u2__abc_44228_n19684) );
  OR2X2 OR2X2_4713 ( .A(u2__abc_44228_n19687), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n19688) );
  OR2X2 OR2X2_4714 ( .A(u2__abc_44228_n19692), .B(u2__abc_44228_n19683), .Y(u2__abc_44228_n19693) );
  OR2X2 OR2X2_4715 ( .A(u2__abc_44228_n19685), .B(sqrto_159_), .Y(u2__abc_44228_n19696) );
  OR2X2 OR2X2_4716 ( .A(u2__abc_44228_n19699), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n19700) );
  OR2X2 OR2X2_4717 ( .A(u2__abc_44228_n19704), .B(u2__abc_44228_n19695), .Y(u2__abc_44228_n19705) );
  OR2X2 OR2X2_4718 ( .A(u2__abc_44228_n19697), .B(sqrto_160_), .Y(u2__abc_44228_n19708) );
  OR2X2 OR2X2_4719 ( .A(u2__abc_44228_n19711), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n19712) );
  OR2X2 OR2X2_472 ( .A(_abc_64468_n1587), .B(_abc_64468_n1588), .Y(_abc_64468_n1589) );
  OR2X2 OR2X2_4720 ( .A(u2__abc_44228_n19716), .B(u2__abc_44228_n19707), .Y(u2__abc_44228_n19717) );
  OR2X2 OR2X2_4721 ( .A(u2__abc_44228_n19709), .B(sqrto_161_), .Y(u2__abc_44228_n19720) );
  OR2X2 OR2X2_4722 ( .A(u2__abc_44228_n19723), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n19724) );
  OR2X2 OR2X2_4723 ( .A(u2__abc_44228_n19728), .B(u2__abc_44228_n19719), .Y(u2__abc_44228_n19729) );
  OR2X2 OR2X2_4724 ( .A(u2__abc_44228_n19721), .B(sqrto_162_), .Y(u2__abc_44228_n19732) );
  OR2X2 OR2X2_4725 ( .A(u2__abc_44228_n19735), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n19736) );
  OR2X2 OR2X2_4726 ( .A(u2__abc_44228_n19740), .B(u2__abc_44228_n19731), .Y(u2__abc_44228_n19741) );
  OR2X2 OR2X2_4727 ( .A(u2__abc_44228_n19733), .B(sqrto_163_), .Y(u2__abc_44228_n19744) );
  OR2X2 OR2X2_4728 ( .A(u2__abc_44228_n19747), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n19748) );
  OR2X2 OR2X2_4729 ( .A(u2__abc_44228_n19752), .B(u2__abc_44228_n19743), .Y(u2__abc_44228_n19753) );
  OR2X2 OR2X2_473 ( .A(_abc_64468_n1590), .B(_abc_64468_n1591), .Y(_auto_iopadmap_cc_313_execute_65414_232_) );
  OR2X2 OR2X2_4730 ( .A(u2__abc_44228_n19745), .B(sqrto_164_), .Y(u2__abc_44228_n19756) );
  OR2X2 OR2X2_4731 ( .A(u2__abc_44228_n19759), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n19760) );
  OR2X2 OR2X2_4732 ( .A(u2__abc_44228_n19764), .B(u2__abc_44228_n19755), .Y(u2__abc_44228_n19765) );
  OR2X2 OR2X2_4733 ( .A(u2__abc_44228_n19757), .B(sqrto_165_), .Y(u2__abc_44228_n19768) );
  OR2X2 OR2X2_4734 ( .A(u2__abc_44228_n19771), .B(u2__abc_44228_n2983_bF_buf1), .Y(u2__abc_44228_n19772) );
  OR2X2 OR2X2_4735 ( .A(u2__abc_44228_n19776), .B(u2__abc_44228_n19767), .Y(u2__abc_44228_n19777) );
  OR2X2 OR2X2_4736 ( .A(u2__abc_44228_n19769), .B(sqrto_166_), .Y(u2__abc_44228_n19780) );
  OR2X2 OR2X2_4737 ( .A(u2__abc_44228_n19783), .B(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n19784) );
  OR2X2 OR2X2_4738 ( .A(u2__abc_44228_n19788), .B(u2__abc_44228_n19779), .Y(u2__abc_44228_n19789) );
  OR2X2 OR2X2_4739 ( .A(u2__abc_44228_n19781), .B(sqrto_167_), .Y(u2__abc_44228_n19792) );
  OR2X2 OR2X2_474 ( .A(_abc_64468_n1596), .B(_abc_64468_n1595), .Y(_abc_64468_n1597) );
  OR2X2 OR2X2_4740 ( .A(u2__abc_44228_n19795), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n19796) );
  OR2X2 OR2X2_4741 ( .A(u2__abc_44228_n19800), .B(u2__abc_44228_n19791), .Y(u2__abc_44228_n19801) );
  OR2X2 OR2X2_4742 ( .A(u2__abc_44228_n19793), .B(sqrto_168_), .Y(u2__abc_44228_n19804) );
  OR2X2 OR2X2_4743 ( .A(u2__abc_44228_n19807), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n19808) );
  OR2X2 OR2X2_4744 ( .A(u2__abc_44228_n19812), .B(u2__abc_44228_n19803), .Y(u2__abc_44228_n19813) );
  OR2X2 OR2X2_4745 ( .A(u2__abc_44228_n19805), .B(sqrto_169_), .Y(u2__abc_44228_n19816) );
  OR2X2 OR2X2_4746 ( .A(u2__abc_44228_n19819), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n19820) );
  OR2X2 OR2X2_4747 ( .A(u2__abc_44228_n19824), .B(u2__abc_44228_n19815), .Y(u2__abc_44228_n19825) );
  OR2X2 OR2X2_4748 ( .A(u2__abc_44228_n19817), .B(sqrto_170_), .Y(u2__abc_44228_n19828) );
  OR2X2 OR2X2_4749 ( .A(u2__abc_44228_n19831), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n19832) );
  OR2X2 OR2X2_475 ( .A(_abc_64468_n1602), .B(_abc_64468_n1603), .Y(_abc_64468_n1604) );
  OR2X2 OR2X2_4750 ( .A(u2__abc_44228_n19836), .B(u2__abc_44228_n19827), .Y(u2__abc_44228_n19837) );
  OR2X2 OR2X2_4751 ( .A(u2__abc_44228_n19829), .B(sqrto_171_), .Y(u2__abc_44228_n19840) );
  OR2X2 OR2X2_4752 ( .A(u2__abc_44228_n19843), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n19844) );
  OR2X2 OR2X2_4753 ( .A(u2__abc_44228_n19848), .B(u2__abc_44228_n19839), .Y(u2__abc_44228_n19849) );
  OR2X2 OR2X2_4754 ( .A(u2__abc_44228_n19841), .B(sqrto_172_), .Y(u2__abc_44228_n19852) );
  OR2X2 OR2X2_4755 ( .A(u2__abc_44228_n19855), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n19856) );
  OR2X2 OR2X2_4756 ( .A(u2__abc_44228_n19860), .B(u2__abc_44228_n19851), .Y(u2__abc_44228_n19861) );
  OR2X2 OR2X2_4757 ( .A(u2__abc_44228_n19853), .B(sqrto_173_), .Y(u2__abc_44228_n19864) );
  OR2X2 OR2X2_4758 ( .A(u2__abc_44228_n19867), .B(u2__abc_44228_n2983_bF_buf127), .Y(u2__abc_44228_n19868) );
  OR2X2 OR2X2_4759 ( .A(u2__abc_44228_n19872), .B(u2__abc_44228_n19863), .Y(u2__abc_44228_n19873) );
  OR2X2 OR2X2_476 ( .A(_abc_64468_n1605), .B(_abc_64468_n1593), .Y(_auto_iopadmap_cc_313_execute_65414_233_) );
  OR2X2 OR2X2_4760 ( .A(u2__abc_44228_n19865), .B(sqrto_174_), .Y(u2__abc_44228_n19876) );
  OR2X2 OR2X2_4761 ( .A(u2__abc_44228_n19879), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n19880) );
  OR2X2 OR2X2_4762 ( .A(u2__abc_44228_n19884), .B(u2__abc_44228_n19875), .Y(u2__abc_44228_n19885) );
  OR2X2 OR2X2_4763 ( .A(u2__abc_44228_n19877), .B(sqrto_175_), .Y(u2__abc_44228_n19888) );
  OR2X2 OR2X2_4764 ( .A(u2__abc_44228_n19891), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n19892) );
  OR2X2 OR2X2_4765 ( .A(u2__abc_44228_n19896), .B(u2__abc_44228_n19887), .Y(u2__abc_44228_n19897) );
  OR2X2 OR2X2_4766 ( .A(u2__abc_44228_n19889), .B(sqrto_176_), .Y(u2__abc_44228_n19900) );
  OR2X2 OR2X2_4767 ( .A(u2__abc_44228_n19903), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n19904) );
  OR2X2 OR2X2_4768 ( .A(u2__abc_44228_n19908), .B(u2__abc_44228_n19899), .Y(u2__abc_44228_n19909) );
  OR2X2 OR2X2_4769 ( .A(u2__abc_44228_n19901), .B(sqrto_177_), .Y(u2__abc_44228_n19912) );
  OR2X2 OR2X2_477 ( .A(_abc_64468_n1609), .B(_abc_64468_n1608), .Y(_abc_64468_n1610) );
  OR2X2 OR2X2_4770 ( .A(u2__abc_44228_n19915), .B(u2__abc_44228_n2983_bF_buf119), .Y(u2__abc_44228_n19916) );
  OR2X2 OR2X2_4771 ( .A(u2__abc_44228_n19920), .B(u2__abc_44228_n19911), .Y(u2__abc_44228_n19921) );
  OR2X2 OR2X2_4772 ( .A(u2__abc_44228_n19913), .B(sqrto_178_), .Y(u2__abc_44228_n19924) );
  OR2X2 OR2X2_4773 ( .A(u2__abc_44228_n19927), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n19928) );
  OR2X2 OR2X2_4774 ( .A(u2__abc_44228_n19932), .B(u2__abc_44228_n19923), .Y(u2__abc_44228_n19933) );
  OR2X2 OR2X2_4775 ( .A(u2__abc_44228_n19925), .B(sqrto_179_), .Y(u2__abc_44228_n19936) );
  OR2X2 OR2X2_4776 ( .A(u2__abc_44228_n19939), .B(u2__abc_44228_n2983_bF_buf115), .Y(u2__abc_44228_n19940) );
  OR2X2 OR2X2_4777 ( .A(u2__abc_44228_n19944), .B(u2__abc_44228_n19935), .Y(u2__abc_44228_n19945) );
  OR2X2 OR2X2_4778 ( .A(u2__abc_44228_n19937), .B(sqrto_180_), .Y(u2__abc_44228_n19948) );
  OR2X2 OR2X2_4779 ( .A(u2__abc_44228_n19951), .B(u2__abc_44228_n2983_bF_buf113), .Y(u2__abc_44228_n19952) );
  OR2X2 OR2X2_478 ( .A(_abc_64468_n1615), .B(_abc_64468_n1616), .Y(_abc_64468_n1617) );
  OR2X2 OR2X2_4780 ( .A(u2__abc_44228_n19956), .B(u2__abc_44228_n19947), .Y(u2__abc_44228_n19957) );
  OR2X2 OR2X2_4781 ( .A(u2__abc_44228_n19949), .B(sqrto_181_), .Y(u2__abc_44228_n19960) );
  OR2X2 OR2X2_4782 ( .A(u2__abc_44228_n19963), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n19964) );
  OR2X2 OR2X2_4783 ( .A(u2__abc_44228_n19968), .B(u2__abc_44228_n19959), .Y(u2__abc_44228_n19969) );
  OR2X2 OR2X2_4784 ( .A(u2__abc_44228_n19961), .B(sqrto_182_), .Y(u2__abc_44228_n19972) );
  OR2X2 OR2X2_4785 ( .A(u2__abc_44228_n19975), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n19976) );
  OR2X2 OR2X2_4786 ( .A(u2__abc_44228_n19980), .B(u2__abc_44228_n19971), .Y(u2__abc_44228_n19981) );
  OR2X2 OR2X2_4787 ( .A(u2__abc_44228_n19973), .B(sqrto_183_), .Y(u2__abc_44228_n19984) );
  OR2X2 OR2X2_4788 ( .A(u2__abc_44228_n19987), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n19988) );
  OR2X2 OR2X2_4789 ( .A(u2__abc_44228_n19992), .B(u2__abc_44228_n19983), .Y(u2__abc_44228_n19993) );
  OR2X2 OR2X2_479 ( .A(_abc_64468_n1618), .B(_abc_64468_n1619), .Y(_auto_iopadmap_cc_313_execute_65414_234_) );
  OR2X2 OR2X2_4790 ( .A(u2__abc_44228_n19985), .B(sqrto_184_), .Y(u2__abc_44228_n19996) );
  OR2X2 OR2X2_4791 ( .A(u2__abc_44228_n19999), .B(u2__abc_44228_n2983_bF_buf105), .Y(u2__abc_44228_n20000) );
  OR2X2 OR2X2_4792 ( .A(u2__abc_44228_n20004), .B(u2__abc_44228_n19995), .Y(u2__abc_44228_n20005) );
  OR2X2 OR2X2_4793 ( .A(u2__abc_44228_n19997), .B(sqrto_185_), .Y(u2__abc_44228_n20008) );
  OR2X2 OR2X2_4794 ( .A(u2__abc_44228_n20011), .B(u2__abc_44228_n2983_bF_buf103), .Y(u2__abc_44228_n20012) );
  OR2X2 OR2X2_4795 ( .A(u2__abc_44228_n20016), .B(u2__abc_44228_n20007), .Y(u2__abc_44228_n20017) );
  OR2X2 OR2X2_4796 ( .A(u2__abc_44228_n20009), .B(sqrto_186_), .Y(u2__abc_44228_n20020) );
  OR2X2 OR2X2_4797 ( .A(u2__abc_44228_n20023), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n20024) );
  OR2X2 OR2X2_4798 ( .A(u2__abc_44228_n20028), .B(u2__abc_44228_n20019), .Y(u2__abc_44228_n20029) );
  OR2X2 OR2X2_4799 ( .A(u2__abc_44228_n20021), .B(sqrto_187_), .Y(u2__abc_44228_n20032) );
  OR2X2 OR2X2_48 ( .A(_abc_64468_n753_bF_buf12), .B(\a[23] ), .Y(_abc_64468_n900) );
  OR2X2 OR2X2_480 ( .A(_abc_64468_n1624), .B(_abc_64468_n1623), .Y(_abc_64468_n1625) );
  OR2X2 OR2X2_4800 ( .A(u2__abc_44228_n20035), .B(u2__abc_44228_n2983_bF_buf99), .Y(u2__abc_44228_n20036) );
  OR2X2 OR2X2_4801 ( .A(u2__abc_44228_n20040), .B(u2__abc_44228_n20031), .Y(u2__abc_44228_n20041) );
  OR2X2 OR2X2_4802 ( .A(u2__abc_44228_n20033), .B(sqrto_188_), .Y(u2__abc_44228_n20044) );
  OR2X2 OR2X2_4803 ( .A(u2__abc_44228_n20047), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n20048) );
  OR2X2 OR2X2_4804 ( .A(u2__abc_44228_n20052), .B(u2__abc_44228_n20043), .Y(u2__abc_44228_n20053) );
  OR2X2 OR2X2_4805 ( .A(u2__abc_44228_n20045), .B(sqrto_189_), .Y(u2__abc_44228_n20056) );
  OR2X2 OR2X2_4806 ( .A(u2__abc_44228_n20059), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n20060) );
  OR2X2 OR2X2_4807 ( .A(u2__abc_44228_n20064), .B(u2__abc_44228_n20055), .Y(u2__abc_44228_n20065) );
  OR2X2 OR2X2_4808 ( .A(u2__abc_44228_n20057), .B(sqrto_190_), .Y(u2__abc_44228_n20068) );
  OR2X2 OR2X2_4809 ( .A(u2__abc_44228_n20071), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n20072) );
  OR2X2 OR2X2_481 ( .A(_abc_64468_n1630), .B(_abc_64468_n1631), .Y(_abc_64468_n1632) );
  OR2X2 OR2X2_4810 ( .A(u2__abc_44228_n20076), .B(u2__abc_44228_n20067), .Y(u2__abc_44228_n20077) );
  OR2X2 OR2X2_4811 ( .A(u2__abc_44228_n20069), .B(sqrto_191_), .Y(u2__abc_44228_n20080) );
  OR2X2 OR2X2_4812 ( .A(u2__abc_44228_n20083), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n20084) );
  OR2X2 OR2X2_4813 ( .A(u2__abc_44228_n20088), .B(u2__abc_44228_n20079), .Y(u2__abc_44228_n20089) );
  OR2X2 OR2X2_4814 ( .A(u2__abc_44228_n20081), .B(sqrto_192_), .Y(u2__abc_44228_n20092) );
  OR2X2 OR2X2_4815 ( .A(u2__abc_44228_n20095), .B(u2__abc_44228_n2983_bF_buf89), .Y(u2__abc_44228_n20096) );
  OR2X2 OR2X2_4816 ( .A(u2__abc_44228_n20100), .B(u2__abc_44228_n20091), .Y(u2__abc_44228_n20101) );
  OR2X2 OR2X2_4817 ( .A(u2__abc_44228_n20093), .B(sqrto_193_), .Y(u2__abc_44228_n20104) );
  OR2X2 OR2X2_4818 ( .A(u2__abc_44228_n20107), .B(u2__abc_44228_n2983_bF_buf87), .Y(u2__abc_44228_n20108) );
  OR2X2 OR2X2_4819 ( .A(u2__abc_44228_n20112), .B(u2__abc_44228_n20103), .Y(u2__abc_44228_n20113) );
  OR2X2 OR2X2_482 ( .A(_abc_64468_n1633), .B(_abc_64468_n1621), .Y(_auto_iopadmap_cc_313_execute_65414_235_) );
  OR2X2 OR2X2_4820 ( .A(u2__abc_44228_n20105), .B(sqrto_194_), .Y(u2__abc_44228_n20116) );
  OR2X2 OR2X2_4821 ( .A(u2__abc_44228_n20119), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n20120) );
  OR2X2 OR2X2_4822 ( .A(u2__abc_44228_n20124), .B(u2__abc_44228_n20115), .Y(u2__abc_44228_n20125) );
  OR2X2 OR2X2_4823 ( .A(u2__abc_44228_n20117), .B(sqrto_195_), .Y(u2__abc_44228_n20128) );
  OR2X2 OR2X2_4824 ( .A(u2__abc_44228_n20131), .B(u2__abc_44228_n2983_bF_buf83), .Y(u2__abc_44228_n20132) );
  OR2X2 OR2X2_4825 ( .A(u2__abc_44228_n20136), .B(u2__abc_44228_n20127), .Y(u2__abc_44228_n20137) );
  OR2X2 OR2X2_4826 ( .A(u2__abc_44228_n20129), .B(sqrto_196_), .Y(u2__abc_44228_n20140) );
  OR2X2 OR2X2_4827 ( .A(u2__abc_44228_n20143), .B(u2__abc_44228_n2983_bF_buf81), .Y(u2__abc_44228_n20144) );
  OR2X2 OR2X2_4828 ( .A(u2__abc_44228_n20148), .B(u2__abc_44228_n20139), .Y(u2__abc_44228_n20149) );
  OR2X2 OR2X2_4829 ( .A(u2__abc_44228_n20141), .B(sqrto_197_), .Y(u2__abc_44228_n20152) );
  OR2X2 OR2X2_483 ( .A(_abc_64468_n1637), .B(_abc_64468_n1636), .Y(_abc_64468_n1638) );
  OR2X2 OR2X2_4830 ( .A(u2__abc_44228_n20155), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n20156) );
  OR2X2 OR2X2_4831 ( .A(u2__abc_44228_n20160), .B(u2__abc_44228_n20151), .Y(u2__abc_44228_n20161) );
  OR2X2 OR2X2_4832 ( .A(u2__abc_44228_n20153), .B(sqrto_198_), .Y(u2__abc_44228_n20164) );
  OR2X2 OR2X2_4833 ( .A(u2__abc_44228_n20167), .B(u2__abc_44228_n2983_bF_buf77), .Y(u2__abc_44228_n20168) );
  OR2X2 OR2X2_4834 ( .A(u2__abc_44228_n20172), .B(u2__abc_44228_n20163), .Y(u2__abc_44228_n20173) );
  OR2X2 OR2X2_4835 ( .A(u2__abc_44228_n20165), .B(sqrto_199_), .Y(u2__abc_44228_n20176) );
  OR2X2 OR2X2_4836 ( .A(u2__abc_44228_n20179), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n20180) );
  OR2X2 OR2X2_4837 ( .A(u2__abc_44228_n20184), .B(u2__abc_44228_n20175), .Y(u2__abc_44228_n20185) );
  OR2X2 OR2X2_4838 ( .A(u2__abc_44228_n20177), .B(sqrto_200_), .Y(u2__abc_44228_n20188) );
  OR2X2 OR2X2_4839 ( .A(u2__abc_44228_n20191), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n20192) );
  OR2X2 OR2X2_484 ( .A(_abc_64468_n1643), .B(_abc_64468_n1644), .Y(_abc_64468_n1645) );
  OR2X2 OR2X2_4840 ( .A(u2__abc_44228_n20196), .B(u2__abc_44228_n20187), .Y(u2__abc_44228_n20197) );
  OR2X2 OR2X2_4841 ( .A(u2__abc_44228_n20189), .B(sqrto_201_), .Y(u2__abc_44228_n20200) );
  OR2X2 OR2X2_4842 ( .A(u2__abc_44228_n20203), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n20204) );
  OR2X2 OR2X2_4843 ( .A(u2__abc_44228_n20208), .B(u2__abc_44228_n20199), .Y(u2__abc_44228_n20209) );
  OR2X2 OR2X2_4844 ( .A(u2__abc_44228_n20201), .B(sqrto_202_), .Y(u2__abc_44228_n20212) );
  OR2X2 OR2X2_4845 ( .A(u2__abc_44228_n20215), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n20216) );
  OR2X2 OR2X2_4846 ( .A(u2__abc_44228_n20220), .B(u2__abc_44228_n20211), .Y(u2__abc_44228_n20221) );
  OR2X2 OR2X2_4847 ( .A(u2__abc_44228_n20213), .B(sqrto_203_), .Y(u2__abc_44228_n20224) );
  OR2X2 OR2X2_4848 ( .A(u2__abc_44228_n20227), .B(u2__abc_44228_n2983_bF_buf67), .Y(u2__abc_44228_n20228) );
  OR2X2 OR2X2_4849 ( .A(u2__abc_44228_n20232), .B(u2__abc_44228_n20223), .Y(u2__abc_44228_n20233) );
  OR2X2 OR2X2_485 ( .A(_abc_64468_n1646), .B(_abc_64468_n1647), .Y(_auto_iopadmap_cc_313_execute_65414_236_) );
  OR2X2 OR2X2_4850 ( .A(u2__abc_44228_n20225), .B(sqrto_204_), .Y(u2__abc_44228_n20236) );
  OR2X2 OR2X2_4851 ( .A(u2__abc_44228_n20239), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n20240) );
  OR2X2 OR2X2_4852 ( .A(u2__abc_44228_n20244), .B(u2__abc_44228_n20235), .Y(u2__abc_44228_n20245) );
  OR2X2 OR2X2_4853 ( .A(u2__abc_44228_n20237), .B(sqrto_205_), .Y(u2__abc_44228_n20248) );
  OR2X2 OR2X2_4854 ( .A(u2__abc_44228_n20251), .B(u2__abc_44228_n2983_bF_buf63), .Y(u2__abc_44228_n20252) );
  OR2X2 OR2X2_4855 ( .A(u2__abc_44228_n20256), .B(u2__abc_44228_n20247), .Y(u2__abc_44228_n20257) );
  OR2X2 OR2X2_4856 ( .A(u2__abc_44228_n20249), .B(sqrto_206_), .Y(u2__abc_44228_n20260) );
  OR2X2 OR2X2_4857 ( .A(u2__abc_44228_n20263), .B(u2__abc_44228_n2983_bF_buf61), .Y(u2__abc_44228_n20264) );
  OR2X2 OR2X2_4858 ( .A(u2__abc_44228_n20268), .B(u2__abc_44228_n20259), .Y(u2__abc_44228_n20269) );
  OR2X2 OR2X2_4859 ( .A(u2__abc_44228_n20261), .B(sqrto_207_), .Y(u2__abc_44228_n20272) );
  OR2X2 OR2X2_486 ( .A(_abc_64468_n1652), .B(_abc_64468_n1651), .Y(_abc_64468_n1653) );
  OR2X2 OR2X2_4860 ( .A(u2__abc_44228_n20275), .B(u2__abc_44228_n2983_bF_buf59), .Y(u2__abc_44228_n20276) );
  OR2X2 OR2X2_4861 ( .A(u2__abc_44228_n20280), .B(u2__abc_44228_n20271), .Y(u2__abc_44228_n20281) );
  OR2X2 OR2X2_4862 ( .A(u2__abc_44228_n20273), .B(sqrto_208_), .Y(u2__abc_44228_n20284) );
  OR2X2 OR2X2_4863 ( .A(u2__abc_44228_n20287), .B(u2__abc_44228_n2983_bF_buf57), .Y(u2__abc_44228_n20288) );
  OR2X2 OR2X2_4864 ( .A(u2__abc_44228_n20292), .B(u2__abc_44228_n20283), .Y(u2__abc_44228_n20293) );
  OR2X2 OR2X2_4865 ( .A(u2__abc_44228_n20285), .B(sqrto_209_), .Y(u2__abc_44228_n20296) );
  OR2X2 OR2X2_4866 ( .A(u2__abc_44228_n20299), .B(u2__abc_44228_n2983_bF_buf55), .Y(u2__abc_44228_n20300) );
  OR2X2 OR2X2_4867 ( .A(u2__abc_44228_n20304), .B(u2__abc_44228_n20295), .Y(u2__abc_44228_n20305) );
  OR2X2 OR2X2_4868 ( .A(u2__abc_44228_n20297), .B(sqrto_210_), .Y(u2__abc_44228_n20308) );
  OR2X2 OR2X2_4869 ( .A(u2__abc_44228_n20311), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n20312) );
  OR2X2 OR2X2_487 ( .A(_abc_64468_n1658), .B(_abc_64468_n1659), .Y(_abc_64468_n1660) );
  OR2X2 OR2X2_4870 ( .A(u2__abc_44228_n20316), .B(u2__abc_44228_n20307), .Y(u2__abc_44228_n20317) );
  OR2X2 OR2X2_4871 ( .A(u2__abc_44228_n20309), .B(sqrto_211_), .Y(u2__abc_44228_n20320) );
  OR2X2 OR2X2_4872 ( .A(u2__abc_44228_n20323), .B(u2__abc_44228_n2983_bF_buf51), .Y(u2__abc_44228_n20324) );
  OR2X2 OR2X2_4873 ( .A(u2__abc_44228_n20328), .B(u2__abc_44228_n20319), .Y(u2__abc_44228_n20329) );
  OR2X2 OR2X2_4874 ( .A(u2__abc_44228_n20321), .B(sqrto_212_), .Y(u2__abc_44228_n20332) );
  OR2X2 OR2X2_4875 ( .A(u2__abc_44228_n20335), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n20336) );
  OR2X2 OR2X2_4876 ( .A(u2__abc_44228_n20340), .B(u2__abc_44228_n20331), .Y(u2__abc_44228_n20341) );
  OR2X2 OR2X2_4877 ( .A(u2__abc_44228_n20333), .B(sqrto_213_), .Y(u2__abc_44228_n20344) );
  OR2X2 OR2X2_4878 ( .A(u2__abc_44228_n20347), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n20348) );
  OR2X2 OR2X2_4879 ( .A(u2__abc_44228_n20352), .B(u2__abc_44228_n20343), .Y(u2__abc_44228_n20353) );
  OR2X2 OR2X2_488 ( .A(_abc_64468_n1661), .B(_abc_64468_n1649), .Y(_auto_iopadmap_cc_313_execute_65414_237_) );
  OR2X2 OR2X2_4880 ( .A(u2__abc_44228_n20345), .B(sqrto_214_), .Y(u2__abc_44228_n20356) );
  OR2X2 OR2X2_4881 ( .A(u2__abc_44228_n20359), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n20360) );
  OR2X2 OR2X2_4882 ( .A(u2__abc_44228_n20364), .B(u2__abc_44228_n20355), .Y(u2__abc_44228_n20365) );
  OR2X2 OR2X2_4883 ( .A(u2__abc_44228_n20357), .B(sqrto_215_), .Y(u2__abc_44228_n20368) );
  OR2X2 OR2X2_4884 ( .A(u2__abc_44228_n20371), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n20372) );
  OR2X2 OR2X2_4885 ( .A(u2__abc_44228_n20376), .B(u2__abc_44228_n20367), .Y(u2__abc_44228_n20377) );
  OR2X2 OR2X2_4886 ( .A(u2__abc_44228_n20369), .B(sqrto_216_), .Y(u2__abc_44228_n20380) );
  OR2X2 OR2X2_4887 ( .A(u2__abc_44228_n20383), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n20384) );
  OR2X2 OR2X2_4888 ( .A(u2__abc_44228_n20388), .B(u2__abc_44228_n20379), .Y(u2__abc_44228_n20389) );
  OR2X2 OR2X2_4889 ( .A(u2__abc_44228_n20381), .B(sqrto_217_), .Y(u2__abc_44228_n20392) );
  OR2X2 OR2X2_489 ( .A(_abc_64468_n1665), .B(_abc_64468_n1664), .Y(_abc_64468_n1666) );
  OR2X2 OR2X2_4890 ( .A(u2__abc_44228_n20395), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n20396) );
  OR2X2 OR2X2_4891 ( .A(u2__abc_44228_n20400), .B(u2__abc_44228_n20391), .Y(u2__abc_44228_n20401) );
  OR2X2 OR2X2_4892 ( .A(u2__abc_44228_n20393), .B(sqrto_218_), .Y(u2__abc_44228_n20404) );
  OR2X2 OR2X2_4893 ( .A(u2__abc_44228_n20407), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n20408) );
  OR2X2 OR2X2_4894 ( .A(u2__abc_44228_n20412), .B(u2__abc_44228_n20403), .Y(u2__abc_44228_n20413) );
  OR2X2 OR2X2_4895 ( .A(u2__abc_44228_n20405), .B(sqrto_219_), .Y(u2__abc_44228_n20416) );
  OR2X2 OR2X2_4896 ( .A(u2__abc_44228_n20419), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n20420) );
  OR2X2 OR2X2_4897 ( .A(u2__abc_44228_n20424), .B(u2__abc_44228_n20415), .Y(u2__abc_44228_n20425) );
  OR2X2 OR2X2_4898 ( .A(u2__abc_44228_n20417), .B(sqrto_220_), .Y(u2__abc_44228_n20428) );
  OR2X2 OR2X2_4899 ( .A(u2__abc_44228_n20431), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n20432) );
  OR2X2 OR2X2_49 ( .A(aNan_bF_buf7), .B(sqrto_100_), .Y(_abc_64468_n902) );
  OR2X2 OR2X2_490 ( .A(_abc_64468_n1671), .B(_abc_64468_n1672), .Y(_abc_64468_n1673) );
  OR2X2 OR2X2_4900 ( .A(u2__abc_44228_n20436), .B(u2__abc_44228_n20427), .Y(u2__abc_44228_n20437) );
  OR2X2 OR2X2_4901 ( .A(u2__abc_44228_n20429), .B(sqrto_221_), .Y(u2__abc_44228_n20440) );
  OR2X2 OR2X2_4902 ( .A(u2__abc_44228_n20443), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n20444) );
  OR2X2 OR2X2_4903 ( .A(u2__abc_44228_n20448), .B(u2__abc_44228_n20439), .Y(u2__abc_44228_n20449) );
  OR2X2 OR2X2_4904 ( .A(u2__abc_44228_n20441), .B(sqrto_222_), .Y(u2__abc_44228_n20452) );
  OR2X2 OR2X2_4905 ( .A(u2__abc_44228_n20455), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n20456) );
  OR2X2 OR2X2_4906 ( .A(u2__abc_44228_n20460), .B(u2__abc_44228_n20451), .Y(u2__abc_44228_n20461) );
  OR2X2 OR2X2_4907 ( .A(u2__abc_44228_n20453), .B(sqrto_223_), .Y(u2__abc_44228_n20464) );
  OR2X2 OR2X2_4908 ( .A(u2__abc_44228_n20467), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n20468) );
  OR2X2 OR2X2_4909 ( .A(u2__abc_44228_n20472), .B(u2__abc_44228_n20463), .Y(u2__abc_44228_n20473) );
  OR2X2 OR2X2_491 ( .A(_abc_64468_n1674), .B(_abc_64468_n1675), .Y(_auto_iopadmap_cc_313_execute_65414_238_) );
  OR2X2 OR2X2_4910 ( .A(u2__abc_44228_n20465), .B(sqrto_224_), .Y(u2__abc_44228_n20476) );
  OR2X2 OR2X2_4911 ( .A(u2__abc_44228_n20479), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n20480) );
  OR2X2 OR2X2_4912 ( .A(u2__abc_44228_n20484), .B(u2__abc_44228_n20475), .Y(u2__abc_44228_n20485) );
  OR2X2 OR2X2_4913 ( .A(u2__abc_44228_n20477), .B(sqrto_225_), .Y(u2__abc_44228_n20488) );
  OR2X2 OR2X2_4914 ( .A(u2__abc_44228_n20491), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n20492) );
  OR2X2 OR2X2_4915 ( .A(u2__abc_44228_n20496), .B(u2__abc_44228_n20487), .Y(u2__abc_44228_n20497) );
  OR2X2 OR2X2_4916 ( .A(u2__abc_44228_n20489), .B(u2_o_226_), .Y(u2__abc_44228_n20500) );
  OR2X2 OR2X2_4917 ( .A(u2__abc_44228_n20503), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n20504) );
  OR2X2 OR2X2_4918 ( .A(u2__abc_44228_n20508), .B(u2__abc_44228_n20499), .Y(u2__abc_44228_n20509) );
  OR2X2 OR2X2_4919 ( .A(u2__abc_44228_n20501), .B(u2_o_227_), .Y(u2__abc_44228_n20512) );
  OR2X2 OR2X2_492 ( .A(_abc_64468_n753_bF_buf6), .B(\a[125] ), .Y(_abc_64468_n1677) );
  OR2X2 OR2X2_4920 ( .A(u2__abc_44228_n20515), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n20516) );
  OR2X2 OR2X2_4921 ( .A(u2__abc_44228_n20520), .B(u2__abc_44228_n20511), .Y(u2__abc_44228_n20521) );
  OR2X2 OR2X2_4922 ( .A(u2__abc_44228_n20513), .B(u2_o_228_), .Y(u2__abc_44228_n20524) );
  OR2X2 OR2X2_4923 ( .A(u2__abc_44228_n20527), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n20528) );
  OR2X2 OR2X2_4924 ( .A(u2__abc_44228_n20532), .B(u2__abc_44228_n20523), .Y(u2__abc_44228_n20533) );
  OR2X2 OR2X2_4925 ( .A(u2__abc_44228_n20525), .B(u2_o_229_), .Y(u2__abc_44228_n20536) );
  OR2X2 OR2X2_4926 ( .A(u2__abc_44228_n20539), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n20540) );
  OR2X2 OR2X2_4927 ( .A(u2__abc_44228_n20544), .B(u2__abc_44228_n20535), .Y(u2__abc_44228_n20545) );
  OR2X2 OR2X2_4928 ( .A(u2__abc_44228_n20537), .B(u2_o_230_), .Y(u2__abc_44228_n20548) );
  OR2X2 OR2X2_4929 ( .A(u2__abc_44228_n20551), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n20552) );
  OR2X2 OR2X2_493 ( .A(_abc_64468_n1679), .B(_abc_64468_n1678), .Y(_abc_64468_n1680) );
  OR2X2 OR2X2_4930 ( .A(u2__abc_44228_n20556), .B(u2__abc_44228_n20547), .Y(u2__abc_44228_n20557) );
  OR2X2 OR2X2_4931 ( .A(u2__abc_44228_n20549), .B(u2_o_231_), .Y(u2__abc_44228_n20560) );
  OR2X2 OR2X2_4932 ( .A(u2__abc_44228_n20563), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n20564) );
  OR2X2 OR2X2_4933 ( .A(u2__abc_44228_n20568), .B(u2__abc_44228_n20559), .Y(u2__abc_44228_n20569) );
  OR2X2 OR2X2_4934 ( .A(u2__abc_44228_n20561), .B(u2_o_232_), .Y(u2__abc_44228_n20572) );
  OR2X2 OR2X2_4935 ( .A(u2__abc_44228_n20575), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n20576) );
  OR2X2 OR2X2_4936 ( .A(u2__abc_44228_n20580), .B(u2__abc_44228_n20571), .Y(u2__abc_44228_n20581) );
  OR2X2 OR2X2_4937 ( .A(u2__abc_44228_n20573), .B(u2_o_233_), .Y(u2__abc_44228_n20584) );
  OR2X2 OR2X2_4938 ( .A(u2__abc_44228_n20587), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n20588) );
  OR2X2 OR2X2_4939 ( .A(u2__abc_44228_n20592), .B(u2__abc_44228_n20583), .Y(u2__abc_44228_n20593) );
  OR2X2 OR2X2_494 ( .A(_abc_64468_n1672), .B(_abc_64468_n1683), .Y(_abc_64468_n1684) );
  OR2X2 OR2X2_4940 ( .A(u2__abc_44228_n20585), .B(u2_o_234_), .Y(u2__abc_44228_n20596) );
  OR2X2 OR2X2_4941 ( .A(u2__abc_44228_n20599), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n20600) );
  OR2X2 OR2X2_4942 ( .A(u2__abc_44228_n20604), .B(u2__abc_44228_n20595), .Y(u2__abc_44228_n20605) );
  OR2X2 OR2X2_4943 ( .A(u2__abc_44228_n20597), .B(u2_o_235_), .Y(u2__abc_44228_n20608) );
  OR2X2 OR2X2_4944 ( .A(u2__abc_44228_n20611), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n20612) );
  OR2X2 OR2X2_4945 ( .A(u2__abc_44228_n20616), .B(u2__abc_44228_n20607), .Y(u2__abc_44228_n20617) );
  OR2X2 OR2X2_4946 ( .A(u2__abc_44228_n20609), .B(u2_o_236_), .Y(u2__abc_44228_n20620) );
  OR2X2 OR2X2_4947 ( .A(u2__abc_44228_n20623), .B(u2__abc_44228_n2983_bF_buf1), .Y(u2__abc_44228_n20624) );
  OR2X2 OR2X2_4948 ( .A(u2__abc_44228_n20628), .B(u2__abc_44228_n20619), .Y(u2__abc_44228_n20629) );
  OR2X2 OR2X2_4949 ( .A(u2__abc_44228_n20621), .B(u2_o_237_), .Y(u2__abc_44228_n20632) );
  OR2X2 OR2X2_495 ( .A(_abc_64468_n1687), .B(aNan_bF_buf5), .Y(_abc_64468_n1688) );
  OR2X2 OR2X2_4950 ( .A(u2__abc_44228_n20635), .B(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n20636) );
  OR2X2 OR2X2_4951 ( .A(u2__abc_44228_n20640), .B(u2__abc_44228_n20631), .Y(u2__abc_44228_n20641) );
  OR2X2 OR2X2_4952 ( .A(u2__abc_44228_n20633), .B(u2_o_238_), .Y(u2__abc_44228_n20644) );
  OR2X2 OR2X2_4953 ( .A(u2__abc_44228_n20647), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n20648) );
  OR2X2 OR2X2_4954 ( .A(u2__abc_44228_n20652), .B(u2__abc_44228_n20643), .Y(u2__abc_44228_n20653) );
  OR2X2 OR2X2_4955 ( .A(u2__abc_44228_n20645), .B(u2_o_239_), .Y(u2__abc_44228_n20656) );
  OR2X2 OR2X2_4956 ( .A(u2__abc_44228_n20659), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n20660) );
  OR2X2 OR2X2_4957 ( .A(u2__abc_44228_n20664), .B(u2__abc_44228_n20655), .Y(u2__abc_44228_n20665) );
  OR2X2 OR2X2_4958 ( .A(u2__abc_44228_n20657), .B(u2_o_240_), .Y(u2__abc_44228_n20668) );
  OR2X2 OR2X2_4959 ( .A(u2__abc_44228_n20671), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n20672) );
  OR2X2 OR2X2_496 ( .A(_abc_64468_n1679), .B(aNan_bF_buf4), .Y(_abc_64468_n1690) );
  OR2X2 OR2X2_4960 ( .A(u2__abc_44228_n20676), .B(u2__abc_44228_n20667), .Y(u2__abc_44228_n20677) );
  OR2X2 OR2X2_4961 ( .A(u2__abc_44228_n20669), .B(u2_o_241_), .Y(u2__abc_44228_n20680) );
  OR2X2 OR2X2_4962 ( .A(u2__abc_44228_n20683), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n20684) );
  OR2X2 OR2X2_4963 ( .A(u2__abc_44228_n20688), .B(u2__abc_44228_n20679), .Y(u2__abc_44228_n20689) );
  OR2X2 OR2X2_4964 ( .A(u2__abc_44228_n20681), .B(u2_o_242_), .Y(u2__abc_44228_n20692) );
  OR2X2 OR2X2_4965 ( .A(u2__abc_44228_n20695), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n20696) );
  OR2X2 OR2X2_4966 ( .A(u2__abc_44228_n20700), .B(u2__abc_44228_n20691), .Y(u2__abc_44228_n20701) );
  OR2X2 OR2X2_4967 ( .A(u2__abc_44228_n20693), .B(u2_o_243_), .Y(u2__abc_44228_n20704) );
  OR2X2 OR2X2_4968 ( .A(u2__abc_44228_n20707), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n20708) );
  OR2X2 OR2X2_4969 ( .A(u2__abc_44228_n20712), .B(u2__abc_44228_n20703), .Y(u2__abc_44228_n20713) );
  OR2X2 OR2X2_497 ( .A(_abc_64468_n1693), .B(_abc_64468_n1691), .Y(_auto_iopadmap_cc_313_execute_65414_240_) );
  OR2X2 OR2X2_4970 ( .A(u2__abc_44228_n20705), .B(u2_o_244_), .Y(u2__abc_44228_n20716) );
  OR2X2 OR2X2_4971 ( .A(u2__abc_44228_n20719), .B(u2__abc_44228_n2983_bF_buf127), .Y(u2__abc_44228_n20720) );
  OR2X2 OR2X2_4972 ( .A(u2__abc_44228_n20724), .B(u2__abc_44228_n20715), .Y(u2__abc_44228_n20725) );
  OR2X2 OR2X2_4973 ( .A(u2__abc_44228_n20717), .B(u2_o_245_), .Y(u2__abc_44228_n20728) );
  OR2X2 OR2X2_4974 ( .A(u2__abc_44228_n20731), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n20732) );
  OR2X2 OR2X2_4975 ( .A(u2__abc_44228_n20736), .B(u2__abc_44228_n20727), .Y(u2__abc_44228_n20737) );
  OR2X2 OR2X2_4976 ( .A(u2__abc_44228_n20729), .B(u2_o_246_), .Y(u2__abc_44228_n20740) );
  OR2X2 OR2X2_4977 ( .A(u2__abc_44228_n20743), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n20744) );
  OR2X2 OR2X2_4978 ( .A(u2__abc_44228_n20748), .B(u2__abc_44228_n20739), .Y(u2__abc_44228_n20749) );
  OR2X2 OR2X2_4979 ( .A(u2__abc_44228_n20741), .B(u2_o_247_), .Y(u2__abc_44228_n20752) );
  OR2X2 OR2X2_498 ( .A(\a[125] ), .B(\a[126] ), .Y(u1__abc_43968_n137) );
  OR2X2 OR2X2_4980 ( .A(u2__abc_44228_n20755), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n20756) );
  OR2X2 OR2X2_4981 ( .A(u2__abc_44228_n20760), .B(u2__abc_44228_n20751), .Y(u2__abc_44228_n20761) );
  OR2X2 OR2X2_4982 ( .A(u2__abc_44228_n20753), .B(u2_o_248_), .Y(u2__abc_44228_n20764) );
  OR2X2 OR2X2_4983 ( .A(u2__abc_44228_n20767), .B(u2__abc_44228_n2983_bF_buf119), .Y(u2__abc_44228_n20768) );
  OR2X2 OR2X2_4984 ( .A(u2__abc_44228_n20772), .B(u2__abc_44228_n20763), .Y(u2__abc_44228_n20773) );
  OR2X2 OR2X2_4985 ( .A(u2__abc_44228_n20765), .B(u2_o_249_), .Y(u2__abc_44228_n20776) );
  OR2X2 OR2X2_4986 ( .A(u2__abc_44228_n20779), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n20780) );
  OR2X2 OR2X2_4987 ( .A(u2__abc_44228_n20784), .B(u2__abc_44228_n20775), .Y(u2__abc_44228_n20785) );
  OR2X2 OR2X2_4988 ( .A(u2__abc_44228_n20777), .B(u2_o_250_), .Y(u2__abc_44228_n20788) );
  OR2X2 OR2X2_4989 ( .A(u2__abc_44228_n20791), .B(u2__abc_44228_n2983_bF_buf115), .Y(u2__abc_44228_n20792) );
  OR2X2 OR2X2_499 ( .A(\a[123] ), .B(\a[124] ), .Y(u1__abc_43968_n138) );
  OR2X2 OR2X2_4990 ( .A(u2__abc_44228_n20796), .B(u2__abc_44228_n20787), .Y(u2__abc_44228_n20797) );
  OR2X2 OR2X2_4991 ( .A(u2__abc_44228_n20789), .B(u2_o_251_), .Y(u2__abc_44228_n20800) );
  OR2X2 OR2X2_4992 ( .A(u2__abc_44228_n20803), .B(u2__abc_44228_n2983_bF_buf113), .Y(u2__abc_44228_n20804) );
  OR2X2 OR2X2_4993 ( .A(u2__abc_44228_n20808), .B(u2__abc_44228_n20799), .Y(u2__abc_44228_n20809) );
  OR2X2 OR2X2_4994 ( .A(u2__abc_44228_n20801), .B(u2_o_252_), .Y(u2__abc_44228_n20812) );
  OR2X2 OR2X2_4995 ( .A(u2__abc_44228_n20815), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n20816) );
  OR2X2 OR2X2_4996 ( .A(u2__abc_44228_n20820), .B(u2__abc_44228_n20811), .Y(u2__abc_44228_n20821) );
  OR2X2 OR2X2_4997 ( .A(u2__abc_44228_n20813), .B(u2_o_253_), .Y(u2__abc_44228_n20824) );
  OR2X2 OR2X2_4998 ( .A(u2__abc_44228_n20827), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n20828) );
  OR2X2 OR2X2_4999 ( .A(u2__abc_44228_n20832), .B(u2__abc_44228_n20823), .Y(u2__abc_44228_n20833) );
  OR2X2 OR2X2_5 ( .A(aNan_bF_buf7), .B(sqrto_78_), .Y(_abc_64468_n836) );
  OR2X2 OR2X2_50 ( .A(_abc_64468_n753_bF_buf11), .B(\a[24] ), .Y(_abc_64468_n903) );
  OR2X2 OR2X2_500 ( .A(u1__abc_43968_n137), .B(u1__abc_43968_n138), .Y(u1__abc_43968_n139_1) );
  OR2X2 OR2X2_5000 ( .A(u2__abc_44228_n20825), .B(u2_o_254_), .Y(u2__abc_44228_n20836) );
  OR2X2 OR2X2_5001 ( .A(u2__abc_44228_n20839), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n20840) );
  OR2X2 OR2X2_5002 ( .A(u2__abc_44228_n20844), .B(u2__abc_44228_n20835), .Y(u2__abc_44228_n20845) );
  OR2X2 OR2X2_5003 ( .A(u2__abc_44228_n20837), .B(u2_o_255_), .Y(u2__abc_44228_n20848) );
  OR2X2 OR2X2_5004 ( .A(u2__abc_44228_n20851), .B(u2__abc_44228_n2983_bF_buf105), .Y(u2__abc_44228_n20852) );
  OR2X2 OR2X2_5005 ( .A(u2__abc_44228_n20856), .B(u2__abc_44228_n20847), .Y(u2__abc_44228_n20857) );
  OR2X2 OR2X2_5006 ( .A(u2__abc_44228_n20849), .B(u2_o_256_), .Y(u2__abc_44228_n20860) );
  OR2X2 OR2X2_5007 ( .A(u2__abc_44228_n20863), .B(u2__abc_44228_n2983_bF_buf103), .Y(u2__abc_44228_n20864) );
  OR2X2 OR2X2_5008 ( .A(u2__abc_44228_n20868), .B(u2__abc_44228_n20859), .Y(u2__abc_44228_n20869) );
  OR2X2 OR2X2_5009 ( .A(u2__abc_44228_n20861), .B(u2_o_257_), .Y(u2__abc_44228_n20872) );
  OR2X2 OR2X2_501 ( .A(\a[121] ), .B(\a[122] ), .Y(u1__abc_43968_n140_1) );
  OR2X2 OR2X2_5010 ( .A(u2__abc_44228_n20875), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n20876) );
  OR2X2 OR2X2_5011 ( .A(u2__abc_44228_n20880), .B(u2__abc_44228_n20871), .Y(u2__abc_44228_n20881) );
  OR2X2 OR2X2_5012 ( .A(u2__abc_44228_n20873), .B(u2_o_258_), .Y(u2__abc_44228_n20884) );
  OR2X2 OR2X2_5013 ( .A(u2__abc_44228_n20887), .B(u2__abc_44228_n2983_bF_buf99), .Y(u2__abc_44228_n20888) );
  OR2X2 OR2X2_5014 ( .A(u2__abc_44228_n20892), .B(u2__abc_44228_n20883), .Y(u2__abc_44228_n20893) );
  OR2X2 OR2X2_5015 ( .A(u2__abc_44228_n20885), .B(u2_o_259_), .Y(u2__abc_44228_n20896) );
  OR2X2 OR2X2_5016 ( .A(u2__abc_44228_n20899), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n20900) );
  OR2X2 OR2X2_5017 ( .A(u2__abc_44228_n20904), .B(u2__abc_44228_n20895), .Y(u2__abc_44228_n20905) );
  OR2X2 OR2X2_5018 ( .A(u2__abc_44228_n20897), .B(u2_o_260_), .Y(u2__abc_44228_n20908) );
  OR2X2 OR2X2_5019 ( .A(u2__abc_44228_n20911), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n20912) );
  OR2X2 OR2X2_502 ( .A(\a[119] ), .B(\a[120] ), .Y(u1__abc_43968_n141) );
  OR2X2 OR2X2_5020 ( .A(u2__abc_44228_n20916), .B(u2__abc_44228_n20907), .Y(u2__abc_44228_n20917) );
  OR2X2 OR2X2_5021 ( .A(u2__abc_44228_n20909), .B(u2_o_261_), .Y(u2__abc_44228_n20920) );
  OR2X2 OR2X2_5022 ( .A(u2__abc_44228_n20923), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n20924) );
  OR2X2 OR2X2_5023 ( .A(u2__abc_44228_n20928), .B(u2__abc_44228_n20919), .Y(u2__abc_44228_n20929) );
  OR2X2 OR2X2_5024 ( .A(u2__abc_44228_n20921), .B(u2_o_262_), .Y(u2__abc_44228_n20932) );
  OR2X2 OR2X2_5025 ( .A(u2__abc_44228_n20935), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n20936) );
  OR2X2 OR2X2_5026 ( .A(u2__abc_44228_n20940), .B(u2__abc_44228_n20931), .Y(u2__abc_44228_n20941) );
  OR2X2 OR2X2_5027 ( .A(u2__abc_44228_n20933), .B(u2_o_263_), .Y(u2__abc_44228_n20944) );
  OR2X2 OR2X2_5028 ( .A(u2__abc_44228_n20947), .B(u2__abc_44228_n2983_bF_buf89), .Y(u2__abc_44228_n20948) );
  OR2X2 OR2X2_5029 ( .A(u2__abc_44228_n20952), .B(u2__abc_44228_n20943), .Y(u2__abc_44228_n20953) );
  OR2X2 OR2X2_503 ( .A(u1__abc_43968_n140_1), .B(u1__abc_43968_n141), .Y(u1__abc_43968_n142_1) );
  OR2X2 OR2X2_5030 ( .A(u2__abc_44228_n20945), .B(u2_o_264_), .Y(u2__abc_44228_n20956) );
  OR2X2 OR2X2_5031 ( .A(u2__abc_44228_n20959), .B(u2__abc_44228_n2983_bF_buf87), .Y(u2__abc_44228_n20960) );
  OR2X2 OR2X2_5032 ( .A(u2__abc_44228_n20964), .B(u2__abc_44228_n20955), .Y(u2__abc_44228_n20965) );
  OR2X2 OR2X2_5033 ( .A(u2__abc_44228_n20957), .B(u2_o_265_), .Y(u2__abc_44228_n20968) );
  OR2X2 OR2X2_5034 ( .A(u2__abc_44228_n20971), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n20972) );
  OR2X2 OR2X2_5035 ( .A(u2__abc_44228_n20976), .B(u2__abc_44228_n20967), .Y(u2__abc_44228_n20977) );
  OR2X2 OR2X2_5036 ( .A(u2__abc_44228_n20969), .B(u2_o_266_), .Y(u2__abc_44228_n20980) );
  OR2X2 OR2X2_5037 ( .A(u2__abc_44228_n20983), .B(u2__abc_44228_n2983_bF_buf83), .Y(u2__abc_44228_n20984) );
  OR2X2 OR2X2_5038 ( .A(u2__abc_44228_n20988), .B(u2__abc_44228_n20979), .Y(u2__abc_44228_n20989) );
  OR2X2 OR2X2_5039 ( .A(u2__abc_44228_n20981), .B(u2_o_267_), .Y(u2__abc_44228_n20992) );
  OR2X2 OR2X2_504 ( .A(u1__abc_43968_n139_1), .B(u1__abc_43968_n142_1), .Y(u1__abc_43968_n143_1) );
  OR2X2 OR2X2_5040 ( .A(u2__abc_44228_n20995), .B(u2__abc_44228_n2983_bF_buf81), .Y(u2__abc_44228_n20996) );
  OR2X2 OR2X2_5041 ( .A(u2__abc_44228_n21000), .B(u2__abc_44228_n20991), .Y(u2__abc_44228_n21001) );
  OR2X2 OR2X2_5042 ( .A(u2__abc_44228_n20993), .B(u2_o_268_), .Y(u2__abc_44228_n21004) );
  OR2X2 OR2X2_5043 ( .A(u2__abc_44228_n21007), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n21008) );
  OR2X2 OR2X2_5044 ( .A(u2__abc_44228_n21012), .B(u2__abc_44228_n21003), .Y(u2__abc_44228_n21013) );
  OR2X2 OR2X2_5045 ( .A(u2__abc_44228_n21005), .B(u2_o_269_), .Y(u2__abc_44228_n21016) );
  OR2X2 OR2X2_5046 ( .A(u2__abc_44228_n21019), .B(u2__abc_44228_n2983_bF_buf77), .Y(u2__abc_44228_n21020) );
  OR2X2 OR2X2_5047 ( .A(u2__abc_44228_n21024), .B(u2__abc_44228_n21015), .Y(u2__abc_44228_n21025) );
  OR2X2 OR2X2_5048 ( .A(u2__abc_44228_n21017), .B(u2_o_270_), .Y(u2__abc_44228_n21028) );
  OR2X2 OR2X2_5049 ( .A(u2__abc_44228_n21031), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n21032) );
  OR2X2 OR2X2_505 ( .A(\a[118] ), .B(\a[115] ), .Y(u1__abc_43968_n144) );
  OR2X2 OR2X2_5050 ( .A(u2__abc_44228_n21036), .B(u2__abc_44228_n21027), .Y(u2__abc_44228_n21037) );
  OR2X2 OR2X2_5051 ( .A(u2__abc_44228_n21029), .B(u2_o_271_), .Y(u2__abc_44228_n21040) );
  OR2X2 OR2X2_5052 ( .A(u2__abc_44228_n21043), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n21044) );
  OR2X2 OR2X2_5053 ( .A(u2__abc_44228_n21048), .B(u2__abc_44228_n21039), .Y(u2__abc_44228_n21049) );
  OR2X2 OR2X2_5054 ( .A(u2__abc_44228_n21041), .B(u2_o_272_), .Y(u2__abc_44228_n21052) );
  OR2X2 OR2X2_5055 ( .A(u2__abc_44228_n21055), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n21056) );
  OR2X2 OR2X2_5056 ( .A(u2__abc_44228_n21060), .B(u2__abc_44228_n21051), .Y(u2__abc_44228_n21061) );
  OR2X2 OR2X2_5057 ( .A(u2__abc_44228_n21053), .B(u2_o_273_), .Y(u2__abc_44228_n21064) );
  OR2X2 OR2X2_5058 ( .A(u2__abc_44228_n21067), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n21068) );
  OR2X2 OR2X2_5059 ( .A(u2__abc_44228_n21072), .B(u2__abc_44228_n21063), .Y(u2__abc_44228_n21073) );
  OR2X2 OR2X2_506 ( .A(u1__abc_43968_n144), .B(\a[116] ), .Y(u1__abc_43968_n145) );
  OR2X2 OR2X2_5060 ( .A(u2__abc_44228_n21065), .B(u2_o_274_), .Y(u2__abc_44228_n21076) );
  OR2X2 OR2X2_5061 ( .A(u2__abc_44228_n21079), .B(u2__abc_44228_n2983_bF_buf67), .Y(u2__abc_44228_n21080) );
  OR2X2 OR2X2_5062 ( .A(u2__abc_44228_n21084), .B(u2__abc_44228_n21075), .Y(u2__abc_44228_n21085) );
  OR2X2 OR2X2_5063 ( .A(u2__abc_44228_n21077), .B(u2_o_275_), .Y(u2__abc_44228_n21088) );
  OR2X2 OR2X2_5064 ( .A(u2__abc_44228_n21091), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n21092) );
  OR2X2 OR2X2_5065 ( .A(u2__abc_44228_n21096), .B(u2__abc_44228_n21087), .Y(u2__abc_44228_n21097) );
  OR2X2 OR2X2_5066 ( .A(u2__abc_44228_n21089), .B(u2_o_276_), .Y(u2__abc_44228_n21100) );
  OR2X2 OR2X2_5067 ( .A(u2__abc_44228_n21103), .B(u2__abc_44228_n2983_bF_buf63), .Y(u2__abc_44228_n21104) );
  OR2X2 OR2X2_5068 ( .A(u2__abc_44228_n21108), .B(u2__abc_44228_n21099), .Y(u2__abc_44228_n21109) );
  OR2X2 OR2X2_5069 ( .A(u2__abc_44228_n21101), .B(u2_o_277_), .Y(u2__abc_44228_n21112) );
  OR2X2 OR2X2_507 ( .A(\a[113] ), .B(\a[114] ), .Y(u1__abc_43968_n146_1) );
  OR2X2 OR2X2_5070 ( .A(u2__abc_44228_n21115), .B(u2__abc_44228_n2983_bF_buf61), .Y(u2__abc_44228_n21116) );
  OR2X2 OR2X2_5071 ( .A(u2__abc_44228_n21120), .B(u2__abc_44228_n21111), .Y(u2__abc_44228_n21121) );
  OR2X2 OR2X2_5072 ( .A(u2__abc_44228_n21113), .B(u2_o_278_), .Y(u2__abc_44228_n21124) );
  OR2X2 OR2X2_5073 ( .A(u2__abc_44228_n21127), .B(u2__abc_44228_n2983_bF_buf59), .Y(u2__abc_44228_n21128) );
  OR2X2 OR2X2_5074 ( .A(u2__abc_44228_n21132), .B(u2__abc_44228_n21123), .Y(u2__abc_44228_n21133) );
  OR2X2 OR2X2_5075 ( .A(u2__abc_44228_n21125), .B(u2_o_279_), .Y(u2__abc_44228_n21136) );
  OR2X2 OR2X2_5076 ( .A(u2__abc_44228_n21139), .B(u2__abc_44228_n2983_bF_buf57), .Y(u2__abc_44228_n21140) );
  OR2X2 OR2X2_5077 ( .A(u2__abc_44228_n21144), .B(u2__abc_44228_n21135), .Y(u2__abc_44228_n21145) );
  OR2X2 OR2X2_5078 ( .A(u2__abc_44228_n21137), .B(u2_o_280_), .Y(u2__abc_44228_n21148) );
  OR2X2 OR2X2_5079 ( .A(u2__abc_44228_n21151), .B(u2__abc_44228_n2983_bF_buf55), .Y(u2__abc_44228_n21152) );
  OR2X2 OR2X2_508 ( .A(a_112_bF_buf2), .B(\a[117] ), .Y(u1__abc_43968_n147_1) );
  OR2X2 OR2X2_5080 ( .A(u2__abc_44228_n21156), .B(u2__abc_44228_n21147), .Y(u2__abc_44228_n21157) );
  OR2X2 OR2X2_5081 ( .A(u2__abc_44228_n21149), .B(u2_o_281_), .Y(u2__abc_44228_n21160) );
  OR2X2 OR2X2_5082 ( .A(u2__abc_44228_n21163), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n21164) );
  OR2X2 OR2X2_5083 ( .A(u2__abc_44228_n21168), .B(u2__abc_44228_n21159), .Y(u2__abc_44228_n21169) );
  OR2X2 OR2X2_5084 ( .A(u2__abc_44228_n21161), .B(u2_o_282_), .Y(u2__abc_44228_n21172) );
  OR2X2 OR2X2_5085 ( .A(u2__abc_44228_n21175), .B(u2__abc_44228_n2983_bF_buf51), .Y(u2__abc_44228_n21176) );
  OR2X2 OR2X2_5086 ( .A(u2__abc_44228_n21180), .B(u2__abc_44228_n21171), .Y(u2__abc_44228_n21181) );
  OR2X2 OR2X2_5087 ( .A(u2__abc_44228_n21173), .B(u2_o_283_), .Y(u2__abc_44228_n21184) );
  OR2X2 OR2X2_5088 ( .A(u2__abc_44228_n21187), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n21188) );
  OR2X2 OR2X2_5089 ( .A(u2__abc_44228_n21192), .B(u2__abc_44228_n21183), .Y(u2__abc_44228_n21193) );
  OR2X2 OR2X2_509 ( .A(u1__abc_43968_n146_1), .B(u1__abc_43968_n147_1), .Y(u1__abc_43968_n148) );
  OR2X2 OR2X2_5090 ( .A(u2__abc_44228_n21185), .B(u2_o_284_), .Y(u2__abc_44228_n21196) );
  OR2X2 OR2X2_5091 ( .A(u2__abc_44228_n21199), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n21200) );
  OR2X2 OR2X2_5092 ( .A(u2__abc_44228_n21204), .B(u2__abc_44228_n21195), .Y(u2__abc_44228_n21205) );
  OR2X2 OR2X2_5093 ( .A(u2__abc_44228_n21197), .B(u2_o_285_), .Y(u2__abc_44228_n21208) );
  OR2X2 OR2X2_5094 ( .A(u2__abc_44228_n21211), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n21212) );
  OR2X2 OR2X2_5095 ( .A(u2__abc_44228_n21216), .B(u2__abc_44228_n21207), .Y(u2__abc_44228_n21217) );
  OR2X2 OR2X2_5096 ( .A(u2__abc_44228_n21209), .B(u2_o_286_), .Y(u2__abc_44228_n21220) );
  OR2X2 OR2X2_5097 ( .A(u2__abc_44228_n21223), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n21224) );
  OR2X2 OR2X2_5098 ( .A(u2__abc_44228_n21228), .B(u2__abc_44228_n21219), .Y(u2__abc_44228_n21229) );
  OR2X2 OR2X2_5099 ( .A(u2__abc_44228_n21221), .B(u2_o_287_), .Y(u2__abc_44228_n21232) );
  OR2X2 OR2X2_51 ( .A(aNan_bF_buf6), .B(sqrto_101_), .Y(_abc_64468_n905) );
  OR2X2 OR2X2_510 ( .A(u1__abc_43968_n148), .B(u1__abc_43968_n145), .Y(u1__abc_43968_n149_1) );
  OR2X2 OR2X2_5100 ( .A(u2__abc_44228_n21235), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n21236) );
  OR2X2 OR2X2_5101 ( .A(u2__abc_44228_n21240), .B(u2__abc_44228_n21231), .Y(u2__abc_44228_n21241) );
  OR2X2 OR2X2_5102 ( .A(u2__abc_44228_n21233), .B(u2_o_288_), .Y(u2__abc_44228_n21244) );
  OR2X2 OR2X2_5103 ( .A(u2__abc_44228_n21247), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n21248) );
  OR2X2 OR2X2_5104 ( .A(u2__abc_44228_n21252), .B(u2__abc_44228_n21243), .Y(u2__abc_44228_n21253) );
  OR2X2 OR2X2_5105 ( .A(u2__abc_44228_n21245), .B(u2_o_289_), .Y(u2__abc_44228_n21256) );
  OR2X2 OR2X2_5106 ( .A(u2__abc_44228_n21259), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n21260) );
  OR2X2 OR2X2_5107 ( .A(u2__abc_44228_n21264), .B(u2__abc_44228_n21255), .Y(u2__abc_44228_n21265) );
  OR2X2 OR2X2_5108 ( .A(u2__abc_44228_n21257), .B(u2_o_290_), .Y(u2__abc_44228_n21268) );
  OR2X2 OR2X2_5109 ( .A(u2__abc_44228_n21271), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n21272) );
  OR2X2 OR2X2_511 ( .A(u1__abc_43968_n143_1), .B(u1__abc_43968_n149_1), .Y(fracta_112_) );
  OR2X2 OR2X2_5110 ( .A(u2__abc_44228_n21276), .B(u2__abc_44228_n21267), .Y(u2__abc_44228_n21277) );
  OR2X2 OR2X2_5111 ( .A(u2__abc_44228_n21269), .B(u2_o_291_), .Y(u2__abc_44228_n21280) );
  OR2X2 OR2X2_5112 ( .A(u2__abc_44228_n21283), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n21284) );
  OR2X2 OR2X2_5113 ( .A(u2__abc_44228_n21288), .B(u2__abc_44228_n21279), .Y(u2__abc_44228_n21289) );
  OR2X2 OR2X2_5114 ( .A(u2__abc_44228_n21281), .B(u2_o_292_), .Y(u2__abc_44228_n21292) );
  OR2X2 OR2X2_5115 ( .A(u2__abc_44228_n21295), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n21296) );
  OR2X2 OR2X2_5116 ( .A(u2__abc_44228_n21300), .B(u2__abc_44228_n21291), .Y(u2__abc_44228_n21301) );
  OR2X2 OR2X2_5117 ( .A(u2__abc_44228_n21293), .B(u2_o_293_), .Y(u2__abc_44228_n21304) );
  OR2X2 OR2X2_5118 ( .A(u2__abc_44228_n21307), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n21308) );
  OR2X2 OR2X2_5119 ( .A(u2__abc_44228_n21312), .B(u2__abc_44228_n21303), .Y(u2__abc_44228_n21313) );
  OR2X2 OR2X2_512 ( .A(u2__abc_44228_n2963), .B(_auto_iopadmap_cc_313_execute_65412), .Y(u2__abc_44228_n2964) );
  OR2X2 OR2X2_5120 ( .A(u2__abc_44228_n21305), .B(u2_o_294_), .Y(u2__abc_44228_n21316) );
  OR2X2 OR2X2_5121 ( .A(u2__abc_44228_n21319), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n21320) );
  OR2X2 OR2X2_5122 ( .A(u2__abc_44228_n21324), .B(u2__abc_44228_n21315), .Y(u2__abc_44228_n21325) );
  OR2X2 OR2X2_5123 ( .A(u2__abc_44228_n21317), .B(u2_o_295_), .Y(u2__abc_44228_n21328) );
  OR2X2 OR2X2_5124 ( .A(u2__abc_44228_n21331), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n21332) );
  OR2X2 OR2X2_5125 ( .A(u2__abc_44228_n21336), .B(u2__abc_44228_n21327), .Y(u2__abc_44228_n21337) );
  OR2X2 OR2X2_5126 ( .A(u2__abc_44228_n21329), .B(u2_o_296_), .Y(u2__abc_44228_n21340) );
  OR2X2 OR2X2_5127 ( .A(u2__abc_44228_n21343), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n21344) );
  OR2X2 OR2X2_5128 ( .A(u2__abc_44228_n21348), .B(u2__abc_44228_n21339), .Y(u2__abc_44228_n21349) );
  OR2X2 OR2X2_5129 ( .A(u2__abc_44228_n21341), .B(u2_o_297_), .Y(u2__abc_44228_n21352) );
  OR2X2 OR2X2_513 ( .A(u2__abc_44228_n2969), .B(rst), .Y(u2__abc_44228_n2970) );
  OR2X2 OR2X2_5130 ( .A(u2__abc_44228_n21355), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n21356) );
  OR2X2 OR2X2_5131 ( .A(u2__abc_44228_n21360), .B(u2__abc_44228_n21351), .Y(u2__abc_44228_n21361) );
  OR2X2 OR2X2_5132 ( .A(u2__abc_44228_n21353), .B(u2_o_298_), .Y(u2__abc_44228_n21364) );
  OR2X2 OR2X2_5133 ( .A(u2__abc_44228_n21367), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n21368) );
  OR2X2 OR2X2_5134 ( .A(u2__abc_44228_n21372), .B(u2__abc_44228_n21363), .Y(u2__abc_44228_n21373) );
  OR2X2 OR2X2_5135 ( .A(u2__abc_44228_n21365), .B(u2_o_299_), .Y(u2__abc_44228_n21376) );
  OR2X2 OR2X2_5136 ( .A(u2__abc_44228_n21379), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n21380) );
  OR2X2 OR2X2_5137 ( .A(u2__abc_44228_n21384), .B(u2__abc_44228_n21375), .Y(u2__abc_44228_n21385) );
  OR2X2 OR2X2_5138 ( .A(u2__abc_44228_n21377), .B(u2_o_300_), .Y(u2__abc_44228_n21388) );
  OR2X2 OR2X2_5139 ( .A(u2__abc_44228_n21391), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n21392) );
  OR2X2 OR2X2_514 ( .A(u2__abc_44228_n2970), .B(u2__abc_44228_n2965), .Y(u2__abc_29664_n1191) );
  OR2X2 OR2X2_5140 ( .A(u2__abc_44228_n21396), .B(u2__abc_44228_n21387), .Y(u2__abc_44228_n21397) );
  OR2X2 OR2X2_5141 ( .A(u2__abc_44228_n21389), .B(u2_o_301_), .Y(u2__abc_44228_n21400) );
  OR2X2 OR2X2_5142 ( .A(u2__abc_44228_n21403), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n21404) );
  OR2X2 OR2X2_5143 ( .A(u2__abc_44228_n21408), .B(u2__abc_44228_n21399), .Y(u2__abc_44228_n21409) );
  OR2X2 OR2X2_5144 ( .A(u2__abc_44228_n21401), .B(u2_o_302_), .Y(u2__abc_44228_n21412) );
  OR2X2 OR2X2_5145 ( .A(u2__abc_44228_n21415), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n21416) );
  OR2X2 OR2X2_5146 ( .A(u2__abc_44228_n21420), .B(u2__abc_44228_n21411), .Y(u2__abc_44228_n21421) );
  OR2X2 OR2X2_5147 ( .A(u2__abc_44228_n21413), .B(u2_o_303_), .Y(u2__abc_44228_n21424) );
  OR2X2 OR2X2_5148 ( .A(u2__abc_44228_n21427), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n21428) );
  OR2X2 OR2X2_5149 ( .A(u2__abc_44228_n21432), .B(u2__abc_44228_n21423), .Y(u2__abc_44228_n21433) );
  OR2X2 OR2X2_515 ( .A(u2_cnt_3_), .B(u2_cnt_2_), .Y(u2__abc_44228_n2976) );
  OR2X2 OR2X2_5150 ( .A(u2__abc_44228_n21425), .B(u2_o_304_), .Y(u2__abc_44228_n21436) );
  OR2X2 OR2X2_5151 ( .A(u2__abc_44228_n21439), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n21440) );
  OR2X2 OR2X2_5152 ( .A(u2__abc_44228_n21444), .B(u2__abc_44228_n21435), .Y(u2__abc_44228_n21445) );
  OR2X2 OR2X2_5153 ( .A(u2__abc_44228_n21437), .B(u2_o_305_), .Y(u2__abc_44228_n21448) );
  OR2X2 OR2X2_5154 ( .A(u2__abc_44228_n21451), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n21452) );
  OR2X2 OR2X2_5155 ( .A(u2__abc_44228_n21456), .B(u2__abc_44228_n21447), .Y(u2__abc_44228_n21457) );
  OR2X2 OR2X2_5156 ( .A(u2__abc_44228_n21449), .B(u2_o_306_), .Y(u2__abc_44228_n21460) );
  OR2X2 OR2X2_5157 ( .A(u2__abc_44228_n21463), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n21464) );
  OR2X2 OR2X2_5158 ( .A(u2__abc_44228_n21468), .B(u2__abc_44228_n21459), .Y(u2__abc_44228_n21469) );
  OR2X2 OR2X2_5159 ( .A(u2__abc_44228_n21461), .B(u2_o_307_), .Y(u2__abc_44228_n21472) );
  OR2X2 OR2X2_516 ( .A(u2__abc_44228_n2986), .B(u2__abc_44228_n2989_bF_buf3), .Y(u2__abc_44228_n2990) );
  OR2X2 OR2X2_5160 ( .A(u2__abc_44228_n21475), .B(u2__abc_44228_n2983_bF_buf1), .Y(u2__abc_44228_n21476) );
  OR2X2 OR2X2_5161 ( .A(u2__abc_44228_n21480), .B(u2__abc_44228_n21471), .Y(u2__abc_44228_n21481) );
  OR2X2 OR2X2_5162 ( .A(u2__abc_44228_n21473), .B(u2_o_308_), .Y(u2__abc_44228_n21484) );
  OR2X2 OR2X2_5163 ( .A(u2__abc_44228_n21487), .B(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n21488) );
  OR2X2 OR2X2_5164 ( .A(u2__abc_44228_n21492), .B(u2__abc_44228_n21483), .Y(u2__abc_44228_n21493) );
  OR2X2 OR2X2_5165 ( .A(u2__abc_44228_n21485), .B(u2_o_309_), .Y(u2__abc_44228_n21496) );
  OR2X2 OR2X2_5166 ( .A(u2__abc_44228_n21499), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n21500) );
  OR2X2 OR2X2_5167 ( .A(u2__abc_44228_n21504), .B(u2__abc_44228_n21495), .Y(u2__abc_44228_n21505) );
  OR2X2 OR2X2_5168 ( .A(u2__abc_44228_n21497), .B(u2_o_310_), .Y(u2__abc_44228_n21508) );
  OR2X2 OR2X2_5169 ( .A(u2__abc_44228_n21511), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n21512) );
  OR2X2 OR2X2_517 ( .A(u2__abc_44228_n2985), .B(u2__abc_44228_n2990), .Y(u2__abc_29664_n3922) );
  OR2X2 OR2X2_5170 ( .A(u2__abc_44228_n21516), .B(u2__abc_44228_n21507), .Y(u2__abc_44228_n21517) );
  OR2X2 OR2X2_5171 ( .A(u2__abc_44228_n21509), .B(u2_o_311_), .Y(u2__abc_44228_n21520) );
  OR2X2 OR2X2_5172 ( .A(u2__abc_44228_n21523), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n21524) );
  OR2X2 OR2X2_5173 ( .A(u2__abc_44228_n21528), .B(u2__abc_44228_n21519), .Y(u2__abc_44228_n21529) );
  OR2X2 OR2X2_5174 ( .A(u2__abc_44228_n21521), .B(u2_o_312_), .Y(u2__abc_44228_n21532) );
  OR2X2 OR2X2_5175 ( .A(u2__abc_44228_n21535), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n21536) );
  OR2X2 OR2X2_5176 ( .A(u2__abc_44228_n21540), .B(u2__abc_44228_n21531), .Y(u2__abc_44228_n21541) );
  OR2X2 OR2X2_5177 ( .A(u2__abc_44228_n21533), .B(u2_o_313_), .Y(u2__abc_44228_n21544) );
  OR2X2 OR2X2_5178 ( .A(u2__abc_44228_n21547), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n21548) );
  OR2X2 OR2X2_5179 ( .A(u2__abc_44228_n21552), .B(u2__abc_44228_n21543), .Y(u2__abc_44228_n21553) );
  OR2X2 OR2X2_518 ( .A(u2__abc_44228_n2993), .B(u2__abc_44228_n2992), .Y(u2__abc_29664_n3927) );
  OR2X2 OR2X2_5180 ( .A(u2__abc_44228_n21545), .B(u2_o_314_), .Y(u2__abc_44228_n21556) );
  OR2X2 OR2X2_5181 ( .A(u2__abc_44228_n21559), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n21560) );
  OR2X2 OR2X2_5182 ( .A(u2__abc_44228_n21564), .B(u2__abc_44228_n21555), .Y(u2__abc_44228_n21565) );
  OR2X2 OR2X2_5183 ( .A(u2__abc_44228_n21557), .B(u2_o_315_), .Y(u2__abc_44228_n21568) );
  OR2X2 OR2X2_5184 ( .A(u2__abc_44228_n21571), .B(u2__abc_44228_n2983_bF_buf127), .Y(u2__abc_44228_n21572) );
  OR2X2 OR2X2_5185 ( .A(u2__abc_44228_n21576), .B(u2__abc_44228_n21567), .Y(u2__abc_44228_n21577) );
  OR2X2 OR2X2_5186 ( .A(u2__abc_44228_n21569), .B(u2_o_316_), .Y(u2__abc_44228_n21580) );
  OR2X2 OR2X2_5187 ( .A(u2__abc_44228_n21583), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n21584) );
  OR2X2 OR2X2_5188 ( .A(u2__abc_44228_n21588), .B(u2__abc_44228_n21579), .Y(u2__abc_44228_n21589) );
  OR2X2 OR2X2_5189 ( .A(u2__abc_44228_n21581), .B(u2_o_317_), .Y(u2__abc_44228_n21592) );
  OR2X2 OR2X2_519 ( .A(u2__abc_44228_n2997), .B(u2_cnt_0_), .Y(u2__abc_44228_n2998) );
  OR2X2 OR2X2_5190 ( .A(u2__abc_44228_n21595), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n21596) );
  OR2X2 OR2X2_5191 ( .A(u2__abc_44228_n21600), .B(u2__abc_44228_n21591), .Y(u2__abc_44228_n21601) );
  OR2X2 OR2X2_5192 ( .A(u2__abc_44228_n21593), .B(u2_o_318_), .Y(u2__abc_44228_n21604) );
  OR2X2 OR2X2_5193 ( .A(u2__abc_44228_n21607), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n21608) );
  OR2X2 OR2X2_5194 ( .A(u2__abc_44228_n21612), .B(u2__abc_44228_n21603), .Y(u2__abc_44228_n21613) );
  OR2X2 OR2X2_5195 ( .A(u2__abc_44228_n21605), .B(u2_o_319_), .Y(u2__abc_44228_n21616) );
  OR2X2 OR2X2_5196 ( .A(u2__abc_44228_n21619), .B(u2__abc_44228_n2983_bF_buf119), .Y(u2__abc_44228_n21620) );
  OR2X2 OR2X2_5197 ( .A(u2__abc_44228_n21624), .B(u2__abc_44228_n21615), .Y(u2__abc_44228_n21625) );
  OR2X2 OR2X2_5198 ( .A(u2__abc_44228_n21617), .B(u2_o_320_), .Y(u2__abc_44228_n21628) );
  OR2X2 OR2X2_5199 ( .A(u2__abc_44228_n21631), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n21632) );
  OR2X2 OR2X2_52 ( .A(_abc_64468_n753_bF_buf10), .B(\a[25] ), .Y(_abc_64468_n906) );
  OR2X2 OR2X2_520 ( .A(u2__abc_44228_n2968), .B(u2__abc_44228_n2974), .Y(u2__abc_44228_n2999) );
  OR2X2 OR2X2_5200 ( .A(u2__abc_44228_n21636), .B(u2__abc_44228_n21627), .Y(u2__abc_44228_n21637) );
  OR2X2 OR2X2_5201 ( .A(u2__abc_44228_n21629), .B(u2_o_321_), .Y(u2__abc_44228_n21640) );
  OR2X2 OR2X2_5202 ( .A(u2__abc_44228_n21643), .B(u2__abc_44228_n2983_bF_buf115), .Y(u2__abc_44228_n21644) );
  OR2X2 OR2X2_5203 ( .A(u2__abc_44228_n21648), .B(u2__abc_44228_n21639), .Y(u2__abc_44228_n21649) );
  OR2X2 OR2X2_5204 ( .A(u2__abc_44228_n21641), .B(u2_o_322_), .Y(u2__abc_44228_n21652) );
  OR2X2 OR2X2_5205 ( .A(u2__abc_44228_n21655), .B(u2__abc_44228_n2983_bF_buf113), .Y(u2__abc_44228_n21656) );
  OR2X2 OR2X2_5206 ( .A(u2__abc_44228_n21660), .B(u2__abc_44228_n21651), .Y(u2__abc_44228_n21661) );
  OR2X2 OR2X2_5207 ( .A(u2__abc_44228_n21653), .B(u2_o_323_), .Y(u2__abc_44228_n21664) );
  OR2X2 OR2X2_5208 ( .A(u2__abc_44228_n21667), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n21668) );
  OR2X2 OR2X2_5209 ( .A(u2__abc_44228_n21672), .B(u2__abc_44228_n21663), .Y(u2__abc_44228_n21673) );
  OR2X2 OR2X2_521 ( .A(u2_cnt_1_), .B(u2_cnt_0_), .Y(u2__abc_44228_n3002) );
  OR2X2 OR2X2_5210 ( .A(u2__abc_44228_n21665), .B(u2_o_324_), .Y(u2__abc_44228_n21676) );
  OR2X2 OR2X2_5211 ( .A(u2__abc_44228_n21679), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n21680) );
  OR2X2 OR2X2_5212 ( .A(u2__abc_44228_n21684), .B(u2__abc_44228_n21675), .Y(u2__abc_44228_n21685) );
  OR2X2 OR2X2_5213 ( .A(u2__abc_44228_n21677), .B(u2_o_325_), .Y(u2__abc_44228_n21688) );
  OR2X2 OR2X2_5214 ( .A(u2__abc_44228_n21691), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n21692) );
  OR2X2 OR2X2_5215 ( .A(u2__abc_44228_n21696), .B(u2__abc_44228_n21687), .Y(u2__abc_44228_n21697) );
  OR2X2 OR2X2_5216 ( .A(u2__abc_44228_n21689), .B(u2_o_326_), .Y(u2__abc_44228_n21700) );
  OR2X2 OR2X2_5217 ( .A(u2__abc_44228_n21703), .B(u2__abc_44228_n2983_bF_buf105), .Y(u2__abc_44228_n21704) );
  OR2X2 OR2X2_5218 ( .A(u2__abc_44228_n21708), .B(u2__abc_44228_n21699), .Y(u2__abc_44228_n21709) );
  OR2X2 OR2X2_5219 ( .A(u2__abc_44228_n21701), .B(u2_o_327_), .Y(u2__abc_44228_n21712) );
  OR2X2 OR2X2_522 ( .A(u2__abc_44228_n3006), .B(u2__abc_44228_n3001), .Y(u2_cnt_1__FF_INPUT) );
  OR2X2 OR2X2_5220 ( .A(u2__abc_44228_n21715), .B(u2__abc_44228_n2983_bF_buf103), .Y(u2__abc_44228_n21716) );
  OR2X2 OR2X2_5221 ( .A(u2__abc_44228_n21720), .B(u2__abc_44228_n21711), .Y(u2__abc_44228_n21721) );
  OR2X2 OR2X2_5222 ( .A(u2__abc_44228_n21713), .B(u2_o_328_), .Y(u2__abc_44228_n21724) );
  OR2X2 OR2X2_5223 ( .A(u2__abc_44228_n21727), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n21728) );
  OR2X2 OR2X2_5224 ( .A(u2__abc_44228_n21732), .B(u2__abc_44228_n21723), .Y(u2__abc_44228_n21733) );
  OR2X2 OR2X2_5225 ( .A(u2__abc_44228_n21725), .B(u2_o_329_), .Y(u2__abc_44228_n21736) );
  OR2X2 OR2X2_5226 ( .A(u2__abc_44228_n21739), .B(u2__abc_44228_n2983_bF_buf99), .Y(u2__abc_44228_n21740) );
  OR2X2 OR2X2_5227 ( .A(u2__abc_44228_n21744), .B(u2__abc_44228_n21735), .Y(u2__abc_44228_n21745) );
  OR2X2 OR2X2_5228 ( .A(u2__abc_44228_n21737), .B(u2_o_330_), .Y(u2__abc_44228_n21748) );
  OR2X2 OR2X2_5229 ( .A(u2__abc_44228_n21751), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n21752) );
  OR2X2 OR2X2_523 ( .A(u2__abc_44228_n3008), .B(u2_cnt_2_), .Y(u2__abc_44228_n3009) );
  OR2X2 OR2X2_5230 ( .A(u2__abc_44228_n21756), .B(u2__abc_44228_n21747), .Y(u2__abc_44228_n21757) );
  OR2X2 OR2X2_5231 ( .A(u2__abc_44228_n21749), .B(u2_o_331_), .Y(u2__abc_44228_n21760) );
  OR2X2 OR2X2_5232 ( .A(u2__abc_44228_n21763), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n21764) );
  OR2X2 OR2X2_5233 ( .A(u2__abc_44228_n21768), .B(u2__abc_44228_n21759), .Y(u2__abc_44228_n21769) );
  OR2X2 OR2X2_5234 ( .A(u2__abc_44228_n21761), .B(u2_o_332_), .Y(u2__abc_44228_n21772) );
  OR2X2 OR2X2_5235 ( .A(u2__abc_44228_n21775), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n21776) );
  OR2X2 OR2X2_5236 ( .A(u2__abc_44228_n21780), .B(u2__abc_44228_n21771), .Y(u2__abc_44228_n21781) );
  OR2X2 OR2X2_5237 ( .A(u2__abc_44228_n21773), .B(u2_o_333_), .Y(u2__abc_44228_n21784) );
  OR2X2 OR2X2_5238 ( .A(u2__abc_44228_n21787), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n21788) );
  OR2X2 OR2X2_5239 ( .A(u2__abc_44228_n21792), .B(u2__abc_44228_n21783), .Y(u2__abc_44228_n21793) );
  OR2X2 OR2X2_524 ( .A(u2__abc_44228_n3003), .B(u2_cnt_2_), .Y(u2__abc_44228_n3013) );
  OR2X2 OR2X2_5240 ( .A(u2__abc_44228_n21785), .B(u2_o_334_), .Y(u2__abc_44228_n21796) );
  OR2X2 OR2X2_5241 ( .A(u2__abc_44228_n21799), .B(u2__abc_44228_n2983_bF_buf89), .Y(u2__abc_44228_n21800) );
  OR2X2 OR2X2_5242 ( .A(u2__abc_44228_n21804), .B(u2__abc_44228_n21795), .Y(u2__abc_44228_n21805) );
  OR2X2 OR2X2_5243 ( .A(u2__abc_44228_n21797), .B(u2_o_335_), .Y(u2__abc_44228_n21808) );
  OR2X2 OR2X2_5244 ( .A(u2__abc_44228_n21811), .B(u2__abc_44228_n2983_bF_buf87), .Y(u2__abc_44228_n21812) );
  OR2X2 OR2X2_5245 ( .A(u2__abc_44228_n21816), .B(u2__abc_44228_n21807), .Y(u2__abc_44228_n21817) );
  OR2X2 OR2X2_5246 ( .A(u2__abc_44228_n21809), .B(u2_o_336_), .Y(u2__abc_44228_n21820) );
  OR2X2 OR2X2_5247 ( .A(u2__abc_44228_n21823), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n21824) );
  OR2X2 OR2X2_5248 ( .A(u2__abc_44228_n21828), .B(u2__abc_44228_n21819), .Y(u2__abc_44228_n21829) );
  OR2X2 OR2X2_5249 ( .A(u2__abc_44228_n21821), .B(u2_o_337_), .Y(u2__abc_44228_n21832) );
  OR2X2 OR2X2_525 ( .A(u2__abc_44228_n3015), .B(u2__abc_44228_n3010), .Y(u2__abc_44228_n3016) );
  OR2X2 OR2X2_5250 ( .A(u2__abc_44228_n21835), .B(u2__abc_44228_n2983_bF_buf83), .Y(u2__abc_44228_n21836) );
  OR2X2 OR2X2_5251 ( .A(u2__abc_44228_n21840), .B(u2__abc_44228_n21831), .Y(u2__abc_44228_n21841) );
  OR2X2 OR2X2_5252 ( .A(u2__abc_44228_n21833), .B(u2_o_338_), .Y(u2__abc_44228_n21844) );
  OR2X2 OR2X2_5253 ( .A(u2__abc_44228_n21847), .B(u2__abc_44228_n2983_bF_buf81), .Y(u2__abc_44228_n21848) );
  OR2X2 OR2X2_5254 ( .A(u2__abc_44228_n21852), .B(u2__abc_44228_n21843), .Y(u2__abc_44228_n21853) );
  OR2X2 OR2X2_5255 ( .A(u2__abc_44228_n21845), .B(u2_o_339_), .Y(u2__abc_44228_n21856) );
  OR2X2 OR2X2_5256 ( .A(u2__abc_44228_n21859), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n21860) );
  OR2X2 OR2X2_5257 ( .A(u2__abc_44228_n21864), .B(u2__abc_44228_n21855), .Y(u2__abc_44228_n21865) );
  OR2X2 OR2X2_5258 ( .A(u2__abc_44228_n21857), .B(u2_o_340_), .Y(u2__abc_44228_n21868) );
  OR2X2 OR2X2_5259 ( .A(u2__abc_44228_n21871), .B(u2__abc_44228_n2983_bF_buf77), .Y(u2__abc_44228_n21872) );
  OR2X2 OR2X2_526 ( .A(u2__abc_44228_n3011), .B(u2_cnt_3_), .Y(u2__abc_44228_n3019) );
  OR2X2 OR2X2_5260 ( .A(u2__abc_44228_n21876), .B(u2__abc_44228_n21867), .Y(u2__abc_44228_n21877) );
  OR2X2 OR2X2_5261 ( .A(u2__abc_44228_n21869), .B(u2_o_341_), .Y(u2__abc_44228_n21880) );
  OR2X2 OR2X2_5262 ( .A(u2__abc_44228_n21883), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n21884) );
  OR2X2 OR2X2_5263 ( .A(u2__abc_44228_n21888), .B(u2__abc_44228_n21879), .Y(u2__abc_44228_n21889) );
  OR2X2 OR2X2_5264 ( .A(u2__abc_44228_n21881), .B(u2_o_342_), .Y(u2__abc_44228_n21892) );
  OR2X2 OR2X2_5265 ( .A(u2__abc_44228_n21895), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n21896) );
  OR2X2 OR2X2_5266 ( .A(u2__abc_44228_n21900), .B(u2__abc_44228_n21891), .Y(u2__abc_44228_n21901) );
  OR2X2 OR2X2_5267 ( .A(u2__abc_44228_n21893), .B(u2_o_343_), .Y(u2__abc_44228_n21904) );
  OR2X2 OR2X2_5268 ( .A(u2__abc_44228_n21907), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n21908) );
  OR2X2 OR2X2_5269 ( .A(u2__abc_44228_n21912), .B(u2__abc_44228_n21903), .Y(u2__abc_44228_n21913) );
  OR2X2 OR2X2_527 ( .A(u2__abc_44228_n3023), .B(u2__abc_44228_n3018), .Y(u2_cnt_3__FF_INPUT) );
  OR2X2 OR2X2_5270 ( .A(u2__abc_44228_n21905), .B(u2_o_344_), .Y(u2__abc_44228_n21916) );
  OR2X2 OR2X2_5271 ( .A(u2__abc_44228_n21919), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n21920) );
  OR2X2 OR2X2_5272 ( .A(u2__abc_44228_n21924), .B(u2__abc_44228_n21915), .Y(u2__abc_44228_n21925) );
  OR2X2 OR2X2_5273 ( .A(u2__abc_44228_n21917), .B(u2_o_345_), .Y(u2__abc_44228_n21928) );
  OR2X2 OR2X2_5274 ( .A(u2__abc_44228_n21931), .B(u2__abc_44228_n2983_bF_buf67), .Y(u2__abc_44228_n21932) );
  OR2X2 OR2X2_5275 ( .A(u2__abc_44228_n21936), .B(u2__abc_44228_n21927), .Y(u2__abc_44228_n21937) );
  OR2X2 OR2X2_5276 ( .A(u2__abc_44228_n21929), .B(u2_o_346_), .Y(u2__abc_44228_n21940) );
  OR2X2 OR2X2_5277 ( .A(u2__abc_44228_n21943), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n21944) );
  OR2X2 OR2X2_5278 ( .A(u2__abc_44228_n21948), .B(u2__abc_44228_n21939), .Y(u2__abc_44228_n21949) );
  OR2X2 OR2X2_5279 ( .A(u2__abc_44228_n21941), .B(u2_o_347_), .Y(u2__abc_44228_n21952) );
  OR2X2 OR2X2_528 ( .A(u2__abc_44228_n3020), .B(u2_cnt_4_), .Y(u2__abc_44228_n3028) );
  OR2X2 OR2X2_5280 ( .A(u2__abc_44228_n21955), .B(u2__abc_44228_n2983_bF_buf63), .Y(u2__abc_44228_n21956) );
  OR2X2 OR2X2_5281 ( .A(u2__abc_44228_n21960), .B(u2__abc_44228_n21951), .Y(u2__abc_44228_n21961) );
  OR2X2 OR2X2_5282 ( .A(u2__abc_44228_n21953), .B(u2_o_348_), .Y(u2__abc_44228_n21964) );
  OR2X2 OR2X2_5283 ( .A(u2__abc_44228_n21967), .B(u2__abc_44228_n2983_bF_buf61), .Y(u2__abc_44228_n21968) );
  OR2X2 OR2X2_5284 ( .A(u2__abc_44228_n21972), .B(u2__abc_44228_n21963), .Y(u2__abc_44228_n21973) );
  OR2X2 OR2X2_5285 ( .A(u2__abc_44228_n21965), .B(u2_o_349_), .Y(u2__abc_44228_n21976) );
  OR2X2 OR2X2_5286 ( .A(u2__abc_44228_n21979), .B(u2__abc_44228_n2983_bF_buf59), .Y(u2__abc_44228_n21980) );
  OR2X2 OR2X2_5287 ( .A(u2__abc_44228_n21984), .B(u2__abc_44228_n21975), .Y(u2__abc_44228_n21985) );
  OR2X2 OR2X2_5288 ( .A(u2__abc_44228_n21977), .B(u2_o_350_), .Y(u2__abc_44228_n21988) );
  OR2X2 OR2X2_5289 ( .A(u2__abc_44228_n21991), .B(u2__abc_44228_n2983_bF_buf57), .Y(u2__abc_44228_n21992) );
  OR2X2 OR2X2_529 ( .A(u2__abc_44228_n3030), .B(u2__abc_44228_n3025), .Y(u2_cnt_4__FF_INPUT) );
  OR2X2 OR2X2_5290 ( .A(u2__abc_44228_n21996), .B(u2__abc_44228_n21987), .Y(u2__abc_44228_n21997) );
  OR2X2 OR2X2_5291 ( .A(u2__abc_44228_n21989), .B(u2_o_351_), .Y(u2__abc_44228_n22000) );
  OR2X2 OR2X2_5292 ( .A(u2__abc_44228_n22003), .B(u2__abc_44228_n2983_bF_buf55), .Y(u2__abc_44228_n22004) );
  OR2X2 OR2X2_5293 ( .A(u2__abc_44228_n22008), .B(u2__abc_44228_n21999), .Y(u2__abc_44228_n22009) );
  OR2X2 OR2X2_5294 ( .A(u2__abc_44228_n22001), .B(u2_o_352_), .Y(u2__abc_44228_n22012) );
  OR2X2 OR2X2_5295 ( .A(u2__abc_44228_n22015), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n22016) );
  OR2X2 OR2X2_5296 ( .A(u2__abc_44228_n22020), .B(u2__abc_44228_n22011), .Y(u2__abc_44228_n22021) );
  OR2X2 OR2X2_5297 ( .A(u2__abc_44228_n22013), .B(u2_o_353_), .Y(u2__abc_44228_n22024) );
  OR2X2 OR2X2_5298 ( .A(u2__abc_44228_n22027), .B(u2__abc_44228_n2983_bF_buf51), .Y(u2__abc_44228_n22028) );
  OR2X2 OR2X2_5299 ( .A(u2__abc_44228_n22032), .B(u2__abc_44228_n22023), .Y(u2__abc_44228_n22033) );
  OR2X2 OR2X2_53 ( .A(aNan_bF_buf5), .B(sqrto_102_), .Y(_abc_64468_n908) );
  OR2X2 OR2X2_530 ( .A(u2__abc_44228_n3026), .B(u2_cnt_5_), .Y(u2__abc_44228_n3033) );
  OR2X2 OR2X2_5300 ( .A(u2__abc_44228_n22025), .B(u2_o_354_), .Y(u2__abc_44228_n22036) );
  OR2X2 OR2X2_5301 ( .A(u2__abc_44228_n22039), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n22040) );
  OR2X2 OR2X2_5302 ( .A(u2__abc_44228_n22044), .B(u2__abc_44228_n22035), .Y(u2__abc_44228_n22045) );
  OR2X2 OR2X2_5303 ( .A(u2__abc_44228_n22037), .B(u2_o_355_), .Y(u2__abc_44228_n22048) );
  OR2X2 OR2X2_5304 ( .A(u2__abc_44228_n22051), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n22052) );
  OR2X2 OR2X2_5305 ( .A(u2__abc_44228_n22056), .B(u2__abc_44228_n22047), .Y(u2__abc_44228_n22057) );
  OR2X2 OR2X2_5306 ( .A(u2__abc_44228_n22049), .B(u2_o_356_), .Y(u2__abc_44228_n22060) );
  OR2X2 OR2X2_5307 ( .A(u2__abc_44228_n22063), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n22064) );
  OR2X2 OR2X2_5308 ( .A(u2__abc_44228_n22068), .B(u2__abc_44228_n22059), .Y(u2__abc_44228_n22069) );
  OR2X2 OR2X2_5309 ( .A(u2__abc_44228_n22061), .B(u2_o_357_), .Y(u2__abc_44228_n22072) );
  OR2X2 OR2X2_531 ( .A(u2__abc_44228_n3037), .B(u2__abc_44228_n3032), .Y(u2_cnt_5__FF_INPUT) );
  OR2X2 OR2X2_5310 ( .A(u2__abc_44228_n22075), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n22076) );
  OR2X2 OR2X2_5311 ( .A(u2__abc_44228_n22080), .B(u2__abc_44228_n22071), .Y(u2__abc_44228_n22081) );
  OR2X2 OR2X2_5312 ( .A(u2__abc_44228_n22073), .B(u2_o_358_), .Y(u2__abc_44228_n22084) );
  OR2X2 OR2X2_5313 ( .A(u2__abc_44228_n22087), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n22088) );
  OR2X2 OR2X2_5314 ( .A(u2__abc_44228_n22092), .B(u2__abc_44228_n22083), .Y(u2__abc_44228_n22093) );
  OR2X2 OR2X2_5315 ( .A(u2__abc_44228_n22085), .B(u2_o_359_), .Y(u2__abc_44228_n22096) );
  OR2X2 OR2X2_5316 ( .A(u2__abc_44228_n22099), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n22100) );
  OR2X2 OR2X2_5317 ( .A(u2__abc_44228_n22104), .B(u2__abc_44228_n22095), .Y(u2__abc_44228_n22105) );
  OR2X2 OR2X2_5318 ( .A(u2__abc_44228_n22097), .B(u2_o_360_), .Y(u2__abc_44228_n22108) );
  OR2X2 OR2X2_5319 ( .A(u2__abc_44228_n22111), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n22112) );
  OR2X2 OR2X2_532 ( .A(u2__abc_44228_n3034), .B(u2__abc_44228_n3010), .Y(u2__abc_44228_n3039) );
  OR2X2 OR2X2_5320 ( .A(u2__abc_44228_n22116), .B(u2__abc_44228_n22107), .Y(u2__abc_44228_n22117) );
  OR2X2 OR2X2_5321 ( .A(u2__abc_44228_n22109), .B(u2_o_361_), .Y(u2__abc_44228_n22120) );
  OR2X2 OR2X2_5322 ( .A(u2__abc_44228_n22123), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n22124) );
  OR2X2 OR2X2_5323 ( .A(u2__abc_44228_n22128), .B(u2__abc_44228_n22119), .Y(u2__abc_44228_n22129) );
  OR2X2 OR2X2_5324 ( .A(u2__abc_44228_n22121), .B(u2_o_362_), .Y(u2__abc_44228_n22132) );
  OR2X2 OR2X2_5325 ( .A(u2__abc_44228_n22135), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n22136) );
  OR2X2 OR2X2_5326 ( .A(u2__abc_44228_n22140), .B(u2__abc_44228_n22131), .Y(u2__abc_44228_n22141) );
  OR2X2 OR2X2_5327 ( .A(u2__abc_44228_n22133), .B(u2_o_363_), .Y(u2__abc_44228_n22144) );
  OR2X2 OR2X2_5328 ( .A(u2__abc_44228_n22147), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n22148) );
  OR2X2 OR2X2_5329 ( .A(u2__abc_44228_n22152), .B(u2__abc_44228_n22143), .Y(u2__abc_44228_n22153) );
  OR2X2 OR2X2_533 ( .A(u2__abc_44228_n3040), .B(u2_cnt_6_), .Y(u2__abc_44228_n3041) );
  OR2X2 OR2X2_5330 ( .A(u2__abc_44228_n22145), .B(u2_o_364_), .Y(u2__abc_44228_n22156) );
  OR2X2 OR2X2_5331 ( .A(u2__abc_44228_n22159), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n22160) );
  OR2X2 OR2X2_5332 ( .A(u2__abc_44228_n22164), .B(u2__abc_44228_n22155), .Y(u2__abc_44228_n22165) );
  OR2X2 OR2X2_5333 ( .A(u2__abc_44228_n22157), .B(u2_o_365_), .Y(u2__abc_44228_n22168) );
  OR2X2 OR2X2_5334 ( .A(u2__abc_44228_n22171), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n22172) );
  OR2X2 OR2X2_5335 ( .A(u2__abc_44228_n22176), .B(u2__abc_44228_n22167), .Y(u2__abc_44228_n22177) );
  OR2X2 OR2X2_5336 ( .A(u2__abc_44228_n22169), .B(u2_o_366_), .Y(u2__abc_44228_n22180) );
  OR2X2 OR2X2_5337 ( .A(u2__abc_44228_n22183), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n22184) );
  OR2X2 OR2X2_5338 ( .A(u2__abc_44228_n22188), .B(u2__abc_44228_n22179), .Y(u2__abc_44228_n22189) );
  OR2X2 OR2X2_5339 ( .A(u2__abc_44228_n22181), .B(u2_o_367_), .Y(u2__abc_44228_n22192) );
  OR2X2 OR2X2_534 ( .A(u2__abc_44228_n3044), .B(u2__abc_44228_n3010), .Y(u2__abc_44228_n3045) );
  OR2X2 OR2X2_5340 ( .A(u2__abc_44228_n22195), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n22196) );
  OR2X2 OR2X2_5341 ( .A(u2__abc_44228_n22200), .B(u2__abc_44228_n22191), .Y(u2__abc_44228_n22201) );
  OR2X2 OR2X2_5342 ( .A(u2__abc_44228_n22193), .B(u2_o_368_), .Y(u2__abc_44228_n22204) );
  OR2X2 OR2X2_5343 ( .A(u2__abc_44228_n22207), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n22208) );
  OR2X2 OR2X2_5344 ( .A(u2__abc_44228_n22212), .B(u2__abc_44228_n22203), .Y(u2__abc_44228_n22213) );
  OR2X2 OR2X2_5345 ( .A(u2__abc_44228_n22205), .B(u2_o_369_), .Y(u2__abc_44228_n22216) );
  OR2X2 OR2X2_5346 ( .A(u2__abc_44228_n22219), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n22220) );
  OR2X2 OR2X2_5347 ( .A(u2__abc_44228_n22224), .B(u2__abc_44228_n22215), .Y(u2__abc_44228_n22225) );
  OR2X2 OR2X2_5348 ( .A(u2__abc_44228_n22217), .B(u2_o_370_), .Y(u2__abc_44228_n22228) );
  OR2X2 OR2X2_5349 ( .A(u2__abc_44228_n22231), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n22232) );
  OR2X2 OR2X2_535 ( .A(u2__abc_44228_n3054), .B(rst), .Y(u2__abc_44228_n3055) );
  OR2X2 OR2X2_5350 ( .A(u2__abc_44228_n22236), .B(u2__abc_44228_n22227), .Y(u2__abc_44228_n22237) );
  OR2X2 OR2X2_5351 ( .A(u2__abc_44228_n22229), .B(u2_o_371_), .Y(u2__abc_44228_n22240) );
  OR2X2 OR2X2_5352 ( .A(u2__abc_44228_n22243), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n22244) );
  OR2X2 OR2X2_5353 ( .A(u2__abc_44228_n22248), .B(u2__abc_44228_n22239), .Y(u2__abc_44228_n22249) );
  OR2X2 OR2X2_5354 ( .A(u2__abc_44228_n22241), .B(u2_o_372_), .Y(u2__abc_44228_n22252) );
  OR2X2 OR2X2_5355 ( .A(u2__abc_44228_n22255), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n22256) );
  OR2X2 OR2X2_5356 ( .A(u2__abc_44228_n22260), .B(u2__abc_44228_n22251), .Y(u2__abc_44228_n22261) );
  OR2X2 OR2X2_5357 ( .A(u2__abc_44228_n22253), .B(u2_o_373_), .Y(u2__abc_44228_n22264) );
  OR2X2 OR2X2_5358 ( .A(u2__abc_44228_n22267), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n22268) );
  OR2X2 OR2X2_5359 ( .A(u2__abc_44228_n22272), .B(u2__abc_44228_n22263), .Y(u2__abc_44228_n22273) );
  OR2X2 OR2X2_536 ( .A(u2__abc_44228_n3055), .B(u2__abc_44228_n3052), .Y(u2__abc_44228_n3056) );
  OR2X2 OR2X2_5360 ( .A(u2__abc_44228_n22265), .B(u2_o_374_), .Y(u2__abc_44228_n22276) );
  OR2X2 OR2X2_5361 ( .A(u2__abc_44228_n22279), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n22280) );
  OR2X2 OR2X2_5362 ( .A(u2__abc_44228_n22284), .B(u2__abc_44228_n22275), .Y(u2__abc_44228_n22285) );
  OR2X2 OR2X2_5363 ( .A(u2__abc_44228_n22277), .B(u2_o_375_), .Y(u2__abc_44228_n22288) );
  OR2X2 OR2X2_5364 ( .A(u2__abc_44228_n22291), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n22292) );
  OR2X2 OR2X2_5365 ( .A(u2__abc_44228_n22296), .B(u2__abc_44228_n22287), .Y(u2__abc_44228_n22297) );
  OR2X2 OR2X2_5366 ( .A(u2__abc_44228_n22289), .B(u2_o_376_), .Y(u2__abc_44228_n22300) );
  OR2X2 OR2X2_5367 ( .A(u2__abc_44228_n22303), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n22304) );
  OR2X2 OR2X2_5368 ( .A(u2__abc_44228_n22308), .B(u2__abc_44228_n22299), .Y(u2__abc_44228_n22309) );
  OR2X2 OR2X2_5369 ( .A(u2__abc_44228_n22301), .B(u2_o_377_), .Y(u2__abc_44228_n22312) );
  OR2X2 OR2X2_537 ( .A(u2__abc_44228_n3061), .B(u2__abc_44228_n2963), .Y(u2__abc_44228_n3062) );
  OR2X2 OR2X2_5370 ( .A(u2__abc_44228_n22315), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n22316) );
  OR2X2 OR2X2_5371 ( .A(u2__abc_44228_n22320), .B(u2__abc_44228_n22311), .Y(u2__abc_44228_n22321) );
  OR2X2 OR2X2_5372 ( .A(u2__abc_44228_n22313), .B(u2_o_378_), .Y(u2__abc_44228_n22324) );
  OR2X2 OR2X2_5373 ( .A(u2__abc_44228_n22327), .B(u2__abc_44228_n2983_bF_buf1), .Y(u2__abc_44228_n22328) );
  OR2X2 OR2X2_5374 ( .A(u2__abc_44228_n22332), .B(u2__abc_44228_n22323), .Y(u2__abc_44228_n22333) );
  OR2X2 OR2X2_5375 ( .A(u2__abc_44228_n22325), .B(u2_o_379_), .Y(u2__abc_44228_n22336) );
  OR2X2 OR2X2_5376 ( .A(u2__abc_44228_n22339), .B(u2__abc_44228_n2983_bF_buf141), .Y(u2__abc_44228_n22340) );
  OR2X2 OR2X2_5377 ( .A(u2__abc_44228_n22344), .B(u2__abc_44228_n22335), .Y(u2__abc_44228_n22345) );
  OR2X2 OR2X2_5378 ( .A(u2__abc_44228_n22337), .B(u2_o_380_), .Y(u2__abc_44228_n22348) );
  OR2X2 OR2X2_5379 ( .A(u2__abc_44228_n22351), .B(u2__abc_44228_n2983_bF_buf139), .Y(u2__abc_44228_n22352) );
  OR2X2 OR2X2_538 ( .A(u2__abc_44228_n3064), .B(u2_root_0_), .Y(u2__abc_44228_n3065) );
  OR2X2 OR2X2_5380 ( .A(u2__abc_44228_n22356), .B(u2__abc_44228_n22347), .Y(u2__abc_44228_n22357) );
  OR2X2 OR2X2_5381 ( .A(u2__abc_44228_n22349), .B(u2_o_381_), .Y(u2__abc_44228_n22360) );
  OR2X2 OR2X2_5382 ( .A(u2__abc_44228_n22363), .B(u2__abc_44228_n2983_bF_buf137), .Y(u2__abc_44228_n22364) );
  OR2X2 OR2X2_5383 ( .A(u2__abc_44228_n22368), .B(u2__abc_44228_n22359), .Y(u2__abc_44228_n22369) );
  OR2X2 OR2X2_5384 ( .A(u2__abc_44228_n22361), .B(u2_o_382_), .Y(u2__abc_44228_n22372) );
  OR2X2 OR2X2_5385 ( .A(u2__abc_44228_n22375), .B(u2__abc_44228_n2983_bF_buf135), .Y(u2__abc_44228_n22376) );
  OR2X2 OR2X2_5386 ( .A(u2__abc_44228_n22380), .B(u2__abc_44228_n22371), .Y(u2__abc_44228_n22381) );
  OR2X2 OR2X2_5387 ( .A(u2__abc_44228_n22373), .B(u2_o_383_), .Y(u2__abc_44228_n22384) );
  OR2X2 OR2X2_5388 ( .A(u2__abc_44228_n22387), .B(u2__abc_44228_n2983_bF_buf133), .Y(u2__abc_44228_n22388) );
  OR2X2 OR2X2_5389 ( .A(u2__abc_44228_n22392), .B(u2__abc_44228_n22383), .Y(u2__abc_44228_n22393) );
  OR2X2 OR2X2_539 ( .A(u2__abc_44228_n3067), .B(u2_remHiShift_1_), .Y(u2__abc_44228_n3068) );
  OR2X2 OR2X2_5390 ( .A(u2__abc_44228_n22385), .B(u2_o_384_), .Y(u2__abc_44228_n22396) );
  OR2X2 OR2X2_5391 ( .A(u2__abc_44228_n22399), .B(u2__abc_44228_n2983_bF_buf131), .Y(u2__abc_44228_n22400) );
  OR2X2 OR2X2_5392 ( .A(u2__abc_44228_n22404), .B(u2__abc_44228_n22395), .Y(u2__abc_44228_n22405) );
  OR2X2 OR2X2_5393 ( .A(u2__abc_44228_n22397), .B(u2_o_385_), .Y(u2__abc_44228_n22408) );
  OR2X2 OR2X2_5394 ( .A(u2__abc_44228_n22411), .B(u2__abc_44228_n2983_bF_buf129), .Y(u2__abc_44228_n22412) );
  OR2X2 OR2X2_5395 ( .A(u2__abc_44228_n22416), .B(u2__abc_44228_n22407), .Y(u2__abc_44228_n22417) );
  OR2X2 OR2X2_5396 ( .A(u2__abc_44228_n22409), .B(u2_o_386_), .Y(u2__abc_44228_n22420) );
  OR2X2 OR2X2_5397 ( .A(u2__abc_44228_n22423), .B(u2__abc_44228_n2983_bF_buf127), .Y(u2__abc_44228_n22424) );
  OR2X2 OR2X2_5398 ( .A(u2__abc_44228_n22428), .B(u2__abc_44228_n22419), .Y(u2__abc_44228_n22429) );
  OR2X2 OR2X2_5399 ( .A(u2__abc_44228_n22421), .B(u2_o_387_), .Y(u2__abc_44228_n22432) );
  OR2X2 OR2X2_54 ( .A(_abc_64468_n753_bF_buf9), .B(\a[26] ), .Y(_abc_64468_n909) );
  OR2X2 OR2X2_540 ( .A(u2__abc_44228_n3070), .B(u2__abc_44228_n3066), .Y(u2__abc_44228_n3071) );
  OR2X2 OR2X2_5400 ( .A(u2__abc_44228_n22435), .B(u2__abc_44228_n2983_bF_buf125), .Y(u2__abc_44228_n22436) );
  OR2X2 OR2X2_5401 ( .A(u2__abc_44228_n22440), .B(u2__abc_44228_n22431), .Y(u2__abc_44228_n22441) );
  OR2X2 OR2X2_5402 ( .A(u2__abc_44228_n22433), .B(u2_o_388_), .Y(u2__abc_44228_n22444) );
  OR2X2 OR2X2_5403 ( .A(u2__abc_44228_n22447), .B(u2__abc_44228_n2983_bF_buf123), .Y(u2__abc_44228_n22448) );
  OR2X2 OR2X2_5404 ( .A(u2__abc_44228_n22452), .B(u2__abc_44228_n22443), .Y(u2__abc_44228_n22453) );
  OR2X2 OR2X2_5405 ( .A(u2__abc_44228_n22445), .B(u2_o_389_), .Y(u2__abc_44228_n22456) );
  OR2X2 OR2X2_5406 ( .A(u2__abc_44228_n22459), .B(u2__abc_44228_n2983_bF_buf121), .Y(u2__abc_44228_n22460) );
  OR2X2 OR2X2_5407 ( .A(u2__abc_44228_n22464), .B(u2__abc_44228_n22455), .Y(u2__abc_44228_n22465) );
  OR2X2 OR2X2_5408 ( .A(u2__abc_44228_n22457), .B(u2_o_390_), .Y(u2__abc_44228_n22468) );
  OR2X2 OR2X2_5409 ( .A(u2__abc_44228_n22471), .B(u2__abc_44228_n2983_bF_buf119), .Y(u2__abc_44228_n22472) );
  OR2X2 OR2X2_541 ( .A(u2__abc_44228_n3072), .B(sqrto_1_), .Y(u2__abc_44228_n3073) );
  OR2X2 OR2X2_5410 ( .A(u2__abc_44228_n22476), .B(u2__abc_44228_n22467), .Y(u2__abc_44228_n22477) );
  OR2X2 OR2X2_5411 ( .A(u2__abc_44228_n22469), .B(u2_o_391_), .Y(u2__abc_44228_n22480) );
  OR2X2 OR2X2_5412 ( .A(u2__abc_44228_n22483), .B(u2__abc_44228_n2983_bF_buf117), .Y(u2__abc_44228_n22484) );
  OR2X2 OR2X2_5413 ( .A(u2__abc_44228_n22488), .B(u2__abc_44228_n22479), .Y(u2__abc_44228_n22489) );
  OR2X2 OR2X2_5414 ( .A(u2__abc_44228_n22481), .B(u2_o_392_), .Y(u2__abc_44228_n22492) );
  OR2X2 OR2X2_5415 ( .A(u2__abc_44228_n22495), .B(u2__abc_44228_n2983_bF_buf115), .Y(u2__abc_44228_n22496) );
  OR2X2 OR2X2_5416 ( .A(u2__abc_44228_n22500), .B(u2__abc_44228_n22491), .Y(u2__abc_44228_n22501) );
  OR2X2 OR2X2_5417 ( .A(u2__abc_44228_n22493), .B(u2_o_393_), .Y(u2__abc_44228_n22504) );
  OR2X2 OR2X2_5418 ( .A(u2__abc_44228_n22507), .B(u2__abc_44228_n2983_bF_buf113), .Y(u2__abc_44228_n22508) );
  OR2X2 OR2X2_5419 ( .A(u2__abc_44228_n22512), .B(u2__abc_44228_n22503), .Y(u2__abc_44228_n22513) );
  OR2X2 OR2X2_542 ( .A(u2__abc_44228_n3074), .B(u2_remHi_1_), .Y(u2__abc_44228_n3075) );
  OR2X2 OR2X2_5420 ( .A(u2__abc_44228_n22505), .B(u2_o_394_), .Y(u2__abc_44228_n22516) );
  OR2X2 OR2X2_5421 ( .A(u2__abc_44228_n22519), .B(u2__abc_44228_n2983_bF_buf111), .Y(u2__abc_44228_n22520) );
  OR2X2 OR2X2_5422 ( .A(u2__abc_44228_n22524), .B(u2__abc_44228_n22515), .Y(u2__abc_44228_n22525) );
  OR2X2 OR2X2_5423 ( .A(u2__abc_44228_n22517), .B(u2_o_395_), .Y(u2__abc_44228_n22528) );
  OR2X2 OR2X2_5424 ( .A(u2__abc_44228_n22531), .B(u2__abc_44228_n2983_bF_buf109), .Y(u2__abc_44228_n22532) );
  OR2X2 OR2X2_5425 ( .A(u2__abc_44228_n22536), .B(u2__abc_44228_n22527), .Y(u2__abc_44228_n22537) );
  OR2X2 OR2X2_5426 ( .A(u2__abc_44228_n22529), .B(u2_o_396_), .Y(u2__abc_44228_n22540) );
  OR2X2 OR2X2_5427 ( .A(u2__abc_44228_n22543), .B(u2__abc_44228_n2983_bF_buf107), .Y(u2__abc_44228_n22544) );
  OR2X2 OR2X2_5428 ( .A(u2__abc_44228_n22548), .B(u2__abc_44228_n22539), .Y(u2__abc_44228_n22549) );
  OR2X2 OR2X2_5429 ( .A(u2__abc_44228_n22541), .B(u2_o_397_), .Y(u2__abc_44228_n22552) );
  OR2X2 OR2X2_543 ( .A(u2__abc_44228_n3077), .B(u2_remHi_0_), .Y(u2__abc_44228_n3080) );
  OR2X2 OR2X2_5430 ( .A(u2__abc_44228_n22555), .B(u2__abc_44228_n2983_bF_buf105), .Y(u2__abc_44228_n22556) );
  OR2X2 OR2X2_5431 ( .A(u2__abc_44228_n22560), .B(u2__abc_44228_n22551), .Y(u2__abc_44228_n22561) );
  OR2X2 OR2X2_5432 ( .A(u2__abc_44228_n22553), .B(u2_o_398_), .Y(u2__abc_44228_n22564) );
  OR2X2 OR2X2_5433 ( .A(u2__abc_44228_n22567), .B(u2__abc_44228_n2983_bF_buf103), .Y(u2__abc_44228_n22568) );
  OR2X2 OR2X2_5434 ( .A(u2__abc_44228_n22572), .B(u2__abc_44228_n22563), .Y(u2__abc_44228_n22573) );
  OR2X2 OR2X2_5435 ( .A(u2__abc_44228_n22565), .B(u2_o_399_), .Y(u2__abc_44228_n22576) );
  OR2X2 OR2X2_5436 ( .A(u2__abc_44228_n22579), .B(u2__abc_44228_n2983_bF_buf101), .Y(u2__abc_44228_n22580) );
  OR2X2 OR2X2_5437 ( .A(u2__abc_44228_n22584), .B(u2__abc_44228_n22575), .Y(u2__abc_44228_n22585) );
  OR2X2 OR2X2_5438 ( .A(u2__abc_44228_n22577), .B(u2_o_400_), .Y(u2__abc_44228_n22588) );
  OR2X2 OR2X2_5439 ( .A(u2__abc_44228_n22591), .B(u2__abc_44228_n2983_bF_buf99), .Y(u2__abc_44228_n22592) );
  OR2X2 OR2X2_544 ( .A(u2__abc_44228_n3085), .B(u2__abc_44228_n3084), .Y(u2__abc_44228_n3086) );
  OR2X2 OR2X2_5440 ( .A(u2__abc_44228_n22596), .B(u2__abc_44228_n22587), .Y(u2__abc_44228_n22597) );
  OR2X2 OR2X2_5441 ( .A(u2__abc_44228_n22589), .B(u2_o_401_), .Y(u2__abc_44228_n22600) );
  OR2X2 OR2X2_5442 ( .A(u2__abc_44228_n22603), .B(u2__abc_44228_n2983_bF_buf97), .Y(u2__abc_44228_n22604) );
  OR2X2 OR2X2_5443 ( .A(u2__abc_44228_n22608), .B(u2__abc_44228_n22599), .Y(u2__abc_44228_n22609) );
  OR2X2 OR2X2_5444 ( .A(u2__abc_44228_n22601), .B(u2_o_402_), .Y(u2__abc_44228_n22612) );
  OR2X2 OR2X2_5445 ( .A(u2__abc_44228_n22615), .B(u2__abc_44228_n2983_bF_buf95), .Y(u2__abc_44228_n22616) );
  OR2X2 OR2X2_5446 ( .A(u2__abc_44228_n22620), .B(u2__abc_44228_n22611), .Y(u2__abc_44228_n22621) );
  OR2X2 OR2X2_5447 ( .A(u2__abc_44228_n22613), .B(u2_o_403_), .Y(u2__abc_44228_n22624) );
  OR2X2 OR2X2_5448 ( .A(u2__abc_44228_n22627), .B(u2__abc_44228_n2983_bF_buf93), .Y(u2__abc_44228_n22628) );
  OR2X2 OR2X2_5449 ( .A(u2__abc_44228_n22632), .B(u2__abc_44228_n22623), .Y(u2__abc_44228_n22633) );
  OR2X2 OR2X2_545 ( .A(u2__abc_44228_n3083), .B(u2__abc_44228_n3086), .Y(u2__abc_44228_n3087) );
  OR2X2 OR2X2_5450 ( .A(u2__abc_44228_n22625), .B(u2_o_404_), .Y(u2__abc_44228_n22636) );
  OR2X2 OR2X2_5451 ( .A(u2__abc_44228_n22639), .B(u2__abc_44228_n2983_bF_buf91), .Y(u2__abc_44228_n22640) );
  OR2X2 OR2X2_5452 ( .A(u2__abc_44228_n22644), .B(u2__abc_44228_n22635), .Y(u2__abc_44228_n22645) );
  OR2X2 OR2X2_5453 ( .A(u2__abc_44228_n22637), .B(u2_o_405_), .Y(u2__abc_44228_n22648) );
  OR2X2 OR2X2_5454 ( .A(u2__abc_44228_n22651), .B(u2__abc_44228_n2983_bF_buf89), .Y(u2__abc_44228_n22652) );
  OR2X2 OR2X2_5455 ( .A(u2__abc_44228_n22656), .B(u2__abc_44228_n22647), .Y(u2__abc_44228_n22657) );
  OR2X2 OR2X2_5456 ( .A(u2__abc_44228_n22649), .B(u2_o_406_), .Y(u2__abc_44228_n22660) );
  OR2X2 OR2X2_5457 ( .A(u2__abc_44228_n22663), .B(u2__abc_44228_n2983_bF_buf87), .Y(u2__abc_44228_n22664) );
  OR2X2 OR2X2_5458 ( .A(u2__abc_44228_n22668), .B(u2__abc_44228_n22659), .Y(u2__abc_44228_n22669) );
  OR2X2 OR2X2_5459 ( .A(u2__abc_44228_n22661), .B(u2_o_407_), .Y(u2__abc_44228_n22672) );
  OR2X2 OR2X2_546 ( .A(u2__abc_44228_n3088), .B(sqrto_5_), .Y(u2__abc_44228_n3089) );
  OR2X2 OR2X2_5460 ( .A(u2__abc_44228_n22675), .B(u2__abc_44228_n2983_bF_buf85), .Y(u2__abc_44228_n22676) );
  OR2X2 OR2X2_5461 ( .A(u2__abc_44228_n22680), .B(u2__abc_44228_n22671), .Y(u2__abc_44228_n22681) );
  OR2X2 OR2X2_5462 ( .A(u2__abc_44228_n22673), .B(u2_o_408_), .Y(u2__abc_44228_n22684) );
  OR2X2 OR2X2_5463 ( .A(u2__abc_44228_n22687), .B(u2__abc_44228_n2983_bF_buf83), .Y(u2__abc_44228_n22688) );
  OR2X2 OR2X2_5464 ( .A(u2__abc_44228_n22692), .B(u2__abc_44228_n22683), .Y(u2__abc_44228_n22693) );
  OR2X2 OR2X2_5465 ( .A(u2__abc_44228_n22685), .B(u2_o_409_), .Y(u2__abc_44228_n22696) );
  OR2X2 OR2X2_5466 ( .A(u2__abc_44228_n22699), .B(u2__abc_44228_n2983_bF_buf81), .Y(u2__abc_44228_n22700) );
  OR2X2 OR2X2_5467 ( .A(u2__abc_44228_n22704), .B(u2__abc_44228_n22695), .Y(u2__abc_44228_n22705) );
  OR2X2 OR2X2_5468 ( .A(u2__abc_44228_n22697), .B(u2_o_410_), .Y(u2__abc_44228_n22708) );
  OR2X2 OR2X2_5469 ( .A(u2__abc_44228_n22711), .B(u2__abc_44228_n2983_bF_buf79), .Y(u2__abc_44228_n22712) );
  OR2X2 OR2X2_547 ( .A(u2__abc_44228_n3090), .B(u2_remHi_5_), .Y(u2__abc_44228_n3091) );
  OR2X2 OR2X2_5470 ( .A(u2__abc_44228_n22716), .B(u2__abc_44228_n22707), .Y(u2__abc_44228_n22717) );
  OR2X2 OR2X2_5471 ( .A(u2__abc_44228_n22709), .B(u2_o_411_), .Y(u2__abc_44228_n22720) );
  OR2X2 OR2X2_5472 ( .A(u2__abc_44228_n22723), .B(u2__abc_44228_n2983_bF_buf77), .Y(u2__abc_44228_n22724) );
  OR2X2 OR2X2_5473 ( .A(u2__abc_44228_n22728), .B(u2__abc_44228_n22719), .Y(u2__abc_44228_n22729) );
  OR2X2 OR2X2_5474 ( .A(u2__abc_44228_n22721), .B(u2_o_412_), .Y(u2__abc_44228_n22732) );
  OR2X2 OR2X2_5475 ( .A(u2__abc_44228_n22735), .B(u2__abc_44228_n2983_bF_buf75), .Y(u2__abc_44228_n22736) );
  OR2X2 OR2X2_5476 ( .A(u2__abc_44228_n22740), .B(u2__abc_44228_n22731), .Y(u2__abc_44228_n22741) );
  OR2X2 OR2X2_5477 ( .A(u2__abc_44228_n22733), .B(u2_o_413_), .Y(u2__abc_44228_n22744) );
  OR2X2 OR2X2_5478 ( .A(u2__abc_44228_n22747), .B(u2__abc_44228_n2983_bF_buf73), .Y(u2__abc_44228_n22748) );
  OR2X2 OR2X2_5479 ( .A(u2__abc_44228_n22752), .B(u2__abc_44228_n22743), .Y(u2__abc_44228_n22753) );
  OR2X2 OR2X2_548 ( .A(u2__abc_44228_n3093), .B(sqrto_4_), .Y(u2__abc_44228_n3094) );
  OR2X2 OR2X2_5480 ( .A(u2__abc_44228_n22745), .B(u2_o_414_), .Y(u2__abc_44228_n22756) );
  OR2X2 OR2X2_5481 ( .A(u2__abc_44228_n22759), .B(u2__abc_44228_n2983_bF_buf71), .Y(u2__abc_44228_n22760) );
  OR2X2 OR2X2_5482 ( .A(u2__abc_44228_n22764), .B(u2__abc_44228_n22755), .Y(u2__abc_44228_n22765) );
  OR2X2 OR2X2_5483 ( .A(u2__abc_44228_n22757), .B(u2_o_415_), .Y(u2__abc_44228_n22768) );
  OR2X2 OR2X2_5484 ( .A(u2__abc_44228_n22771), .B(u2__abc_44228_n2983_bF_buf69), .Y(u2__abc_44228_n22772) );
  OR2X2 OR2X2_5485 ( .A(u2__abc_44228_n22776), .B(u2__abc_44228_n22767), .Y(u2__abc_44228_n22777) );
  OR2X2 OR2X2_5486 ( .A(u2__abc_44228_n22769), .B(u2_o_416_), .Y(u2__abc_44228_n22780) );
  OR2X2 OR2X2_5487 ( .A(u2__abc_44228_n22783), .B(u2__abc_44228_n2983_bF_buf67), .Y(u2__abc_44228_n22784) );
  OR2X2 OR2X2_5488 ( .A(u2__abc_44228_n22788), .B(u2__abc_44228_n22779), .Y(u2__abc_44228_n22789) );
  OR2X2 OR2X2_5489 ( .A(u2__abc_44228_n22781), .B(u2_o_417_), .Y(u2__abc_44228_n22792) );
  OR2X2 OR2X2_549 ( .A(u2__abc_44228_n3095), .B(u2_remHi_4_), .Y(u2__abc_44228_n3096) );
  OR2X2 OR2X2_5490 ( .A(u2__abc_44228_n22795), .B(u2__abc_44228_n2983_bF_buf65), .Y(u2__abc_44228_n22796) );
  OR2X2 OR2X2_5491 ( .A(u2__abc_44228_n22800), .B(u2__abc_44228_n22791), .Y(u2__abc_44228_n22801) );
  OR2X2 OR2X2_5492 ( .A(u2__abc_44228_n22793), .B(u2_o_418_), .Y(u2__abc_44228_n22804) );
  OR2X2 OR2X2_5493 ( .A(u2__abc_44228_n22807), .B(u2__abc_44228_n2983_bF_buf63), .Y(u2__abc_44228_n22808) );
  OR2X2 OR2X2_5494 ( .A(u2__abc_44228_n22812), .B(u2__abc_44228_n22803), .Y(u2__abc_44228_n22813) );
  OR2X2 OR2X2_5495 ( .A(u2__abc_44228_n22805), .B(u2_o_419_), .Y(u2__abc_44228_n22816) );
  OR2X2 OR2X2_5496 ( .A(u2__abc_44228_n22819), .B(u2__abc_44228_n2983_bF_buf61), .Y(u2__abc_44228_n22820) );
  OR2X2 OR2X2_5497 ( .A(u2__abc_44228_n22824), .B(u2__abc_44228_n22815), .Y(u2__abc_44228_n22825) );
  OR2X2 OR2X2_5498 ( .A(u2__abc_44228_n22817), .B(u2_o_420_), .Y(u2__abc_44228_n22828) );
  OR2X2 OR2X2_5499 ( .A(u2__abc_44228_n22831), .B(u2__abc_44228_n2983_bF_buf59), .Y(u2__abc_44228_n22832) );
  OR2X2 OR2X2_55 ( .A(aNan_bF_buf4), .B(sqrto_103_), .Y(_abc_64468_n911) );
  OR2X2 OR2X2_550 ( .A(u2__abc_44228_n3099), .B(u2_remHi_3_), .Y(u2__abc_44228_n3102) );
  OR2X2 OR2X2_5500 ( .A(u2__abc_44228_n22836), .B(u2__abc_44228_n22827), .Y(u2__abc_44228_n22837) );
  OR2X2 OR2X2_5501 ( .A(u2__abc_44228_n22829), .B(u2_o_421_), .Y(u2__abc_44228_n22840) );
  OR2X2 OR2X2_5502 ( .A(u2__abc_44228_n22843), .B(u2__abc_44228_n2983_bF_buf57), .Y(u2__abc_44228_n22844) );
  OR2X2 OR2X2_5503 ( .A(u2__abc_44228_n22848), .B(u2__abc_44228_n22839), .Y(u2__abc_44228_n22849) );
  OR2X2 OR2X2_5504 ( .A(u2__abc_44228_n22841), .B(u2_o_422_), .Y(u2__abc_44228_n22852) );
  OR2X2 OR2X2_5505 ( .A(u2__abc_44228_n22855), .B(u2__abc_44228_n2983_bF_buf55), .Y(u2__abc_44228_n22856) );
  OR2X2 OR2X2_5506 ( .A(u2__abc_44228_n22860), .B(u2__abc_44228_n22851), .Y(u2__abc_44228_n22861) );
  OR2X2 OR2X2_5507 ( .A(u2__abc_44228_n22853), .B(u2_o_423_), .Y(u2__abc_44228_n22864) );
  OR2X2 OR2X2_5508 ( .A(u2__abc_44228_n22867), .B(u2__abc_44228_n2983_bF_buf53), .Y(u2__abc_44228_n22868) );
  OR2X2 OR2X2_5509 ( .A(u2__abc_44228_n22872), .B(u2__abc_44228_n22863), .Y(u2__abc_44228_n22873) );
  OR2X2 OR2X2_551 ( .A(u2__abc_44228_n3104), .B(u2_remHi_2_), .Y(u2__abc_44228_n3107) );
  OR2X2 OR2X2_5510 ( .A(u2__abc_44228_n22865), .B(u2_o_424_), .Y(u2__abc_44228_n22876) );
  OR2X2 OR2X2_5511 ( .A(u2__abc_44228_n22879), .B(u2__abc_44228_n2983_bF_buf51), .Y(u2__abc_44228_n22880) );
  OR2X2 OR2X2_5512 ( .A(u2__abc_44228_n22884), .B(u2__abc_44228_n22875), .Y(u2__abc_44228_n22885) );
  OR2X2 OR2X2_5513 ( .A(u2__abc_44228_n22877), .B(u2_o_425_), .Y(u2__abc_44228_n22888) );
  OR2X2 OR2X2_5514 ( .A(u2__abc_44228_n22891), .B(u2__abc_44228_n2983_bF_buf49), .Y(u2__abc_44228_n22892) );
  OR2X2 OR2X2_5515 ( .A(u2__abc_44228_n22896), .B(u2__abc_44228_n22887), .Y(u2__abc_44228_n22897) );
  OR2X2 OR2X2_5516 ( .A(u2__abc_44228_n22889), .B(u2_o_426_), .Y(u2__abc_44228_n22900) );
  OR2X2 OR2X2_5517 ( .A(u2__abc_44228_n22903), .B(u2__abc_44228_n2983_bF_buf47), .Y(u2__abc_44228_n22904) );
  OR2X2 OR2X2_5518 ( .A(u2__abc_44228_n22908), .B(u2__abc_44228_n22899), .Y(u2__abc_44228_n22909) );
  OR2X2 OR2X2_5519 ( .A(u2__abc_44228_n22901), .B(u2_o_427_), .Y(u2__abc_44228_n22912) );
  OR2X2 OR2X2_552 ( .A(u2__abc_44228_n3100), .B(u2__abc_44228_n3105), .Y(u2__abc_44228_n3112) );
  OR2X2 OR2X2_5520 ( .A(u2__abc_44228_n22915), .B(u2__abc_44228_n2983_bF_buf45), .Y(u2__abc_44228_n22916) );
  OR2X2 OR2X2_5521 ( .A(u2__abc_44228_n22920), .B(u2__abc_44228_n22911), .Y(u2__abc_44228_n22921) );
  OR2X2 OR2X2_5522 ( .A(u2__abc_44228_n22913), .B(u2_o_428_), .Y(u2__abc_44228_n22924) );
  OR2X2 OR2X2_5523 ( .A(u2__abc_44228_n22927), .B(u2__abc_44228_n2983_bF_buf43), .Y(u2__abc_44228_n22928) );
  OR2X2 OR2X2_5524 ( .A(u2__abc_44228_n22932), .B(u2__abc_44228_n22923), .Y(u2__abc_44228_n22933) );
  OR2X2 OR2X2_5525 ( .A(u2__abc_44228_n22925), .B(u2_o_429_), .Y(u2__abc_44228_n22936) );
  OR2X2 OR2X2_5526 ( .A(u2__abc_44228_n22939), .B(u2__abc_44228_n2983_bF_buf41), .Y(u2__abc_44228_n22940) );
  OR2X2 OR2X2_5527 ( .A(u2__abc_44228_n22944), .B(u2__abc_44228_n22935), .Y(u2__abc_44228_n22945) );
  OR2X2 OR2X2_5528 ( .A(u2__abc_44228_n22937), .B(u2_o_430_), .Y(u2__abc_44228_n22948) );
  OR2X2 OR2X2_5529 ( .A(u2__abc_44228_n22951), .B(u2__abc_44228_n2983_bF_buf39), .Y(u2__abc_44228_n22952) );
  OR2X2 OR2X2_553 ( .A(u2__abc_44228_n3117), .B(u2__abc_44228_n3115), .Y(u2__abc_44228_n3118) );
  OR2X2 OR2X2_5530 ( .A(u2__abc_44228_n22956), .B(u2__abc_44228_n22947), .Y(u2__abc_44228_n22957) );
  OR2X2 OR2X2_5531 ( .A(u2__abc_44228_n22949), .B(u2_o_431_), .Y(u2__abc_44228_n22960) );
  OR2X2 OR2X2_5532 ( .A(u2__abc_44228_n22963), .B(u2__abc_44228_n2983_bF_buf37), .Y(u2__abc_44228_n22964) );
  OR2X2 OR2X2_5533 ( .A(u2__abc_44228_n22968), .B(u2__abc_44228_n22959), .Y(u2__abc_44228_n22969) );
  OR2X2 OR2X2_5534 ( .A(u2__abc_44228_n22961), .B(u2_o_432_), .Y(u2__abc_44228_n22972) );
  OR2X2 OR2X2_5535 ( .A(u2__abc_44228_n22975), .B(u2__abc_44228_n2983_bF_buf35), .Y(u2__abc_44228_n22976) );
  OR2X2 OR2X2_5536 ( .A(u2__abc_44228_n22980), .B(u2__abc_44228_n22971), .Y(u2__abc_44228_n22981) );
  OR2X2 OR2X2_5537 ( .A(u2__abc_44228_n22973), .B(u2_o_433_), .Y(u2__abc_44228_n22984) );
  OR2X2 OR2X2_5538 ( .A(u2__abc_44228_n22987), .B(u2__abc_44228_n2983_bF_buf33), .Y(u2__abc_44228_n22988) );
  OR2X2 OR2X2_5539 ( .A(u2__abc_44228_n22992), .B(u2__abc_44228_n22983), .Y(u2__abc_44228_n22993) );
  OR2X2 OR2X2_554 ( .A(u2__abc_44228_n3114), .B(u2__abc_44228_n3118), .Y(u2__abc_44228_n3119) );
  OR2X2 OR2X2_5540 ( .A(u2__abc_44228_n22985), .B(u2_o_434_), .Y(u2__abc_44228_n22996) );
  OR2X2 OR2X2_5541 ( .A(u2__abc_44228_n22999), .B(u2__abc_44228_n2983_bF_buf31), .Y(u2__abc_44228_n23000) );
  OR2X2 OR2X2_5542 ( .A(u2__abc_44228_n23004), .B(u2__abc_44228_n22995), .Y(u2__abc_44228_n23005) );
  OR2X2 OR2X2_5543 ( .A(u2__abc_44228_n22997), .B(u2_o_435_), .Y(u2__abc_44228_n23008) );
  OR2X2 OR2X2_5544 ( .A(u2__abc_44228_n23011), .B(u2__abc_44228_n2983_bF_buf29), .Y(u2__abc_44228_n23012) );
  OR2X2 OR2X2_5545 ( .A(u2__abc_44228_n23016), .B(u2__abc_44228_n23007), .Y(u2__abc_44228_n23017) );
  OR2X2 OR2X2_5546 ( .A(u2__abc_44228_n23009), .B(u2_o_436_), .Y(u2__abc_44228_n23020) );
  OR2X2 OR2X2_5547 ( .A(u2__abc_44228_n23023), .B(u2__abc_44228_n2983_bF_buf27), .Y(u2__abc_44228_n23024) );
  OR2X2 OR2X2_5548 ( .A(u2__abc_44228_n23028), .B(u2__abc_44228_n23019), .Y(u2__abc_44228_n23029) );
  OR2X2 OR2X2_5549 ( .A(u2__abc_44228_n23021), .B(u2_o_437_), .Y(u2__abc_44228_n23032) );
  OR2X2 OR2X2_555 ( .A(u2__abc_44228_n3111), .B(u2__abc_44228_n3119), .Y(u2__abc_44228_n3120) );
  OR2X2 OR2X2_5550 ( .A(u2__abc_44228_n23035), .B(u2__abc_44228_n2983_bF_buf25), .Y(u2__abc_44228_n23036) );
  OR2X2 OR2X2_5551 ( .A(u2__abc_44228_n23040), .B(u2__abc_44228_n23031), .Y(u2__abc_44228_n23041) );
  OR2X2 OR2X2_5552 ( .A(u2__abc_44228_n23033), .B(u2_o_438_), .Y(u2__abc_44228_n23044) );
  OR2X2 OR2X2_5553 ( .A(u2__abc_44228_n23047), .B(u2__abc_44228_n2983_bF_buf23), .Y(u2__abc_44228_n23048) );
  OR2X2 OR2X2_5554 ( .A(u2__abc_44228_n23052), .B(u2__abc_44228_n23043), .Y(u2__abc_44228_n23053) );
  OR2X2 OR2X2_5555 ( .A(u2__abc_44228_n23045), .B(u2_o_439_), .Y(u2__abc_44228_n23056) );
  OR2X2 OR2X2_5556 ( .A(u2__abc_44228_n23059), .B(u2__abc_44228_n2983_bF_buf21), .Y(u2__abc_44228_n23060) );
  OR2X2 OR2X2_5557 ( .A(u2__abc_44228_n23064), .B(u2__abc_44228_n23055), .Y(u2__abc_44228_n23065) );
  OR2X2 OR2X2_5558 ( .A(u2__abc_44228_n23057), .B(u2_o_440_), .Y(u2__abc_44228_n23068) );
  OR2X2 OR2X2_5559 ( .A(u2__abc_44228_n23071), .B(u2__abc_44228_n2983_bF_buf19), .Y(u2__abc_44228_n23072) );
  OR2X2 OR2X2_556 ( .A(u2__abc_44228_n3129), .B(u2__abc_44228_n3131), .Y(u2__abc_44228_n3132) );
  OR2X2 OR2X2_5560 ( .A(u2__abc_44228_n23076), .B(u2__abc_44228_n23067), .Y(u2__abc_44228_n23077) );
  OR2X2 OR2X2_5561 ( .A(u2__abc_44228_n23069), .B(u2_o_441_), .Y(u2__abc_44228_n23080) );
  OR2X2 OR2X2_5562 ( .A(u2__abc_44228_n23083), .B(u2__abc_44228_n2983_bF_buf17), .Y(u2__abc_44228_n23084) );
  OR2X2 OR2X2_5563 ( .A(u2__abc_44228_n23088), .B(u2__abc_44228_n23079), .Y(u2__abc_44228_n23089) );
  OR2X2 OR2X2_5564 ( .A(u2__abc_44228_n23081), .B(u2_o_442_), .Y(u2__abc_44228_n23092) );
  OR2X2 OR2X2_5565 ( .A(u2__abc_44228_n23095), .B(u2__abc_44228_n2983_bF_buf15), .Y(u2__abc_44228_n23096) );
  OR2X2 OR2X2_5566 ( .A(u2__abc_44228_n23100), .B(u2__abc_44228_n23091), .Y(u2__abc_44228_n23101) );
  OR2X2 OR2X2_5567 ( .A(u2__abc_44228_n23093), .B(u2_o_443_), .Y(u2__abc_44228_n23104) );
  OR2X2 OR2X2_5568 ( .A(u2__abc_44228_n23107), .B(u2__abc_44228_n2983_bF_buf13), .Y(u2__abc_44228_n23108) );
  OR2X2 OR2X2_5569 ( .A(u2__abc_44228_n23112), .B(u2__abc_44228_n23103), .Y(u2__abc_44228_n23113) );
  OR2X2 OR2X2_557 ( .A(u2__abc_44228_n3143), .B(u2__abc_44228_n3145), .Y(u2__abc_44228_n3146) );
  OR2X2 OR2X2_5570 ( .A(u2__abc_44228_n23105), .B(u2_o_444_), .Y(u2__abc_44228_n23116) );
  OR2X2 OR2X2_5571 ( .A(u2__abc_44228_n23119), .B(u2__abc_44228_n2983_bF_buf11), .Y(u2__abc_44228_n23120) );
  OR2X2 OR2X2_5572 ( .A(u2__abc_44228_n23124), .B(u2__abc_44228_n23115), .Y(u2__abc_44228_n23125) );
  OR2X2 OR2X2_5573 ( .A(u2__abc_44228_n23117), .B(u2_o_445_), .Y(u2__abc_44228_n23128) );
  OR2X2 OR2X2_5574 ( .A(u2__abc_44228_n23131), .B(u2__abc_44228_n2983_bF_buf9), .Y(u2__abc_44228_n23132) );
  OR2X2 OR2X2_5575 ( .A(u2__abc_44228_n23136), .B(u2__abc_44228_n23127), .Y(u2__abc_44228_n23137) );
  OR2X2 OR2X2_5576 ( .A(u2__abc_44228_n23129), .B(u2_o_446_), .Y(u2__abc_44228_n23140) );
  OR2X2 OR2X2_5577 ( .A(u2__abc_44228_n23143), .B(u2__abc_44228_n2983_bF_buf7), .Y(u2__abc_44228_n23144) );
  OR2X2 OR2X2_5578 ( .A(u2__abc_44228_n23148), .B(u2__abc_44228_n23139), .Y(u2__abc_44228_n23149) );
  OR2X2 OR2X2_5579 ( .A(u2__abc_44228_n23141), .B(u2_o_447_), .Y(u2__abc_44228_n23152) );
  OR2X2 OR2X2_558 ( .A(u2__abc_44228_n3150), .B(sqrto_9_), .Y(u2__abc_44228_n3151) );
  OR2X2 OR2X2_5580 ( .A(u2__abc_44228_n23155), .B(u2__abc_44228_n2983_bF_buf5), .Y(u2__abc_44228_n23156) );
  OR2X2 OR2X2_5581 ( .A(u2__abc_44228_n23160), .B(u2__abc_44228_n23151), .Y(u2__abc_44228_n23161) );
  OR2X2 OR2X2_5582 ( .A(u2__abc_44228_n23153), .B(u2_o_448_), .Y(u2__abc_44228_n23164) );
  OR2X2 OR2X2_5583 ( .A(u2__abc_44228_n23167), .B(u2__abc_44228_n2983_bF_buf3), .Y(u2__abc_44228_n23168) );
  OR2X2 OR2X2_5584 ( .A(u2__abc_44228_n23172), .B(u2__abc_44228_n23163), .Y(u2__abc_44228_n23173) );
  OR2X2 OR2X2_559 ( .A(u2__abc_44228_n3152), .B(u2_remHi_9_), .Y(u2__abc_44228_n3153) );
  OR2X2 OR2X2_56 ( .A(_abc_64468_n753_bF_buf8), .B(\a[27] ), .Y(_abc_64468_n912) );
  OR2X2 OR2X2_560 ( .A(u2__abc_44228_n3155), .B(sqrto_8_), .Y(u2__abc_44228_n3156) );
  OR2X2 OR2X2_561 ( .A(u2__abc_44228_n3157), .B(u2_remHi_8_), .Y(u2__abc_44228_n3158) );
  OR2X2 OR2X2_562 ( .A(u2__abc_44228_n3162), .B(u2__abc_44228_n3164), .Y(u2__abc_44228_n3165) );
  OR2X2 OR2X2_563 ( .A(u2__abc_44228_n3162), .B(u2__abc_44228_n3168), .Y(u2__abc_44228_n3178) );
  OR2X2 OR2X2_564 ( .A(u2__abc_44228_n3183), .B(u2__abc_44228_n3181), .Y(u2__abc_44228_n3184) );
  OR2X2 OR2X2_565 ( .A(u2__abc_44228_n3180), .B(u2__abc_44228_n3184), .Y(u2__abc_44228_n3185) );
  OR2X2 OR2X2_566 ( .A(u2__abc_44228_n3136), .B(u2__abc_44228_n3143), .Y(u2__abc_44228_n3187) );
  OR2X2 OR2X2_567 ( .A(u2__abc_44228_n3190), .B(u2__abc_44228_n3122), .Y(u2__abc_44228_n3191) );
  OR2X2 OR2X2_568 ( .A(u2__abc_44228_n3189), .B(u2__abc_44228_n3191), .Y(u2__abc_44228_n3192) );
  OR2X2 OR2X2_569 ( .A(u2__abc_44228_n3186), .B(u2__abc_44228_n3192), .Y(u2__abc_44228_n3193) );
  OR2X2 OR2X2_57 ( .A(aNan_bF_buf3), .B(sqrto_104_), .Y(_abc_64468_n914) );
  OR2X2 OR2X2_570 ( .A(u2__abc_44228_n3177), .B(u2__abc_44228_n3193), .Y(u2__abc_44228_n3194) );
  OR2X2 OR2X2_571 ( .A(u2__abc_44228_n3203), .B(u2__abc_44228_n3205), .Y(u2__abc_44228_n3206) );
  OR2X2 OR2X2_572 ( .A(u2__abc_44228_n3210), .B(u2__abc_44228_n3212), .Y(u2__abc_44228_n3213) );
  OR2X2 OR2X2_573 ( .A(u2__abc_44228_n3232), .B(u2__abc_44228_n3234), .Y(u2__abc_44228_n3235) );
  OR2X2 OR2X2_574 ( .A(u2__abc_44228_n3246), .B(u2__abc_44228_n3248), .Y(u2__abc_44228_n3249) );
  OR2X2 OR2X2_575 ( .A(u2__abc_44228_n3262), .B(u2__abc_44228_n3264), .Y(u2__abc_44228_n3265) );
  OR2X2 OR2X2_576 ( .A(u2__abc_44228_n3269), .B(u2__abc_44228_n3271), .Y(u2__abc_44228_n3272) );
  OR2X2 OR2X2_577 ( .A(u2__abc_44228_n3283), .B(sqrto_17_), .Y(u2__abc_44228_n3284) );
  OR2X2 OR2X2_578 ( .A(u2__abc_44228_n3285), .B(u2_remHi_17_), .Y(u2__abc_44228_n3286) );
  OR2X2 OR2X2_579 ( .A(u2__abc_44228_n3288), .B(sqrto_16_), .Y(u2__abc_44228_n3289) );
  OR2X2 OR2X2_58 ( .A(_abc_64468_n753_bF_buf7), .B(\a[28] ), .Y(_abc_64468_n915) );
  OR2X2 OR2X2_580 ( .A(u2__abc_44228_n3290), .B(u2_remHi_16_), .Y(u2__abc_44228_n3291) );
  OR2X2 OR2X2_581 ( .A(u2__abc_44228_n3302), .B(u2__abc_44228_n3304), .Y(u2__abc_44228_n3305) );
  OR2X2 OR2X2_582 ( .A(u2__abc_44228_n3295), .B(u2__abc_44228_n3302), .Y(u2__abc_44228_n3312) );
  OR2X2 OR2X2_583 ( .A(u2__abc_44228_n3317), .B(u2__abc_44228_n3315), .Y(u2__abc_44228_n3318) );
  OR2X2 OR2X2_584 ( .A(u2__abc_44228_n3314), .B(u2__abc_44228_n3318), .Y(u2__abc_44228_n3319) );
  OR2X2 OR2X2_585 ( .A(u2__abc_44228_n3269), .B(u2__abc_44228_n3275), .Y(u2__abc_44228_n3321) );
  OR2X2 OR2X2_586 ( .A(u2__abc_44228_n3324), .B(u2__abc_44228_n3255), .Y(u2__abc_44228_n3325) );
  OR2X2 OR2X2_587 ( .A(u2__abc_44228_n3323), .B(u2__abc_44228_n3325), .Y(u2__abc_44228_n3326) );
  OR2X2 OR2X2_588 ( .A(u2__abc_44228_n3320), .B(u2__abc_44228_n3326), .Y(u2__abc_44228_n3327) );
  OR2X2 OR2X2_589 ( .A(u2__abc_44228_n3225), .B(u2__abc_44228_n3232), .Y(u2__abc_44228_n3329) );
  OR2X2 OR2X2_59 ( .A(aNan_bF_buf2), .B(sqrto_105_), .Y(_abc_64468_n917) );
  OR2X2 OR2X2_590 ( .A(u2__abc_44228_n3331), .B(u2__abc_44228_n3335), .Y(u2__abc_44228_n3336) );
  OR2X2 OR2X2_591 ( .A(u2__abc_44228_n3343), .B(u2__abc_44228_n3196), .Y(u2__abc_44228_n3344) );
  OR2X2 OR2X2_592 ( .A(u2__abc_44228_n3342), .B(u2__abc_44228_n3344), .Y(u2__abc_44228_n3345) );
  OR2X2 OR2X2_593 ( .A(u2__abc_44228_n3337), .B(u2__abc_44228_n3345), .Y(u2__abc_44228_n3346) );
  OR2X2 OR2X2_594 ( .A(u2__abc_44228_n3328), .B(u2__abc_44228_n3346), .Y(u2__abc_44228_n3347) );
  OR2X2 OR2X2_595 ( .A(u2__abc_44228_n3311), .B(u2__abc_44228_n3347), .Y(u2__abc_44228_n3348) );
  OR2X2 OR2X2_596 ( .A(u2__abc_44228_n3357), .B(u2__abc_44228_n3359), .Y(u2__abc_44228_n3360) );
  OR2X2 OR2X2_597 ( .A(u2__abc_44228_n3364), .B(u2__abc_44228_n3366), .Y(u2__abc_44228_n3367) );
  OR2X2 OR2X2_598 ( .A(u2__abc_44228_n3386), .B(u2__abc_44228_n3388), .Y(u2__abc_44228_n3389) );
  OR2X2 OR2X2_599 ( .A(u2__abc_44228_n3400), .B(u2__abc_44228_n3402), .Y(u2__abc_44228_n3403) );
  OR2X2 OR2X2_6 ( .A(_abc_64468_n753_bF_buf5), .B(\a[2] ), .Y(_abc_64468_n837) );
  OR2X2 OR2X2_60 ( .A(_abc_64468_n753_bF_buf6), .B(\a[29] ), .Y(_abc_64468_n918) );
  OR2X2 OR2X2_600 ( .A(u2__abc_44228_n3416), .B(u2__abc_44228_n3418), .Y(u2__abc_44228_n3419) );
  OR2X2 OR2X2_601 ( .A(u2__abc_44228_n3423), .B(u2__abc_44228_n3425), .Y(u2__abc_44228_n3426) );
  OR2X2 OR2X2_602 ( .A(u2__abc_44228_n3445), .B(u2__abc_44228_n3447), .Y(u2__abc_44228_n3448) );
  OR2X2 OR2X2_603 ( .A(u2__abc_44228_n3459), .B(u2__abc_44228_n3461), .Y(u2__abc_44228_n3462) );
  OR2X2 OR2X2_604 ( .A(u2__abc_44228_n3476), .B(u2__abc_44228_n3478), .Y(u2__abc_44228_n3479) );
  OR2X2 OR2X2_605 ( .A(u2__abc_44228_n3483), .B(u2__abc_44228_n3485), .Y(u2__abc_44228_n3486) );
  OR2X2 OR2X2_606 ( .A(u2__abc_44228_n3505_1), .B(u2__abc_44228_n3507), .Y(u2__abc_44228_n3508) );
  OR2X2 OR2X2_607 ( .A(u2__abc_44228_n3519), .B(u2__abc_44228_n3521), .Y(u2__abc_44228_n3522) );
  OR2X2 OR2X2_608 ( .A(u2__abc_44228_n3535), .B(u2__abc_44228_n3537), .Y(u2__abc_44228_n3538) );
  OR2X2 OR2X2_609 ( .A(u2__abc_44228_n3542), .B(u2__abc_44228_n3544), .Y(u2__abc_44228_n3545) );
  OR2X2 OR2X2_61 ( .A(aNan_bF_buf1), .B(sqrto_106_), .Y(_abc_64468_n920) );
  OR2X2 OR2X2_610 ( .A(u2__abc_44228_n3556), .B(sqrto_33_), .Y(u2__abc_44228_n3557) );
  OR2X2 OR2X2_611 ( .A(u2__abc_44228_n3558), .B(u2_remHi_33_), .Y(u2__abc_44228_n3559) );
  OR2X2 OR2X2_612 ( .A(u2__abc_44228_n3561), .B(sqrto_32_), .Y(u2__abc_44228_n3562_1) );
  OR2X2 OR2X2_613 ( .A(u2__abc_44228_n3563), .B(u2_remHi_32_), .Y(u2__abc_44228_n3564) );
  OR2X2 OR2X2_614 ( .A(u2__abc_44228_n3568), .B(u2__abc_44228_n3570), .Y(u2__abc_44228_n3571_1) );
  OR2X2 OR2X2_615 ( .A(u2__abc_44228_n3568), .B(u2__abc_44228_n3574), .Y(u2__abc_44228_n3586) );
  OR2X2 OR2X2_616 ( .A(u2__abc_44228_n3591), .B(u2__abc_44228_n3589), .Y(u2__abc_44228_n3592) );
  OR2X2 OR2X2_617 ( .A(u2__abc_44228_n3588_1), .B(u2__abc_44228_n3592), .Y(u2__abc_44228_n3593) );
  OR2X2 OR2X2_618 ( .A(u2__abc_44228_n3528), .B(u2__abc_44228_n3535), .Y(u2__abc_44228_n3600) );
  OR2X2 OR2X2_619 ( .A(u2__abc_44228_n3599), .B(u2__abc_44228_n3601), .Y(u2__abc_44228_n3602) );
  OR2X2 OR2X2_62 ( .A(_abc_64468_n753_bF_buf5), .B(\a[30] ), .Y(_abc_64468_n921) );
  OR2X2 OR2X2_620 ( .A(u2__abc_44228_n3594), .B(u2__abc_44228_n3602), .Y(u2__abc_44228_n3603) );
  OR2X2 OR2X2_621 ( .A(u2__abc_44228_n3498), .B(u2__abc_44228_n3505_1), .Y(u2__abc_44228_n3605) );
  OR2X2 OR2X2_622 ( .A(u2__abc_44228_n3607), .B(u2__abc_44228_n3611), .Y(u2__abc_44228_n3612) );
  OR2X2 OR2X2_623 ( .A(u2__abc_44228_n3614), .B(u2__abc_44228_n3469), .Y(u2__abc_44228_n3615) );
  OR2X2 OR2X2_624 ( .A(u2__abc_44228_n3620), .B(u2__abc_44228_n3615), .Y(u2__abc_44228_n3621) );
  OR2X2 OR2X2_625 ( .A(u2__abc_44228_n3613), .B(u2__abc_44228_n3621), .Y(u2__abc_44228_n3622) );
  OR2X2 OR2X2_626 ( .A(u2__abc_44228_n3604), .B(u2__abc_44228_n3622), .Y(u2__abc_44228_n3623) );
  OR2X2 OR2X2_627 ( .A(u2__abc_44228_n3452), .B(u2__abc_44228_n3459), .Y(u2__abc_44228_n3625) );
  OR2X2 OR2X2_628 ( .A(u2__abc_44228_n3628), .B(u2__abc_44228_n3438), .Y(u2__abc_44228_n3629) );
  OR2X2 OR2X2_629 ( .A(u2__abc_44228_n3627_1), .B(u2__abc_44228_n3629), .Y(u2__abc_44228_n3630) );
  OR2X2 OR2X2_63 ( .A(aNan_bF_buf0), .B(sqrto_107_), .Y(_abc_64468_n923) );
  OR2X2 OR2X2_630 ( .A(u2__abc_44228_n3637_1), .B(u2__abc_44228_n3409), .Y(u2__abc_44228_n3638) );
  OR2X2 OR2X2_631 ( .A(u2__abc_44228_n3636), .B(u2__abc_44228_n3638), .Y(u2__abc_44228_n3639) );
  OR2X2 OR2X2_632 ( .A(u2__abc_44228_n3631), .B(u2__abc_44228_n3639), .Y(u2__abc_44228_n3640) );
  OR2X2 OR2X2_633 ( .A(u2__abc_44228_n3642), .B(u2__abc_44228_n3396), .Y(u2__abc_44228_n3643) );
  OR2X2 OR2X2_634 ( .A(u2__abc_44228_n3646), .B(u2__abc_44228_n3650), .Y(u2__abc_44228_n3651) );
  OR2X2 OR2X2_635 ( .A(u2__abc_44228_n3653), .B(u2__abc_44228_n3350), .Y(u2__abc_44228_n3654) );
  OR2X2 OR2X2_636 ( .A(u2__abc_44228_n3659), .B(u2__abc_44228_n3654), .Y(u2__abc_44228_n3660) );
  OR2X2 OR2X2_637 ( .A(u2__abc_44228_n3652), .B(u2__abc_44228_n3660), .Y(u2__abc_44228_n3661) );
  OR2X2 OR2X2_638 ( .A(u2__abc_44228_n3641), .B(u2__abc_44228_n3661), .Y(u2__abc_44228_n3662) );
  OR2X2 OR2X2_639 ( .A(u2__abc_44228_n3624), .B(u2__abc_44228_n3662), .Y(u2__abc_44228_n3663) );
  OR2X2 OR2X2_64 ( .A(_abc_64468_n753_bF_buf4), .B(\a[31] ), .Y(_abc_64468_n924) );
  OR2X2 OR2X2_640 ( .A(u2__abc_44228_n3585), .B(u2__abc_44228_n3663), .Y(u2__abc_44228_n3664) );
  OR2X2 OR2X2_641 ( .A(u2__abc_44228_n3673), .B(u2__abc_44228_n3675_1), .Y(u2__abc_44228_n3676) );
  OR2X2 OR2X2_642 ( .A(u2__abc_44228_n3680), .B(u2__abc_44228_n3682), .Y(u2__abc_44228_n3683) );
  OR2X2 OR2X2_643 ( .A(u2__abc_44228_n3702), .B(u2__abc_44228_n3704_1), .Y(u2__abc_44228_n3705) );
  OR2X2 OR2X2_644 ( .A(u2__abc_44228_n3716), .B(u2__abc_44228_n3718), .Y(u2__abc_44228_n3719) );
  OR2X2 OR2X2_645 ( .A(u2__abc_44228_n3732_1), .B(u2__abc_44228_n3734), .Y(u2__abc_44228_n3735) );
  OR2X2 OR2X2_646 ( .A(u2__abc_44228_n3746), .B(u2__abc_44228_n3748), .Y(u2__abc_44228_n3749) );
  OR2X2 OR2X2_647 ( .A(u2__abc_44228_n3761), .B(u2__abc_44228_n3763), .Y(u2__abc_44228_n3764) );
  OR2X2 OR2X2_648 ( .A(u2__abc_44228_n3768_1), .B(u2__abc_44228_n3770), .Y(u2__abc_44228_n3771) );
  OR2X2 OR2X2_649 ( .A(u2__abc_44228_n3792), .B(u2__abc_44228_n3794), .Y(u2__abc_44228_n3795) );
  OR2X2 OR2X2_65 ( .A(aNan_bF_buf10), .B(sqrto_108_), .Y(_abc_64468_n926) );
  OR2X2 OR2X2_650 ( .A(u2__abc_44228_n3799), .B(u2__abc_44228_n3801), .Y(u2__abc_44228_n3802) );
  OR2X2 OR2X2_651 ( .A(u2__abc_44228_n3821), .B(u2__abc_44228_n3823), .Y(u2__abc_44228_n3824) );
  OR2X2 OR2X2_652 ( .A(u2__abc_44228_n3835_1), .B(u2__abc_44228_n3837), .Y(u2__abc_44228_n3838) );
  OR2X2 OR2X2_653 ( .A(u2__abc_44228_n3851), .B(u2__abc_44228_n3853), .Y(u2__abc_44228_n3854_1) );
  OR2X2 OR2X2_654 ( .A(u2__abc_44228_n3858), .B(u2__abc_44228_n3860), .Y(u2__abc_44228_n3861) );
  OR2X2 OR2X2_655 ( .A(u2__abc_44228_n3880), .B(u2__abc_44228_n3882_1), .Y(u2__abc_44228_n3883) );
  OR2X2 OR2X2_656 ( .A(u2__abc_44228_n3887), .B(u2__abc_44228_n3889), .Y(u2__abc_44228_n3890) );
  OR2X2 OR2X2_657 ( .A(u2__abc_44228_n3912_1), .B(u2__abc_44228_n3914), .Y(u2__abc_44228_n3915) );
  OR2X2 OR2X2_658 ( .A(u2__abc_44228_n3919), .B(u2__abc_44228_n3921_1), .Y(u2__abc_44228_n3922) );
  OR2X2 OR2X2_659 ( .A(u2__abc_44228_n3941), .B(u2__abc_44228_n3943), .Y(u2__abc_44228_n3944) );
  OR2X2 OR2X2_66 ( .A(_abc_64468_n753_bF_buf3), .B(\a[32] ), .Y(_abc_64468_n927) );
  OR2X2 OR2X2_660 ( .A(u2__abc_44228_n3948), .B(u2__abc_44228_n3950), .Y(u2__abc_44228_n3951) );
  OR2X2 OR2X2_661 ( .A(u2__abc_44228_n3971), .B(u2__abc_44228_n3973), .Y(u2__abc_44228_n3974) );
  OR2X2 OR2X2_662 ( .A(u2__abc_44228_n3978), .B(u2__abc_44228_n3980), .Y(u2__abc_44228_n3981) );
  OR2X2 OR2X2_663 ( .A(u2__abc_44228_n4000), .B(u2__abc_44228_n4002), .Y(u2__abc_44228_n4003) );
  OR2X2 OR2X2_664 ( .A(u2__abc_44228_n4007), .B(u2__abc_44228_n4009), .Y(u2__abc_44228_n4010) );
  OR2X2 OR2X2_665 ( .A(u2__abc_44228_n4031), .B(u2__abc_44228_n4033_1), .Y(u2__abc_44228_n4034) );
  OR2X2 OR2X2_666 ( .A(u2__abc_44228_n4038), .B(u2__abc_44228_n4040), .Y(u2__abc_44228_n4041_1) );
  OR2X2 OR2X2_667 ( .A(u2__abc_44228_n4060), .B(u2__abc_44228_n4062), .Y(u2__abc_44228_n4063) );
  OR2X2 OR2X2_668 ( .A(u2__abc_44228_n4074), .B(u2__abc_44228_n4076), .Y(u2__abc_44228_n4077) );
  OR2X2 OR2X2_669 ( .A(u2__abc_44228_n4090_1), .B(u2__abc_44228_n4092), .Y(u2__abc_44228_n4093) );
  OR2X2 OR2X2_67 ( .A(aNan_bF_buf9), .B(sqrto_109_), .Y(_abc_64468_n929) );
  OR2X2 OR2X2_670 ( .A(u2__abc_44228_n4104), .B(u2__abc_44228_n4106), .Y(u2__abc_44228_n4107) );
  OR2X2 OR2X2_671 ( .A(u2__abc_44228_n4111), .B(sqrto_65_), .Y(u2__abc_44228_n4112) );
  OR2X2 OR2X2_672 ( .A(u2__abc_44228_n4113), .B(u2_remHi_65_), .Y(u2__abc_44228_n4114) );
  OR2X2 OR2X2_673 ( .A(u2__abc_44228_n4116), .B(sqrto_64_), .Y(u2__abc_44228_n4117) );
  OR2X2 OR2X2_674 ( .A(u2__abc_44228_n4118), .B(u2_remHi_64_), .Y(u2__abc_44228_n4119_1) );
  OR2X2 OR2X2_675 ( .A(u2__abc_44228_n4130), .B(u2__abc_44228_n4132), .Y(u2__abc_44228_n4133) );
  OR2X2 OR2X2_676 ( .A(u2__abc_44228_n4123), .B(u2__abc_44228_n4130), .Y(u2__abc_44228_n4142) );
  OR2X2 OR2X2_677 ( .A(u2__abc_44228_n4147_1), .B(u2__abc_44228_n4145), .Y(u2__abc_44228_n4148) );
  OR2X2 OR2X2_678 ( .A(u2__abc_44228_n4144), .B(u2__abc_44228_n4148), .Y(u2__abc_44228_n4149) );
  OR2X2 OR2X2_679 ( .A(u2__abc_44228_n4097), .B(u2__abc_44228_n4104), .Y(u2__abc_44228_n4151) );
  OR2X2 OR2X2_68 ( .A(_abc_64468_n753_bF_buf2), .B(\a[33] ), .Y(_abc_64468_n930) );
  OR2X2 OR2X2_680 ( .A(u2__abc_44228_n4154), .B(u2__abc_44228_n4083), .Y(u2__abc_44228_n4155) );
  OR2X2 OR2X2_681 ( .A(u2__abc_44228_n4153), .B(u2__abc_44228_n4155), .Y(u2__abc_44228_n4156) );
  OR2X2 OR2X2_682 ( .A(u2__abc_44228_n4150), .B(u2__abc_44228_n4156), .Y(u2__abc_44228_n4157_1) );
  OR2X2 OR2X2_683 ( .A(u2__abc_44228_n4053), .B(u2__abc_44228_n4060), .Y(u2__abc_44228_n4159) );
  OR2X2 OR2X2_684 ( .A(u2__abc_44228_n4161), .B(u2__abc_44228_n4165), .Y(u2__abc_44228_n4166) );
  OR2X2 OR2X2_685 ( .A(u2__abc_44228_n4173), .B(u2__abc_44228_n4024_1), .Y(u2__abc_44228_n4174) );
  OR2X2 OR2X2_686 ( .A(u2__abc_44228_n4174), .B(u2__abc_44228_n4168), .Y(u2__abc_44228_n4175) );
  OR2X2 OR2X2_687 ( .A(u2__abc_44228_n4175), .B(u2__abc_44228_n4167_1), .Y(u2__abc_44228_n4176_1) );
  OR2X2 OR2X2_688 ( .A(u2__abc_44228_n4176_1), .B(u2__abc_44228_n4158), .Y(u2__abc_44228_n4177) );
  OR2X2 OR2X2_689 ( .A(u2__abc_44228_n4184), .B(u2__abc_44228_n3993), .Y(u2__abc_44228_n4185_1) );
  OR2X2 OR2X2_69 ( .A(aNan_bF_buf8), .B(sqrto_110_), .Y(_abc_64468_n932) );
  OR2X2 OR2X2_690 ( .A(u2__abc_44228_n4183), .B(u2__abc_44228_n4185_1), .Y(u2__abc_44228_n4186) );
  OR2X2 OR2X2_691 ( .A(u2__abc_44228_n4188), .B(u2__abc_44228_n3987), .Y(u2__abc_44228_n4189) );
  OR2X2 OR2X2_692 ( .A(u2__abc_44228_n4193), .B(u2__abc_44228_n3964), .Y(u2__abc_44228_n4194) );
  OR2X2 OR2X2_693 ( .A(u2__abc_44228_n4192), .B(u2__abc_44228_n4194), .Y(u2__abc_44228_n4195_1) );
  OR2X2 OR2X2_694 ( .A(u2__abc_44228_n4187), .B(u2__abc_44228_n4195_1), .Y(u2__abc_44228_n4196) );
  OR2X2 OR2X2_695 ( .A(u2__abc_44228_n4203), .B(u2__abc_44228_n3934), .Y(u2__abc_44228_n4204) );
  OR2X2 OR2X2_696 ( .A(u2__abc_44228_n4202), .B(u2__abc_44228_n4204), .Y(u2__abc_44228_n4205_1) );
  OR2X2 OR2X2_697 ( .A(u2__abc_44228_n4212), .B(u2__abc_44228_n3905), .Y(u2__abc_44228_n4213) );
  OR2X2 OR2X2_698 ( .A(u2__abc_44228_n4211), .B(u2__abc_44228_n4213), .Y(u2__abc_44228_n4214) );
  OR2X2 OR2X2_699 ( .A(u2__abc_44228_n4206), .B(u2__abc_44228_n4214), .Y(u2__abc_44228_n4215_1) );
  OR2X2 OR2X2_7 ( .A(aNan_bF_buf6), .B(sqrto_79_), .Y(_abc_64468_n839_1) );
  OR2X2 OR2X2_70 ( .A(_abc_64468_n753_bF_buf1), .B(\a[34] ), .Y(_abc_64468_n933) );
  OR2X2 OR2X2_700 ( .A(u2__abc_44228_n4197), .B(u2__abc_44228_n4215_1), .Y(u2__abc_44228_n4216) );
  OR2X2 OR2X2_701 ( .A(u2__abc_44228_n4178), .B(u2__abc_44228_n4216), .Y(u2__abc_44228_n4217) );
  OR2X2 OR2X2_702 ( .A(u2__abc_44228_n4224_1), .B(u2__abc_44228_n3873_1), .Y(u2__abc_44228_n4225) );
  OR2X2 OR2X2_703 ( .A(u2__abc_44228_n4223), .B(u2__abc_44228_n4225), .Y(u2__abc_44228_n4226) );
  OR2X2 OR2X2_704 ( .A(u2__abc_44228_n4228), .B(u2__abc_44228_n3867), .Y(u2__abc_44228_n4229) );
  OR2X2 OR2X2_705 ( .A(u2__abc_44228_n4233_1), .B(u2__abc_44228_n3844_1), .Y(u2__abc_44228_n4234) );
  OR2X2 OR2X2_706 ( .A(u2__abc_44228_n4232), .B(u2__abc_44228_n4234), .Y(u2__abc_44228_n4235) );
  OR2X2 OR2X2_707 ( .A(u2__abc_44228_n4227), .B(u2__abc_44228_n4235), .Y(u2__abc_44228_n4236) );
  OR2X2 OR2X2_708 ( .A(u2__abc_44228_n4238), .B(u2__abc_44228_n3817), .Y(u2__abc_44228_n4239) );
  OR2X2 OR2X2_709 ( .A(u2__abc_44228_n4242), .B(u2__abc_44228_n4246), .Y(u2__abc_44228_n4247) );
  OR2X2 OR2X2_71 ( .A(aNan_bF_buf7), .B(sqrto_111_), .Y(_abc_64468_n935) );
  OR2X2 OR2X2_710 ( .A(u2__abc_44228_n4254), .B(u2__abc_44228_n3785), .Y(u2__abc_44228_n4255) );
  OR2X2 OR2X2_711 ( .A(u2__abc_44228_n4253_1), .B(u2__abc_44228_n4255), .Y(u2__abc_44228_n4256) );
  OR2X2 OR2X2_712 ( .A(u2__abc_44228_n4248), .B(u2__abc_44228_n4256), .Y(u2__abc_44228_n4257) );
  OR2X2 OR2X2_713 ( .A(u2__abc_44228_n4237), .B(u2__abc_44228_n4257), .Y(u2__abc_44228_n4258) );
  OR2X2 OR2X2_714 ( .A(u2__abc_44228_n4260), .B(u2__abc_44228_n3698), .Y(u2__abc_44228_n4261) );
  OR2X2 OR2X2_715 ( .A(u2__abc_44228_n3709), .B(u2__abc_44228_n3716), .Y(u2__abc_44228_n4265) );
  OR2X2 OR2X2_716 ( .A(u2__abc_44228_n4264), .B(u2__abc_44228_n4266), .Y(u2__abc_44228_n4267) );
  OR2X2 OR2X2_717 ( .A(u2__abc_44228_n4274), .B(u2__abc_44228_n3666_1), .Y(u2__abc_44228_n4275) );
  OR2X2 OR2X2_718 ( .A(u2__abc_44228_n4273), .B(u2__abc_44228_n4275), .Y(u2__abc_44228_n4276) );
  OR2X2 OR2X2_719 ( .A(u2__abc_44228_n4268), .B(u2__abc_44228_n4276), .Y(u2__abc_44228_n4277) );
  OR2X2 OR2X2_72 ( .A(_abc_64468_n753_bF_buf0), .B(\a[35] ), .Y(_abc_64468_n936) );
  OR2X2 OR2X2_720 ( .A(u2__abc_44228_n4283), .B(u2__abc_44228_n3754), .Y(u2__abc_44228_n4284) );
  OR2X2 OR2X2_721 ( .A(u2__abc_44228_n4282), .B(u2__abc_44228_n4284), .Y(u2__abc_44228_n4285) );
  OR2X2 OR2X2_722 ( .A(u2__abc_44228_n4287), .B(u2__abc_44228_n3742), .Y(u2__abc_44228_n4288) );
  OR2X2 OR2X2_723 ( .A(u2__abc_44228_n4292), .B(u2__abc_44228_n3725), .Y(u2__abc_44228_n4293) );
  OR2X2 OR2X2_724 ( .A(u2__abc_44228_n4291_1), .B(u2__abc_44228_n4293), .Y(u2__abc_44228_n4294) );
  OR2X2 OR2X2_725 ( .A(u2__abc_44228_n4286), .B(u2__abc_44228_n4294), .Y(u2__abc_44228_n4295) );
  OR2X2 OR2X2_726 ( .A(u2__abc_44228_n4296), .B(u2__abc_44228_n4277), .Y(u2__abc_44228_n4297) );
  OR2X2 OR2X2_727 ( .A(u2__abc_44228_n4259), .B(u2__abc_44228_n4297), .Y(u2__abc_44228_n4298) );
  OR2X2 OR2X2_728 ( .A(u2__abc_44228_n4218), .B(u2__abc_44228_n4298), .Y(u2__abc_44228_n4299) );
  OR2X2 OR2X2_729 ( .A(u2__abc_44228_n4141), .B(u2__abc_44228_n4299), .Y(u2__abc_44228_n4300_1) );
  OR2X2 OR2X2_73 ( .A(aNan_bF_buf6), .B(sqrto_112_), .Y(_abc_64468_n938) );
  OR2X2 OR2X2_730 ( .A(u2__abc_44228_n4309), .B(u2__abc_44228_n4311), .Y(u2__abc_44228_n4312) );
  OR2X2 OR2X2_731 ( .A(u2__abc_44228_n4316), .B(u2__abc_44228_n4318), .Y(u2__abc_44228_n4319) );
  OR2X2 OR2X2_732 ( .A(u2__abc_44228_n4338_1), .B(u2__abc_44228_n4340), .Y(u2__abc_44228_n4341) );
  OR2X2 OR2X2_733 ( .A(u2__abc_44228_n4345), .B(u2__abc_44228_n4347), .Y(u2__abc_44228_n4348) );
  OR2X2 OR2X2_734 ( .A(u2__abc_44228_n4368_1), .B(u2__abc_44228_n4370), .Y(u2__abc_44228_n4371) );
  OR2X2 OR2X2_735 ( .A(u2__abc_44228_n4375), .B(u2__abc_44228_n4377_1), .Y(u2__abc_44228_n4378) );
  OR2X2 OR2X2_736 ( .A(u2__abc_44228_n4397), .B(u2__abc_44228_n4399), .Y(u2__abc_44228_n4400) );
  OR2X2 OR2X2_737 ( .A(u2__abc_44228_n4404), .B(u2__abc_44228_n4406), .Y(u2__abc_44228_n4407) );
  OR2X2 OR2X2_738 ( .A(u2__abc_44228_n4428), .B(u2__abc_44228_n4430), .Y(u2__abc_44228_n4431) );
  OR2X2 OR2X2_739 ( .A(u2__abc_44228_n4435), .B(u2__abc_44228_n4437), .Y(u2__abc_44228_n4438) );
  OR2X2 OR2X2_74 ( .A(_abc_64468_n753_bF_buf13), .B(\a[36] ), .Y(_abc_64468_n939) );
  OR2X2 OR2X2_740 ( .A(u2__abc_44228_n4457), .B(u2__abc_44228_n4459), .Y(u2__abc_44228_n4460) );
  OR2X2 OR2X2_741 ( .A(u2__abc_44228_n4471_1), .B(u2__abc_44228_n4473), .Y(u2__abc_44228_n4474) );
  OR2X2 OR2X2_742 ( .A(u2__abc_44228_n4487), .B(u2__abc_44228_n4489_1), .Y(u2__abc_44228_n4490) );
  OR2X2 OR2X2_743 ( .A(u2__abc_44228_n4494), .B(u2__abc_44228_n4496), .Y(u2__abc_44228_n4497) );
  OR2X2 OR2X2_744 ( .A(u2__abc_44228_n4516), .B(u2__abc_44228_n4518), .Y(u2__abc_44228_n4519) );
  OR2X2 OR2X2_745 ( .A(u2__abc_44228_n4523), .B(u2__abc_44228_n4525), .Y(u2__abc_44228_n4526_1) );
  OR2X2 OR2X2_746 ( .A(u2__abc_44228_n4548), .B(u2__abc_44228_n4550), .Y(u2__abc_44228_n4551) );
  OR2X2 OR2X2_747 ( .A(u2__abc_44228_n4555), .B(u2__abc_44228_n4557), .Y(u2__abc_44228_n4558) );
  OR2X2 OR2X2_748 ( .A(u2__abc_44228_n4577), .B(u2__abc_44228_n4579), .Y(u2__abc_44228_n4580) );
  OR2X2 OR2X2_749 ( .A(u2__abc_44228_n4584), .B(u2__abc_44228_n4586), .Y(u2__abc_44228_n4587) );
  OR2X2 OR2X2_75 ( .A(aNan_bF_buf5), .B(sqrto_113_), .Y(_abc_64468_n941) );
  OR2X2 OR2X2_750 ( .A(u2__abc_44228_n4607), .B(u2__abc_44228_n4609), .Y(u2__abc_44228_n4610_1) );
  OR2X2 OR2X2_751 ( .A(u2__abc_44228_n4614), .B(u2__abc_44228_n4616), .Y(u2__abc_44228_n4617) );
  OR2X2 OR2X2_752 ( .A(u2__abc_44228_n4636), .B(u2__abc_44228_n4638_1), .Y(u2__abc_44228_n4639) );
  OR2X2 OR2X2_753 ( .A(u2__abc_44228_n4650), .B(u2__abc_44228_n4652), .Y(u2__abc_44228_n4653) );
  OR2X2 OR2X2_754 ( .A(u2__abc_44228_n4667), .B(u2__abc_44228_n4669), .Y(u2__abc_44228_n4670) );
  OR2X2 OR2X2_755 ( .A(u2__abc_44228_n4681), .B(u2__abc_44228_n4683), .Y(u2__abc_44228_n4684) );
  OR2X2 OR2X2_756 ( .A(u2__abc_44228_n4696), .B(u2__abc_44228_n4698), .Y(u2__abc_44228_n4699) );
  OR2X2 OR2X2_757 ( .A(u2__abc_44228_n4703), .B(u2__abc_44228_n4705), .Y(u2__abc_44228_n4706) );
  OR2X2 OR2X2_758 ( .A(u2__abc_44228_n4726), .B(u2__abc_44228_n4728), .Y(u2__abc_44228_n4729) );
  OR2X2 OR2X2_759 ( .A(u2__abc_44228_n4740), .B(u2__abc_44228_n4742), .Y(u2__abc_44228_n4743) );
  OR2X2 OR2X2_76 ( .A(_abc_64468_n753_bF_buf12), .B(\a[37] ), .Y(_abc_64468_n942) );
  OR2X2 OR2X2_760 ( .A(u2__abc_44228_n4755), .B(u2__abc_44228_n4757), .Y(u2__abc_44228_n4758) );
  OR2X2 OR2X2_761 ( .A(u2__abc_44228_n4762), .B(u2__abc_44228_n4764), .Y(u2__abc_44228_n4765) );
  OR2X2 OR2X2_762 ( .A(u2__abc_44228_n4788_1), .B(u2__abc_44228_n4790), .Y(u2__abc_44228_n4791) );
  OR2X2 OR2X2_763 ( .A(u2__abc_44228_n4802), .B(u2__abc_44228_n4804), .Y(u2__abc_44228_n4805) );
  OR2X2 OR2X2_764 ( .A(u2__abc_44228_n4817), .B(u2__abc_44228_n4819), .Y(u2__abc_44228_n4820) );
  OR2X2 OR2X2_765 ( .A(u2__abc_44228_n4831), .B(u2__abc_44228_n4833), .Y(u2__abc_44228_n4834) );
  OR2X2 OR2X2_766 ( .A(u2__abc_44228_n4847), .B(u2__abc_44228_n4849), .Y(u2__abc_44228_n4850) );
  OR2X2 OR2X2_767 ( .A(u2__abc_44228_n4861), .B(u2__abc_44228_n4863), .Y(u2__abc_44228_n4864_1) );
  OR2X2 OR2X2_768 ( .A(u2__abc_44228_n4876), .B(u2__abc_44228_n4878), .Y(u2__abc_44228_n4879) );
  OR2X2 OR2X2_769 ( .A(u2__abc_44228_n4890), .B(u2__abc_44228_n4892_1), .Y(u2__abc_44228_n4893) );
  OR2X2 OR2X2_77 ( .A(aNan_bF_buf4), .B(sqrto_114_), .Y(_abc_64468_n944) );
  OR2X2 OR2X2_770 ( .A(u2__abc_44228_n4907), .B(u2__abc_44228_n4909), .Y(u2__abc_44228_n4910) );
  OR2X2 OR2X2_771 ( .A(u2__abc_44228_n4914), .B(u2__abc_44228_n4916), .Y(u2__abc_44228_n4917) );
  OR2X2 OR2X2_772 ( .A(u2__abc_44228_n4936), .B(u2__abc_44228_n4938), .Y(u2__abc_44228_n4939_1) );
  OR2X2 OR2X2_773 ( .A(u2__abc_44228_n4943), .B(u2__abc_44228_n4945), .Y(u2__abc_44228_n4946) );
  OR2X2 OR2X2_774 ( .A(u2__abc_44228_n4966), .B(u2__abc_44228_n4968), .Y(u2__abc_44228_n4969) );
  OR2X2 OR2X2_775 ( .A(u2__abc_44228_n4973), .B(u2__abc_44228_n4975), .Y(u2__abc_44228_n4976_1) );
  OR2X2 OR2X2_776 ( .A(u2__abc_44228_n4995), .B(u2__abc_44228_n4997), .Y(u2__abc_44228_n4998) );
  OR2X2 OR2X2_777 ( .A(u2__abc_44228_n5002), .B(u2__abc_44228_n5004), .Y(u2__abc_44228_n5005_1) );
  OR2X2 OR2X2_778 ( .A(u2__abc_44228_n5027), .B(u2__abc_44228_n5029), .Y(u2__abc_44228_n5030) );
  OR2X2 OR2X2_779 ( .A(u2__abc_44228_n5041), .B(u2__abc_44228_n5043), .Y(u2__abc_44228_n5044) );
  OR2X2 OR2X2_78 ( .A(_abc_64468_n753_bF_buf11), .B(\a[38] ), .Y(_abc_64468_n945) );
  OR2X2 OR2X2_780 ( .A(u2__abc_44228_n5056), .B(u2__abc_44228_n5058), .Y(u2__abc_44228_n5059) );
  OR2X2 OR2X2_781 ( .A(u2__abc_44228_n5063), .B(u2__abc_44228_n5065), .Y(u2__abc_44228_n5066) );
  OR2X2 OR2X2_782 ( .A(u2__abc_44228_n5086), .B(u2__abc_44228_n5088), .Y(u2__abc_44228_n5089_1) );
  OR2X2 OR2X2_783 ( .A(u2__abc_44228_n5093), .B(u2__abc_44228_n5095), .Y(u2__abc_44228_n5096) );
  OR2X2 OR2X2_784 ( .A(u2__abc_44228_n5115), .B(u2__abc_44228_n5117), .Y(u2__abc_44228_n5118_1) );
  OR2X2 OR2X2_785 ( .A(u2__abc_44228_n5129), .B(u2__abc_44228_n5131), .Y(u2__abc_44228_n5132) );
  OR2X2 OR2X2_786 ( .A(u2__abc_44228_n5146_1), .B(u2__abc_44228_n5148), .Y(u2__abc_44228_n5149) );
  OR2X2 OR2X2_787 ( .A(u2__abc_44228_n5160), .B(u2__abc_44228_n5162), .Y(u2__abc_44228_n5163) );
  OR2X2 OR2X2_788 ( .A(u2__abc_44228_n5175), .B(u2__abc_44228_n5177), .Y(u2__abc_44228_n5178) );
  OR2X2 OR2X2_789 ( .A(u2__abc_44228_n5189), .B(u2__abc_44228_n5191), .Y(u2__abc_44228_n5192_1) );
  OR2X2 OR2X2_79 ( .A(aNan_bF_buf3), .B(sqrto_115_), .Y(_abc_64468_n947) );
  OR2X2 OR2X2_790 ( .A(u2__abc_44228_n5205), .B(u2__abc_44228_n5207), .Y(u2__abc_44228_n5208) );
  OR2X2 OR2X2_791 ( .A(u2__abc_44228_n5219), .B(u2__abc_44228_n5221_1), .Y(u2__abc_44228_n5222) );
  OR2X2 OR2X2_792 ( .A(u2__abc_44228_n5226), .B(sqrto_129_), .Y(u2__abc_44228_n5227) );
  OR2X2 OR2X2_793 ( .A(u2__abc_44228_n5228), .B(u2_remHi_129_), .Y(u2__abc_44228_n5229) );
  OR2X2 OR2X2_794 ( .A(u2__abc_44228_n5231), .B(sqrto_128_), .Y(u2__abc_44228_n5232) );
  OR2X2 OR2X2_795 ( .A(u2__abc_44228_n5233), .B(u2_remHi_128_), .Y(u2__abc_44228_n5234) );
  OR2X2 OR2X2_796 ( .A(u2__abc_44228_n5245), .B(u2__abc_44228_n5247), .Y(u2__abc_44228_n5248) );
  OR2X2 OR2X2_797 ( .A(u2__abc_44228_n5238), .B(u2__abc_44228_n5245), .Y(u2__abc_44228_n5258) );
  OR2X2 OR2X2_798 ( .A(u2__abc_44228_n5263), .B(u2__abc_44228_n5261), .Y(u2__abc_44228_n5264) );
  OR2X2 OR2X2_799 ( .A(u2__abc_44228_n5260_1), .B(u2__abc_44228_n5264), .Y(u2__abc_44228_n5265) );
  OR2X2 OR2X2_8 ( .A(_abc_64468_n753_bF_buf4), .B(\a[3] ), .Y(_abc_64468_n840_1) );
  OR2X2 OR2X2_80 ( .A(_abc_64468_n753_bF_buf10), .B(\a[39] ), .Y(_abc_64468_n948) );
  OR2X2 OR2X2_800 ( .A(u2__abc_44228_n5212), .B(u2__abc_44228_n5219), .Y(u2__abc_44228_n5267) );
  OR2X2 OR2X2_801 ( .A(u2__abc_44228_n5270), .B(u2__abc_44228_n5198), .Y(u2__abc_44228_n5271) );
  OR2X2 OR2X2_802 ( .A(u2__abc_44228_n5269_1), .B(u2__abc_44228_n5271), .Y(u2__abc_44228_n5272) );
  OR2X2 OR2X2_803 ( .A(u2__abc_44228_n5266), .B(u2__abc_44228_n5272), .Y(u2__abc_44228_n5273) );
  OR2X2 OR2X2_804 ( .A(u2__abc_44228_n5168), .B(u2__abc_44228_n5175), .Y(u2__abc_44228_n5275) );
  OR2X2 OR2X2_805 ( .A(u2__abc_44228_n5182_1), .B(u2__abc_44228_n5189), .Y(u2__abc_44228_n5278_1) );
  OR2X2 OR2X2_806 ( .A(u2__abc_44228_n5277), .B(u2__abc_44228_n5279), .Y(u2__abc_44228_n5280) );
  OR2X2 OR2X2_807 ( .A(u2__abc_44228_n5139), .B(u2__abc_44228_n5146_1), .Y(u2__abc_44228_n5287_1) );
  OR2X2 OR2X2_808 ( .A(u2__abc_44228_n5286), .B(u2__abc_44228_n5288), .Y(u2__abc_44228_n5289) );
  OR2X2 OR2X2_809 ( .A(u2__abc_44228_n5281), .B(u2__abc_44228_n5289), .Y(u2__abc_44228_n5290) );
  OR2X2 OR2X2_81 ( .A(aNan_bF_buf2), .B(sqrto_116_), .Y(_abc_64468_n950) );
  OR2X2 OR2X2_810 ( .A(u2__abc_44228_n5274), .B(u2__abc_44228_n5290), .Y(u2__abc_44228_n5291) );
  OR2X2 OR2X2_811 ( .A(u2__abc_44228_n5122), .B(u2__abc_44228_n5129), .Y(u2__abc_44228_n5293) );
  OR2X2 OR2X2_812 ( .A(u2__abc_44228_n5295), .B(u2__abc_44228_n5299), .Y(u2__abc_44228_n5300) );
  OR2X2 OR2X2_813 ( .A(u2__abc_44228_n5307), .B(u2__abc_44228_n5079), .Y(u2__abc_44228_n5308) );
  OR2X2 OR2X2_814 ( .A(u2__abc_44228_n5306_1), .B(u2__abc_44228_n5308), .Y(u2__abc_44228_n5309) );
  OR2X2 OR2X2_815 ( .A(u2__abc_44228_n5301), .B(u2__abc_44228_n5309), .Y(u2__abc_44228_n5310) );
  OR2X2 OR2X2_816 ( .A(u2__abc_44228_n5049), .B(u2__abc_44228_n5056), .Y(u2__abc_44228_n5312) );
  OR2X2 OR2X2_817 ( .A(u2__abc_44228_n5318), .B(u2__abc_44228_n5313), .Y(u2__abc_44228_n5319) );
  OR2X2 OR2X2_818 ( .A(u2__abc_44228_n5321), .B(u2__abc_44228_n5020), .Y(u2__abc_44228_n5322) );
  OR2X2 OR2X2_819 ( .A(u2__abc_44228_n5323), .B(u2__abc_44228_n5037), .Y(u2__abc_44228_n5324_1) );
  OR2X2 OR2X2_82 ( .A(_abc_64468_n753_bF_buf9), .B(\a[40] ), .Y(_abc_64468_n951) );
  OR2X2 OR2X2_820 ( .A(u2__abc_44228_n5327), .B(u2__abc_44228_n5322), .Y(u2__abc_44228_n5328) );
  OR2X2 OR2X2_821 ( .A(u2__abc_44228_n5320), .B(u2__abc_44228_n5328), .Y(u2__abc_44228_n5329) );
  OR2X2 OR2X2_822 ( .A(u2__abc_44228_n5311), .B(u2__abc_44228_n5329), .Y(u2__abc_44228_n5330) );
  OR2X2 OR2X2_823 ( .A(u2__abc_44228_n5292), .B(u2__abc_44228_n5330), .Y(u2__abc_44228_n5331) );
  OR2X2 OR2X2_824 ( .A(u2__abc_44228_n5002), .B(u2__abc_44228_n5008), .Y(u2__abc_44228_n5333_1) );
  OR2X2 OR2X2_825 ( .A(u2__abc_44228_n5336), .B(u2__abc_44228_n4988), .Y(u2__abc_44228_n5337) );
  OR2X2 OR2X2_826 ( .A(u2__abc_44228_n5335), .B(u2__abc_44228_n5337), .Y(u2__abc_44228_n5338) );
  OR2X2 OR2X2_827 ( .A(u2__abc_44228_n5345), .B(u2__abc_44228_n4959), .Y(u2__abc_44228_n5346) );
  OR2X2 OR2X2_828 ( .A(u2__abc_44228_n5344), .B(u2__abc_44228_n5346), .Y(u2__abc_44228_n5347) );
  OR2X2 OR2X2_829 ( .A(u2__abc_44228_n5339), .B(u2__abc_44228_n5347), .Y(u2__abc_44228_n5348) );
  OR2X2 OR2X2_83 ( .A(aNan_bF_buf1), .B(sqrto_117_), .Y(_abc_64468_n953) );
  OR2X2 OR2X2_830 ( .A(u2__abc_44228_n4929), .B(u2__abc_44228_n4936), .Y(u2__abc_44228_n5350) );
  OR2X2 OR2X2_831 ( .A(u2__abc_44228_n5356), .B(u2__abc_44228_n5351), .Y(u2__abc_44228_n5357) );
  OR2X2 OR2X2_832 ( .A(u2__abc_44228_n5364), .B(u2__abc_44228_n4900), .Y(u2__abc_44228_n5365) );
  OR2X2 OR2X2_833 ( .A(u2__abc_44228_n5363), .B(u2__abc_44228_n5365), .Y(u2__abc_44228_n5366) );
  OR2X2 OR2X2_834 ( .A(u2__abc_44228_n5358), .B(u2__abc_44228_n5366), .Y(u2__abc_44228_n5367) );
  OR2X2 OR2X2_835 ( .A(u2__abc_44228_n5349), .B(u2__abc_44228_n5367), .Y(u2__abc_44228_n5368) );
  OR2X2 OR2X2_836 ( .A(u2__abc_44228_n5370), .B(u2__abc_44228_n4886), .Y(u2__abc_44228_n5371) );
  OR2X2 OR2X2_837 ( .A(u2__abc_44228_n5375), .B(u2__abc_44228_n4869), .Y(u2__abc_44228_n5376) );
  OR2X2 OR2X2_838 ( .A(u2__abc_44228_n5374), .B(u2__abc_44228_n5376), .Y(u2__abc_44228_n5377) );
  OR2X2 OR2X2_839 ( .A(u2__abc_44228_n5379), .B(u2__abc_44228_n4857), .Y(u2__abc_44228_n5380) );
  OR2X2 OR2X2_84 ( .A(_abc_64468_n753_bF_buf8), .B(\a[41] ), .Y(_abc_64468_n954) );
  OR2X2 OR2X2_840 ( .A(u2__abc_44228_n5384), .B(u2__abc_44228_n4840), .Y(u2__abc_44228_n5385) );
  OR2X2 OR2X2_841 ( .A(u2__abc_44228_n5383), .B(u2__abc_44228_n5385), .Y(u2__abc_44228_n5386) );
  OR2X2 OR2X2_842 ( .A(u2__abc_44228_n5378), .B(u2__abc_44228_n5386), .Y(u2__abc_44228_n5387) );
  OR2X2 OR2X2_843 ( .A(u2__abc_44228_n5389), .B(u2__abc_44228_n4798), .Y(u2__abc_44228_n5390_1) );
  OR2X2 OR2X2_844 ( .A(u2__abc_44228_n5394), .B(u2__abc_44228_n4781), .Y(u2__abc_44228_n5395) );
  OR2X2 OR2X2_845 ( .A(u2__abc_44228_n5393), .B(u2__abc_44228_n5395), .Y(u2__abc_44228_n5396) );
  OR2X2 OR2X2_846 ( .A(u2__abc_44228_n5397), .B(u2__abc_44228_n4813), .Y(u2__abc_44228_n5398) );
  OR2X2 OR2X2_847 ( .A(u2__abc_44228_n5401), .B(u2__abc_44228_n5405), .Y(u2__abc_44228_n5406) );
  OR2X2 OR2X2_848 ( .A(u2__abc_44228_n5407), .B(u2__abc_44228_n5396), .Y(u2__abc_44228_n5408) );
  OR2X2 OR2X2_849 ( .A(u2__abc_44228_n5388), .B(u2__abc_44228_n5408), .Y(u2__abc_44228_n5409) );
  OR2X2 OR2X2_85 ( .A(aNan_bF_buf0), .B(sqrto_118_), .Y(_abc_64468_n956) );
  OR2X2 OR2X2_850 ( .A(u2__abc_44228_n5369), .B(u2__abc_44228_n5409), .Y(u2__abc_44228_n5410_1) );
  OR2X2 OR2X2_851 ( .A(u2__abc_44228_n5332), .B(u2__abc_44228_n5410_1), .Y(u2__abc_44228_n5411) );
  OR2X2 OR2X2_852 ( .A(u2__abc_44228_n4762), .B(u2__abc_44228_n4768), .Y(u2__abc_44228_n5413) );
  OR2X2 OR2X2_853 ( .A(u2__abc_44228_n5416), .B(u2__abc_44228_n4748), .Y(u2__abc_44228_n5417) );
  OR2X2 OR2X2_854 ( .A(u2__abc_44228_n5415), .B(u2__abc_44228_n5417), .Y(u2__abc_44228_n5418) );
  OR2X2 OR2X2_855 ( .A(u2__abc_44228_n5420), .B(u2__abc_44228_n4736), .Y(u2__abc_44228_n5421) );
  OR2X2 OR2X2_856 ( .A(u2__abc_44228_n5425), .B(u2__abc_44228_n4719), .Y(u2__abc_44228_n5426) );
  OR2X2 OR2X2_857 ( .A(u2__abc_44228_n5424), .B(u2__abc_44228_n5426), .Y(u2__abc_44228_n5427) );
  OR2X2 OR2X2_858 ( .A(u2__abc_44228_n5419_1), .B(u2__abc_44228_n5427), .Y(u2__abc_44228_n5428_1) );
  OR2X2 OR2X2_859 ( .A(u2__abc_44228_n5435), .B(u2__abc_44228_n4689), .Y(u2__abc_44228_n5436) );
  OR2X2 OR2X2_86 ( .A(_abc_64468_n753_bF_buf7), .B(\a[42] ), .Y(_abc_64468_n957) );
  OR2X2 OR2X2_860 ( .A(u2__abc_44228_n5434), .B(u2__abc_44228_n5436), .Y(u2__abc_44228_n5437_1) );
  OR2X2 OR2X2_861 ( .A(u2__abc_44228_n5439), .B(u2__abc_44228_n4677), .Y(u2__abc_44228_n5440) );
  OR2X2 OR2X2_862 ( .A(u2__abc_44228_n5444), .B(u2__abc_44228_n4660), .Y(u2__abc_44228_n5445) );
  OR2X2 OR2X2_863 ( .A(u2__abc_44228_n5443), .B(u2__abc_44228_n5445), .Y(u2__abc_44228_n5446) );
  OR2X2 OR2X2_864 ( .A(u2__abc_44228_n5438), .B(u2__abc_44228_n5446), .Y(u2__abc_44228_n5447_1) );
  OR2X2 OR2X2_865 ( .A(u2__abc_44228_n5429), .B(u2__abc_44228_n5447_1), .Y(u2__abc_44228_n5448) );
  OR2X2 OR2X2_866 ( .A(u2__abc_44228_n5450), .B(u2__abc_44228_n4646_1), .Y(u2__abc_44228_n5451) );
  OR2X2 OR2X2_867 ( .A(u2__abc_44228_n5455), .B(u2__abc_44228_n4629_1), .Y(u2__abc_44228_n5456_1) );
  OR2X2 OR2X2_868 ( .A(u2__abc_44228_n5454), .B(u2__abc_44228_n5456_1), .Y(u2__abc_44228_n5457) );
  OR2X2 OR2X2_869 ( .A(u2__abc_44228_n5464), .B(u2__abc_44228_n4600_1), .Y(u2__abc_44228_n5465_1) );
  OR2X2 OR2X2_87 ( .A(aNan_bF_buf10), .B(sqrto_119_), .Y(_abc_64468_n959) );
  OR2X2 OR2X2_870 ( .A(u2__abc_44228_n5463), .B(u2__abc_44228_n5465_1), .Y(u2__abc_44228_n5466) );
  OR2X2 OR2X2_871 ( .A(u2__abc_44228_n5458), .B(u2__abc_44228_n5466), .Y(u2__abc_44228_n5467) );
  OR2X2 OR2X2_872 ( .A(u2__abc_44228_n5474_1), .B(u2__abc_44228_n4570), .Y(u2__abc_44228_n5475) );
  OR2X2 OR2X2_873 ( .A(u2__abc_44228_n5473), .B(u2__abc_44228_n5475), .Y(u2__abc_44228_n5476) );
  OR2X2 OR2X2_874 ( .A(u2__abc_44228_n5478), .B(u2__abc_44228_n4541), .Y(u2__abc_44228_n5479) );
  OR2X2 OR2X2_875 ( .A(u2__abc_44228_n5484), .B(u2__abc_44228_n5479), .Y(u2__abc_44228_n5485) );
  OR2X2 OR2X2_876 ( .A(u2__abc_44228_n5477), .B(u2__abc_44228_n5485), .Y(u2__abc_44228_n5486) );
  OR2X2 OR2X2_877 ( .A(u2__abc_44228_n5468), .B(u2__abc_44228_n5486), .Y(u2__abc_44228_n5487) );
  OR2X2 OR2X2_878 ( .A(u2__abc_44228_n5449), .B(u2__abc_44228_n5487), .Y(u2__abc_44228_n5488) );
  OR2X2 OR2X2_879 ( .A(u2__abc_44228_n5490), .B(u2__abc_44228_n4532), .Y(u2__abc_44228_n5491) );
  OR2X2 OR2X2_88 ( .A(_abc_64468_n753_bF_buf6), .B(\a[43] ), .Y(_abc_64468_n960) );
  OR2X2 OR2X2_880 ( .A(u2__abc_44228_n5495), .B(u2__abc_44228_n4509), .Y(u2__abc_44228_n5496) );
  OR2X2 OR2X2_881 ( .A(u2__abc_44228_n5494), .B(u2__abc_44228_n5496), .Y(u2__abc_44228_n5497) );
  OR2X2 OR2X2_882 ( .A(u2__abc_44228_n5504), .B(u2__abc_44228_n4480_1), .Y(u2__abc_44228_n5505) );
  OR2X2 OR2X2_883 ( .A(u2__abc_44228_n5503), .B(u2__abc_44228_n5505), .Y(u2__abc_44228_n5506) );
  OR2X2 OR2X2_884 ( .A(u2__abc_44228_n5498), .B(u2__abc_44228_n5506), .Y(u2__abc_44228_n5507) );
  OR2X2 OR2X2_885 ( .A(u2__abc_44228_n5509), .B(u2__abc_44228_n4453), .Y(u2__abc_44228_n5510) );
  OR2X2 OR2X2_886 ( .A(u2__abc_44228_n5513), .B(u2__abc_44228_n5517), .Y(u2__abc_44228_n5518) );
  OR2X2 OR2X2_887 ( .A(u2__abc_44228_n5525), .B(u2__abc_44228_n4421), .Y(u2__abc_44228_n5526) );
  OR2X2 OR2X2_888 ( .A(u2__abc_44228_n5524), .B(u2__abc_44228_n5526), .Y(u2__abc_44228_n5527) );
  OR2X2 OR2X2_889 ( .A(u2__abc_44228_n5519), .B(u2__abc_44228_n5527), .Y(u2__abc_44228_n5528) );
  OR2X2 OR2X2_89 ( .A(aNan_bF_buf9), .B(sqrto_120_), .Y(_abc_64468_n962) );
  OR2X2 OR2X2_890 ( .A(u2__abc_44228_n5508), .B(u2__abc_44228_n5528), .Y(u2__abc_44228_n5529) );
  OR2X2 OR2X2_891 ( .A(u2__abc_44228_n5536), .B(u2__abc_44228_n4331), .Y(u2__abc_44228_n5537) );
  OR2X2 OR2X2_892 ( .A(u2__abc_44228_n5535), .B(u2__abc_44228_n5537), .Y(u2__abc_44228_n5538) );
  OR2X2 OR2X2_893 ( .A(u2__abc_44228_n4302), .B(u2__abc_44228_n4309), .Y(u2__abc_44228_n5540_1) );
  OR2X2 OR2X2_894 ( .A(u2__abc_44228_n5546), .B(u2__abc_44228_n5541), .Y(u2__abc_44228_n5547) );
  OR2X2 OR2X2_895 ( .A(u2__abc_44228_n5539), .B(u2__abc_44228_n5547), .Y(u2__abc_44228_n5548) );
  OR2X2 OR2X2_896 ( .A(u2__abc_44228_n5554), .B(u2__abc_44228_n4390), .Y(u2__abc_44228_n5555) );
  OR2X2 OR2X2_897 ( .A(u2__abc_44228_n5553), .B(u2__abc_44228_n5555), .Y(u2__abc_44228_n5556) );
  OR2X2 OR2X2_898 ( .A(u2__abc_44228_n5563), .B(u2__abc_44228_n4361), .Y(u2__abc_44228_n5564) );
  OR2X2 OR2X2_899 ( .A(u2__abc_44228_n5562), .B(u2__abc_44228_n5564), .Y(u2__abc_44228_n5565) );
  OR2X2 OR2X2_9 ( .A(aNan_bF_buf5), .B(sqrto_80_), .Y(_abc_64468_n842) );
  OR2X2 OR2X2_90 ( .A(_abc_64468_n753_bF_buf5), .B(\a[44] ), .Y(_abc_64468_n963) );
  OR2X2 OR2X2_900 ( .A(u2__abc_44228_n5557), .B(u2__abc_44228_n5565), .Y(u2__abc_44228_n5566) );
  OR2X2 OR2X2_901 ( .A(u2__abc_44228_n5567), .B(u2__abc_44228_n5548), .Y(u2__abc_44228_n5568_1) );
  OR2X2 OR2X2_902 ( .A(u2__abc_44228_n5530), .B(u2__abc_44228_n5568_1), .Y(u2__abc_44228_n5569) );
  OR2X2 OR2X2_903 ( .A(u2__abc_44228_n5489), .B(u2__abc_44228_n5569), .Y(u2__abc_44228_n5570) );
  OR2X2 OR2X2_904 ( .A(u2__abc_44228_n5412), .B(u2__abc_44228_n5570), .Y(u2__abc_44228_n5571) );
  OR2X2 OR2X2_905 ( .A(u2__abc_44228_n5257), .B(u2__abc_44228_n5571), .Y(u2__abc_44228_n5572) );
  OR2X2 OR2X2_906 ( .A(u2__abc_44228_n5581), .B(u2__abc_44228_n5583), .Y(u2__abc_44228_n5584) );
  OR2X2 OR2X2_907 ( .A(u2__abc_44228_n5595), .B(u2__abc_44228_n5597_1), .Y(u2__abc_44228_n5598) );
  OR2X2 OR2X2_908 ( .A(u2__abc_44228_n5610), .B(u2__abc_44228_n5612), .Y(u2__abc_44228_n5613) );
  OR2X2 OR2X2_909 ( .A(u2__abc_44228_n5624_1), .B(u2__abc_44228_n5626), .Y(u2__abc_44228_n5627) );
  OR2X2 OR2X2_91 ( .A(aNan_bF_buf8), .B(sqrto_121_), .Y(_abc_64468_n965) );
  OR2X2 OR2X2_910 ( .A(u2__abc_44228_n5640), .B(u2__abc_44228_n5642), .Y(u2__abc_44228_n5643_1) );
  OR2X2 OR2X2_911 ( .A(u2__abc_44228_n5647), .B(u2__abc_44228_n5649), .Y(u2__abc_44228_n5650) );
  OR2X2 OR2X2_912 ( .A(u2__abc_44228_n5669), .B(u2__abc_44228_n5671), .Y(u2__abc_44228_n5672_1) );
  OR2X2 OR2X2_913 ( .A(u2__abc_44228_n5683), .B(u2__abc_44228_n5685), .Y(u2__abc_44228_n5686) );
  OR2X2 OR2X2_914 ( .A(u2__abc_44228_n5700_1), .B(u2__abc_44228_n5702), .Y(u2__abc_44228_n5703) );
  OR2X2 OR2X2_915 ( .A(u2__abc_44228_n5714), .B(u2__abc_44228_n5716), .Y(u2__abc_44228_n5717) );
  OR2X2 OR2X2_916 ( .A(u2__abc_44228_n5729), .B(u2__abc_44228_n5731), .Y(u2__abc_44228_n5732) );
  OR2X2 OR2X2_917 ( .A(u2__abc_44228_n5743), .B(u2__abc_44228_n5745), .Y(u2__abc_44228_n5746) );
  OR2X2 OR2X2_918 ( .A(u2__abc_44228_n5759), .B(u2__abc_44228_n5761), .Y(u2__abc_44228_n5762) );
  OR2X2 OR2X2_919 ( .A(u2__abc_44228_n5766), .B(u2__abc_44228_n5768), .Y(u2__abc_44228_n5769) );
  OR2X2 OR2X2_92 ( .A(_abc_64468_n753_bF_buf4), .B(\a[45] ), .Y(_abc_64468_n966) );
  OR2X2 OR2X2_920 ( .A(u2__abc_44228_n5788), .B(u2__abc_44228_n5790), .Y(u2__abc_44228_n5791) );
  OR2X2 OR2X2_921 ( .A(u2__abc_44228_n5802_1), .B(u2__abc_44228_n5804), .Y(u2__abc_44228_n5805) );
  OR2X2 OR2X2_922 ( .A(u2__abc_44228_n5820), .B(u2__abc_44228_n5822_1), .Y(u2__abc_44228_n5823) );
  OR2X2 OR2X2_923 ( .A(u2__abc_44228_n5827), .B(u2__abc_44228_n5829), .Y(u2__abc_44228_n5830_1) );
  OR2X2 OR2X2_924 ( .A(u2__abc_44228_n5849), .B(u2__abc_44228_n5851), .Y(u2__abc_44228_n5852) );
  OR2X2 OR2X2_925 ( .A(u2__abc_44228_n5863_1), .B(u2__abc_44228_n5865), .Y(u2__abc_44228_n5866) );
  OR2X2 OR2X2_926 ( .A(u2__abc_44228_n5879), .B(u2__abc_44228_n5881), .Y(u2__abc_44228_n5882) );
  OR2X2 OR2X2_927 ( .A(u2__abc_44228_n5886), .B(u2__abc_44228_n5888), .Y(u2__abc_44228_n5889) );
  OR2X2 OR2X2_928 ( .A(u2__abc_44228_n5908), .B(u2__abc_44228_n5910), .Y(u2__abc_44228_n5911_1) );
  OR2X2 OR2X2_929 ( .A(u2__abc_44228_n5922), .B(u2__abc_44228_n5924), .Y(u2__abc_44228_n5925) );
  OR2X2 OR2X2_93 ( .A(aNan_bF_buf7), .B(sqrto_122_), .Y(_abc_64468_n968) );
  OR2X2 OR2X2_930 ( .A(u2__abc_44228_n5939), .B(u2__abc_44228_n5941), .Y(u2__abc_44228_n5942) );
  OR2X2 OR2X2_931 ( .A(u2__abc_44228_n5953), .B(u2__abc_44228_n5955), .Y(u2__abc_44228_n5956) );
  OR2X2 OR2X2_932 ( .A(u2__abc_44228_n5968), .B(u2__abc_44228_n5970), .Y(u2__abc_44228_n5971) );
  OR2X2 OR2X2_933 ( .A(u2__abc_44228_n5982), .B(u2__abc_44228_n5984), .Y(u2__abc_44228_n5985_1) );
  OR2X2 OR2X2_934 ( .A(u2__abc_44228_n5998), .B(u2__abc_44228_n6000), .Y(u2__abc_44228_n6001) );
  OR2X2 OR2X2_935 ( .A(u2__abc_44228_n6005), .B(u2__abc_44228_n6007), .Y(u2__abc_44228_n6008) );
  OR2X2 OR2X2_936 ( .A(u2__abc_44228_n6027), .B(u2__abc_44228_n6029), .Y(u2__abc_44228_n6030) );
  OR2X2 OR2X2_937 ( .A(u2__abc_44228_n6034), .B(u2__abc_44228_n6036), .Y(u2__abc_44228_n6037) );
  OR2X2 OR2X2_938 ( .A(u2__abc_44228_n6060), .B(u2__abc_44228_n6062), .Y(u2__abc_44228_n6063) );
  OR2X2 OR2X2_939 ( .A(u2__abc_44228_n6074), .B(u2__abc_44228_n6076), .Y(u2__abc_44228_n6077) );
  OR2X2 OR2X2_94 ( .A(_abc_64468_n753_bF_buf3), .B(\a[46] ), .Y(_abc_64468_n969) );
  OR2X2 OR2X2_940 ( .A(u2__abc_44228_n6089), .B(u2__abc_44228_n6091), .Y(u2__abc_44228_n6092) );
  OR2X2 OR2X2_941 ( .A(u2__abc_44228_n6103), .B(u2__abc_44228_n6105), .Y(u2__abc_44228_n6106) );
  OR2X2 OR2X2_942 ( .A(u2__abc_44228_n6119), .B(u2__abc_44228_n6121), .Y(u2__abc_44228_n6122_1) );
  OR2X2 OR2X2_943 ( .A(u2__abc_44228_n6126), .B(u2__abc_44228_n6128), .Y(u2__abc_44228_n6129) );
  OR2X2 OR2X2_944 ( .A(u2__abc_44228_n6148), .B(u2__abc_44228_n6150), .Y(u2__abc_44228_n6151_1) );
  OR2X2 OR2X2_945 ( .A(u2__abc_44228_n6155), .B(u2__abc_44228_n6157), .Y(u2__abc_44228_n6158) );
  OR2X2 OR2X2_946 ( .A(u2__abc_44228_n6179), .B(u2__abc_44228_n6181), .Y(u2__abc_44228_n6182) );
  OR2X2 OR2X2_947 ( .A(u2__abc_44228_n6193), .B(u2__abc_44228_n6195), .Y(u2__abc_44228_n6196_1) );
  OR2X2 OR2X2_948 ( .A(u2__abc_44228_n6208), .B(u2__abc_44228_n6210), .Y(u2__abc_44228_n6211) );
  OR2X2 OR2X2_949 ( .A(u2__abc_44228_n6222), .B(u2__abc_44228_n6224_1), .Y(u2__abc_44228_n6225) );
  OR2X2 OR2X2_95 ( .A(aNan_bF_buf6), .B(sqrto_123_), .Y(_abc_64468_n971) );
  OR2X2 OR2X2_950 ( .A(u2__abc_44228_n6238), .B(u2__abc_44228_n6240), .Y(u2__abc_44228_n6241) );
  OR2X2 OR2X2_951 ( .A(u2__abc_44228_n6252), .B(u2__abc_44228_n6254), .Y(u2__abc_44228_n6255) );
  OR2X2 OR2X2_952 ( .A(u2__abc_44228_n6267), .B(u2__abc_44228_n6269_1), .Y(u2__abc_44228_n6270) );
  OR2X2 OR2X2_953 ( .A(u2__abc_44228_n6281), .B(u2__abc_44228_n6283), .Y(u2__abc_44228_n6284) );
  OR2X2 OR2X2_954 ( .A(u2__abc_44228_n6299), .B(u2__abc_44228_n6301), .Y(u2__abc_44228_n6302) );
  OR2X2 OR2X2_955 ( .A(u2__abc_44228_n6313), .B(u2__abc_44228_n6315_1), .Y(u2__abc_44228_n6316) );
  OR2X2 OR2X2_956 ( .A(u2__abc_44228_n6328), .B(u2__abc_44228_n6330), .Y(u2__abc_44228_n6331) );
  OR2X2 OR2X2_957 ( .A(u2__abc_44228_n6342_1), .B(u2__abc_44228_n6344), .Y(u2__abc_44228_n6345) );
  OR2X2 OR2X2_958 ( .A(u2__abc_44228_n6358), .B(u2__abc_44228_n6360), .Y(u2__abc_44228_n6361_1) );
  OR2X2 OR2X2_959 ( .A(u2__abc_44228_n6372), .B(u2__abc_44228_n6374), .Y(u2__abc_44228_n6375) );
  OR2X2 OR2X2_96 ( .A(_abc_64468_n753_bF_buf2), .B(\a[47] ), .Y(_abc_64468_n972) );
  OR2X2 OR2X2_960 ( .A(u2__abc_44228_n6387), .B(u2__abc_44228_n6389_1), .Y(u2__abc_44228_n6390) );
  OR2X2 OR2X2_961 ( .A(u2__abc_44228_n6394), .B(u2__abc_44228_n6396), .Y(u2__abc_44228_n6397_1) );
  OR2X2 OR2X2_962 ( .A(u2__abc_44228_n6418), .B(u2__abc_44228_n6420), .Y(u2__abc_44228_n6421) );
  OR2X2 OR2X2_963 ( .A(u2__abc_44228_n6432), .B(u2__abc_44228_n6434), .Y(u2__abc_44228_n6435_1) );
  OR2X2 OR2X2_964 ( .A(u2__abc_44228_n6447), .B(u2__abc_44228_n6449), .Y(u2__abc_44228_n6450) );
  OR2X2 OR2X2_965 ( .A(u2__abc_44228_n6461), .B(u2__abc_44228_n6463_1), .Y(u2__abc_44228_n6464) );
  OR2X2 OR2X2_966 ( .A(u2__abc_44228_n6477), .B(u2__abc_44228_n6479), .Y(u2__abc_44228_n6480_1) );
  OR2X2 OR2X2_967 ( .A(u2__abc_44228_n6491), .B(u2__abc_44228_n6493), .Y(u2__abc_44228_n6494) );
  OR2X2 OR2X2_968 ( .A(u2__abc_44228_n6506), .B(u2__abc_44228_n6508), .Y(u2__abc_44228_n6509) );
  OR2X2 OR2X2_969 ( .A(u2__abc_44228_n6520), .B(u2__abc_44228_n6522), .Y(u2__abc_44228_n6523) );
  OR2X2 OR2X2_97 ( .A(aNan_bF_buf5), .B(sqrto_124_), .Y(_abc_64468_n974) );
  OR2X2 OR2X2_970 ( .A(u2__abc_44228_n6533), .B(u2__abc_44228_n6516), .Y(u2__abc_44228_n6534) );
  OR2X2 OR2X2_971 ( .A(u2__abc_44228_n6538), .B(u2__abc_44228_n6499_1), .Y(u2__abc_44228_n6539) );
  OR2X2 OR2X2_972 ( .A(u2__abc_44228_n6537), .B(u2__abc_44228_n6539), .Y(u2__abc_44228_n6540) );
  OR2X2 OR2X2_973 ( .A(u2__abc_44228_n6542), .B(u2__abc_44228_n6487), .Y(u2__abc_44228_n6543_1) );
  OR2X2 OR2X2_974 ( .A(u2__abc_44228_n6547), .B(u2__abc_44228_n6470), .Y(u2__abc_44228_n6548) );
  OR2X2 OR2X2_975 ( .A(u2__abc_44228_n6546), .B(u2__abc_44228_n6548), .Y(u2__abc_44228_n6549) );
  OR2X2 OR2X2_976 ( .A(u2__abc_44228_n6541), .B(u2__abc_44228_n6549), .Y(u2__abc_44228_n6550) );
  OR2X2 OR2X2_977 ( .A(u2__abc_44228_n6440), .B(u2__abc_44228_n6447), .Y(u2__abc_44228_n6552_1) );
  OR2X2 OR2X2_978 ( .A(u2__abc_44228_n6558), .B(u2__abc_44228_n6553), .Y(u2__abc_44228_n6559) );
  OR2X2 OR2X2_979 ( .A(u2__abc_44228_n6561_1), .B(u2__abc_44228_n6428), .Y(u2__abc_44228_n6562) );
  OR2X2 OR2X2_98 ( .A(_abc_64468_n753_bF_buf1), .B(\a[48] ), .Y(_abc_64468_n975) );
  OR2X2 OR2X2_980 ( .A(u2__abc_44228_n6566), .B(u2__abc_44228_n6411), .Y(u2__abc_44228_n6567) );
  OR2X2 OR2X2_981 ( .A(u2__abc_44228_n6565), .B(u2__abc_44228_n6567), .Y(u2__abc_44228_n6568) );
  OR2X2 OR2X2_982 ( .A(u2__abc_44228_n6560), .B(u2__abc_44228_n6568), .Y(u2__abc_44228_n6569) );
  OR2X2 OR2X2_983 ( .A(u2__abc_44228_n6551), .B(u2__abc_44228_n6569), .Y(u2__abc_44228_n6570) );
  OR2X2 OR2X2_984 ( .A(u2__abc_44228_n6577), .B(u2__abc_44228_n6380), .Y(u2__abc_44228_n6578) );
  OR2X2 OR2X2_985 ( .A(u2__abc_44228_n6576), .B(u2__abc_44228_n6578), .Y(u2__abc_44228_n6579_1) );
  OR2X2 OR2X2_986 ( .A(u2__abc_44228_n6581), .B(u2__abc_44228_n6368), .Y(u2__abc_44228_n6582) );
  OR2X2 OR2X2_987 ( .A(u2__abc_44228_n6586), .B(u2__abc_44228_n6351), .Y(u2__abc_44228_n6587) );
  OR2X2 OR2X2_988 ( .A(u2__abc_44228_n6585), .B(u2__abc_44228_n6587), .Y(u2__abc_44228_n6588_1) );
  OR2X2 OR2X2_989 ( .A(u2__abc_44228_n6580), .B(u2__abc_44228_n6588_1), .Y(u2__abc_44228_n6589) );
  OR2X2 OR2X2_99 ( .A(aNan_bF_buf4), .B(sqrto_125_), .Y(_abc_64468_n977) );
  OR2X2 OR2X2_990 ( .A(u2__abc_44228_n6591), .B(u2__abc_44228_n6324_1), .Y(u2__abc_44228_n6592) );
  OR2X2 OR2X2_991 ( .A(u2__abc_44228_n6595), .B(u2__abc_44228_n6599), .Y(u2__abc_44228_n6600) );
  OR2X2 OR2X2_992 ( .A(u2__abc_44228_n6602), .B(u2__abc_44228_n6292), .Y(u2__abc_44228_n6603) );
  OR2X2 OR2X2_993 ( .A(u2__abc_44228_n6608), .B(u2__abc_44228_n6603), .Y(u2__abc_44228_n6609) );
  OR2X2 OR2X2_994 ( .A(u2__abc_44228_n6601), .B(u2__abc_44228_n6609), .Y(u2__abc_44228_n6610) );
  OR2X2 OR2X2_995 ( .A(u2__abc_44228_n6590), .B(u2__abc_44228_n6610), .Y(u2__abc_44228_n6611) );
  OR2X2 OR2X2_996 ( .A(u2__abc_44228_n6571_1), .B(u2__abc_44228_n6611), .Y(u2__abc_44228_n6612) );
  OR2X2 OR2X2_997 ( .A(u2__abc_44228_n6614), .B(u2__abc_44228_n6277), .Y(u2__abc_44228_n6615) );
  OR2X2 OR2X2_998 ( .A(u2__abc_44228_n6619), .B(u2__abc_44228_n6260_1), .Y(u2__abc_44228_n6620) );
  OR2X2 OR2X2_999 ( .A(u2__abc_44228_n6618), .B(u2__abc_44228_n6620), .Y(u2__abc_44228_n6621) );
endmodule
