module siphash(clk, reset_n, cs, we, \addr[0] , \addr[1] , \addr[2] , \addr[3] , \addr[4] , \addr[5] , \addr[6] , \addr[7] , \write_data[0] , \write_data[1] , \write_data[2] , \write_data[3] , \write_data[4] , \write_data[5] , \write_data[6] , \write_data[7] , \write_data[8] , \write_data[9] , \write_data[10] , \write_data[11] , \write_data[12] , \write_data[13] , \write_data[14] , \write_data[15] , \write_data[16] , \write_data[17] , \write_data[18] , \write_data[19] , \write_data[20] , \write_data[21] , \write_data[22] , \write_data[23] , \write_data[24] , \write_data[25] , \write_data[26] , \write_data[27] , \write_data[28] , \write_data[29] , \write_data[30] , \write_data[31] , \read_data[0] , \read_data[1] , \read_data[2] , \read_data[3] , \read_data[4] , \read_data[5] , \read_data[6] , \read_data[7] , \read_data[8] , \read_data[9] , \read_data[10] , \read_data[11] , \read_data[12] , \read_data[13] , \read_data[14] , \read_data[15] , \read_data[16] , \read_data[17] , \read_data[18] , \read_data[19] , \read_data[20] , \read_data[21] , \read_data[22] , \read_data[23] , \read_data[24] , \read_data[25] , \read_data[26] , \read_data[27] , \read_data[28] , \read_data[29] , \read_data[30] , \read_data[31] );

wire _0ctrl_reg_2_0__0_; 
wire _0ctrl_reg_2_0__1_; 
wire _0ctrl_reg_2_0__2_; 
wire _0key0_reg_31_0__0_; 
wire _0key0_reg_31_0__10_; 
wire _0key0_reg_31_0__11_; 
wire _0key0_reg_31_0__12_; 
wire _0key0_reg_31_0__13_; 
wire _0key0_reg_31_0__14_; 
wire _0key0_reg_31_0__15_; 
wire _0key0_reg_31_0__16_; 
wire _0key0_reg_31_0__17_; 
wire _0key0_reg_31_0__18_; 
wire _0key0_reg_31_0__19_; 
wire _0key0_reg_31_0__1_; 
wire _0key0_reg_31_0__20_; 
wire _0key0_reg_31_0__21_; 
wire _0key0_reg_31_0__22_; 
wire _0key0_reg_31_0__23_; 
wire _0key0_reg_31_0__24_; 
wire _0key0_reg_31_0__25_; 
wire _0key0_reg_31_0__26_; 
wire _0key0_reg_31_0__27_; 
wire _0key0_reg_31_0__28_; 
wire _0key0_reg_31_0__29_; 
wire _0key0_reg_31_0__2_; 
wire _0key0_reg_31_0__30_; 
wire _0key0_reg_31_0__31_; 
wire _0key0_reg_31_0__3_; 
wire _0key0_reg_31_0__4_; 
wire _0key0_reg_31_0__5_; 
wire _0key0_reg_31_0__6_; 
wire _0key0_reg_31_0__7_; 
wire _0key0_reg_31_0__8_; 
wire _0key0_reg_31_0__9_; 
wire _0key1_reg_31_0__0_; 
wire _0key1_reg_31_0__10_; 
wire _0key1_reg_31_0__11_; 
wire _0key1_reg_31_0__12_; 
wire _0key1_reg_31_0__13_; 
wire _0key1_reg_31_0__14_; 
wire _0key1_reg_31_0__15_; 
wire _0key1_reg_31_0__16_; 
wire _0key1_reg_31_0__17_; 
wire _0key1_reg_31_0__18_; 
wire _0key1_reg_31_0__19_; 
wire _0key1_reg_31_0__1_; 
wire _0key1_reg_31_0__20_; 
wire _0key1_reg_31_0__21_; 
wire _0key1_reg_31_0__22_; 
wire _0key1_reg_31_0__23_; 
wire _0key1_reg_31_0__24_; 
wire _0key1_reg_31_0__25_; 
wire _0key1_reg_31_0__26_; 
wire _0key1_reg_31_0__27_; 
wire _0key1_reg_31_0__28_; 
wire _0key1_reg_31_0__29_; 
wire _0key1_reg_31_0__2_; 
wire _0key1_reg_31_0__30_; 
wire _0key1_reg_31_0__31_; 
wire _0key1_reg_31_0__3_; 
wire _0key1_reg_31_0__4_; 
wire _0key1_reg_31_0__5_; 
wire _0key1_reg_31_0__6_; 
wire _0key1_reg_31_0__7_; 
wire _0key1_reg_31_0__8_; 
wire _0key1_reg_31_0__9_; 
wire _0key2_reg_31_0__0_; 
wire _0key2_reg_31_0__10_; 
wire _0key2_reg_31_0__11_; 
wire _0key2_reg_31_0__12_; 
wire _0key2_reg_31_0__13_; 
wire _0key2_reg_31_0__14_; 
wire _0key2_reg_31_0__15_; 
wire _0key2_reg_31_0__16_; 
wire _0key2_reg_31_0__17_; 
wire _0key2_reg_31_0__18_; 
wire _0key2_reg_31_0__19_; 
wire _0key2_reg_31_0__1_; 
wire _0key2_reg_31_0__20_; 
wire _0key2_reg_31_0__21_; 
wire _0key2_reg_31_0__22_; 
wire _0key2_reg_31_0__23_; 
wire _0key2_reg_31_0__24_; 
wire _0key2_reg_31_0__25_; 
wire _0key2_reg_31_0__26_; 
wire _0key2_reg_31_0__27_; 
wire _0key2_reg_31_0__28_; 
wire _0key2_reg_31_0__29_; 
wire _0key2_reg_31_0__2_; 
wire _0key2_reg_31_0__30_; 
wire _0key2_reg_31_0__31_; 
wire _0key2_reg_31_0__3_; 
wire _0key2_reg_31_0__4_; 
wire _0key2_reg_31_0__5_; 
wire _0key2_reg_31_0__6_; 
wire _0key2_reg_31_0__7_; 
wire _0key2_reg_31_0__8_; 
wire _0key2_reg_31_0__9_; 
wire _0key3_reg_31_0__0_; 
wire _0key3_reg_31_0__10_; 
wire _0key3_reg_31_0__11_; 
wire _0key3_reg_31_0__12_; 
wire _0key3_reg_31_0__13_; 
wire _0key3_reg_31_0__14_; 
wire _0key3_reg_31_0__15_; 
wire _0key3_reg_31_0__16_; 
wire _0key3_reg_31_0__17_; 
wire _0key3_reg_31_0__18_; 
wire _0key3_reg_31_0__19_; 
wire _0key3_reg_31_0__1_; 
wire _0key3_reg_31_0__20_; 
wire _0key3_reg_31_0__21_; 
wire _0key3_reg_31_0__22_; 
wire _0key3_reg_31_0__23_; 
wire _0key3_reg_31_0__24_; 
wire _0key3_reg_31_0__25_; 
wire _0key3_reg_31_0__26_; 
wire _0key3_reg_31_0__27_; 
wire _0key3_reg_31_0__28_; 
wire _0key3_reg_31_0__29_; 
wire _0key3_reg_31_0__2_; 
wire _0key3_reg_31_0__30_; 
wire _0key3_reg_31_0__31_; 
wire _0key3_reg_31_0__3_; 
wire _0key3_reg_31_0__4_; 
wire _0key3_reg_31_0__5_; 
wire _0key3_reg_31_0__6_; 
wire _0key3_reg_31_0__7_; 
wire _0key3_reg_31_0__8_; 
wire _0key3_reg_31_0__9_; 
wire _0long_reg_0_0_; 
wire _0mi0_reg_31_0__0_; 
wire _0mi0_reg_31_0__10_; 
wire _0mi0_reg_31_0__11_; 
wire _0mi0_reg_31_0__12_; 
wire _0mi0_reg_31_0__13_; 
wire _0mi0_reg_31_0__14_; 
wire _0mi0_reg_31_0__15_; 
wire _0mi0_reg_31_0__16_; 
wire _0mi0_reg_31_0__17_; 
wire _0mi0_reg_31_0__18_; 
wire _0mi0_reg_31_0__19_; 
wire _0mi0_reg_31_0__1_; 
wire _0mi0_reg_31_0__20_; 
wire _0mi0_reg_31_0__21_; 
wire _0mi0_reg_31_0__22_; 
wire _0mi0_reg_31_0__23_; 
wire _0mi0_reg_31_0__24_; 
wire _0mi0_reg_31_0__25_; 
wire _0mi0_reg_31_0__26_; 
wire _0mi0_reg_31_0__27_; 
wire _0mi0_reg_31_0__28_; 
wire _0mi0_reg_31_0__29_; 
wire _0mi0_reg_31_0__2_; 
wire _0mi0_reg_31_0__30_; 
wire _0mi0_reg_31_0__31_; 
wire _0mi0_reg_31_0__3_; 
wire _0mi0_reg_31_0__4_; 
wire _0mi0_reg_31_0__5_; 
wire _0mi0_reg_31_0__6_; 
wire _0mi0_reg_31_0__7_; 
wire _0mi0_reg_31_0__8_; 
wire _0mi0_reg_31_0__9_; 
wire _0mi1_reg_31_0__0_; 
wire _0mi1_reg_31_0__10_; 
wire _0mi1_reg_31_0__11_; 
wire _0mi1_reg_31_0__12_; 
wire _0mi1_reg_31_0__13_; 
wire _0mi1_reg_31_0__14_; 
wire _0mi1_reg_31_0__15_; 
wire _0mi1_reg_31_0__16_; 
wire _0mi1_reg_31_0__17_; 
wire _0mi1_reg_31_0__18_; 
wire _0mi1_reg_31_0__19_; 
wire _0mi1_reg_31_0__1_; 
wire _0mi1_reg_31_0__20_; 
wire _0mi1_reg_31_0__21_; 
wire _0mi1_reg_31_0__22_; 
wire _0mi1_reg_31_0__23_; 
wire _0mi1_reg_31_0__24_; 
wire _0mi1_reg_31_0__25_; 
wire _0mi1_reg_31_0__26_; 
wire _0mi1_reg_31_0__27_; 
wire _0mi1_reg_31_0__28_; 
wire _0mi1_reg_31_0__29_; 
wire _0mi1_reg_31_0__2_; 
wire _0mi1_reg_31_0__30_; 
wire _0mi1_reg_31_0__31_; 
wire _0mi1_reg_31_0__3_; 
wire _0mi1_reg_31_0__4_; 
wire _0mi1_reg_31_0__5_; 
wire _0mi1_reg_31_0__6_; 
wire _0mi1_reg_31_0__7_; 
wire _0mi1_reg_31_0__8_; 
wire _0mi1_reg_31_0__9_; 
wire _0param_reg_7_0__0_; 
wire _0param_reg_7_0__1_; 
wire _0param_reg_7_0__2_; 
wire _0param_reg_7_0__3_; 
wire _0param_reg_7_0__4_; 
wire _0param_reg_7_0__5_; 
wire _0param_reg_7_0__6_; 
wire _0param_reg_7_0__7_; 
wire _0word0_reg_31_0__0_; 
wire _0word0_reg_31_0__10_; 
wire _0word0_reg_31_0__11_; 
wire _0word0_reg_31_0__12_; 
wire _0word0_reg_31_0__13_; 
wire _0word0_reg_31_0__14_; 
wire _0word0_reg_31_0__15_; 
wire _0word0_reg_31_0__16_; 
wire _0word0_reg_31_0__17_; 
wire _0word0_reg_31_0__18_; 
wire _0word0_reg_31_0__19_; 
wire _0word0_reg_31_0__1_; 
wire _0word0_reg_31_0__20_; 
wire _0word0_reg_31_0__21_; 
wire _0word0_reg_31_0__22_; 
wire _0word0_reg_31_0__23_; 
wire _0word0_reg_31_0__24_; 
wire _0word0_reg_31_0__25_; 
wire _0word0_reg_31_0__26_; 
wire _0word0_reg_31_0__27_; 
wire _0word0_reg_31_0__28_; 
wire _0word0_reg_31_0__29_; 
wire _0word0_reg_31_0__2_; 
wire _0word0_reg_31_0__30_; 
wire _0word0_reg_31_0__31_; 
wire _0word0_reg_31_0__3_; 
wire _0word0_reg_31_0__4_; 
wire _0word0_reg_31_0__5_; 
wire _0word0_reg_31_0__6_; 
wire _0word0_reg_31_0__7_; 
wire _0word0_reg_31_0__8_; 
wire _0word0_reg_31_0__9_; 
wire _0word1_reg_31_0__0_; 
wire _0word1_reg_31_0__10_; 
wire _0word1_reg_31_0__11_; 
wire _0word1_reg_31_0__12_; 
wire _0word1_reg_31_0__13_; 
wire _0word1_reg_31_0__14_; 
wire _0word1_reg_31_0__15_; 
wire _0word1_reg_31_0__16_; 
wire _0word1_reg_31_0__17_; 
wire _0word1_reg_31_0__18_; 
wire _0word1_reg_31_0__19_; 
wire _0word1_reg_31_0__1_; 
wire _0word1_reg_31_0__20_; 
wire _0word1_reg_31_0__21_; 
wire _0word1_reg_31_0__22_; 
wire _0word1_reg_31_0__23_; 
wire _0word1_reg_31_0__24_; 
wire _0word1_reg_31_0__25_; 
wire _0word1_reg_31_0__26_; 
wire _0word1_reg_31_0__27_; 
wire _0word1_reg_31_0__28_; 
wire _0word1_reg_31_0__29_; 
wire _0word1_reg_31_0__2_; 
wire _0word1_reg_31_0__30_; 
wire _0word1_reg_31_0__31_; 
wire _0word1_reg_31_0__3_; 
wire _0word1_reg_31_0__4_; 
wire _0word1_reg_31_0__5_; 
wire _0word1_reg_31_0__6_; 
wire _0word1_reg_31_0__7_; 
wire _0word1_reg_31_0__8_; 
wire _0word1_reg_31_0__9_; 
wire _0word2_reg_31_0__0_; 
wire _0word2_reg_31_0__10_; 
wire _0word2_reg_31_0__11_; 
wire _0word2_reg_31_0__12_; 
wire _0word2_reg_31_0__13_; 
wire _0word2_reg_31_0__14_; 
wire _0word2_reg_31_0__15_; 
wire _0word2_reg_31_0__16_; 
wire _0word2_reg_31_0__17_; 
wire _0word2_reg_31_0__18_; 
wire _0word2_reg_31_0__19_; 
wire _0word2_reg_31_0__1_; 
wire _0word2_reg_31_0__20_; 
wire _0word2_reg_31_0__21_; 
wire _0word2_reg_31_0__22_; 
wire _0word2_reg_31_0__23_; 
wire _0word2_reg_31_0__24_; 
wire _0word2_reg_31_0__25_; 
wire _0word2_reg_31_0__26_; 
wire _0word2_reg_31_0__27_; 
wire _0word2_reg_31_0__28_; 
wire _0word2_reg_31_0__29_; 
wire _0word2_reg_31_0__2_; 
wire _0word2_reg_31_0__30_; 
wire _0word2_reg_31_0__31_; 
wire _0word2_reg_31_0__3_; 
wire _0word2_reg_31_0__4_; 
wire _0word2_reg_31_0__5_; 
wire _0word2_reg_31_0__6_; 
wire _0word2_reg_31_0__7_; 
wire _0word2_reg_31_0__8_; 
wire _0word2_reg_31_0__9_; 
wire _0word3_reg_31_0__0_; 
wire _0word3_reg_31_0__10_; 
wire _0word3_reg_31_0__11_; 
wire _0word3_reg_31_0__12_; 
wire _0word3_reg_31_0__13_; 
wire _0word3_reg_31_0__14_; 
wire _0word3_reg_31_0__15_; 
wire _0word3_reg_31_0__16_; 
wire _0word3_reg_31_0__17_; 
wire _0word3_reg_31_0__18_; 
wire _0word3_reg_31_0__19_; 
wire _0word3_reg_31_0__1_; 
wire _0word3_reg_31_0__20_; 
wire _0word3_reg_31_0__21_; 
wire _0word3_reg_31_0__22_; 
wire _0word3_reg_31_0__23_; 
wire _0word3_reg_31_0__24_; 
wire _0word3_reg_31_0__25_; 
wire _0word3_reg_31_0__26_; 
wire _0word3_reg_31_0__27_; 
wire _0word3_reg_31_0__28_; 
wire _0word3_reg_31_0__29_; 
wire _0word3_reg_31_0__2_; 
wire _0word3_reg_31_0__30_; 
wire _0word3_reg_31_0__31_; 
wire _0word3_reg_31_0__3_; 
wire _0word3_reg_31_0__4_; 
wire _0word3_reg_31_0__5_; 
wire _0word3_reg_31_0__6_; 
wire _0word3_reg_31_0__7_; 
wire _0word3_reg_31_0__8_; 
wire _0word3_reg_31_0__9_; 
wire _abc_19873_new_n1000_; 
wire _abc_19873_new_n1001_; 
wire _abc_19873_new_n1002_; 
wire _abc_19873_new_n1003_; 
wire _abc_19873_new_n1004_; 
wire _abc_19873_new_n1005_; 
wire _abc_19873_new_n1006_; 
wire _abc_19873_new_n1007_; 
wire _abc_19873_new_n1008_; 
wire _abc_19873_new_n1009_; 
wire _abc_19873_new_n1010_; 
wire _abc_19873_new_n1011_; 
wire _abc_19873_new_n1012_; 
wire _abc_19873_new_n1013_; 
wire _abc_19873_new_n1014_; 
wire _abc_19873_new_n1015_; 
wire _abc_19873_new_n1016_; 
wire _abc_19873_new_n1018_; 
wire _abc_19873_new_n1019_; 
wire _abc_19873_new_n1020_; 
wire _abc_19873_new_n1021_; 
wire _abc_19873_new_n1022_; 
wire _abc_19873_new_n1023_; 
wire _abc_19873_new_n1024_; 
wire _abc_19873_new_n1025_; 
wire _abc_19873_new_n1026_; 
wire _abc_19873_new_n1027_; 
wire _abc_19873_new_n1028_; 
wire _abc_19873_new_n1029_; 
wire _abc_19873_new_n1030_; 
wire _abc_19873_new_n1031_; 
wire _abc_19873_new_n1032_; 
wire _abc_19873_new_n1033_; 
wire _abc_19873_new_n1034_; 
wire _abc_19873_new_n1035_; 
wire _abc_19873_new_n1036_; 
wire _abc_19873_new_n1037_; 
wire _abc_19873_new_n1039_; 
wire _abc_19873_new_n1040_; 
wire _abc_19873_new_n1041_; 
wire _abc_19873_new_n1042_; 
wire _abc_19873_new_n1043_; 
wire _abc_19873_new_n1044_; 
wire _abc_19873_new_n1045_; 
wire _abc_19873_new_n1046_; 
wire _abc_19873_new_n1047_; 
wire _abc_19873_new_n1048_; 
wire _abc_19873_new_n1049_; 
wire _abc_19873_new_n1050_; 
wire _abc_19873_new_n1051_; 
wire _abc_19873_new_n1052_; 
wire _abc_19873_new_n1053_; 
wire _abc_19873_new_n1054_; 
wire _abc_19873_new_n1055_; 
wire _abc_19873_new_n1056_; 
wire _abc_19873_new_n1057_; 
wire _abc_19873_new_n1059_; 
wire _abc_19873_new_n1060_; 
wire _abc_19873_new_n1061_; 
wire _abc_19873_new_n1062_; 
wire _abc_19873_new_n1063_; 
wire _abc_19873_new_n1064_; 
wire _abc_19873_new_n1064__bF_buf0; 
wire _abc_19873_new_n1064__bF_buf1; 
wire _abc_19873_new_n1064__bF_buf2; 
wire _abc_19873_new_n1064__bF_buf3; 
wire _abc_19873_new_n1065_; 
wire _abc_19873_new_n1066_; 
wire _abc_19873_new_n1067_; 
wire _abc_19873_new_n1068_; 
wire _abc_19873_new_n1069_; 
wire _abc_19873_new_n1070_; 
wire _abc_19873_new_n1071_; 
wire _abc_19873_new_n1072_; 
wire _abc_19873_new_n1073_; 
wire _abc_19873_new_n1074_; 
wire _abc_19873_new_n1075_; 
wire _abc_19873_new_n1076_; 
wire _abc_19873_new_n1077_; 
wire _abc_19873_new_n1079_; 
wire _abc_19873_new_n1080_; 
wire _abc_19873_new_n1081_; 
wire _abc_19873_new_n1082_; 
wire _abc_19873_new_n1083_; 
wire _abc_19873_new_n1084_; 
wire _abc_19873_new_n1085_; 
wire _abc_19873_new_n1086_; 
wire _abc_19873_new_n1087_; 
wire _abc_19873_new_n1088_; 
wire _abc_19873_new_n1089_; 
wire _abc_19873_new_n1090_; 
wire _abc_19873_new_n1091_; 
wire _abc_19873_new_n1092_; 
wire _abc_19873_new_n1093_; 
wire _abc_19873_new_n1094_; 
wire _abc_19873_new_n1095_; 
wire _abc_19873_new_n1096_; 
wire _abc_19873_new_n1098_; 
wire _abc_19873_new_n1099_; 
wire _abc_19873_new_n1100_; 
wire _abc_19873_new_n1101_; 
wire _abc_19873_new_n1102_; 
wire _abc_19873_new_n1103_; 
wire _abc_19873_new_n1104_; 
wire _abc_19873_new_n1105_; 
wire _abc_19873_new_n1106_; 
wire _abc_19873_new_n1107_; 
wire _abc_19873_new_n1108_; 
wire _abc_19873_new_n1109_; 
wire _abc_19873_new_n1110_; 
wire _abc_19873_new_n1111_; 
wire _abc_19873_new_n1112_; 
wire _abc_19873_new_n1113_; 
wire _abc_19873_new_n1114_; 
wire _abc_19873_new_n1115_; 
wire _abc_19873_new_n1117_; 
wire _abc_19873_new_n1118_; 
wire _abc_19873_new_n1119_; 
wire _abc_19873_new_n1120_; 
wire _abc_19873_new_n1121_; 
wire _abc_19873_new_n1122_; 
wire _abc_19873_new_n1123_; 
wire _abc_19873_new_n1124_; 
wire _abc_19873_new_n1125_; 
wire _abc_19873_new_n1126_; 
wire _abc_19873_new_n1127_; 
wire _abc_19873_new_n1128_; 
wire _abc_19873_new_n1129_; 
wire _abc_19873_new_n1130_; 
wire _abc_19873_new_n1131_; 
wire _abc_19873_new_n1132_; 
wire _abc_19873_new_n1133_; 
wire _abc_19873_new_n1134_; 
wire _abc_19873_new_n1136_; 
wire _abc_19873_new_n1137_; 
wire _abc_19873_new_n1138_; 
wire _abc_19873_new_n1139_; 
wire _abc_19873_new_n1140_; 
wire _abc_19873_new_n1141_; 
wire _abc_19873_new_n1142_; 
wire _abc_19873_new_n1143_; 
wire _abc_19873_new_n1144_; 
wire _abc_19873_new_n1145_; 
wire _abc_19873_new_n1146_; 
wire _abc_19873_new_n1147_; 
wire _abc_19873_new_n1148_; 
wire _abc_19873_new_n1149_; 
wire _abc_19873_new_n1150_; 
wire _abc_19873_new_n1151_; 
wire _abc_19873_new_n1152_; 
wire _abc_19873_new_n1153_; 
wire _abc_19873_new_n1155_; 
wire _abc_19873_new_n1156_; 
wire _abc_19873_new_n1157_; 
wire _abc_19873_new_n1158_; 
wire _abc_19873_new_n1159_; 
wire _abc_19873_new_n1160_; 
wire _abc_19873_new_n1161_; 
wire _abc_19873_new_n1162_; 
wire _abc_19873_new_n1163_; 
wire _abc_19873_new_n1164_; 
wire _abc_19873_new_n1165_; 
wire _abc_19873_new_n1166_; 
wire _abc_19873_new_n1167_; 
wire _abc_19873_new_n1168_; 
wire _abc_19873_new_n1169_; 
wire _abc_19873_new_n1170_; 
wire _abc_19873_new_n1171_; 
wire _abc_19873_new_n1172_; 
wire _abc_19873_new_n1174_; 
wire _abc_19873_new_n1175_; 
wire _abc_19873_new_n1176_; 
wire _abc_19873_new_n1177_; 
wire _abc_19873_new_n1178_; 
wire _abc_19873_new_n1179_; 
wire _abc_19873_new_n1180_; 
wire _abc_19873_new_n1181_; 
wire _abc_19873_new_n1182_; 
wire _abc_19873_new_n1183_; 
wire _abc_19873_new_n1184_; 
wire _abc_19873_new_n1185_; 
wire _abc_19873_new_n1186_; 
wire _abc_19873_new_n1187_; 
wire _abc_19873_new_n1188_; 
wire _abc_19873_new_n1189_; 
wire _abc_19873_new_n1190_; 
wire _abc_19873_new_n1192_; 
wire _abc_19873_new_n1193_; 
wire _abc_19873_new_n1194_; 
wire _abc_19873_new_n1195_; 
wire _abc_19873_new_n1196_; 
wire _abc_19873_new_n1197_; 
wire _abc_19873_new_n1198_; 
wire _abc_19873_new_n1199_; 
wire _abc_19873_new_n1200_; 
wire _abc_19873_new_n1201_; 
wire _abc_19873_new_n1202_; 
wire _abc_19873_new_n1203_; 
wire _abc_19873_new_n1204_; 
wire _abc_19873_new_n1205_; 
wire _abc_19873_new_n1206_; 
wire _abc_19873_new_n1207_; 
wire _abc_19873_new_n1208_; 
wire _abc_19873_new_n1210_; 
wire _abc_19873_new_n1211_; 
wire _abc_19873_new_n1212_; 
wire _abc_19873_new_n1213_; 
wire _abc_19873_new_n1214_; 
wire _abc_19873_new_n1215_; 
wire _abc_19873_new_n1216_; 
wire _abc_19873_new_n1217_; 
wire _abc_19873_new_n1218_; 
wire _abc_19873_new_n1219_; 
wire _abc_19873_new_n1220_; 
wire _abc_19873_new_n1221_; 
wire _abc_19873_new_n1222_; 
wire _abc_19873_new_n1223_; 
wire _abc_19873_new_n1224_; 
wire _abc_19873_new_n1225_; 
wire _abc_19873_new_n1226_; 
wire _abc_19873_new_n1227_; 
wire _abc_19873_new_n1229_; 
wire _abc_19873_new_n1230_; 
wire _abc_19873_new_n1231_; 
wire _abc_19873_new_n1232_; 
wire _abc_19873_new_n1233_; 
wire _abc_19873_new_n1234_; 
wire _abc_19873_new_n1235_; 
wire _abc_19873_new_n1236_; 
wire _abc_19873_new_n1237_; 
wire _abc_19873_new_n1238_; 
wire _abc_19873_new_n1239_; 
wire _abc_19873_new_n1240_; 
wire _abc_19873_new_n1241_; 
wire _abc_19873_new_n1242_; 
wire _abc_19873_new_n1243_; 
wire _abc_19873_new_n1244_; 
wire _abc_19873_new_n1245_; 
wire _abc_19873_new_n1247_; 
wire _abc_19873_new_n1248_; 
wire _abc_19873_new_n1249_; 
wire _abc_19873_new_n1250_; 
wire _abc_19873_new_n1251_; 
wire _abc_19873_new_n1252_; 
wire _abc_19873_new_n1253_; 
wire _abc_19873_new_n1254_; 
wire _abc_19873_new_n1255_; 
wire _abc_19873_new_n1256_; 
wire _abc_19873_new_n1257_; 
wire _abc_19873_new_n1258_; 
wire _abc_19873_new_n1259_; 
wire _abc_19873_new_n1260_; 
wire _abc_19873_new_n1261_; 
wire _abc_19873_new_n1262_; 
wire _abc_19873_new_n1263_; 
wire _abc_19873_new_n1264_; 
wire _abc_19873_new_n1266_; 
wire _abc_19873_new_n1267_; 
wire _abc_19873_new_n1268_; 
wire _abc_19873_new_n1269_; 
wire _abc_19873_new_n1270_; 
wire _abc_19873_new_n1271_; 
wire _abc_19873_new_n1272_; 
wire _abc_19873_new_n1273_; 
wire _abc_19873_new_n1274_; 
wire _abc_19873_new_n1275_; 
wire _abc_19873_new_n1276_; 
wire _abc_19873_new_n1277_; 
wire _abc_19873_new_n1278_; 
wire _abc_19873_new_n1279_; 
wire _abc_19873_new_n1280_; 
wire _abc_19873_new_n1281_; 
wire _abc_19873_new_n1282_; 
wire _abc_19873_new_n1284_; 
wire _abc_19873_new_n1285_; 
wire _abc_19873_new_n1286_; 
wire _abc_19873_new_n1287_; 
wire _abc_19873_new_n1288_; 
wire _abc_19873_new_n1289_; 
wire _abc_19873_new_n1290_; 
wire _abc_19873_new_n1291_; 
wire _abc_19873_new_n1292_; 
wire _abc_19873_new_n1293_; 
wire _abc_19873_new_n1294_; 
wire _abc_19873_new_n1295_; 
wire _abc_19873_new_n1296_; 
wire _abc_19873_new_n1297_; 
wire _abc_19873_new_n1298_; 
wire _abc_19873_new_n1299_; 
wire _abc_19873_new_n1300_; 
wire _abc_19873_new_n1302_; 
wire _abc_19873_new_n1303_; 
wire _abc_19873_new_n1304_; 
wire _abc_19873_new_n1305_; 
wire _abc_19873_new_n1306_; 
wire _abc_19873_new_n1307_; 
wire _abc_19873_new_n1308_; 
wire _abc_19873_new_n1309_; 
wire _abc_19873_new_n1310_; 
wire _abc_19873_new_n1311_; 
wire _abc_19873_new_n1312_; 
wire _abc_19873_new_n1313_; 
wire _abc_19873_new_n1314_; 
wire _abc_19873_new_n1315_; 
wire _abc_19873_new_n1316_; 
wire _abc_19873_new_n1317_; 
wire _abc_19873_new_n1318_; 
wire _abc_19873_new_n1320_; 
wire _abc_19873_new_n1321_; 
wire _abc_19873_new_n1322_; 
wire _abc_19873_new_n1323_; 
wire _abc_19873_new_n1324_; 
wire _abc_19873_new_n1325_; 
wire _abc_19873_new_n1326_; 
wire _abc_19873_new_n1327_; 
wire _abc_19873_new_n1328_; 
wire _abc_19873_new_n1329_; 
wire _abc_19873_new_n1330_; 
wire _abc_19873_new_n1331_; 
wire _abc_19873_new_n1332_; 
wire _abc_19873_new_n1333_; 
wire _abc_19873_new_n1334_; 
wire _abc_19873_new_n1335_; 
wire _abc_19873_new_n1336_; 
wire _abc_19873_new_n1338_; 
wire _abc_19873_new_n1339_; 
wire _abc_19873_new_n1340_; 
wire _abc_19873_new_n1341_; 
wire _abc_19873_new_n1342_; 
wire _abc_19873_new_n1343_; 
wire _abc_19873_new_n1344_; 
wire _abc_19873_new_n1345_; 
wire _abc_19873_new_n1346_; 
wire _abc_19873_new_n1347_; 
wire _abc_19873_new_n1348_; 
wire _abc_19873_new_n1349_; 
wire _abc_19873_new_n1350_; 
wire _abc_19873_new_n1351_; 
wire _abc_19873_new_n1352_; 
wire _abc_19873_new_n1353_; 
wire _abc_19873_new_n1354_; 
wire _abc_19873_new_n1356_; 
wire _abc_19873_new_n1357_; 
wire _abc_19873_new_n1358_; 
wire _abc_19873_new_n1359_; 
wire _abc_19873_new_n1360_; 
wire _abc_19873_new_n1361_; 
wire _abc_19873_new_n1362_; 
wire _abc_19873_new_n1363_; 
wire _abc_19873_new_n1364_; 
wire _abc_19873_new_n1365_; 
wire _abc_19873_new_n1366_; 
wire _abc_19873_new_n1367_; 
wire _abc_19873_new_n1368_; 
wire _abc_19873_new_n1369_; 
wire _abc_19873_new_n1370_; 
wire _abc_19873_new_n1371_; 
wire _abc_19873_new_n1372_; 
wire _abc_19873_new_n1373_; 
wire _abc_19873_new_n1375_; 
wire _abc_19873_new_n1376_; 
wire _abc_19873_new_n1377_; 
wire _abc_19873_new_n1378_; 
wire _abc_19873_new_n1379_; 
wire _abc_19873_new_n1380_; 
wire _abc_19873_new_n1381_; 
wire _abc_19873_new_n1382_; 
wire _abc_19873_new_n1383_; 
wire _abc_19873_new_n1384_; 
wire _abc_19873_new_n1385_; 
wire _abc_19873_new_n1386_; 
wire _abc_19873_new_n1387_; 
wire _abc_19873_new_n1388_; 
wire _abc_19873_new_n1389_; 
wire _abc_19873_new_n1390_; 
wire _abc_19873_new_n1391_; 
wire _abc_19873_new_n1393_; 
wire _abc_19873_new_n1394_; 
wire _abc_19873_new_n1395_; 
wire _abc_19873_new_n1396_; 
wire _abc_19873_new_n1397_; 
wire _abc_19873_new_n1398_; 
wire _abc_19873_new_n1399_; 
wire _abc_19873_new_n1400_; 
wire _abc_19873_new_n1401_; 
wire _abc_19873_new_n1402_; 
wire _abc_19873_new_n1403_; 
wire _abc_19873_new_n1404_; 
wire _abc_19873_new_n1405_; 
wire _abc_19873_new_n1406_; 
wire _abc_19873_new_n1407_; 
wire _abc_19873_new_n1408_; 
wire _abc_19873_new_n1409_; 
wire _abc_19873_new_n1411_; 
wire _abc_19873_new_n1412_; 
wire _abc_19873_new_n1413_; 
wire _abc_19873_new_n1414_; 
wire _abc_19873_new_n1415_; 
wire _abc_19873_new_n1416_; 
wire _abc_19873_new_n1417_; 
wire _abc_19873_new_n1418_; 
wire _abc_19873_new_n1419_; 
wire _abc_19873_new_n1420_; 
wire _abc_19873_new_n1421_; 
wire _abc_19873_new_n1422_; 
wire _abc_19873_new_n1423_; 
wire _abc_19873_new_n1424_; 
wire _abc_19873_new_n1425_; 
wire _abc_19873_new_n1426_; 
wire _abc_19873_new_n1427_; 
wire _abc_19873_new_n1428_; 
wire _abc_19873_new_n1430_; 
wire _abc_19873_new_n1431_; 
wire _abc_19873_new_n1432_; 
wire _abc_19873_new_n1433_; 
wire _abc_19873_new_n1434_; 
wire _abc_19873_new_n1435_; 
wire _abc_19873_new_n1436_; 
wire _abc_19873_new_n1437_; 
wire _abc_19873_new_n1438_; 
wire _abc_19873_new_n1439_; 
wire _abc_19873_new_n1440_; 
wire _abc_19873_new_n1441_; 
wire _abc_19873_new_n1442_; 
wire _abc_19873_new_n1443_; 
wire _abc_19873_new_n1444_; 
wire _abc_19873_new_n1445_; 
wire _abc_19873_new_n1446_; 
wire _abc_19873_new_n1447_; 
wire _abc_19873_new_n1449_; 
wire _abc_19873_new_n1450_; 
wire _abc_19873_new_n1451_; 
wire _abc_19873_new_n1452_; 
wire _abc_19873_new_n1453_; 
wire _abc_19873_new_n1454_; 
wire _abc_19873_new_n1455_; 
wire _abc_19873_new_n1456_; 
wire _abc_19873_new_n1457_; 
wire _abc_19873_new_n1458_; 
wire _abc_19873_new_n1459_; 
wire _abc_19873_new_n1460_; 
wire _abc_19873_new_n1461_; 
wire _abc_19873_new_n1462_; 
wire _abc_19873_new_n1463_; 
wire _abc_19873_new_n1464_; 
wire _abc_19873_new_n1465_; 
wire _abc_19873_new_n1467_; 
wire _abc_19873_new_n1468_; 
wire _abc_19873_new_n1469_; 
wire _abc_19873_new_n1470_; 
wire _abc_19873_new_n1471_; 
wire _abc_19873_new_n1472_; 
wire _abc_19873_new_n1473_; 
wire _abc_19873_new_n1474_; 
wire _abc_19873_new_n1475_; 
wire _abc_19873_new_n1476_; 
wire _abc_19873_new_n1477_; 
wire _abc_19873_new_n1478_; 
wire _abc_19873_new_n1479_; 
wire _abc_19873_new_n1480_; 
wire _abc_19873_new_n1481_; 
wire _abc_19873_new_n1482_; 
wire _abc_19873_new_n1483_; 
wire _abc_19873_new_n1484_; 
wire _abc_19873_new_n1485_; 
wire _abc_19873_new_n1487_; 
wire _abc_19873_new_n1488_; 
wire _abc_19873_new_n1489_; 
wire _abc_19873_new_n1490_; 
wire _abc_19873_new_n1491_; 
wire _abc_19873_new_n1492_; 
wire _abc_19873_new_n1493_; 
wire _abc_19873_new_n1494_; 
wire _abc_19873_new_n1495_; 
wire _abc_19873_new_n1496_; 
wire _abc_19873_new_n1497_; 
wire _abc_19873_new_n1498_; 
wire _abc_19873_new_n1499_; 
wire _abc_19873_new_n1500_; 
wire _abc_19873_new_n1501_; 
wire _abc_19873_new_n1502_; 
wire _abc_19873_new_n1503_; 
wire _abc_19873_new_n1505_; 
wire _abc_19873_new_n1506_; 
wire _abc_19873_new_n1507_; 
wire _abc_19873_new_n1508_; 
wire _abc_19873_new_n1509_; 
wire _abc_19873_new_n1510_; 
wire _abc_19873_new_n1511_; 
wire _abc_19873_new_n1512_; 
wire _abc_19873_new_n1513_; 
wire _abc_19873_new_n1514_; 
wire _abc_19873_new_n1515_; 
wire _abc_19873_new_n1516_; 
wire _abc_19873_new_n1517_; 
wire _abc_19873_new_n1518_; 
wire _abc_19873_new_n1519_; 
wire _abc_19873_new_n1520_; 
wire _abc_19873_new_n1521_; 
wire _abc_19873_new_n1522_; 
wire _abc_19873_new_n1524_; 
wire _abc_19873_new_n1524__bF_buf0; 
wire _abc_19873_new_n1524__bF_buf1; 
wire _abc_19873_new_n1524__bF_buf10; 
wire _abc_19873_new_n1524__bF_buf11; 
wire _abc_19873_new_n1524__bF_buf12; 
wire _abc_19873_new_n1524__bF_buf13; 
wire _abc_19873_new_n1524__bF_buf14; 
wire _abc_19873_new_n1524__bF_buf15; 
wire _abc_19873_new_n1524__bF_buf2; 
wire _abc_19873_new_n1524__bF_buf3; 
wire _abc_19873_new_n1524__bF_buf4; 
wire _abc_19873_new_n1524__bF_buf5; 
wire _abc_19873_new_n1524__bF_buf6; 
wire _abc_19873_new_n1524__bF_buf7; 
wire _abc_19873_new_n1524__bF_buf8; 
wire _abc_19873_new_n1524__bF_buf9; 
wire _abc_19873_new_n1525_; 
wire _abc_19873_new_n1527_; 
wire _abc_19873_new_n1529_; 
wire _abc_19873_new_n1530_; 
wire _abc_19873_new_n1532_; 
wire _abc_19873_new_n1534_; 
wire _abc_19873_new_n1536_; 
wire _abc_19873_new_n1538_; 
wire _abc_19873_new_n1540_; 
wire _abc_19873_new_n1541_; 
wire _abc_19873_new_n1543_; 
wire _abc_19873_new_n1545_; 
wire _abc_19873_new_n1547_; 
wire _abc_19873_new_n1549_; 
wire _abc_19873_new_n1550_; 
wire _abc_19873_new_n1552_; 
wire _abc_19873_new_n1553_; 
wire _abc_19873_new_n1555_; 
wire _abc_19873_new_n1556_; 
wire _abc_19873_new_n1558_; 
wire _abc_19873_new_n1559_; 
wire _abc_19873_new_n1561_; 
wire _abc_19873_new_n1563_; 
wire _abc_19873_new_n1564_; 
wire _abc_19873_new_n1566_; 
wire _abc_19873_new_n1567_; 
wire _abc_19873_new_n1569_; 
wire _abc_19873_new_n1570_; 
wire _abc_19873_new_n1572_; 
wire _abc_19873_new_n1573_; 
wire _abc_19873_new_n1575_; 
wire _abc_19873_new_n1576_; 
wire _abc_19873_new_n1578_; 
wire _abc_19873_new_n1579_; 
wire _abc_19873_new_n1581_; 
wire _abc_19873_new_n1582_; 
wire _abc_19873_new_n1584_; 
wire _abc_19873_new_n1586_; 
wire _abc_19873_new_n1587_; 
wire _abc_19873_new_n1589_; 
wire _abc_19873_new_n1590_; 
wire _abc_19873_new_n1592_; 
wire _abc_19873_new_n1594_; 
wire _abc_19873_new_n1596_; 
wire _abc_19873_new_n1597_; 
wire _abc_19873_new_n1599_; 
wire _abc_19873_new_n1601_; 
wire _abc_19873_new_n1602_; 
wire _abc_19873_new_n1604_; 
wire _abc_19873_new_n1606_; 
wire _abc_19873_new_n1607_; 
wire _abc_19873_new_n1609_; 
wire _abc_19873_new_n1610_; 
wire _abc_19873_new_n1612_; 
wire _abc_19873_new_n1614_; 
wire _abc_19873_new_n1615_; 
wire _abc_19873_new_n1617_; 
wire _abc_19873_new_n1618_; 
wire _abc_19873_new_n1620_; 
wire _abc_19873_new_n1621_; 
wire _abc_19873_new_n1623_; 
wire _abc_19873_new_n1624_; 
wire _abc_19873_new_n1626_; 
wire _abc_19873_new_n1627_; 
wire _abc_19873_new_n1629_; 
wire _abc_19873_new_n1631_; 
wire _abc_19873_new_n1633_; 
wire _abc_19873_new_n1635_; 
wire _abc_19873_new_n1636_; 
wire _abc_19873_new_n1638_; 
wire _abc_19873_new_n1639_; 
wire _abc_19873_new_n1641_; 
wire _abc_19873_new_n1643_; 
wire _abc_19873_new_n1644_; 
wire _abc_19873_new_n1646_; 
wire _abc_19873_new_n1648_; 
wire _abc_19873_new_n1649_; 
wire _abc_19873_new_n1651_; 
wire _abc_19873_new_n1652_; 
wire _abc_19873_new_n1654_; 
wire _abc_19873_new_n1655_; 
wire _abc_19873_new_n1657_; 
wire _abc_19873_new_n1658_; 
wire _abc_19873_new_n1660_; 
wire _abc_19873_new_n1661_; 
wire _abc_19873_new_n1663_; 
wire _abc_19873_new_n1665_; 
wire _abc_19873_new_n1666_; 
wire _abc_19873_new_n1668_; 
wire _abc_19873_new_n1670_; 
wire _abc_19873_new_n1671_; 
wire _abc_19873_new_n1673_; 
wire _abc_19873_new_n1674_; 
wire _abc_19873_new_n1676_; 
wire _abc_19873_new_n1678_; 
wire _abc_19873_new_n1680_; 
wire _abc_19873_new_n1681_; 
wire _abc_19873_new_n1683_; 
wire _abc_19873_new_n1685_; 
wire _abc_19873_new_n1686_; 
wire _abc_19873_new_n1688_; 
wire _abc_19873_new_n1690_; 
wire _abc_19873_new_n1692_; 
wire _abc_19873_new_n1694_; 
wire _abc_19873_new_n1695_; 
wire _abc_19873_new_n1697_; 
wire _abc_19873_new_n1698_; 
wire _abc_19873_new_n1700_; 
wire _abc_19873_new_n1701_; 
wire _abc_19873_new_n1703_; 
wire _abc_19873_new_n1705_; 
wire _abc_19873_new_n1706_; 
wire _abc_19873_new_n1708_; 
wire _abc_19873_new_n1709_; 
wire _abc_19873_new_n1711_; 
wire _abc_19873_new_n1713_; 
wire _abc_19873_new_n1715_; 
wire _abc_19873_new_n1717_; 
wire _abc_19873_new_n1718_; 
wire _abc_19873_new_n1720_; 
wire _abc_19873_new_n1721_; 
wire _abc_19873_new_n1723_; 
wire _abc_19873_new_n1724_; 
wire _abc_19873_new_n1726_; 
wire _abc_19873_new_n1727_; 
wire _abc_19873_new_n1729_; 
wire _abc_19873_new_n1731_; 
wire _abc_19873_new_n1732_; 
wire _abc_19873_new_n1734_; 
wire _abc_19873_new_n1735_; 
wire _abc_19873_new_n1737_; 
wire _abc_19873_new_n1738_; 
wire _abc_19873_new_n1740_; 
wire _abc_19873_new_n1741_; 
wire _abc_19873_new_n1743_; 
wire _abc_19873_new_n1744_; 
wire _abc_19873_new_n1746_; 
wire _abc_19873_new_n1747_; 
wire _abc_19873_new_n1749_; 
wire _abc_19873_new_n1750_; 
wire _abc_19873_new_n1752_; 
wire _abc_19873_new_n1754_; 
wire _abc_19873_new_n1755_; 
wire _abc_19873_new_n1757_; 
wire _abc_19873_new_n1758_; 
wire _abc_19873_new_n1760_; 
wire _abc_19873_new_n1762_; 
wire _abc_19873_new_n1764_; 
wire _abc_19873_new_n1765_; 
wire _abc_19873_new_n1767_; 
wire _abc_19873_new_n1769_; 
wire _abc_19873_new_n1770_; 
wire _abc_19873_new_n1772_; 
wire _abc_19873_new_n1774_; 
wire _abc_19873_new_n1775_; 
wire _abc_19873_new_n1777_; 
wire _abc_19873_new_n1778_; 
wire _abc_19873_new_n1780_; 
wire _abc_19873_new_n1781_; 
wire _abc_19873_new_n1783_; 
wire _abc_19873_new_n1784_; 
wire _abc_19873_new_n1786_; 
wire _abc_19873_new_n1787_; 
wire _abc_19873_new_n1789_; 
wire _abc_19873_new_n1790_; 
wire _abc_19873_new_n1792_; 
wire _abc_19873_new_n1793_; 
wire _abc_19873_new_n1795_; 
wire _abc_19873_new_n1797_; 
wire _abc_19873_new_n1799_; 
wire _abc_19873_new_n1801_; 
wire _abc_19873_new_n1803_; 
wire _abc_19873_new_n1805_; 
wire _abc_19873_new_n1807_; 
wire _abc_19873_new_n1808_; 
wire _abc_19873_new_n1810_; 
wire _abc_19873_new_n1812_; 
wire _abc_19873_new_n1814_; 
wire _abc_19873_new_n1816_; 
wire _abc_19873_new_n1818_; 
wire _abc_19873_new_n1820_; 
wire _abc_19873_new_n1822_; 
wire _abc_19873_new_n1824_; 
wire _abc_19873_new_n1825_; 
wire _abc_19873_new_n1827_; 
wire _abc_19873_new_n1829_; 
wire _abc_19873_new_n1831_; 
wire _abc_19873_new_n1833_; 
wire _abc_19873_new_n1835_; 
wire _abc_19873_new_n1837_; 
wire _abc_19873_new_n1839_; 
wire _abc_19873_new_n1841_; 
wire _abc_19873_new_n1843_; 
wire _abc_19873_new_n1845_; 
wire _abc_19873_new_n1847_; 
wire _abc_19873_new_n1848_; 
wire _abc_19873_new_n1849_; 
wire _abc_19873_new_n1849__bF_buf0; 
wire _abc_19873_new_n1849__bF_buf1; 
wire _abc_19873_new_n1849__bF_buf2; 
wire _abc_19873_new_n1849__bF_buf3; 
wire _abc_19873_new_n1849__bF_buf4; 
wire _abc_19873_new_n1849__bF_buf5; 
wire _abc_19873_new_n1849__bF_buf6; 
wire _abc_19873_new_n1849__bF_buf7; 
wire _abc_19873_new_n1850_; 
wire _abc_19873_new_n1852_; 
wire _abc_19873_new_n1853_; 
wire _abc_19873_new_n1855_; 
wire _abc_19873_new_n1857_; 
wire _abc_19873_new_n1859_; 
wire _abc_19873_new_n1861_; 
wire _abc_19873_new_n1862_; 
wire _abc_19873_new_n1864_; 
wire _abc_19873_new_n1866_; 
wire _abc_19873_new_n1868_; 
wire _abc_19873_new_n1870_; 
wire _abc_19873_new_n1872_; 
wire _abc_19873_new_n1874_; 
wire _abc_19873_new_n1876_; 
wire _abc_19873_new_n1878_; 
wire _abc_19873_new_n1880_; 
wire _abc_19873_new_n1881_; 
wire _abc_19873_new_n1883_; 
wire _abc_19873_new_n1885_; 
wire _abc_19873_new_n1886_; 
wire _abc_19873_new_n1888_; 
wire _abc_19873_new_n1890_; 
wire _abc_19873_new_n1892_; 
wire _abc_19873_new_n1893_; 
wire _abc_19873_new_n1895_; 
wire _abc_19873_new_n1897_; 
wire _abc_19873_new_n1899_; 
wire _abc_19873_new_n1900_; 
wire _abc_19873_new_n1902_; 
wire _abc_19873_new_n1904_; 
wire _abc_19873_new_n1905_; 
wire _abc_19873_new_n1907_; 
wire _abc_19873_new_n1908_; 
wire _abc_19873_new_n1910_; 
wire _abc_19873_new_n1912_; 
wire _abc_19873_new_n1914_; 
wire _abc_19873_new_n1915_; 
wire _abc_19873_new_n1917_; 
wire _abc_19873_new_n1918_; 
wire _abc_19873_new_n1920_; 
wire _abc_19873_new_n1921_; 
wire _abc_19873_new_n1923_; 
wire _abc_19873_new_n1925_; 
wire _abc_19873_new_n1925__bF_buf0; 
wire _abc_19873_new_n1925__bF_buf1; 
wire _abc_19873_new_n1925__bF_buf2; 
wire _abc_19873_new_n1925__bF_buf3; 
wire _abc_19873_new_n1925__bF_buf4; 
wire _abc_19873_new_n1925__bF_buf5; 
wire _abc_19873_new_n1925__bF_buf6; 
wire _abc_19873_new_n1925__bF_buf7; 
wire _abc_19873_new_n1926_; 
wire _abc_19873_new_n1928_; 
wire _abc_19873_new_n1930_; 
wire _abc_19873_new_n1932_; 
wire _abc_19873_new_n1934_; 
wire _abc_19873_new_n1936_; 
wire _abc_19873_new_n1938_; 
wire _abc_19873_new_n1940_; 
wire _abc_19873_new_n1942_; 
wire _abc_19873_new_n1944_; 
wire _abc_19873_new_n1946_; 
wire _abc_19873_new_n1948_; 
wire _abc_19873_new_n1950_; 
wire _abc_19873_new_n1952_; 
wire _abc_19873_new_n1954_; 
wire _abc_19873_new_n1956_; 
wire _abc_19873_new_n1958_; 
wire _abc_19873_new_n1960_; 
wire _abc_19873_new_n1961_; 
wire _abc_19873_new_n1963_; 
wire _abc_19873_new_n1965_; 
wire _abc_19873_new_n1967_; 
wire _abc_19873_new_n1969_; 
wire _abc_19873_new_n1971_; 
wire _abc_19873_new_n1973_; 
wire _abc_19873_new_n1975_; 
wire _abc_19873_new_n1977_; 
wire _abc_19873_new_n1979_; 
wire _abc_19873_new_n1981_; 
wire _abc_19873_new_n1983_; 
wire _abc_19873_new_n1985_; 
wire _abc_19873_new_n1986_; 
wire _abc_19873_new_n1988_; 
wire _abc_19873_new_n1990_; 
wire _abc_19873_new_n1992_; 
wire _abc_19873_new_n1992__bF_buf0; 
wire _abc_19873_new_n1992__bF_buf1; 
wire _abc_19873_new_n1992__bF_buf2; 
wire _abc_19873_new_n1992__bF_buf3; 
wire _abc_19873_new_n1992__bF_buf4; 
wire _abc_19873_new_n1992__bF_buf5; 
wire _abc_19873_new_n1992__bF_buf6; 
wire _abc_19873_new_n1992__bF_buf7; 
wire _abc_19873_new_n1993_; 
wire _abc_19873_new_n1995_; 
wire _abc_19873_new_n1997_; 
wire _abc_19873_new_n1999_; 
wire _abc_19873_new_n2001_; 
wire _abc_19873_new_n2003_; 
wire _abc_19873_new_n2005_; 
wire _abc_19873_new_n2007_; 
wire _abc_19873_new_n2009_; 
wire _abc_19873_new_n2011_; 
wire _abc_19873_new_n2013_; 
wire _abc_19873_new_n2015_; 
wire _abc_19873_new_n2017_; 
wire _abc_19873_new_n2019_; 
wire _abc_19873_new_n2021_; 
wire _abc_19873_new_n2023_; 
wire _abc_19873_new_n2025_; 
wire _abc_19873_new_n2027_; 
wire _abc_19873_new_n2029_; 
wire _abc_19873_new_n2031_; 
wire _abc_19873_new_n2033_; 
wire _abc_19873_new_n2035_; 
wire _abc_19873_new_n2037_; 
wire _abc_19873_new_n2039_; 
wire _abc_19873_new_n2041_; 
wire _abc_19873_new_n2043_; 
wire _abc_19873_new_n2045_; 
wire _abc_19873_new_n2047_; 
wire _abc_19873_new_n2049_; 
wire _abc_19873_new_n2051_; 
wire _abc_19873_new_n2052_; 
wire _abc_19873_new_n2054_; 
wire _abc_19873_new_n2056_; 
wire _abc_19873_new_n2058_; 
wire _abc_19873_new_n2058__bF_buf0; 
wire _abc_19873_new_n2058__bF_buf1; 
wire _abc_19873_new_n2058__bF_buf2; 
wire _abc_19873_new_n2058__bF_buf3; 
wire _abc_19873_new_n2058__bF_buf4; 
wire _abc_19873_new_n2058__bF_buf5; 
wire _abc_19873_new_n2058__bF_buf6; 
wire _abc_19873_new_n2058__bF_buf7; 
wire _abc_19873_new_n2059_; 
wire _abc_19873_new_n2061_; 
wire _abc_19873_new_n2063_; 
wire _abc_19873_new_n2065_; 
wire _abc_19873_new_n2067_; 
wire _abc_19873_new_n2069_; 
wire _abc_19873_new_n2071_; 
wire _abc_19873_new_n2072_; 
wire _abc_19873_new_n2074_; 
wire _abc_19873_new_n2075_; 
wire _abc_19873_new_n2077_; 
wire _abc_19873_new_n2079_; 
wire _abc_19873_new_n2081_; 
wire _abc_19873_new_n2083_; 
wire _abc_19873_new_n2085_; 
wire _abc_19873_new_n2087_; 
wire _abc_19873_new_n2089_; 
wire _abc_19873_new_n2091_; 
wire _abc_19873_new_n2093_; 
wire _abc_19873_new_n2095_; 
wire _abc_19873_new_n2097_; 
wire _abc_19873_new_n2099_; 
wire _abc_19873_new_n2101_; 
wire _abc_19873_new_n2103_; 
wire _abc_19873_new_n2105_; 
wire _abc_19873_new_n2107_; 
wire _abc_19873_new_n2109_; 
wire _abc_19873_new_n2111_; 
wire _abc_19873_new_n2113_; 
wire _abc_19873_new_n2115_; 
wire _abc_19873_new_n2117_; 
wire _abc_19873_new_n2119_; 
wire _abc_19873_new_n2121_; 
wire _abc_19873_new_n2123_; 
wire _abc_19873_new_n2125_; 
wire _abc_19873_new_n2125__bF_buf0; 
wire _abc_19873_new_n2125__bF_buf1; 
wire _abc_19873_new_n2125__bF_buf2; 
wire _abc_19873_new_n2125__bF_buf3; 
wire _abc_19873_new_n2125__bF_buf4; 
wire _abc_19873_new_n2125__bF_buf5; 
wire _abc_19873_new_n2125__bF_buf6; 
wire _abc_19873_new_n2125__bF_buf7; 
wire _abc_19873_new_n2126_; 
wire _abc_19873_new_n2128_; 
wire _abc_19873_new_n2130_; 
wire _abc_19873_new_n2132_; 
wire _abc_19873_new_n2133_; 
wire _abc_19873_new_n2135_; 
wire _abc_19873_new_n2136_; 
wire _abc_19873_new_n2138_; 
wire _abc_19873_new_n2139_; 
wire _abc_19873_new_n2141_; 
wire _abc_19873_new_n2143_; 
wire _abc_19873_new_n2145_; 
wire _abc_19873_new_n2147_; 
wire _abc_19873_new_n2149_; 
wire _abc_19873_new_n2151_; 
wire _abc_19873_new_n2152_; 
wire _abc_19873_new_n2154_; 
wire _abc_19873_new_n2155_; 
wire _abc_19873_new_n2157_; 
wire _abc_19873_new_n2159_; 
wire _abc_19873_new_n2161_; 
wire _abc_19873_new_n2163_; 
wire _abc_19873_new_n2165_; 
wire _abc_19873_new_n2167_; 
wire _abc_19873_new_n2168_; 
wire _abc_19873_new_n2170_; 
wire _abc_19873_new_n2172_; 
wire _abc_19873_new_n2173_; 
wire _abc_19873_new_n2175_; 
wire _abc_19873_new_n2177_; 
wire _abc_19873_new_n2179_; 
wire _abc_19873_new_n2181_; 
wire _abc_19873_new_n2183_; 
wire _abc_19873_new_n2185_; 
wire _abc_19873_new_n2187_; 
wire _abc_19873_new_n2189_; 
wire _abc_19873_new_n2191_; 
wire _abc_19873_new_n2193_; 
wire _abc_19873_new_n2195_; 
wire _abc_19873_new_n2197_; 
wire _abc_19873_new_n2198_; 
wire _abc_19873_new_n2198__bF_buf0; 
wire _abc_19873_new_n2198__bF_buf1; 
wire _abc_19873_new_n2198__bF_buf2; 
wire _abc_19873_new_n2198__bF_buf3; 
wire _abc_19873_new_n2198__bF_buf4; 
wire _abc_19873_new_n2198__bF_buf5; 
wire _abc_19873_new_n2198__bF_buf6; 
wire _abc_19873_new_n2198__bF_buf7; 
wire _abc_19873_new_n2199_; 
wire _abc_19873_new_n2201_; 
wire _abc_19873_new_n2202_; 
wire _abc_19873_new_n2204_; 
wire _abc_19873_new_n2206_; 
wire _abc_19873_new_n2208_; 
wire _abc_19873_new_n2210_; 
wire _abc_19873_new_n2212_; 
wire _abc_19873_new_n2214_; 
wire _abc_19873_new_n2216_; 
wire _abc_19873_new_n2218_; 
wire _abc_19873_new_n2220_; 
wire _abc_19873_new_n2222_; 
wire _abc_19873_new_n2224_; 
wire _abc_19873_new_n2226_; 
wire _abc_19873_new_n2228_; 
wire _abc_19873_new_n2230_; 
wire _abc_19873_new_n2232_; 
wire _abc_19873_new_n2234_; 
wire _abc_19873_new_n2236_; 
wire _abc_19873_new_n2238_; 
wire _abc_19873_new_n2240_; 
wire _abc_19873_new_n2242_; 
wire _abc_19873_new_n2244_; 
wire _abc_19873_new_n2246_; 
wire _abc_19873_new_n2248_; 
wire _abc_19873_new_n2250_; 
wire _abc_19873_new_n2252_; 
wire _abc_19873_new_n2254_; 
wire _abc_19873_new_n2256_; 
wire _abc_19873_new_n2258_; 
wire _abc_19873_new_n2259_; 
wire _abc_19873_new_n2261_; 
wire _abc_19873_new_n2263_; 
wire _abc_19873_new_n2265_; 
wire _abc_19873_new_n2266_; 
wire _abc_19873_new_n2267_; 
wire _abc_19873_new_n2269_; 
wire _abc_19873_new_n2270_; 
wire _abc_19873_new_n2272_; 
wire _abc_19873_new_n2274_; 
wire _abc_19873_new_n2276_; 
wire _abc_19873_new_n2278_; 
wire _abc_19873_new_n2280_; 
wire _abc_19873_new_n2282_; 
wire _abc_19873_new_n2284_; 
wire _abc_19873_new_n2285_; 
wire _abc_19873_new_n2286_; 
wire _abc_19873_new_n2287_; 
wire _abc_19873_new_n2289_; 
wire _abc_19873_new_n2291_; 
wire _abc_19873_new_n2293_; 
wire _abc_19873_new_n2294_; 
wire _abc_19873_new_n2295_; 
wire _abc_19873_new_n2296_; 
wire _abc_19873_new_n870_; 
wire _abc_19873_new_n871_; 
wire _abc_19873_new_n872_; 
wire _abc_19873_new_n873_; 
wire _abc_19873_new_n874_; 
wire _abc_19873_new_n875_; 
wire _abc_19873_new_n876_; 
wire _abc_19873_new_n877_; 
wire _abc_19873_new_n878_; 
wire _abc_19873_new_n879_; 
wire _abc_19873_new_n880_; 
wire _abc_19873_new_n881_; 
wire _abc_19873_new_n882_; 
wire _abc_19873_new_n883_; 
wire _abc_19873_new_n884_; 
wire _abc_19873_new_n885_; 
wire _abc_19873_new_n886_; 
wire _abc_19873_new_n887_; 
wire _abc_19873_new_n888_; 
wire _abc_19873_new_n889_; 
wire _abc_19873_new_n889__bF_buf0; 
wire _abc_19873_new_n889__bF_buf1; 
wire _abc_19873_new_n889__bF_buf2; 
wire _abc_19873_new_n889__bF_buf3; 
wire _abc_19873_new_n889__bF_buf4; 
wire _abc_19873_new_n890_; 
wire _abc_19873_new_n891_; 
wire _abc_19873_new_n892_; 
wire _abc_19873_new_n893_; 
wire _abc_19873_new_n893__bF_buf0; 
wire _abc_19873_new_n893__bF_buf1; 
wire _abc_19873_new_n893__bF_buf2; 
wire _abc_19873_new_n893__bF_buf3; 
wire _abc_19873_new_n893__bF_buf4; 
wire _abc_19873_new_n894_; 
wire _abc_19873_new_n894__bF_buf0; 
wire _abc_19873_new_n894__bF_buf1; 
wire _abc_19873_new_n894__bF_buf2; 
wire _abc_19873_new_n894__bF_buf3; 
wire _abc_19873_new_n894__bF_buf4; 
wire _abc_19873_new_n895_; 
wire _abc_19873_new_n895__bF_buf0; 
wire _abc_19873_new_n895__bF_buf1; 
wire _abc_19873_new_n895__bF_buf2; 
wire _abc_19873_new_n895__bF_buf3; 
wire _abc_19873_new_n895__bF_buf4; 
wire _abc_19873_new_n896_; 
wire _abc_19873_new_n896__bF_buf0; 
wire _abc_19873_new_n896__bF_buf1; 
wire _abc_19873_new_n896__bF_buf2; 
wire _abc_19873_new_n896__bF_buf3; 
wire _abc_19873_new_n896__bF_buf4; 
wire _abc_19873_new_n897_; 
wire _abc_19873_new_n898_; 
wire _abc_19873_new_n899_; 
wire _abc_19873_new_n900_; 
wire _abc_19873_new_n901_; 
wire _abc_19873_new_n901__bF_buf0; 
wire _abc_19873_new_n901__bF_buf1; 
wire _abc_19873_new_n901__bF_buf2; 
wire _abc_19873_new_n901__bF_buf3; 
wire _abc_19873_new_n901__bF_buf4; 
wire _abc_19873_new_n901__bF_buf5; 
wire _abc_19873_new_n901__bF_buf6; 
wire _abc_19873_new_n901__bF_buf7; 
wire _abc_19873_new_n902_; 
wire _abc_19873_new_n903_; 
wire _abc_19873_new_n904_; 
wire _abc_19873_new_n905_; 
wire _abc_19873_new_n905__bF_buf0; 
wire _abc_19873_new_n905__bF_buf1; 
wire _abc_19873_new_n905__bF_buf2; 
wire _abc_19873_new_n905__bF_buf3; 
wire _abc_19873_new_n906_; 
wire _abc_19873_new_n907_; 
wire _abc_19873_new_n908_; 
wire _abc_19873_new_n909_; 
wire _abc_19873_new_n910_; 
wire _abc_19873_new_n911_; 
wire _abc_19873_new_n912_; 
wire _abc_19873_new_n912__bF_buf0; 
wire _abc_19873_new_n912__bF_buf1; 
wire _abc_19873_new_n912__bF_buf2; 
wire _abc_19873_new_n912__bF_buf3; 
wire _abc_19873_new_n913_; 
wire _abc_19873_new_n913__bF_buf0; 
wire _abc_19873_new_n913__bF_buf1; 
wire _abc_19873_new_n913__bF_buf2; 
wire _abc_19873_new_n913__bF_buf3; 
wire _abc_19873_new_n913__bF_buf4; 
wire _abc_19873_new_n914_; 
wire _abc_19873_new_n914__bF_buf0; 
wire _abc_19873_new_n914__bF_buf1; 
wire _abc_19873_new_n914__bF_buf2; 
wire _abc_19873_new_n914__bF_buf3; 
wire _abc_19873_new_n914__bF_buf4; 
wire _abc_19873_new_n915_; 
wire _abc_19873_new_n916_; 
wire _abc_19873_new_n917_; 
wire _abc_19873_new_n918_; 
wire _abc_19873_new_n919_; 
wire _abc_19873_new_n920_; 
wire _abc_19873_new_n921_; 
wire _abc_19873_new_n922_; 
wire _abc_19873_new_n923_; 
wire _abc_19873_new_n924_; 
wire _abc_19873_new_n925_; 
wire _abc_19873_new_n926_; 
wire _abc_19873_new_n927_; 
wire _abc_19873_new_n928_; 
wire _abc_19873_new_n928__bF_buf0; 
wire _abc_19873_new_n928__bF_buf1; 
wire _abc_19873_new_n928__bF_buf2; 
wire _abc_19873_new_n928__bF_buf3; 
wire _abc_19873_new_n928__bF_buf4; 
wire _abc_19873_new_n930_; 
wire _abc_19873_new_n931_; 
wire _abc_19873_new_n932_; 
wire _abc_19873_new_n933_; 
wire _abc_19873_new_n934_; 
wire _abc_19873_new_n935_; 
wire _abc_19873_new_n936_; 
wire _abc_19873_new_n937_; 
wire _abc_19873_new_n938_; 
wire _abc_19873_new_n939_; 
wire _abc_19873_new_n940_; 
wire _abc_19873_new_n941_; 
wire _abc_19873_new_n942_; 
wire _abc_19873_new_n943_; 
wire _abc_19873_new_n944_; 
wire _abc_19873_new_n945_; 
wire _abc_19873_new_n946_; 
wire _abc_19873_new_n947_; 
wire _abc_19873_new_n948_; 
wire _abc_19873_new_n949_; 
wire _abc_19873_new_n950_; 
wire _abc_19873_new_n952_; 
wire _abc_19873_new_n953_; 
wire _abc_19873_new_n954_; 
wire _abc_19873_new_n955_; 
wire _abc_19873_new_n956_; 
wire _abc_19873_new_n957_; 
wire _abc_19873_new_n958_; 
wire _abc_19873_new_n959_; 
wire _abc_19873_new_n960_; 
wire _abc_19873_new_n960__bF_buf0; 
wire _abc_19873_new_n960__bF_buf1; 
wire _abc_19873_new_n960__bF_buf2; 
wire _abc_19873_new_n960__bF_buf3; 
wire _abc_19873_new_n960__bF_buf4; 
wire _abc_19873_new_n961_; 
wire _abc_19873_new_n962_; 
wire _abc_19873_new_n963_; 
wire _abc_19873_new_n964_; 
wire _abc_19873_new_n965_; 
wire _abc_19873_new_n966_; 
wire _abc_19873_new_n967_; 
wire _abc_19873_new_n968_; 
wire _abc_19873_new_n969_; 
wire _abc_19873_new_n969__bF_buf0; 
wire _abc_19873_new_n969__bF_buf1; 
wire _abc_19873_new_n969__bF_buf2; 
wire _abc_19873_new_n969__bF_buf3; 
wire _abc_19873_new_n970_; 
wire _abc_19873_new_n971_; 
wire _abc_19873_new_n972_; 
wire _abc_19873_new_n973_; 
wire _abc_19873_new_n974_; 
wire _abc_19873_new_n976_; 
wire _abc_19873_new_n977_; 
wire _abc_19873_new_n978_; 
wire _abc_19873_new_n979_; 
wire _abc_19873_new_n980_; 
wire _abc_19873_new_n981_; 
wire _abc_19873_new_n982_; 
wire _abc_19873_new_n983_; 
wire _abc_19873_new_n984_; 
wire _abc_19873_new_n985_; 
wire _abc_19873_new_n986_; 
wire _abc_19873_new_n987_; 
wire _abc_19873_new_n988_; 
wire _abc_19873_new_n989_; 
wire _abc_19873_new_n990_; 
wire _abc_19873_new_n991_; 
wire _abc_19873_new_n992_; 
wire _abc_19873_new_n993_; 
wire _abc_19873_new_n994_; 
wire _abc_19873_new_n995_; 
wire _abc_19873_new_n997_; 
wire _abc_19873_new_n998_; 
wire _abc_19873_new_n999_; 
wire _auto_iopadmap_cc_368_execute_27087_0_; 
wire _auto_iopadmap_cc_368_execute_27087_10_; 
wire _auto_iopadmap_cc_368_execute_27087_11_; 
wire _auto_iopadmap_cc_368_execute_27087_12_; 
wire _auto_iopadmap_cc_368_execute_27087_13_; 
wire _auto_iopadmap_cc_368_execute_27087_14_; 
wire _auto_iopadmap_cc_368_execute_27087_15_; 
wire _auto_iopadmap_cc_368_execute_27087_16_; 
wire _auto_iopadmap_cc_368_execute_27087_17_; 
wire _auto_iopadmap_cc_368_execute_27087_18_; 
wire _auto_iopadmap_cc_368_execute_27087_19_; 
wire _auto_iopadmap_cc_368_execute_27087_1_; 
wire _auto_iopadmap_cc_368_execute_27087_20_; 
wire _auto_iopadmap_cc_368_execute_27087_21_; 
wire _auto_iopadmap_cc_368_execute_27087_22_; 
wire _auto_iopadmap_cc_368_execute_27087_23_; 
wire _auto_iopadmap_cc_368_execute_27087_24_; 
wire _auto_iopadmap_cc_368_execute_27087_25_; 
wire _auto_iopadmap_cc_368_execute_27087_26_; 
wire _auto_iopadmap_cc_368_execute_27087_27_; 
wire _auto_iopadmap_cc_368_execute_27087_28_; 
wire _auto_iopadmap_cc_368_execute_27087_29_; 
wire _auto_iopadmap_cc_368_execute_27087_2_; 
wire _auto_iopadmap_cc_368_execute_27087_30_; 
wire _auto_iopadmap_cc_368_execute_27087_31_; 
wire _auto_iopadmap_cc_368_execute_27087_3_; 
wire _auto_iopadmap_cc_368_execute_27087_4_; 
wire _auto_iopadmap_cc_368_execute_27087_5_; 
wire _auto_iopadmap_cc_368_execute_27087_6_; 
wire _auto_iopadmap_cc_368_execute_27087_7_; 
wire _auto_iopadmap_cc_368_execute_27087_8_; 
wire _auto_iopadmap_cc_368_execute_27087_9_; 
input \addr[0] ;
input \addr[1] ;
input \addr[2] ;
input \addr[3] ;
input \addr[4] ;
input \addr[5] ;
input \addr[6] ;
input \addr[7] ;
input clk;
wire clk_bF_buf0; 
wire clk_bF_buf1; 
wire clk_bF_buf10; 
wire clk_bF_buf11; 
wire clk_bF_buf12; 
wire clk_bF_buf13; 
wire clk_bF_buf14; 
wire clk_bF_buf15; 
wire clk_bF_buf16; 
wire clk_bF_buf17; 
wire clk_bF_buf18; 
wire clk_bF_buf19; 
wire clk_bF_buf2; 
wire clk_bF_buf20; 
wire clk_bF_buf21; 
wire clk_bF_buf22; 
wire clk_bF_buf23; 
wire clk_bF_buf24; 
wire clk_bF_buf25; 
wire clk_bF_buf26; 
wire clk_bF_buf27; 
wire clk_bF_buf28; 
wire clk_bF_buf29; 
wire clk_bF_buf3; 
wire clk_bF_buf30; 
wire clk_bF_buf31; 
wire clk_bF_buf32; 
wire clk_bF_buf33; 
wire clk_bF_buf34; 
wire clk_bF_buf35; 
wire clk_bF_buf36; 
wire clk_bF_buf37; 
wire clk_bF_buf38; 
wire clk_bF_buf39; 
wire clk_bF_buf4; 
wire clk_bF_buf40; 
wire clk_bF_buf41; 
wire clk_bF_buf42; 
wire clk_bF_buf43; 
wire clk_bF_buf44; 
wire clk_bF_buf45; 
wire clk_bF_buf46; 
wire clk_bF_buf47; 
wire clk_bF_buf48; 
wire clk_bF_buf49; 
wire clk_bF_buf5; 
wire clk_bF_buf50; 
wire clk_bF_buf51; 
wire clk_bF_buf52; 
wire clk_bF_buf53; 
wire clk_bF_buf54; 
wire clk_bF_buf55; 
wire clk_bF_buf56; 
wire clk_bF_buf57; 
wire clk_bF_buf58; 
wire clk_bF_buf59; 
wire clk_bF_buf6; 
wire clk_bF_buf60; 
wire clk_bF_buf61; 
wire clk_bF_buf62; 
wire clk_bF_buf63; 
wire clk_bF_buf64; 
wire clk_bF_buf65; 
wire clk_bF_buf66; 
wire clk_bF_buf67; 
wire clk_bF_buf68; 
wire clk_bF_buf69; 
wire clk_bF_buf7; 
wire clk_bF_buf70; 
wire clk_bF_buf71; 
wire clk_bF_buf72; 
wire clk_bF_buf73; 
wire clk_bF_buf74; 
wire clk_bF_buf75; 
wire clk_bF_buf76; 
wire clk_bF_buf77; 
wire clk_bF_buf78; 
wire clk_bF_buf79; 
wire clk_bF_buf8; 
wire clk_bF_buf80; 
wire clk_bF_buf81; 
wire clk_bF_buf82; 
wire clk_bF_buf83; 
wire clk_bF_buf84; 
wire clk_bF_buf9; 
wire clk_hier0_bF_buf0; 
wire clk_hier0_bF_buf1; 
wire clk_hier0_bF_buf2; 
wire clk_hier0_bF_buf3; 
wire clk_hier0_bF_buf4; 
wire clk_hier0_bF_buf5; 
wire clk_hier0_bF_buf6; 
wire clk_hier0_bF_buf7; 
wire clk_hier0_bF_buf8; 
wire core__0loop_ctr_reg_3_0__0_; 
wire core__0loop_ctr_reg_3_0__1_; 
wire core__0loop_ctr_reg_3_0__2_; 
wire core__0loop_ctr_reg_3_0__3_; 
wire core__0mi_reg_63_0__0_; 
wire core__0mi_reg_63_0__10_; 
wire core__0mi_reg_63_0__11_; 
wire core__0mi_reg_63_0__12_; 
wire core__0mi_reg_63_0__13_; 
wire core__0mi_reg_63_0__14_; 
wire core__0mi_reg_63_0__15_; 
wire core__0mi_reg_63_0__16_; 
wire core__0mi_reg_63_0__17_; 
wire core__0mi_reg_63_0__18_; 
wire core__0mi_reg_63_0__19_; 
wire core__0mi_reg_63_0__1_; 
wire core__0mi_reg_63_0__20_; 
wire core__0mi_reg_63_0__21_; 
wire core__0mi_reg_63_0__22_; 
wire core__0mi_reg_63_0__23_; 
wire core__0mi_reg_63_0__24_; 
wire core__0mi_reg_63_0__25_; 
wire core__0mi_reg_63_0__26_; 
wire core__0mi_reg_63_0__27_; 
wire core__0mi_reg_63_0__28_; 
wire core__0mi_reg_63_0__29_; 
wire core__0mi_reg_63_0__2_; 
wire core__0mi_reg_63_0__30_; 
wire core__0mi_reg_63_0__31_; 
wire core__0mi_reg_63_0__32_; 
wire core__0mi_reg_63_0__33_; 
wire core__0mi_reg_63_0__34_; 
wire core__0mi_reg_63_0__35_; 
wire core__0mi_reg_63_0__36_; 
wire core__0mi_reg_63_0__37_; 
wire core__0mi_reg_63_0__38_; 
wire core__0mi_reg_63_0__39_; 
wire core__0mi_reg_63_0__3_; 
wire core__0mi_reg_63_0__40_; 
wire core__0mi_reg_63_0__41_; 
wire core__0mi_reg_63_0__42_; 
wire core__0mi_reg_63_0__43_; 
wire core__0mi_reg_63_0__44_; 
wire core__0mi_reg_63_0__45_; 
wire core__0mi_reg_63_0__46_; 
wire core__0mi_reg_63_0__47_; 
wire core__0mi_reg_63_0__48_; 
wire core__0mi_reg_63_0__49_; 
wire core__0mi_reg_63_0__4_; 
wire core__0mi_reg_63_0__50_; 
wire core__0mi_reg_63_0__51_; 
wire core__0mi_reg_63_0__52_; 
wire core__0mi_reg_63_0__53_; 
wire core__0mi_reg_63_0__54_; 
wire core__0mi_reg_63_0__55_; 
wire core__0mi_reg_63_0__56_; 
wire core__0mi_reg_63_0__57_; 
wire core__0mi_reg_63_0__58_; 
wire core__0mi_reg_63_0__59_; 
wire core__0mi_reg_63_0__5_; 
wire core__0mi_reg_63_0__60_; 
wire core__0mi_reg_63_0__61_; 
wire core__0mi_reg_63_0__62_; 
wire core__0mi_reg_63_0__63_; 
wire core__0mi_reg_63_0__6_; 
wire core__0mi_reg_63_0__7_; 
wire core__0mi_reg_63_0__8_; 
wire core__0mi_reg_63_0__9_; 
wire core__0ready_reg_0_0_; 
wire core__0siphash_valid_reg_0_0_; 
wire core__0siphash_word0_reg_63_0__0_; 
wire core__0siphash_word0_reg_63_0__10_; 
wire core__0siphash_word0_reg_63_0__11_; 
wire core__0siphash_word0_reg_63_0__12_; 
wire core__0siphash_word0_reg_63_0__13_; 
wire core__0siphash_word0_reg_63_0__14_; 
wire core__0siphash_word0_reg_63_0__15_; 
wire core__0siphash_word0_reg_63_0__16_; 
wire core__0siphash_word0_reg_63_0__17_; 
wire core__0siphash_word0_reg_63_0__18_; 
wire core__0siphash_word0_reg_63_0__19_; 
wire core__0siphash_word0_reg_63_0__1_; 
wire core__0siphash_word0_reg_63_0__20_; 
wire core__0siphash_word0_reg_63_0__21_; 
wire core__0siphash_word0_reg_63_0__22_; 
wire core__0siphash_word0_reg_63_0__23_; 
wire core__0siphash_word0_reg_63_0__24_; 
wire core__0siphash_word0_reg_63_0__25_; 
wire core__0siphash_word0_reg_63_0__26_; 
wire core__0siphash_word0_reg_63_0__27_; 
wire core__0siphash_word0_reg_63_0__28_; 
wire core__0siphash_word0_reg_63_0__29_; 
wire core__0siphash_word0_reg_63_0__2_; 
wire core__0siphash_word0_reg_63_0__30_; 
wire core__0siphash_word0_reg_63_0__31_; 
wire core__0siphash_word0_reg_63_0__32_; 
wire core__0siphash_word0_reg_63_0__33_; 
wire core__0siphash_word0_reg_63_0__34_; 
wire core__0siphash_word0_reg_63_0__35_; 
wire core__0siphash_word0_reg_63_0__36_; 
wire core__0siphash_word0_reg_63_0__37_; 
wire core__0siphash_word0_reg_63_0__38_; 
wire core__0siphash_word0_reg_63_0__39_; 
wire core__0siphash_word0_reg_63_0__3_; 
wire core__0siphash_word0_reg_63_0__40_; 
wire core__0siphash_word0_reg_63_0__41_; 
wire core__0siphash_word0_reg_63_0__42_; 
wire core__0siphash_word0_reg_63_0__43_; 
wire core__0siphash_word0_reg_63_0__44_; 
wire core__0siphash_word0_reg_63_0__45_; 
wire core__0siphash_word0_reg_63_0__46_; 
wire core__0siphash_word0_reg_63_0__47_; 
wire core__0siphash_word0_reg_63_0__48_; 
wire core__0siphash_word0_reg_63_0__49_; 
wire core__0siphash_word0_reg_63_0__4_; 
wire core__0siphash_word0_reg_63_0__50_; 
wire core__0siphash_word0_reg_63_0__51_; 
wire core__0siphash_word0_reg_63_0__52_; 
wire core__0siphash_word0_reg_63_0__53_; 
wire core__0siphash_word0_reg_63_0__54_; 
wire core__0siphash_word0_reg_63_0__55_; 
wire core__0siphash_word0_reg_63_0__56_; 
wire core__0siphash_word0_reg_63_0__57_; 
wire core__0siphash_word0_reg_63_0__58_; 
wire core__0siphash_word0_reg_63_0__59_; 
wire core__0siphash_word0_reg_63_0__5_; 
wire core__0siphash_word0_reg_63_0__60_; 
wire core__0siphash_word0_reg_63_0__61_; 
wire core__0siphash_word0_reg_63_0__62_; 
wire core__0siphash_word0_reg_63_0__63_; 
wire core__0siphash_word0_reg_63_0__6_; 
wire core__0siphash_word0_reg_63_0__7_; 
wire core__0siphash_word0_reg_63_0__8_; 
wire core__0siphash_word0_reg_63_0__9_; 
wire core__0siphash_word1_reg_63_0__0_; 
wire core__0siphash_word1_reg_63_0__10_; 
wire core__0siphash_word1_reg_63_0__11_; 
wire core__0siphash_word1_reg_63_0__12_; 
wire core__0siphash_word1_reg_63_0__13_; 
wire core__0siphash_word1_reg_63_0__14_; 
wire core__0siphash_word1_reg_63_0__15_; 
wire core__0siphash_word1_reg_63_0__16_; 
wire core__0siphash_word1_reg_63_0__17_; 
wire core__0siphash_word1_reg_63_0__18_; 
wire core__0siphash_word1_reg_63_0__19_; 
wire core__0siphash_word1_reg_63_0__1_; 
wire core__0siphash_word1_reg_63_0__20_; 
wire core__0siphash_word1_reg_63_0__21_; 
wire core__0siphash_word1_reg_63_0__22_; 
wire core__0siphash_word1_reg_63_0__23_; 
wire core__0siphash_word1_reg_63_0__24_; 
wire core__0siphash_word1_reg_63_0__25_; 
wire core__0siphash_word1_reg_63_0__26_; 
wire core__0siphash_word1_reg_63_0__27_; 
wire core__0siphash_word1_reg_63_0__28_; 
wire core__0siphash_word1_reg_63_0__29_; 
wire core__0siphash_word1_reg_63_0__2_; 
wire core__0siphash_word1_reg_63_0__30_; 
wire core__0siphash_word1_reg_63_0__31_; 
wire core__0siphash_word1_reg_63_0__32_; 
wire core__0siphash_word1_reg_63_0__33_; 
wire core__0siphash_word1_reg_63_0__34_; 
wire core__0siphash_word1_reg_63_0__35_; 
wire core__0siphash_word1_reg_63_0__36_; 
wire core__0siphash_word1_reg_63_0__37_; 
wire core__0siphash_word1_reg_63_0__38_; 
wire core__0siphash_word1_reg_63_0__39_; 
wire core__0siphash_word1_reg_63_0__3_; 
wire core__0siphash_word1_reg_63_0__40_; 
wire core__0siphash_word1_reg_63_0__41_; 
wire core__0siphash_word1_reg_63_0__42_; 
wire core__0siphash_word1_reg_63_0__43_; 
wire core__0siphash_word1_reg_63_0__44_; 
wire core__0siphash_word1_reg_63_0__45_; 
wire core__0siphash_word1_reg_63_0__46_; 
wire core__0siphash_word1_reg_63_0__47_; 
wire core__0siphash_word1_reg_63_0__48_; 
wire core__0siphash_word1_reg_63_0__49_; 
wire core__0siphash_word1_reg_63_0__4_; 
wire core__0siphash_word1_reg_63_0__50_; 
wire core__0siphash_word1_reg_63_0__51_; 
wire core__0siphash_word1_reg_63_0__52_; 
wire core__0siphash_word1_reg_63_0__53_; 
wire core__0siphash_word1_reg_63_0__54_; 
wire core__0siphash_word1_reg_63_0__55_; 
wire core__0siphash_word1_reg_63_0__56_; 
wire core__0siphash_word1_reg_63_0__57_; 
wire core__0siphash_word1_reg_63_0__58_; 
wire core__0siphash_word1_reg_63_0__59_; 
wire core__0siphash_word1_reg_63_0__5_; 
wire core__0siphash_word1_reg_63_0__60_; 
wire core__0siphash_word1_reg_63_0__61_; 
wire core__0siphash_word1_reg_63_0__62_; 
wire core__0siphash_word1_reg_63_0__63_; 
wire core__0siphash_word1_reg_63_0__6_; 
wire core__0siphash_word1_reg_63_0__7_; 
wire core__0siphash_word1_reg_63_0__8_; 
wire core__0siphash_word1_reg_63_0__9_; 
wire core__0v0_reg_63_0__0_; 
wire core__0v0_reg_63_0__10_; 
wire core__0v0_reg_63_0__11_; 
wire core__0v0_reg_63_0__12_; 
wire core__0v0_reg_63_0__13_; 
wire core__0v0_reg_63_0__14_; 
wire core__0v0_reg_63_0__15_; 
wire core__0v0_reg_63_0__16_; 
wire core__0v0_reg_63_0__17_; 
wire core__0v0_reg_63_0__18_; 
wire core__0v0_reg_63_0__19_; 
wire core__0v0_reg_63_0__1_; 
wire core__0v0_reg_63_0__20_; 
wire core__0v0_reg_63_0__21_; 
wire core__0v0_reg_63_0__22_; 
wire core__0v0_reg_63_0__23_; 
wire core__0v0_reg_63_0__24_; 
wire core__0v0_reg_63_0__25_; 
wire core__0v0_reg_63_0__26_; 
wire core__0v0_reg_63_0__27_; 
wire core__0v0_reg_63_0__28_; 
wire core__0v0_reg_63_0__29_; 
wire core__0v0_reg_63_0__2_; 
wire core__0v0_reg_63_0__30_; 
wire core__0v0_reg_63_0__31_; 
wire core__0v0_reg_63_0__32_; 
wire core__0v0_reg_63_0__33_; 
wire core__0v0_reg_63_0__34_; 
wire core__0v0_reg_63_0__35_; 
wire core__0v0_reg_63_0__36_; 
wire core__0v0_reg_63_0__37_; 
wire core__0v0_reg_63_0__38_; 
wire core__0v0_reg_63_0__39_; 
wire core__0v0_reg_63_0__3_; 
wire core__0v0_reg_63_0__40_; 
wire core__0v0_reg_63_0__41_; 
wire core__0v0_reg_63_0__42_; 
wire core__0v0_reg_63_0__43_; 
wire core__0v0_reg_63_0__44_; 
wire core__0v0_reg_63_0__45_; 
wire core__0v0_reg_63_0__46_; 
wire core__0v0_reg_63_0__47_; 
wire core__0v0_reg_63_0__48_; 
wire core__0v0_reg_63_0__49_; 
wire core__0v0_reg_63_0__4_; 
wire core__0v0_reg_63_0__50_; 
wire core__0v0_reg_63_0__51_; 
wire core__0v0_reg_63_0__52_; 
wire core__0v0_reg_63_0__53_; 
wire core__0v0_reg_63_0__54_; 
wire core__0v0_reg_63_0__55_; 
wire core__0v0_reg_63_0__56_; 
wire core__0v0_reg_63_0__57_; 
wire core__0v0_reg_63_0__58_; 
wire core__0v0_reg_63_0__59_; 
wire core__0v0_reg_63_0__5_; 
wire core__0v0_reg_63_0__60_; 
wire core__0v0_reg_63_0__61_; 
wire core__0v0_reg_63_0__62_; 
wire core__0v0_reg_63_0__63_; 
wire core__0v0_reg_63_0__6_; 
wire core__0v0_reg_63_0__7_; 
wire core__0v0_reg_63_0__8_; 
wire core__0v0_reg_63_0__9_; 
wire core__0v1_reg_63_0__0_; 
wire core__0v1_reg_63_0__10_; 
wire core__0v1_reg_63_0__11_; 
wire core__0v1_reg_63_0__12_; 
wire core__0v1_reg_63_0__13_; 
wire core__0v1_reg_63_0__14_; 
wire core__0v1_reg_63_0__15_; 
wire core__0v1_reg_63_0__16_; 
wire core__0v1_reg_63_0__17_; 
wire core__0v1_reg_63_0__18_; 
wire core__0v1_reg_63_0__19_; 
wire core__0v1_reg_63_0__1_; 
wire core__0v1_reg_63_0__20_; 
wire core__0v1_reg_63_0__21_; 
wire core__0v1_reg_63_0__22_; 
wire core__0v1_reg_63_0__23_; 
wire core__0v1_reg_63_0__24_; 
wire core__0v1_reg_63_0__25_; 
wire core__0v1_reg_63_0__26_; 
wire core__0v1_reg_63_0__27_; 
wire core__0v1_reg_63_0__28_; 
wire core__0v1_reg_63_0__29_; 
wire core__0v1_reg_63_0__2_; 
wire core__0v1_reg_63_0__30_; 
wire core__0v1_reg_63_0__31_; 
wire core__0v1_reg_63_0__32_; 
wire core__0v1_reg_63_0__33_; 
wire core__0v1_reg_63_0__34_; 
wire core__0v1_reg_63_0__35_; 
wire core__0v1_reg_63_0__36_; 
wire core__0v1_reg_63_0__37_; 
wire core__0v1_reg_63_0__38_; 
wire core__0v1_reg_63_0__39_; 
wire core__0v1_reg_63_0__3_; 
wire core__0v1_reg_63_0__40_; 
wire core__0v1_reg_63_0__41_; 
wire core__0v1_reg_63_0__42_; 
wire core__0v1_reg_63_0__43_; 
wire core__0v1_reg_63_0__44_; 
wire core__0v1_reg_63_0__45_; 
wire core__0v1_reg_63_0__46_; 
wire core__0v1_reg_63_0__47_; 
wire core__0v1_reg_63_0__48_; 
wire core__0v1_reg_63_0__49_; 
wire core__0v1_reg_63_0__4_; 
wire core__0v1_reg_63_0__50_; 
wire core__0v1_reg_63_0__51_; 
wire core__0v1_reg_63_0__52_; 
wire core__0v1_reg_63_0__53_; 
wire core__0v1_reg_63_0__54_; 
wire core__0v1_reg_63_0__55_; 
wire core__0v1_reg_63_0__56_; 
wire core__0v1_reg_63_0__57_; 
wire core__0v1_reg_63_0__58_; 
wire core__0v1_reg_63_0__59_; 
wire core__0v1_reg_63_0__5_; 
wire core__0v1_reg_63_0__60_; 
wire core__0v1_reg_63_0__61_; 
wire core__0v1_reg_63_0__62_; 
wire core__0v1_reg_63_0__63_; 
wire core__0v1_reg_63_0__6_; 
wire core__0v1_reg_63_0__7_; 
wire core__0v1_reg_63_0__8_; 
wire core__0v1_reg_63_0__9_; 
wire core__0v2_reg_63_0__0_; 
wire core__0v2_reg_63_0__10_; 
wire core__0v2_reg_63_0__11_; 
wire core__0v2_reg_63_0__12_; 
wire core__0v2_reg_63_0__13_; 
wire core__0v2_reg_63_0__14_; 
wire core__0v2_reg_63_0__15_; 
wire core__0v2_reg_63_0__16_; 
wire core__0v2_reg_63_0__17_; 
wire core__0v2_reg_63_0__18_; 
wire core__0v2_reg_63_0__19_; 
wire core__0v2_reg_63_0__1_; 
wire core__0v2_reg_63_0__20_; 
wire core__0v2_reg_63_0__21_; 
wire core__0v2_reg_63_0__22_; 
wire core__0v2_reg_63_0__23_; 
wire core__0v2_reg_63_0__24_; 
wire core__0v2_reg_63_0__25_; 
wire core__0v2_reg_63_0__26_; 
wire core__0v2_reg_63_0__27_; 
wire core__0v2_reg_63_0__28_; 
wire core__0v2_reg_63_0__29_; 
wire core__0v2_reg_63_0__2_; 
wire core__0v2_reg_63_0__30_; 
wire core__0v2_reg_63_0__31_; 
wire core__0v2_reg_63_0__32_; 
wire core__0v2_reg_63_0__33_; 
wire core__0v2_reg_63_0__34_; 
wire core__0v2_reg_63_0__35_; 
wire core__0v2_reg_63_0__36_; 
wire core__0v2_reg_63_0__37_; 
wire core__0v2_reg_63_0__38_; 
wire core__0v2_reg_63_0__39_; 
wire core__0v2_reg_63_0__3_; 
wire core__0v2_reg_63_0__40_; 
wire core__0v2_reg_63_0__41_; 
wire core__0v2_reg_63_0__42_; 
wire core__0v2_reg_63_0__43_; 
wire core__0v2_reg_63_0__44_; 
wire core__0v2_reg_63_0__45_; 
wire core__0v2_reg_63_0__46_; 
wire core__0v2_reg_63_0__47_; 
wire core__0v2_reg_63_0__48_; 
wire core__0v2_reg_63_0__49_; 
wire core__0v2_reg_63_0__4_; 
wire core__0v2_reg_63_0__50_; 
wire core__0v2_reg_63_0__51_; 
wire core__0v2_reg_63_0__52_; 
wire core__0v2_reg_63_0__53_; 
wire core__0v2_reg_63_0__54_; 
wire core__0v2_reg_63_0__55_; 
wire core__0v2_reg_63_0__56_; 
wire core__0v2_reg_63_0__57_; 
wire core__0v2_reg_63_0__58_; 
wire core__0v2_reg_63_0__59_; 
wire core__0v2_reg_63_0__5_; 
wire core__0v2_reg_63_0__60_; 
wire core__0v2_reg_63_0__61_; 
wire core__0v2_reg_63_0__62_; 
wire core__0v2_reg_63_0__63_; 
wire core__0v2_reg_63_0__6_; 
wire core__0v2_reg_63_0__7_; 
wire core__0v2_reg_63_0__8_; 
wire core__0v2_reg_63_0__9_; 
wire core__0v3_reg_63_0__0_; 
wire core__0v3_reg_63_0__10_; 
wire core__0v3_reg_63_0__11_; 
wire core__0v3_reg_63_0__12_; 
wire core__0v3_reg_63_0__13_; 
wire core__0v3_reg_63_0__14_; 
wire core__0v3_reg_63_0__15_; 
wire core__0v3_reg_63_0__16_; 
wire core__0v3_reg_63_0__17_; 
wire core__0v3_reg_63_0__18_; 
wire core__0v3_reg_63_0__19_; 
wire core__0v3_reg_63_0__1_; 
wire core__0v3_reg_63_0__20_; 
wire core__0v3_reg_63_0__21_; 
wire core__0v3_reg_63_0__22_; 
wire core__0v3_reg_63_0__23_; 
wire core__0v3_reg_63_0__24_; 
wire core__0v3_reg_63_0__25_; 
wire core__0v3_reg_63_0__26_; 
wire core__0v3_reg_63_0__27_; 
wire core__0v3_reg_63_0__28_; 
wire core__0v3_reg_63_0__29_; 
wire core__0v3_reg_63_0__2_; 
wire core__0v3_reg_63_0__30_; 
wire core__0v3_reg_63_0__31_; 
wire core__0v3_reg_63_0__32_; 
wire core__0v3_reg_63_0__33_; 
wire core__0v3_reg_63_0__34_; 
wire core__0v3_reg_63_0__35_; 
wire core__0v3_reg_63_0__36_; 
wire core__0v3_reg_63_0__37_; 
wire core__0v3_reg_63_0__38_; 
wire core__0v3_reg_63_0__39_; 
wire core__0v3_reg_63_0__3_; 
wire core__0v3_reg_63_0__40_; 
wire core__0v3_reg_63_0__41_; 
wire core__0v3_reg_63_0__42_; 
wire core__0v3_reg_63_0__43_; 
wire core__0v3_reg_63_0__44_; 
wire core__0v3_reg_63_0__45_; 
wire core__0v3_reg_63_0__46_; 
wire core__0v3_reg_63_0__47_; 
wire core__0v3_reg_63_0__48_; 
wire core__0v3_reg_63_0__49_; 
wire core__0v3_reg_63_0__4_; 
wire core__0v3_reg_63_0__50_; 
wire core__0v3_reg_63_0__51_; 
wire core__0v3_reg_63_0__52_; 
wire core__0v3_reg_63_0__53_; 
wire core__0v3_reg_63_0__54_; 
wire core__0v3_reg_63_0__55_; 
wire core__0v3_reg_63_0__56_; 
wire core__0v3_reg_63_0__57_; 
wire core__0v3_reg_63_0__58_; 
wire core__0v3_reg_63_0__59_; 
wire core__0v3_reg_63_0__5_; 
wire core__0v3_reg_63_0__60_; 
wire core__0v3_reg_63_0__61_; 
wire core__0v3_reg_63_0__62_; 
wire core__0v3_reg_63_0__63_; 
wire core__0v3_reg_63_0__6_; 
wire core__0v3_reg_63_0__7_; 
wire core__0v3_reg_63_0__8_; 
wire core__0v3_reg_63_0__9_; 
wire core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1470; 
wire core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1474; 
wire core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1496; 
wire core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1509; 
wire core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_0_; 
wire core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_3_; 
wire core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_4_; 
wire core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_6_; 
wire core__abc_21302_new_n1130_; 
wire core__abc_21302_new_n1131_; 
wire core__abc_21302_new_n1132_; 
wire core__abc_21302_new_n1133_; 
wire core__abc_21302_new_n1134_; 
wire core__abc_21302_new_n1135_; 
wire core__abc_21302_new_n1136_; 
wire core__abc_21302_new_n1137_; 
wire core__abc_21302_new_n1138_; 
wire core__abc_21302_new_n1139_; 
wire core__abc_21302_new_n1140_; 
wire core__abc_21302_new_n1141_; 
wire core__abc_21302_new_n1142_; 
wire core__abc_21302_new_n1143_; 
wire core__abc_21302_new_n1144_; 
wire core__abc_21302_new_n1145_; 
wire core__abc_21302_new_n1146_; 
wire core__abc_21302_new_n1147_; 
wire core__abc_21302_new_n1148_; 
wire core__abc_21302_new_n1149_; 
wire core__abc_21302_new_n1150_; 
wire core__abc_21302_new_n1151_; 
wire core__abc_21302_new_n1152_; 
wire core__abc_21302_new_n1153_; 
wire core__abc_21302_new_n1154_; 
wire core__abc_21302_new_n1155_; 
wire core__abc_21302_new_n1156_; 
wire core__abc_21302_new_n1157_; 
wire core__abc_21302_new_n1158_; 
wire core__abc_21302_new_n1159_; 
wire core__abc_21302_new_n1160_; 
wire core__abc_21302_new_n1161_; 
wire core__abc_21302_new_n1162_; 
wire core__abc_21302_new_n1163_; 
wire core__abc_21302_new_n1164_; 
wire core__abc_21302_new_n1165_; 
wire core__abc_21302_new_n1166_; 
wire core__abc_21302_new_n1167_; 
wire core__abc_21302_new_n1168_; 
wire core__abc_21302_new_n1169_; 
wire core__abc_21302_new_n1170_; 
wire core__abc_21302_new_n1171_; 
wire core__abc_21302_new_n1172_; 
wire core__abc_21302_new_n1173_; 
wire core__abc_21302_new_n1174_; 
wire core__abc_21302_new_n1175_; 
wire core__abc_21302_new_n1176_; 
wire core__abc_21302_new_n1177_; 
wire core__abc_21302_new_n1178_; 
wire core__abc_21302_new_n1179_; 
wire core__abc_21302_new_n1180_; 
wire core__abc_21302_new_n1181_; 
wire core__abc_21302_new_n1182_; 
wire core__abc_21302_new_n1183_; 
wire core__abc_21302_new_n1184_; 
wire core__abc_21302_new_n1185_; 
wire core__abc_21302_new_n1185__bF_buf0; 
wire core__abc_21302_new_n1185__bF_buf1; 
wire core__abc_21302_new_n1185__bF_buf10; 
wire core__abc_21302_new_n1185__bF_buf11; 
wire core__abc_21302_new_n1185__bF_buf12; 
wire core__abc_21302_new_n1185__bF_buf13; 
wire core__abc_21302_new_n1185__bF_buf2; 
wire core__abc_21302_new_n1185__bF_buf3; 
wire core__abc_21302_new_n1185__bF_buf4; 
wire core__abc_21302_new_n1185__bF_buf5; 
wire core__abc_21302_new_n1185__bF_buf6; 
wire core__abc_21302_new_n1185__bF_buf7; 
wire core__abc_21302_new_n1185__bF_buf8; 
wire core__abc_21302_new_n1185__bF_buf9; 
wire core__abc_21302_new_n1186_; 
wire core__abc_21302_new_n1187_; 
wire core__abc_21302_new_n1188_; 
wire core__abc_21302_new_n1189_; 
wire core__abc_21302_new_n1190_; 
wire core__abc_21302_new_n1191_; 
wire core__abc_21302_new_n1192_; 
wire core__abc_21302_new_n1194_; 
wire core__abc_21302_new_n1195_; 
wire core__abc_21302_new_n1196_; 
wire core__abc_21302_new_n1198_; 
wire core__abc_21302_new_n1199_; 
wire core__abc_21302_new_n1200_; 
wire core__abc_21302_new_n1201_; 
wire core__abc_21302_new_n1203_; 
wire core__abc_21302_new_n1204_; 
wire core__abc_21302_new_n1205_; 
wire core__abc_21302_new_n1206_; 
wire core__abc_21302_new_n1208_; 
wire core__abc_21302_new_n1209_; 
wire core__abc_21302_new_n1210_; 
wire core__abc_21302_new_n1211_; 
wire core__abc_21302_new_n1212_; 
wire core__abc_21302_new_n1213_; 
wire core__abc_21302_new_n1214_; 
wire core__abc_21302_new_n1215_; 
wire core__abc_21302_new_n1216_; 
wire core__abc_21302_new_n1217_; 
wire core__abc_21302_new_n1218_; 
wire core__abc_21302_new_n1220_; 
wire core__abc_21302_new_n1221_; 
wire core__abc_21302_new_n1222_; 
wire core__abc_21302_new_n1223_; 
wire core__abc_21302_new_n1224_; 
wire core__abc_21302_new_n1225_; 
wire core__abc_21302_new_n1226_; 
wire core__abc_21302_new_n1227_; 
wire core__abc_21302_new_n1228_; 
wire core__abc_21302_new_n1229_; 
wire core__abc_21302_new_n1230_; 
wire core__abc_21302_new_n1232_; 
wire core__abc_21302_new_n1233_; 
wire core__abc_21302_new_n1234_; 
wire core__abc_21302_new_n1235_; 
wire core__abc_21302_new_n1236_; 
wire core__abc_21302_new_n1237_; 
wire core__abc_21302_new_n1238_; 
wire core__abc_21302_new_n1239_; 
wire core__abc_21302_new_n1241_; 
wire core__abc_21302_new_n1242_; 
wire core__abc_21302_new_n1243_; 
wire core__abc_21302_new_n1244_; 
wire core__abc_21302_new_n1245_; 
wire core__abc_21302_new_n1246_; 
wire core__abc_21302_new_n1247_; 
wire core__abc_21302_new_n1248_; 
wire core__abc_21302_new_n1249_; 
wire core__abc_21302_new_n1251_; 
wire core__abc_21302_new_n1252_; 
wire core__abc_21302_new_n1253_; 
wire core__abc_21302_new_n1254_; 
wire core__abc_21302_new_n1255_; 
wire core__abc_21302_new_n1256_; 
wire core__abc_21302_new_n1257_; 
wire core__abc_21302_new_n1258_; 
wire core__abc_21302_new_n1259_; 
wire core__abc_21302_new_n1261_; 
wire core__abc_21302_new_n1262_; 
wire core__abc_21302_new_n1263_; 
wire core__abc_21302_new_n1264_; 
wire core__abc_21302_new_n1265_; 
wire core__abc_21302_new_n1266_; 
wire core__abc_21302_new_n1267_; 
wire core__abc_21302_new_n1268_; 
wire core__abc_21302_new_n1269_; 
wire core__abc_21302_new_n1270_; 
wire core__abc_21302_new_n1271_; 
wire core__abc_21302_new_n1273_; 
wire core__abc_21302_new_n1274_; 
wire core__abc_21302_new_n1275_; 
wire core__abc_21302_new_n1276_; 
wire core__abc_21302_new_n1277_; 
wire core__abc_21302_new_n1278_; 
wire core__abc_21302_new_n1279_; 
wire core__abc_21302_new_n1280_; 
wire core__abc_21302_new_n1281_; 
wire core__abc_21302_new_n1283_; 
wire core__abc_21302_new_n1284_; 
wire core__abc_21302_new_n1285_; 
wire core__abc_21302_new_n1286_; 
wire core__abc_21302_new_n1287_; 
wire core__abc_21302_new_n1288_; 
wire core__abc_21302_new_n1289_; 
wire core__abc_21302_new_n1290_; 
wire core__abc_21302_new_n1291_; 
wire core__abc_21302_new_n1293_; 
wire core__abc_21302_new_n1294_; 
wire core__abc_21302_new_n1295_; 
wire core__abc_21302_new_n1296_; 
wire core__abc_21302_new_n1297_; 
wire core__abc_21302_new_n1298_; 
wire core__abc_21302_new_n1299_; 
wire core__abc_21302_new_n1301_; 
wire core__abc_21302_new_n1302_; 
wire core__abc_21302_new_n1303_; 
wire core__abc_21302_new_n1304_; 
wire core__abc_21302_new_n1305_; 
wire core__abc_21302_new_n1306_; 
wire core__abc_21302_new_n1307_; 
wire core__abc_21302_new_n1308_; 
wire core__abc_21302_new_n1309_; 
wire core__abc_21302_new_n1310_; 
wire core__abc_21302_new_n1312_; 
wire core__abc_21302_new_n1313_; 
wire core__abc_21302_new_n1314_; 
wire core__abc_21302_new_n1315_; 
wire core__abc_21302_new_n1316_; 
wire core__abc_21302_new_n1317_; 
wire core__abc_21302_new_n1318_; 
wire core__abc_21302_new_n1319_; 
wire core__abc_21302_new_n1320_; 
wire core__abc_21302_new_n1321_; 
wire core__abc_21302_new_n1322_; 
wire core__abc_21302_new_n1324_; 
wire core__abc_21302_new_n1325_; 
wire core__abc_21302_new_n1326_; 
wire core__abc_21302_new_n1327_; 
wire core__abc_21302_new_n1328_; 
wire core__abc_21302_new_n1329_; 
wire core__abc_21302_new_n1330_; 
wire core__abc_21302_new_n1331_; 
wire core__abc_21302_new_n1332_; 
wire core__abc_21302_new_n1333_; 
wire core__abc_21302_new_n1334_; 
wire core__abc_21302_new_n1336_; 
wire core__abc_21302_new_n1337_; 
wire core__abc_21302_new_n1338_; 
wire core__abc_21302_new_n1339_; 
wire core__abc_21302_new_n1340_; 
wire core__abc_21302_new_n1341_; 
wire core__abc_21302_new_n1342_; 
wire core__abc_21302_new_n1343_; 
wire core__abc_21302_new_n1344_; 
wire core__abc_21302_new_n1346_; 
wire core__abc_21302_new_n1347_; 
wire core__abc_21302_new_n1348_; 
wire core__abc_21302_new_n1349_; 
wire core__abc_21302_new_n1350_; 
wire core__abc_21302_new_n1351_; 
wire core__abc_21302_new_n1352_; 
wire core__abc_21302_new_n1353_; 
wire core__abc_21302_new_n1354_; 
wire core__abc_21302_new_n1355_; 
wire core__abc_21302_new_n1356_; 
wire core__abc_21302_new_n1358_; 
wire core__abc_21302_new_n1359_; 
wire core__abc_21302_new_n1360_; 
wire core__abc_21302_new_n1361_; 
wire core__abc_21302_new_n1362_; 
wire core__abc_21302_new_n1363_; 
wire core__abc_21302_new_n1364_; 
wire core__abc_21302_new_n1365_; 
wire core__abc_21302_new_n1366_; 
wire core__abc_21302_new_n1367_; 
wire core__abc_21302_new_n1368_; 
wire core__abc_21302_new_n1370_; 
wire core__abc_21302_new_n1371_; 
wire core__abc_21302_new_n1372_; 
wire core__abc_21302_new_n1373_; 
wire core__abc_21302_new_n1374_; 
wire core__abc_21302_new_n1375_; 
wire core__abc_21302_new_n1376_; 
wire core__abc_21302_new_n1377_; 
wire core__abc_21302_new_n1378_; 
wire core__abc_21302_new_n1379_; 
wire core__abc_21302_new_n1380_; 
wire core__abc_21302_new_n1382_; 
wire core__abc_21302_new_n1383_; 
wire core__abc_21302_new_n1384_; 
wire core__abc_21302_new_n1385_; 
wire core__abc_21302_new_n1386_; 
wire core__abc_21302_new_n1387_; 
wire core__abc_21302_new_n1388_; 
wire core__abc_21302_new_n1389_; 
wire core__abc_21302_new_n1390_; 
wire core__abc_21302_new_n1391_; 
wire core__abc_21302_new_n1393_; 
wire core__abc_21302_new_n1394_; 
wire core__abc_21302_new_n1395_; 
wire core__abc_21302_new_n1396_; 
wire core__abc_21302_new_n1397_; 
wire core__abc_21302_new_n1398_; 
wire core__abc_21302_new_n1399_; 
wire core__abc_21302_new_n1400_; 
wire core__abc_21302_new_n1401_; 
wire core__abc_21302_new_n1402_; 
wire core__abc_21302_new_n1403_; 
wire core__abc_21302_new_n1405_; 
wire core__abc_21302_new_n1406_; 
wire core__abc_21302_new_n1407_; 
wire core__abc_21302_new_n1408_; 
wire core__abc_21302_new_n1409_; 
wire core__abc_21302_new_n1410_; 
wire core__abc_21302_new_n1411_; 
wire core__abc_21302_new_n1412_; 
wire core__abc_21302_new_n1413_; 
wire core__abc_21302_new_n1414_; 
wire core__abc_21302_new_n1415_; 
wire core__abc_21302_new_n1417_; 
wire core__abc_21302_new_n1418_; 
wire core__abc_21302_new_n1419_; 
wire core__abc_21302_new_n1420_; 
wire core__abc_21302_new_n1421_; 
wire core__abc_21302_new_n1422_; 
wire core__abc_21302_new_n1423_; 
wire core__abc_21302_new_n1424_; 
wire core__abc_21302_new_n1425_; 
wire core__abc_21302_new_n1426_; 
wire core__abc_21302_new_n1427_; 
wire core__abc_21302_new_n1429_; 
wire core__abc_21302_new_n1430_; 
wire core__abc_21302_new_n1431_; 
wire core__abc_21302_new_n1432_; 
wire core__abc_21302_new_n1433_; 
wire core__abc_21302_new_n1434_; 
wire core__abc_21302_new_n1435_; 
wire core__abc_21302_new_n1436_; 
wire core__abc_21302_new_n1437_; 
wire core__abc_21302_new_n1438_; 
wire core__abc_21302_new_n1439_; 
wire core__abc_21302_new_n1441_; 
wire core__abc_21302_new_n1442_; 
wire core__abc_21302_new_n1443_; 
wire core__abc_21302_new_n1444_; 
wire core__abc_21302_new_n1445_; 
wire core__abc_21302_new_n1446_; 
wire core__abc_21302_new_n1447_; 
wire core__abc_21302_new_n1448_; 
wire core__abc_21302_new_n1449_; 
wire core__abc_21302_new_n1450_; 
wire core__abc_21302_new_n1451_; 
wire core__abc_21302_new_n1453_; 
wire core__abc_21302_new_n1454_; 
wire core__abc_21302_new_n1455_; 
wire core__abc_21302_new_n1456_; 
wire core__abc_21302_new_n1457_; 
wire core__abc_21302_new_n1458_; 
wire core__abc_21302_new_n1459_; 
wire core__abc_21302_new_n1460_; 
wire core__abc_21302_new_n1461_; 
wire core__abc_21302_new_n1462_; 
wire core__abc_21302_new_n1463_; 
wire core__abc_21302_new_n1465_; 
wire core__abc_21302_new_n1466_; 
wire core__abc_21302_new_n1467_; 
wire core__abc_21302_new_n1468_; 
wire core__abc_21302_new_n1469_; 
wire core__abc_21302_new_n1470_; 
wire core__abc_21302_new_n1471_; 
wire core__abc_21302_new_n1473_; 
wire core__abc_21302_new_n1474_; 
wire core__abc_21302_new_n1475_; 
wire core__abc_21302_new_n1476_; 
wire core__abc_21302_new_n1477_; 
wire core__abc_21302_new_n1478_; 
wire core__abc_21302_new_n1479_; 
wire core__abc_21302_new_n1480_; 
wire core__abc_21302_new_n1481_; 
wire core__abc_21302_new_n1482_; 
wire core__abc_21302_new_n1483_; 
wire core__abc_21302_new_n1485_; 
wire core__abc_21302_new_n1486_; 
wire core__abc_21302_new_n1487_; 
wire core__abc_21302_new_n1488_; 
wire core__abc_21302_new_n1489_; 
wire core__abc_21302_new_n1490_; 
wire core__abc_21302_new_n1491_; 
wire core__abc_21302_new_n1492_; 
wire core__abc_21302_new_n1493_; 
wire core__abc_21302_new_n1495_; 
wire core__abc_21302_new_n1496_; 
wire core__abc_21302_new_n1497_; 
wire core__abc_21302_new_n1498_; 
wire core__abc_21302_new_n1499_; 
wire core__abc_21302_new_n1500_; 
wire core__abc_21302_new_n1501_; 
wire core__abc_21302_new_n1502_; 
wire core__abc_21302_new_n1503_; 
wire core__abc_21302_new_n1504_; 
wire core__abc_21302_new_n1505_; 
wire core__abc_21302_new_n1507_; 
wire core__abc_21302_new_n1508_; 
wire core__abc_21302_new_n1509_; 
wire core__abc_21302_new_n1510_; 
wire core__abc_21302_new_n1511_; 
wire core__abc_21302_new_n1512_; 
wire core__abc_21302_new_n1513_; 
wire core__abc_21302_new_n1514_; 
wire core__abc_21302_new_n1515_; 
wire core__abc_21302_new_n1516_; 
wire core__abc_21302_new_n1517_; 
wire core__abc_21302_new_n1519_; 
wire core__abc_21302_new_n1520_; 
wire core__abc_21302_new_n1521_; 
wire core__abc_21302_new_n1522_; 
wire core__abc_21302_new_n1523_; 
wire core__abc_21302_new_n1524_; 
wire core__abc_21302_new_n1525_; 
wire core__abc_21302_new_n1526_; 
wire core__abc_21302_new_n1527_; 
wire core__abc_21302_new_n1528_; 
wire core__abc_21302_new_n1529_; 
wire core__abc_21302_new_n1531_; 
wire core__abc_21302_new_n1532_; 
wire core__abc_21302_new_n1533_; 
wire core__abc_21302_new_n1534_; 
wire core__abc_21302_new_n1535_; 
wire core__abc_21302_new_n1536_; 
wire core__abc_21302_new_n1537_; 
wire core__abc_21302_new_n1538_; 
wire core__abc_21302_new_n1539_; 
wire core__abc_21302_new_n1540_; 
wire core__abc_21302_new_n1541_; 
wire core__abc_21302_new_n1542_; 
wire core__abc_21302_new_n1544_; 
wire core__abc_21302_new_n1545_; 
wire core__abc_21302_new_n1546_; 
wire core__abc_21302_new_n1547_; 
wire core__abc_21302_new_n1548_; 
wire core__abc_21302_new_n1549_; 
wire core__abc_21302_new_n1550_; 
wire core__abc_21302_new_n1551_; 
wire core__abc_21302_new_n1552_; 
wire core__abc_21302_new_n1553_; 
wire core__abc_21302_new_n1554_; 
wire core__abc_21302_new_n1556_; 
wire core__abc_21302_new_n1557_; 
wire core__abc_21302_new_n1558_; 
wire core__abc_21302_new_n1559_; 
wire core__abc_21302_new_n1560_; 
wire core__abc_21302_new_n1561_; 
wire core__abc_21302_new_n1562_; 
wire core__abc_21302_new_n1564_; 
wire core__abc_21302_new_n1565_; 
wire core__abc_21302_new_n1566_; 
wire core__abc_21302_new_n1567_; 
wire core__abc_21302_new_n1568_; 
wire core__abc_21302_new_n1569_; 
wire core__abc_21302_new_n1570_; 
wire core__abc_21302_new_n1571_; 
wire core__abc_21302_new_n1572_; 
wire core__abc_21302_new_n1573_; 
wire core__abc_21302_new_n1574_; 
wire core__abc_21302_new_n1576_; 
wire core__abc_21302_new_n1577_; 
wire core__abc_21302_new_n1578_; 
wire core__abc_21302_new_n1579_; 
wire core__abc_21302_new_n1580_; 
wire core__abc_21302_new_n1581_; 
wire core__abc_21302_new_n1582_; 
wire core__abc_21302_new_n1583_; 
wire core__abc_21302_new_n1584_; 
wire core__abc_21302_new_n1585_; 
wire core__abc_21302_new_n1586_; 
wire core__abc_21302_new_n1588_; 
wire core__abc_21302_new_n1589_; 
wire core__abc_21302_new_n1590_; 
wire core__abc_21302_new_n1591_; 
wire core__abc_21302_new_n1592_; 
wire core__abc_21302_new_n1593_; 
wire core__abc_21302_new_n1594_; 
wire core__abc_21302_new_n1595_; 
wire core__abc_21302_new_n1596_; 
wire core__abc_21302_new_n1597_; 
wire core__abc_21302_new_n1598_; 
wire core__abc_21302_new_n1599_; 
wire core__abc_21302_new_n1600_; 
wire core__abc_21302_new_n1602_; 
wire core__abc_21302_new_n1603_; 
wire core__abc_21302_new_n1604_; 
wire core__abc_21302_new_n1605_; 
wire core__abc_21302_new_n1606_; 
wire core__abc_21302_new_n1607_; 
wire core__abc_21302_new_n1608_; 
wire core__abc_21302_new_n1609_; 
wire core__abc_21302_new_n1610_; 
wire core__abc_21302_new_n1611_; 
wire core__abc_21302_new_n1612_; 
wire core__abc_21302_new_n1614_; 
wire core__abc_21302_new_n1615_; 
wire core__abc_21302_new_n1616_; 
wire core__abc_21302_new_n1617_; 
wire core__abc_21302_new_n1618_; 
wire core__abc_21302_new_n1619_; 
wire core__abc_21302_new_n1620_; 
wire core__abc_21302_new_n1621_; 
wire core__abc_21302_new_n1622_; 
wire core__abc_21302_new_n1623_; 
wire core__abc_21302_new_n1625_; 
wire core__abc_21302_new_n1626_; 
wire core__abc_21302_new_n1627_; 
wire core__abc_21302_new_n1628_; 
wire core__abc_21302_new_n1629_; 
wire core__abc_21302_new_n1630_; 
wire core__abc_21302_new_n1631_; 
wire core__abc_21302_new_n1632_; 
wire core__abc_21302_new_n1633_; 
wire core__abc_21302_new_n1634_; 
wire core__abc_21302_new_n1635_; 
wire core__abc_21302_new_n1636_; 
wire core__abc_21302_new_n1638_; 
wire core__abc_21302_new_n1639_; 
wire core__abc_21302_new_n1640_; 
wire core__abc_21302_new_n1641_; 
wire core__abc_21302_new_n1642_; 
wire core__abc_21302_new_n1643_; 
wire core__abc_21302_new_n1644_; 
wire core__abc_21302_new_n1645_; 
wire core__abc_21302_new_n1647_; 
wire core__abc_21302_new_n1648_; 
wire core__abc_21302_new_n1649_; 
wire core__abc_21302_new_n1650_; 
wire core__abc_21302_new_n1651_; 
wire core__abc_21302_new_n1652_; 
wire core__abc_21302_new_n1653_; 
wire core__abc_21302_new_n1654_; 
wire core__abc_21302_new_n1655_; 
wire core__abc_21302_new_n1656_; 
wire core__abc_21302_new_n1658_; 
wire core__abc_21302_new_n1659_; 
wire core__abc_21302_new_n1660_; 
wire core__abc_21302_new_n1661_; 
wire core__abc_21302_new_n1662_; 
wire core__abc_21302_new_n1663_; 
wire core__abc_21302_new_n1664_; 
wire core__abc_21302_new_n1665_; 
wire core__abc_21302_new_n1666_; 
wire core__abc_21302_new_n1667_; 
wire core__abc_21302_new_n1669_; 
wire core__abc_21302_new_n1670_; 
wire core__abc_21302_new_n1671_; 
wire core__abc_21302_new_n1672_; 
wire core__abc_21302_new_n1673_; 
wire core__abc_21302_new_n1674_; 
wire core__abc_21302_new_n1675_; 
wire core__abc_21302_new_n1676_; 
wire core__abc_21302_new_n1677_; 
wire core__abc_21302_new_n1678_; 
wire core__abc_21302_new_n1680_; 
wire core__abc_21302_new_n1681_; 
wire core__abc_21302_new_n1682_; 
wire core__abc_21302_new_n1683_; 
wire core__abc_21302_new_n1684_; 
wire core__abc_21302_new_n1685_; 
wire core__abc_21302_new_n1686_; 
wire core__abc_21302_new_n1687_; 
wire core__abc_21302_new_n1688_; 
wire core__abc_21302_new_n1689_; 
wire core__abc_21302_new_n1691_; 
wire core__abc_21302_new_n1692_; 
wire core__abc_21302_new_n1693_; 
wire core__abc_21302_new_n1694_; 
wire core__abc_21302_new_n1695_; 
wire core__abc_21302_new_n1696_; 
wire core__abc_21302_new_n1697_; 
wire core__abc_21302_new_n1698_; 
wire core__abc_21302_new_n1699_; 
wire core__abc_21302_new_n1700_; 
wire core__abc_21302_new_n1702_; 
wire core__abc_21302_new_n1703_; 
wire core__abc_21302_new_n1704_; 
wire core__abc_21302_new_n1705_; 
wire core__abc_21302_new_n1706_; 
wire core__abc_21302_new_n1707_; 
wire core__abc_21302_new_n1708_; 
wire core__abc_21302_new_n1709_; 
wire core__abc_21302_new_n1710_; 
wire core__abc_21302_new_n1711_; 
wire core__abc_21302_new_n1712_; 
wire core__abc_21302_new_n1714_; 
wire core__abc_21302_new_n1715_; 
wire core__abc_21302_new_n1716_; 
wire core__abc_21302_new_n1717_; 
wire core__abc_21302_new_n1718_; 
wire core__abc_21302_new_n1719_; 
wire core__abc_21302_new_n1720_; 
wire core__abc_21302_new_n1721_; 
wire core__abc_21302_new_n1722_; 
wire core__abc_21302_new_n1723_; 
wire core__abc_21302_new_n1725_; 
wire core__abc_21302_new_n1726_; 
wire core__abc_21302_new_n1727_; 
wire core__abc_21302_new_n1728_; 
wire core__abc_21302_new_n1729_; 
wire core__abc_21302_new_n1730_; 
wire core__abc_21302_new_n1731_; 
wire core__abc_21302_new_n1732_; 
wire core__abc_21302_new_n1733_; 
wire core__abc_21302_new_n1734_; 
wire core__abc_21302_new_n1735_; 
wire core__abc_21302_new_n1737_; 
wire core__abc_21302_new_n1738_; 
wire core__abc_21302_new_n1739_; 
wire core__abc_21302_new_n1740_; 
wire core__abc_21302_new_n1741_; 
wire core__abc_21302_new_n1742_; 
wire core__abc_21302_new_n1743_; 
wire core__abc_21302_new_n1744_; 
wire core__abc_21302_new_n1745_; 
wire core__abc_21302_new_n1746_; 
wire core__abc_21302_new_n1748_; 
wire core__abc_21302_new_n1749_; 
wire core__abc_21302_new_n1750_; 
wire core__abc_21302_new_n1751_; 
wire core__abc_21302_new_n1752_; 
wire core__abc_21302_new_n1753_; 
wire core__abc_21302_new_n1754_; 
wire core__abc_21302_new_n1755_; 
wire core__abc_21302_new_n1756_; 
wire core__abc_21302_new_n1757_; 
wire core__abc_21302_new_n1758_; 
wire core__abc_21302_new_n1759_; 
wire core__abc_21302_new_n1761_; 
wire core__abc_21302_new_n1762_; 
wire core__abc_21302_new_n1763_; 
wire core__abc_21302_new_n1764_; 
wire core__abc_21302_new_n1765_; 
wire core__abc_21302_new_n1766_; 
wire core__abc_21302_new_n1767_; 
wire core__abc_21302_new_n1768_; 
wire core__abc_21302_new_n1770_; 
wire core__abc_21302_new_n1771_; 
wire core__abc_21302_new_n1772_; 
wire core__abc_21302_new_n1773_; 
wire core__abc_21302_new_n1774_; 
wire core__abc_21302_new_n1775_; 
wire core__abc_21302_new_n1776_; 
wire core__abc_21302_new_n1777_; 
wire core__abc_21302_new_n1778_; 
wire core__abc_21302_new_n1779_; 
wire core__abc_21302_new_n1780_; 
wire core__abc_21302_new_n1782_; 
wire core__abc_21302_new_n1783_; 
wire core__abc_21302_new_n1784_; 
wire core__abc_21302_new_n1785_; 
wire core__abc_21302_new_n1786_; 
wire core__abc_21302_new_n1787_; 
wire core__abc_21302_new_n1788_; 
wire core__abc_21302_new_n1789_; 
wire core__abc_21302_new_n1790_; 
wire core__abc_21302_new_n1791_; 
wire core__abc_21302_new_n1793_; 
wire core__abc_21302_new_n1794_; 
wire core__abc_21302_new_n1795_; 
wire core__abc_21302_new_n1796_; 
wire core__abc_21302_new_n1797_; 
wire core__abc_21302_new_n1798_; 
wire core__abc_21302_new_n1799_; 
wire core__abc_21302_new_n1800_; 
wire core__abc_21302_new_n1801_; 
wire core__abc_21302_new_n1802_; 
wire core__abc_21302_new_n1803_; 
wire core__abc_21302_new_n1804_; 
wire core__abc_21302_new_n1805_; 
wire core__abc_21302_new_n1807_; 
wire core__abc_21302_new_n1808_; 
wire core__abc_21302_new_n1809_; 
wire core__abc_21302_new_n1810_; 
wire core__abc_21302_new_n1811_; 
wire core__abc_21302_new_n1812_; 
wire core__abc_21302_new_n1813_; 
wire core__abc_21302_new_n1814_; 
wire core__abc_21302_new_n1815_; 
wire core__abc_21302_new_n1816_; 
wire core__abc_21302_new_n1818_; 
wire core__abc_21302_new_n1819_; 
wire core__abc_21302_new_n1820_; 
wire core__abc_21302_new_n1821_; 
wire core__abc_21302_new_n1822_; 
wire core__abc_21302_new_n1823_; 
wire core__abc_21302_new_n1824_; 
wire core__abc_21302_new_n1825_; 
wire core__abc_21302_new_n1826_; 
wire core__abc_21302_new_n1827_; 
wire core__abc_21302_new_n1828_; 
wire core__abc_21302_new_n1829_; 
wire core__abc_21302_new_n1831_; 
wire core__abc_21302_new_n1832_; 
wire core__abc_21302_new_n1833_; 
wire core__abc_21302_new_n1834_; 
wire core__abc_21302_new_n1835_; 
wire core__abc_21302_new_n1836_; 
wire core__abc_21302_new_n1837_; 
wire core__abc_21302_new_n1838_; 
wire core__abc_21302_new_n1839_; 
wire core__abc_21302_new_n1840_; 
wire core__abc_21302_new_n1841_; 
wire core__abc_21302_new_n1842_; 
wire core__abc_21302_new_n1844_; 
wire core__abc_21302_new_n1845_; 
wire core__abc_21302_new_n1846_; 
wire core__abc_21302_new_n1847_; 
wire core__abc_21302_new_n1848_; 
wire core__abc_21302_new_n1849_; 
wire core__abc_21302_new_n1850_; 
wire core__abc_21302_new_n1851_; 
wire core__abc_21302_new_n1852_; 
wire core__abc_21302_new_n1853_; 
wire core__abc_21302_new_n1854_; 
wire core__abc_21302_new_n1855_; 
wire core__abc_21302_new_n1856_; 
wire core__abc_21302_new_n1858_; 
wire core__abc_21302_new_n1859_; 
wire core__abc_21302_new_n1860_; 
wire core__abc_21302_new_n1861_; 
wire core__abc_21302_new_n1862_; 
wire core__abc_21302_new_n1863_; 
wire core__abc_21302_new_n1864_; 
wire core__abc_21302_new_n1865_; 
wire core__abc_21302_new_n1866_; 
wire core__abc_21302_new_n1867_; 
wire core__abc_21302_new_n1868_; 
wire core__abc_21302_new_n1870_; 
wire core__abc_21302_new_n1871_; 
wire core__abc_21302_new_n1872_; 
wire core__abc_21302_new_n1873_; 
wire core__abc_21302_new_n1874_; 
wire core__abc_21302_new_n1875_; 
wire core__abc_21302_new_n1876_; 
wire core__abc_21302_new_n1877_; 
wire core__abc_21302_new_n1878_; 
wire core__abc_21302_new_n1879_; 
wire core__abc_21302_new_n1880_; 
wire core__abc_21302_new_n1881_; 
wire core__abc_21302_new_n1882_; 
wire core__abc_21302_new_n1884_; 
wire core__abc_21302_new_n1885_; 
wire core__abc_21302_new_n1886_; 
wire core__abc_21302_new_n1887_; 
wire core__abc_21302_new_n1888_; 
wire core__abc_21302_new_n1889_; 
wire core__abc_21302_new_n1890_; 
wire core__abc_21302_new_n1891_; 
wire core__abc_21302_new_n1892_; 
wire core__abc_21302_new_n1893_; 
wire core__abc_21302_new_n1894_; 
wire core__abc_21302_new_n1896_; 
wire core__abc_21302_new_n1897_; 
wire core__abc_21302_new_n1898_; 
wire core__abc_21302_new_n1899_; 
wire core__abc_21302_new_n1900_; 
wire core__abc_21302_new_n1901_; 
wire core__abc_21302_new_n1902_; 
wire core__abc_21302_new_n1903_; 
wire core__abc_21302_new_n1904_; 
wire core__abc_21302_new_n1905_; 
wire core__abc_21302_new_n1906_; 
wire core__abc_21302_new_n1907_; 
wire core__abc_21302_new_n1908_; 
wire core__abc_21302_new_n1910_; 
wire core__abc_21302_new_n1911_; 
wire core__abc_21302_new_n1912_; 
wire core__abc_21302_new_n1913_; 
wire core__abc_21302_new_n1914_; 
wire core__abc_21302_new_n1915_; 
wire core__abc_21302_new_n1916_; 
wire core__abc_21302_new_n1917_; 
wire core__abc_21302_new_n1918_; 
wire core__abc_21302_new_n1919_; 
wire core__abc_21302_new_n1920_; 
wire core__abc_21302_new_n1921_; 
wire core__abc_21302_new_n1922_; 
wire core__abc_21302_new_n1924_; 
wire core__abc_21302_new_n1925_; 
wire core__abc_21302_new_n1926_; 
wire core__abc_21302_new_n1927_; 
wire core__abc_21302_new_n1928_; 
wire core__abc_21302_new_n1929_; 
wire core__abc_21302_new_n1930_; 
wire core__abc_21302_new_n1931_; 
wire core__abc_21302_new_n1932_; 
wire core__abc_21302_new_n1933_; 
wire core__abc_21302_new_n1934_; 
wire core__abc_21302_new_n1935_; 
wire core__abc_21302_new_n1937_; 
wire core__abc_21302_new_n1938_; 
wire core__abc_21302_new_n1939_; 
wire core__abc_21302_new_n1940_; 
wire core__abc_21302_new_n1941_; 
wire core__abc_21302_new_n1943_; 
wire core__abc_21302_new_n1944_; 
wire core__abc_21302_new_n1945_; 
wire core__abc_21302_new_n1945__bF_buf0; 
wire core__abc_21302_new_n1945__bF_buf1; 
wire core__abc_21302_new_n1945__bF_buf10; 
wire core__abc_21302_new_n1945__bF_buf2; 
wire core__abc_21302_new_n1945__bF_buf3; 
wire core__abc_21302_new_n1945__bF_buf4; 
wire core__abc_21302_new_n1945__bF_buf5; 
wire core__abc_21302_new_n1945__bF_buf6; 
wire core__abc_21302_new_n1945__bF_buf7; 
wire core__abc_21302_new_n1945__bF_buf8; 
wire core__abc_21302_new_n1945__bF_buf9; 
wire core__abc_21302_new_n1946_; 
wire core__abc_21302_new_n1947_; 
wire core__abc_21302_new_n1949_; 
wire core__abc_21302_new_n1950_; 
wire core__abc_21302_new_n1952_; 
wire core__abc_21302_new_n1953_; 
wire core__abc_21302_new_n1955_; 
wire core__abc_21302_new_n1956_; 
wire core__abc_21302_new_n1958_; 
wire core__abc_21302_new_n1959_; 
wire core__abc_21302_new_n1961_; 
wire core__abc_21302_new_n1962_; 
wire core__abc_21302_new_n1964_; 
wire core__abc_21302_new_n1965_; 
wire core__abc_21302_new_n1967_; 
wire core__abc_21302_new_n1968_; 
wire core__abc_21302_new_n1970_; 
wire core__abc_21302_new_n1971_; 
wire core__abc_21302_new_n1973_; 
wire core__abc_21302_new_n1974_; 
wire core__abc_21302_new_n1976_; 
wire core__abc_21302_new_n1977_; 
wire core__abc_21302_new_n1979_; 
wire core__abc_21302_new_n1980_; 
wire core__abc_21302_new_n1982_; 
wire core__abc_21302_new_n1983_; 
wire core__abc_21302_new_n1985_; 
wire core__abc_21302_new_n1986_; 
wire core__abc_21302_new_n1988_; 
wire core__abc_21302_new_n1989_; 
wire core__abc_21302_new_n1991_; 
wire core__abc_21302_new_n1992_; 
wire core__abc_21302_new_n1994_; 
wire core__abc_21302_new_n1995_; 
wire core__abc_21302_new_n1997_; 
wire core__abc_21302_new_n1998_; 
wire core__abc_21302_new_n2000_; 
wire core__abc_21302_new_n2001_; 
wire core__abc_21302_new_n2003_; 
wire core__abc_21302_new_n2004_; 
wire core__abc_21302_new_n2006_; 
wire core__abc_21302_new_n2007_; 
wire core__abc_21302_new_n2009_; 
wire core__abc_21302_new_n2010_; 
wire core__abc_21302_new_n2012_; 
wire core__abc_21302_new_n2013_; 
wire core__abc_21302_new_n2015_; 
wire core__abc_21302_new_n2016_; 
wire core__abc_21302_new_n2018_; 
wire core__abc_21302_new_n2019_; 
wire core__abc_21302_new_n2021_; 
wire core__abc_21302_new_n2022_; 
wire core__abc_21302_new_n2024_; 
wire core__abc_21302_new_n2025_; 
wire core__abc_21302_new_n2027_; 
wire core__abc_21302_new_n2028_; 
wire core__abc_21302_new_n2030_; 
wire core__abc_21302_new_n2031_; 
wire core__abc_21302_new_n2033_; 
wire core__abc_21302_new_n2034_; 
wire core__abc_21302_new_n2036_; 
wire core__abc_21302_new_n2037_; 
wire core__abc_21302_new_n2039_; 
wire core__abc_21302_new_n2040_; 
wire core__abc_21302_new_n2042_; 
wire core__abc_21302_new_n2043_; 
wire core__abc_21302_new_n2045_; 
wire core__abc_21302_new_n2046_; 
wire core__abc_21302_new_n2048_; 
wire core__abc_21302_new_n2049_; 
wire core__abc_21302_new_n2051_; 
wire core__abc_21302_new_n2052_; 
wire core__abc_21302_new_n2054_; 
wire core__abc_21302_new_n2055_; 
wire core__abc_21302_new_n2057_; 
wire core__abc_21302_new_n2058_; 
wire core__abc_21302_new_n2060_; 
wire core__abc_21302_new_n2061_; 
wire core__abc_21302_new_n2063_; 
wire core__abc_21302_new_n2064_; 
wire core__abc_21302_new_n2066_; 
wire core__abc_21302_new_n2067_; 
wire core__abc_21302_new_n2069_; 
wire core__abc_21302_new_n2070_; 
wire core__abc_21302_new_n2072_; 
wire core__abc_21302_new_n2073_; 
wire core__abc_21302_new_n2075_; 
wire core__abc_21302_new_n2076_; 
wire core__abc_21302_new_n2078_; 
wire core__abc_21302_new_n2079_; 
wire core__abc_21302_new_n2081_; 
wire core__abc_21302_new_n2082_; 
wire core__abc_21302_new_n2084_; 
wire core__abc_21302_new_n2085_; 
wire core__abc_21302_new_n2087_; 
wire core__abc_21302_new_n2088_; 
wire core__abc_21302_new_n2090_; 
wire core__abc_21302_new_n2091_; 
wire core__abc_21302_new_n2093_; 
wire core__abc_21302_new_n2094_; 
wire core__abc_21302_new_n2096_; 
wire core__abc_21302_new_n2097_; 
wire core__abc_21302_new_n2099_; 
wire core__abc_21302_new_n2100_; 
wire core__abc_21302_new_n2102_; 
wire core__abc_21302_new_n2103_; 
wire core__abc_21302_new_n2105_; 
wire core__abc_21302_new_n2106_; 
wire core__abc_21302_new_n2108_; 
wire core__abc_21302_new_n2109_; 
wire core__abc_21302_new_n2111_; 
wire core__abc_21302_new_n2112_; 
wire core__abc_21302_new_n2114_; 
wire core__abc_21302_new_n2115_; 
wire core__abc_21302_new_n2117_; 
wire core__abc_21302_new_n2118_; 
wire core__abc_21302_new_n2120_; 
wire core__abc_21302_new_n2121_; 
wire core__abc_21302_new_n2123_; 
wire core__abc_21302_new_n2124_; 
wire core__abc_21302_new_n2126_; 
wire core__abc_21302_new_n2127_; 
wire core__abc_21302_new_n2129_; 
wire core__abc_21302_new_n2130_; 
wire core__abc_21302_new_n2132_; 
wire core__abc_21302_new_n2133_; 
wire core__abc_21302_new_n2135_; 
wire core__abc_21302_new_n2136_; 
wire core__abc_21302_new_n2138_; 
wire core__abc_21302_new_n2139_; 
wire core__abc_21302_new_n2140_; 
wire core__abc_21302_new_n2142_; 
wire core__abc_21302_new_n2143_; 
wire core__abc_21302_new_n2144_; 
wire core__abc_21302_new_n2145_; 
wire core__abc_21302_new_n2146_; 
wire core__abc_21302_new_n2147_; 
wire core__abc_21302_new_n2149_; 
wire core__abc_21302_new_n2150_; 
wire core__abc_21302_new_n2151_; 
wire core__abc_21302_new_n2152_; 
wire core__abc_21302_new_n2154_; 
wire core__abc_21302_new_n2155_; 
wire core__abc_21302_new_n2156_; 
wire core__abc_21302_new_n2157_; 
wire core__abc_21302_new_n2158_; 
wire core__abc_21302_new_n2159_; 
wire core__abc_21302_new_n2161_; 
wire core__abc_21302_new_n2162_; 
wire core__abc_21302_new_n2164_; 
wire core__abc_21302_new_n2165_; 
wire core__abc_21302_new_n2166_; 
wire core__abc_21302_new_n2167_; 
wire core__abc_21302_new_n2168_; 
wire core__abc_21302_new_n2168__bF_buf0; 
wire core__abc_21302_new_n2168__bF_buf1; 
wire core__abc_21302_new_n2168__bF_buf10; 
wire core__abc_21302_new_n2168__bF_buf11; 
wire core__abc_21302_new_n2168__bF_buf12; 
wire core__abc_21302_new_n2168__bF_buf2; 
wire core__abc_21302_new_n2168__bF_buf3; 
wire core__abc_21302_new_n2168__bF_buf4; 
wire core__abc_21302_new_n2168__bF_buf5; 
wire core__abc_21302_new_n2168__bF_buf6; 
wire core__abc_21302_new_n2168__bF_buf7; 
wire core__abc_21302_new_n2168__bF_buf8; 
wire core__abc_21302_new_n2168__bF_buf9; 
wire core__abc_21302_new_n2169_; 
wire core__abc_21302_new_n2171_; 
wire core__abc_21302_new_n2172_; 
wire core__abc_21302_new_n2174_; 
wire core__abc_21302_new_n2175_; 
wire core__abc_21302_new_n2177_; 
wire core__abc_21302_new_n2178_; 
wire core__abc_21302_new_n2180_; 
wire core__abc_21302_new_n2181_; 
wire core__abc_21302_new_n2183_; 
wire core__abc_21302_new_n2184_; 
wire core__abc_21302_new_n2186_; 
wire core__abc_21302_new_n2187_; 
wire core__abc_21302_new_n2189_; 
wire core__abc_21302_new_n2190_; 
wire core__abc_21302_new_n2192_; 
wire core__abc_21302_new_n2193_; 
wire core__abc_21302_new_n2195_; 
wire core__abc_21302_new_n2196_; 
wire core__abc_21302_new_n2198_; 
wire core__abc_21302_new_n2199_; 
wire core__abc_21302_new_n2201_; 
wire core__abc_21302_new_n2202_; 
wire core__abc_21302_new_n2204_; 
wire core__abc_21302_new_n2205_; 
wire core__abc_21302_new_n2207_; 
wire core__abc_21302_new_n2208_; 
wire core__abc_21302_new_n2210_; 
wire core__abc_21302_new_n2211_; 
wire core__abc_21302_new_n2213_; 
wire core__abc_21302_new_n2214_; 
wire core__abc_21302_new_n2216_; 
wire core__abc_21302_new_n2217_; 
wire core__abc_21302_new_n2219_; 
wire core__abc_21302_new_n2220_; 
wire core__abc_21302_new_n2222_; 
wire core__abc_21302_new_n2223_; 
wire core__abc_21302_new_n2225_; 
wire core__abc_21302_new_n2226_; 
wire core__abc_21302_new_n2228_; 
wire core__abc_21302_new_n2229_; 
wire core__abc_21302_new_n2231_; 
wire core__abc_21302_new_n2232_; 
wire core__abc_21302_new_n2234_; 
wire core__abc_21302_new_n2235_; 
wire core__abc_21302_new_n2237_; 
wire core__abc_21302_new_n2238_; 
wire core__abc_21302_new_n2240_; 
wire core__abc_21302_new_n2241_; 
wire core__abc_21302_new_n2243_; 
wire core__abc_21302_new_n2244_; 
wire core__abc_21302_new_n2246_; 
wire core__abc_21302_new_n2247_; 
wire core__abc_21302_new_n2249_; 
wire core__abc_21302_new_n2250_; 
wire core__abc_21302_new_n2252_; 
wire core__abc_21302_new_n2253_; 
wire core__abc_21302_new_n2255_; 
wire core__abc_21302_new_n2256_; 
wire core__abc_21302_new_n2258_; 
wire core__abc_21302_new_n2259_; 
wire core__abc_21302_new_n2261_; 
wire core__abc_21302_new_n2262_; 
wire core__abc_21302_new_n2264_; 
wire core__abc_21302_new_n2265_; 
wire core__abc_21302_new_n2267_; 
wire core__abc_21302_new_n2268_; 
wire core__abc_21302_new_n2270_; 
wire core__abc_21302_new_n2271_; 
wire core__abc_21302_new_n2273_; 
wire core__abc_21302_new_n2274_; 
wire core__abc_21302_new_n2276_; 
wire core__abc_21302_new_n2277_; 
wire core__abc_21302_new_n2279_; 
wire core__abc_21302_new_n2280_; 
wire core__abc_21302_new_n2282_; 
wire core__abc_21302_new_n2283_; 
wire core__abc_21302_new_n2285_; 
wire core__abc_21302_new_n2286_; 
wire core__abc_21302_new_n2288_; 
wire core__abc_21302_new_n2289_; 
wire core__abc_21302_new_n2291_; 
wire core__abc_21302_new_n2292_; 
wire core__abc_21302_new_n2294_; 
wire core__abc_21302_new_n2295_; 
wire core__abc_21302_new_n2297_; 
wire core__abc_21302_new_n2298_; 
wire core__abc_21302_new_n2300_; 
wire core__abc_21302_new_n2301_; 
wire core__abc_21302_new_n2303_; 
wire core__abc_21302_new_n2304_; 
wire core__abc_21302_new_n2306_; 
wire core__abc_21302_new_n2307_; 
wire core__abc_21302_new_n2309_; 
wire core__abc_21302_new_n2310_; 
wire core__abc_21302_new_n2312_; 
wire core__abc_21302_new_n2313_; 
wire core__abc_21302_new_n2315_; 
wire core__abc_21302_new_n2316_; 
wire core__abc_21302_new_n2318_; 
wire core__abc_21302_new_n2319_; 
wire core__abc_21302_new_n2321_; 
wire core__abc_21302_new_n2322_; 
wire core__abc_21302_new_n2324_; 
wire core__abc_21302_new_n2325_; 
wire core__abc_21302_new_n2327_; 
wire core__abc_21302_new_n2328_; 
wire core__abc_21302_new_n2330_; 
wire core__abc_21302_new_n2331_; 
wire core__abc_21302_new_n2333_; 
wire core__abc_21302_new_n2334_; 
wire core__abc_21302_new_n2336_; 
wire core__abc_21302_new_n2337_; 
wire core__abc_21302_new_n2339_; 
wire core__abc_21302_new_n2340_; 
wire core__abc_21302_new_n2342_; 
wire core__abc_21302_new_n2343_; 
wire core__abc_21302_new_n2345_; 
wire core__abc_21302_new_n2346_; 
wire core__abc_21302_new_n2348_; 
wire core__abc_21302_new_n2349_; 
wire core__abc_21302_new_n2351_; 
wire core__abc_21302_new_n2352_; 
wire core__abc_21302_new_n2354_; 
wire core__abc_21302_new_n2355_; 
wire core__abc_21302_new_n2357_; 
wire core__abc_21302_new_n2358_; 
wire core__abc_21302_new_n2360_; 
wire core__abc_21302_new_n2361_; 
wire core__abc_21302_new_n2362_; 
wire core__abc_21302_new_n2362__bF_buf0; 
wire core__abc_21302_new_n2362__bF_buf1; 
wire core__abc_21302_new_n2362__bF_buf10; 
wire core__abc_21302_new_n2362__bF_buf11; 
wire core__abc_21302_new_n2362__bF_buf2; 
wire core__abc_21302_new_n2362__bF_buf3; 
wire core__abc_21302_new_n2362__bF_buf4; 
wire core__abc_21302_new_n2362__bF_buf5; 
wire core__abc_21302_new_n2362__bF_buf6; 
wire core__abc_21302_new_n2362__bF_buf7; 
wire core__abc_21302_new_n2362__bF_buf8; 
wire core__abc_21302_new_n2362__bF_buf9; 
wire core__abc_21302_new_n2363_; 
wire core__abc_21302_new_n2363__bF_buf0; 
wire core__abc_21302_new_n2363__bF_buf1; 
wire core__abc_21302_new_n2363__bF_buf2; 
wire core__abc_21302_new_n2363__bF_buf3; 
wire core__abc_21302_new_n2363__bF_buf4; 
wire core__abc_21302_new_n2363__bF_buf5; 
wire core__abc_21302_new_n2364_; 
wire core__abc_21302_new_n2364__bF_buf0; 
wire core__abc_21302_new_n2364__bF_buf1; 
wire core__abc_21302_new_n2364__bF_buf2; 
wire core__abc_21302_new_n2364__bF_buf3; 
wire core__abc_21302_new_n2364__bF_buf4; 
wire core__abc_21302_new_n2364__bF_buf5; 
wire core__abc_21302_new_n2365_; 
wire core__abc_21302_new_n2365__bF_buf0; 
wire core__abc_21302_new_n2365__bF_buf1; 
wire core__abc_21302_new_n2365__bF_buf2; 
wire core__abc_21302_new_n2365__bF_buf3; 
wire core__abc_21302_new_n2365__bF_buf4; 
wire core__abc_21302_new_n2366_; 
wire core__abc_21302_new_n2367_; 
wire core__abc_21302_new_n2368_; 
wire core__abc_21302_new_n2368__bF_buf0; 
wire core__abc_21302_new_n2368__bF_buf1; 
wire core__abc_21302_new_n2368__bF_buf2; 
wire core__abc_21302_new_n2368__bF_buf3; 
wire core__abc_21302_new_n2368__bF_buf4; 
wire core__abc_21302_new_n2369_; 
wire core__abc_21302_new_n2369__bF_buf0; 
wire core__abc_21302_new_n2369__bF_buf1; 
wire core__abc_21302_new_n2369__bF_buf2; 
wire core__abc_21302_new_n2369__bF_buf3; 
wire core__abc_21302_new_n2369__bF_buf4; 
wire core__abc_21302_new_n2369__bF_buf5; 
wire core__abc_21302_new_n2369__bF_buf6; 
wire core__abc_21302_new_n2369__bF_buf7; 
wire core__abc_21302_new_n2370_; 
wire core__abc_21302_new_n2371_; 
wire core__abc_21302_new_n2372_; 
wire core__abc_21302_new_n2373_; 
wire core__abc_21302_new_n2374_; 
wire core__abc_21302_new_n2375_; 
wire core__abc_21302_new_n2376_; 
wire core__abc_21302_new_n2377_; 
wire core__abc_21302_new_n2378_; 
wire core__abc_21302_new_n2379_; 
wire core__abc_21302_new_n2380_; 
wire core__abc_21302_new_n2381_; 
wire core__abc_21302_new_n2382_; 
wire core__abc_21302_new_n2383_; 
wire core__abc_21302_new_n2384_; 
wire core__abc_21302_new_n2385_; 
wire core__abc_21302_new_n2386_; 
wire core__abc_21302_new_n2387_; 
wire core__abc_21302_new_n2388_; 
wire core__abc_21302_new_n2389_; 
wire core__abc_21302_new_n2390_; 
wire core__abc_21302_new_n2391_; 
wire core__abc_21302_new_n2392_; 
wire core__abc_21302_new_n2393_; 
wire core__abc_21302_new_n2394_; 
wire core__abc_21302_new_n2395_; 
wire core__abc_21302_new_n2396_; 
wire core__abc_21302_new_n2397_; 
wire core__abc_21302_new_n2398_; 
wire core__abc_21302_new_n2399_; 
wire core__abc_21302_new_n2400_; 
wire core__abc_21302_new_n2401_; 
wire core__abc_21302_new_n2402_; 
wire core__abc_21302_new_n2403_; 
wire core__abc_21302_new_n2404_; 
wire core__abc_21302_new_n2405_; 
wire core__abc_21302_new_n2406_; 
wire core__abc_21302_new_n2407_; 
wire core__abc_21302_new_n2408_; 
wire core__abc_21302_new_n2409_; 
wire core__abc_21302_new_n2410_; 
wire core__abc_21302_new_n2411_; 
wire core__abc_21302_new_n2412_; 
wire core__abc_21302_new_n2413_; 
wire core__abc_21302_new_n2414_; 
wire core__abc_21302_new_n2415_; 
wire core__abc_21302_new_n2416_; 
wire core__abc_21302_new_n2417_; 
wire core__abc_21302_new_n2418_; 
wire core__abc_21302_new_n2419_; 
wire core__abc_21302_new_n2420_; 
wire core__abc_21302_new_n2421_; 
wire core__abc_21302_new_n2422_; 
wire core__abc_21302_new_n2423_; 
wire core__abc_21302_new_n2424_; 
wire core__abc_21302_new_n2425_; 
wire core__abc_21302_new_n2426_; 
wire core__abc_21302_new_n2427_; 
wire core__abc_21302_new_n2428_; 
wire core__abc_21302_new_n2429_; 
wire core__abc_21302_new_n2430_; 
wire core__abc_21302_new_n2431_; 
wire core__abc_21302_new_n2432_; 
wire core__abc_21302_new_n2433_; 
wire core__abc_21302_new_n2434_; 
wire core__abc_21302_new_n2435_; 
wire core__abc_21302_new_n2436_; 
wire core__abc_21302_new_n2437_; 
wire core__abc_21302_new_n2438_; 
wire core__abc_21302_new_n2439_; 
wire core__abc_21302_new_n2440_; 
wire core__abc_21302_new_n2441_; 
wire core__abc_21302_new_n2442_; 
wire core__abc_21302_new_n2443_; 
wire core__abc_21302_new_n2444_; 
wire core__abc_21302_new_n2445_; 
wire core__abc_21302_new_n2446_; 
wire core__abc_21302_new_n2447_; 
wire core__abc_21302_new_n2448_; 
wire core__abc_21302_new_n2449_; 
wire core__abc_21302_new_n2450_; 
wire core__abc_21302_new_n2451_; 
wire core__abc_21302_new_n2452_; 
wire core__abc_21302_new_n2453_; 
wire core__abc_21302_new_n2454_; 
wire core__abc_21302_new_n2455_; 
wire core__abc_21302_new_n2456_; 
wire core__abc_21302_new_n2457_; 
wire core__abc_21302_new_n2458_; 
wire core__abc_21302_new_n2459_; 
wire core__abc_21302_new_n2460_; 
wire core__abc_21302_new_n2461_; 
wire core__abc_21302_new_n2462_; 
wire core__abc_21302_new_n2463_; 
wire core__abc_21302_new_n2464_; 
wire core__abc_21302_new_n2465_; 
wire core__abc_21302_new_n2466_; 
wire core__abc_21302_new_n2467_; 
wire core__abc_21302_new_n2468_; 
wire core__abc_21302_new_n2469_; 
wire core__abc_21302_new_n2470_; 
wire core__abc_21302_new_n2471_; 
wire core__abc_21302_new_n2472_; 
wire core__abc_21302_new_n2473_; 
wire core__abc_21302_new_n2474_; 
wire core__abc_21302_new_n2475_; 
wire core__abc_21302_new_n2476_; 
wire core__abc_21302_new_n2477_; 
wire core__abc_21302_new_n2478_; 
wire core__abc_21302_new_n2479_; 
wire core__abc_21302_new_n2480_; 
wire core__abc_21302_new_n2481_; 
wire core__abc_21302_new_n2482_; 
wire core__abc_21302_new_n2483_; 
wire core__abc_21302_new_n2484_; 
wire core__abc_21302_new_n2485_; 
wire core__abc_21302_new_n2486_; 
wire core__abc_21302_new_n2487_; 
wire core__abc_21302_new_n2488_; 
wire core__abc_21302_new_n2489_; 
wire core__abc_21302_new_n2490_; 
wire core__abc_21302_new_n2491_; 
wire core__abc_21302_new_n2492_; 
wire core__abc_21302_new_n2493_; 
wire core__abc_21302_new_n2494_; 
wire core__abc_21302_new_n2495_; 
wire core__abc_21302_new_n2496_; 
wire core__abc_21302_new_n2497_; 
wire core__abc_21302_new_n2498_; 
wire core__abc_21302_new_n2499_; 
wire core__abc_21302_new_n2500_; 
wire core__abc_21302_new_n2501_; 
wire core__abc_21302_new_n2502_; 
wire core__abc_21302_new_n2503_; 
wire core__abc_21302_new_n2504_; 
wire core__abc_21302_new_n2505_; 
wire core__abc_21302_new_n2506_; 
wire core__abc_21302_new_n2507_; 
wire core__abc_21302_new_n2508_; 
wire core__abc_21302_new_n2509_; 
wire core__abc_21302_new_n2510_; 
wire core__abc_21302_new_n2511_; 
wire core__abc_21302_new_n2512_; 
wire core__abc_21302_new_n2513_; 
wire core__abc_21302_new_n2514_; 
wire core__abc_21302_new_n2515_; 
wire core__abc_21302_new_n2516_; 
wire core__abc_21302_new_n2517_; 
wire core__abc_21302_new_n2518_; 
wire core__abc_21302_new_n2519_; 
wire core__abc_21302_new_n2520_; 
wire core__abc_21302_new_n2521_; 
wire core__abc_21302_new_n2522_; 
wire core__abc_21302_new_n2523_; 
wire core__abc_21302_new_n2524_; 
wire core__abc_21302_new_n2525_; 
wire core__abc_21302_new_n2526_; 
wire core__abc_21302_new_n2527_; 
wire core__abc_21302_new_n2528_; 
wire core__abc_21302_new_n2529_; 
wire core__abc_21302_new_n2530_; 
wire core__abc_21302_new_n2531_; 
wire core__abc_21302_new_n2532_; 
wire core__abc_21302_new_n2533_; 
wire core__abc_21302_new_n2534_; 
wire core__abc_21302_new_n2535_; 
wire core__abc_21302_new_n2536_; 
wire core__abc_21302_new_n2537_; 
wire core__abc_21302_new_n2538_; 
wire core__abc_21302_new_n2539_; 
wire core__abc_21302_new_n2540_; 
wire core__abc_21302_new_n2541_; 
wire core__abc_21302_new_n2542_; 
wire core__abc_21302_new_n2543_; 
wire core__abc_21302_new_n2544_; 
wire core__abc_21302_new_n2545_; 
wire core__abc_21302_new_n2546_; 
wire core__abc_21302_new_n2547_; 
wire core__abc_21302_new_n2548_; 
wire core__abc_21302_new_n2549_; 
wire core__abc_21302_new_n2550_; 
wire core__abc_21302_new_n2551_; 
wire core__abc_21302_new_n2552_; 
wire core__abc_21302_new_n2553_; 
wire core__abc_21302_new_n2554_; 
wire core__abc_21302_new_n2555_; 
wire core__abc_21302_new_n2556_; 
wire core__abc_21302_new_n2557_; 
wire core__abc_21302_new_n2558_; 
wire core__abc_21302_new_n2559_; 
wire core__abc_21302_new_n2560_; 
wire core__abc_21302_new_n2561_; 
wire core__abc_21302_new_n2562_; 
wire core__abc_21302_new_n2563_; 
wire core__abc_21302_new_n2564_; 
wire core__abc_21302_new_n2565_; 
wire core__abc_21302_new_n2566_; 
wire core__abc_21302_new_n2567_; 
wire core__abc_21302_new_n2568_; 
wire core__abc_21302_new_n2569_; 
wire core__abc_21302_new_n2570_; 
wire core__abc_21302_new_n2571_; 
wire core__abc_21302_new_n2572_; 
wire core__abc_21302_new_n2573_; 
wire core__abc_21302_new_n2574_; 
wire core__abc_21302_new_n2575_; 
wire core__abc_21302_new_n2576_; 
wire core__abc_21302_new_n2577_; 
wire core__abc_21302_new_n2578_; 
wire core__abc_21302_new_n2579_; 
wire core__abc_21302_new_n2580_; 
wire core__abc_21302_new_n2581_; 
wire core__abc_21302_new_n2582_; 
wire core__abc_21302_new_n2583_; 
wire core__abc_21302_new_n2584_; 
wire core__abc_21302_new_n2585_; 
wire core__abc_21302_new_n2586_; 
wire core__abc_21302_new_n2587_; 
wire core__abc_21302_new_n2588_; 
wire core__abc_21302_new_n2589_; 
wire core__abc_21302_new_n2590_; 
wire core__abc_21302_new_n2591_; 
wire core__abc_21302_new_n2592_; 
wire core__abc_21302_new_n2593_; 
wire core__abc_21302_new_n2594_; 
wire core__abc_21302_new_n2595_; 
wire core__abc_21302_new_n2596_; 
wire core__abc_21302_new_n2597_; 
wire core__abc_21302_new_n2598_; 
wire core__abc_21302_new_n2599_; 
wire core__abc_21302_new_n2600_; 
wire core__abc_21302_new_n2601_; 
wire core__abc_21302_new_n2602_; 
wire core__abc_21302_new_n2603_; 
wire core__abc_21302_new_n2604_; 
wire core__abc_21302_new_n2605_; 
wire core__abc_21302_new_n2606_; 
wire core__abc_21302_new_n2607_; 
wire core__abc_21302_new_n2608_; 
wire core__abc_21302_new_n2609_; 
wire core__abc_21302_new_n2610_; 
wire core__abc_21302_new_n2611_; 
wire core__abc_21302_new_n2612_; 
wire core__abc_21302_new_n2613_; 
wire core__abc_21302_new_n2614_; 
wire core__abc_21302_new_n2615_; 
wire core__abc_21302_new_n2616_; 
wire core__abc_21302_new_n2617_; 
wire core__abc_21302_new_n2618_; 
wire core__abc_21302_new_n2619_; 
wire core__abc_21302_new_n2620_; 
wire core__abc_21302_new_n2621_; 
wire core__abc_21302_new_n2622_; 
wire core__abc_21302_new_n2623_; 
wire core__abc_21302_new_n2624_; 
wire core__abc_21302_new_n2625_; 
wire core__abc_21302_new_n2626_; 
wire core__abc_21302_new_n2627_; 
wire core__abc_21302_new_n2628_; 
wire core__abc_21302_new_n2629_; 
wire core__abc_21302_new_n2630_; 
wire core__abc_21302_new_n2631_; 
wire core__abc_21302_new_n2632_; 
wire core__abc_21302_new_n2633_; 
wire core__abc_21302_new_n2634_; 
wire core__abc_21302_new_n2634__bF_buf0; 
wire core__abc_21302_new_n2634__bF_buf1; 
wire core__abc_21302_new_n2634__bF_buf2; 
wire core__abc_21302_new_n2634__bF_buf3; 
wire core__abc_21302_new_n2634__bF_buf4; 
wire core__abc_21302_new_n2634__bF_buf5; 
wire core__abc_21302_new_n2634__bF_buf6; 
wire core__abc_21302_new_n2634__bF_buf7; 
wire core__abc_21302_new_n2634__bF_buf8; 
wire core__abc_21302_new_n2635_; 
wire core__abc_21302_new_n2636_; 
wire core__abc_21302_new_n2637_; 
wire core__abc_21302_new_n2638_; 
wire core__abc_21302_new_n2639_; 
wire core__abc_21302_new_n2639__bF_buf0; 
wire core__abc_21302_new_n2639__bF_buf1; 
wire core__abc_21302_new_n2639__bF_buf2; 
wire core__abc_21302_new_n2639__bF_buf3; 
wire core__abc_21302_new_n2639__bF_buf4; 
wire core__abc_21302_new_n2639__bF_buf5; 
wire core__abc_21302_new_n2639__bF_buf6; 
wire core__abc_21302_new_n2640_; 
wire core__abc_21302_new_n2640__bF_buf0; 
wire core__abc_21302_new_n2640__bF_buf1; 
wire core__abc_21302_new_n2640__bF_buf10; 
wire core__abc_21302_new_n2640__bF_buf11; 
wire core__abc_21302_new_n2640__bF_buf2; 
wire core__abc_21302_new_n2640__bF_buf3; 
wire core__abc_21302_new_n2640__bF_buf4; 
wire core__abc_21302_new_n2640__bF_buf5; 
wire core__abc_21302_new_n2640__bF_buf6; 
wire core__abc_21302_new_n2640__bF_buf7; 
wire core__abc_21302_new_n2640__bF_buf8; 
wire core__abc_21302_new_n2640__bF_buf9; 
wire core__abc_21302_new_n2641_; 
wire core__abc_21302_new_n2642_; 
wire core__abc_21302_new_n2643_; 
wire core__abc_21302_new_n2644_; 
wire core__abc_21302_new_n2645_; 
wire core__abc_21302_new_n2647_; 
wire core__abc_21302_new_n2648_; 
wire core__abc_21302_new_n2649_; 
wire core__abc_21302_new_n2650_; 
wire core__abc_21302_new_n2651_; 
wire core__abc_21302_new_n2652_; 
wire core__abc_21302_new_n2653_; 
wire core__abc_21302_new_n2654_; 
wire core__abc_21302_new_n2655_; 
wire core__abc_21302_new_n2656_; 
wire core__abc_21302_new_n2657_; 
wire core__abc_21302_new_n2658_; 
wire core__abc_21302_new_n2659_; 
wire core__abc_21302_new_n2660_; 
wire core__abc_21302_new_n2661_; 
wire core__abc_21302_new_n2662_; 
wire core__abc_21302_new_n2663_; 
wire core__abc_21302_new_n2664_; 
wire core__abc_21302_new_n2665_; 
wire core__abc_21302_new_n2666_; 
wire core__abc_21302_new_n2667_; 
wire core__abc_21302_new_n2668_; 
wire core__abc_21302_new_n2669_; 
wire core__abc_21302_new_n2670_; 
wire core__abc_21302_new_n2671_; 
wire core__abc_21302_new_n2672_; 
wire core__abc_21302_new_n2673_; 
wire core__abc_21302_new_n2673__bF_buf0; 
wire core__abc_21302_new_n2673__bF_buf1; 
wire core__abc_21302_new_n2673__bF_buf10; 
wire core__abc_21302_new_n2673__bF_buf11; 
wire core__abc_21302_new_n2673__bF_buf2; 
wire core__abc_21302_new_n2673__bF_buf3; 
wire core__abc_21302_new_n2673__bF_buf4; 
wire core__abc_21302_new_n2673__bF_buf5; 
wire core__abc_21302_new_n2673__bF_buf6; 
wire core__abc_21302_new_n2673__bF_buf7; 
wire core__abc_21302_new_n2673__bF_buf8; 
wire core__abc_21302_new_n2673__bF_buf9; 
wire core__abc_21302_new_n2674_; 
wire core__abc_21302_new_n2675_; 
wire core__abc_21302_new_n2676_; 
wire core__abc_21302_new_n2677_; 
wire core__abc_21302_new_n2678_; 
wire core__abc_21302_new_n2679_; 
wire core__abc_21302_new_n2681_; 
wire core__abc_21302_new_n2682_; 
wire core__abc_21302_new_n2683_; 
wire core__abc_21302_new_n2684_; 
wire core__abc_21302_new_n2685_; 
wire core__abc_21302_new_n2686_; 
wire core__abc_21302_new_n2687_; 
wire core__abc_21302_new_n2688_; 
wire core__abc_21302_new_n2689_; 
wire core__abc_21302_new_n2690_; 
wire core__abc_21302_new_n2691_; 
wire core__abc_21302_new_n2692_; 
wire core__abc_21302_new_n2693_; 
wire core__abc_21302_new_n2694_; 
wire core__abc_21302_new_n2695_; 
wire core__abc_21302_new_n2696_; 
wire core__abc_21302_new_n2697_; 
wire core__abc_21302_new_n2698_; 
wire core__abc_21302_new_n2699_; 
wire core__abc_21302_new_n2700_; 
wire core__abc_21302_new_n2701_; 
wire core__abc_21302_new_n2702_; 
wire core__abc_21302_new_n2703_; 
wire core__abc_21302_new_n2704_; 
wire core__abc_21302_new_n2705_; 
wire core__abc_21302_new_n2706_; 
wire core__abc_21302_new_n2707_; 
wire core__abc_21302_new_n2708_; 
wire core__abc_21302_new_n2709_; 
wire core__abc_21302_new_n2710_; 
wire core__abc_21302_new_n2711_; 
wire core__abc_21302_new_n2712_; 
wire core__abc_21302_new_n2713_; 
wire core__abc_21302_new_n2714_; 
wire core__abc_21302_new_n2715_; 
wire core__abc_21302_new_n2716_; 
wire core__abc_21302_new_n2717_; 
wire core__abc_21302_new_n2719_; 
wire core__abc_21302_new_n2720_; 
wire core__abc_21302_new_n2721_; 
wire core__abc_21302_new_n2722_; 
wire core__abc_21302_new_n2723_; 
wire core__abc_21302_new_n2724_; 
wire core__abc_21302_new_n2725_; 
wire core__abc_21302_new_n2726_; 
wire core__abc_21302_new_n2727_; 
wire core__abc_21302_new_n2728_; 
wire core__abc_21302_new_n2729_; 
wire core__abc_21302_new_n2730_; 
wire core__abc_21302_new_n2731_; 
wire core__abc_21302_new_n2732_; 
wire core__abc_21302_new_n2733_; 
wire core__abc_21302_new_n2734_; 
wire core__abc_21302_new_n2735_; 
wire core__abc_21302_new_n2736_; 
wire core__abc_21302_new_n2737_; 
wire core__abc_21302_new_n2738_; 
wire core__abc_21302_new_n2739_; 
wire core__abc_21302_new_n2740_; 
wire core__abc_21302_new_n2741_; 
wire core__abc_21302_new_n2742_; 
wire core__abc_21302_new_n2743_; 
wire core__abc_21302_new_n2744_; 
wire core__abc_21302_new_n2745_; 
wire core__abc_21302_new_n2746_; 
wire core__abc_21302_new_n2747_; 
wire core__abc_21302_new_n2748_; 
wire core__abc_21302_new_n2749_; 
wire core__abc_21302_new_n2750_; 
wire core__abc_21302_new_n2751_; 
wire core__abc_21302_new_n2752_; 
wire core__abc_21302_new_n2753_; 
wire core__abc_21302_new_n2754_; 
wire core__abc_21302_new_n2755_; 
wire core__abc_21302_new_n2756_; 
wire core__abc_21302_new_n2757_; 
wire core__abc_21302_new_n2758_; 
wire core__abc_21302_new_n2759_; 
wire core__abc_21302_new_n2760_; 
wire core__abc_21302_new_n2762_; 
wire core__abc_21302_new_n2763_; 
wire core__abc_21302_new_n2764_; 
wire core__abc_21302_new_n2765_; 
wire core__abc_21302_new_n2766_; 
wire core__abc_21302_new_n2767_; 
wire core__abc_21302_new_n2768_; 
wire core__abc_21302_new_n2769_; 
wire core__abc_21302_new_n2770_; 
wire core__abc_21302_new_n2771_; 
wire core__abc_21302_new_n2772_; 
wire core__abc_21302_new_n2773_; 
wire core__abc_21302_new_n2774_; 
wire core__abc_21302_new_n2775_; 
wire core__abc_21302_new_n2776_; 
wire core__abc_21302_new_n2777_; 
wire core__abc_21302_new_n2778_; 
wire core__abc_21302_new_n2779_; 
wire core__abc_21302_new_n2780_; 
wire core__abc_21302_new_n2781_; 
wire core__abc_21302_new_n2782_; 
wire core__abc_21302_new_n2783_; 
wire core__abc_21302_new_n2784_; 
wire core__abc_21302_new_n2785_; 
wire core__abc_21302_new_n2786_; 
wire core__abc_21302_new_n2787_; 
wire core__abc_21302_new_n2788_; 
wire core__abc_21302_new_n2789_; 
wire core__abc_21302_new_n2790_; 
wire core__abc_21302_new_n2791_; 
wire core__abc_21302_new_n2792_; 
wire core__abc_21302_new_n2793_; 
wire core__abc_21302_new_n2794_; 
wire core__abc_21302_new_n2795_; 
wire core__abc_21302_new_n2796_; 
wire core__abc_21302_new_n2798_; 
wire core__abc_21302_new_n2799_; 
wire core__abc_21302_new_n2800_; 
wire core__abc_21302_new_n2801_; 
wire core__abc_21302_new_n2802_; 
wire core__abc_21302_new_n2803_; 
wire core__abc_21302_new_n2804_; 
wire core__abc_21302_new_n2805_; 
wire core__abc_21302_new_n2806_; 
wire core__abc_21302_new_n2807_; 
wire core__abc_21302_new_n2808_; 
wire core__abc_21302_new_n2809_; 
wire core__abc_21302_new_n2810_; 
wire core__abc_21302_new_n2811_; 
wire core__abc_21302_new_n2812_; 
wire core__abc_21302_new_n2813_; 
wire core__abc_21302_new_n2814_; 
wire core__abc_21302_new_n2815_; 
wire core__abc_21302_new_n2816_; 
wire core__abc_21302_new_n2817_; 
wire core__abc_21302_new_n2818_; 
wire core__abc_21302_new_n2819_; 
wire core__abc_21302_new_n2820_; 
wire core__abc_21302_new_n2821_; 
wire core__abc_21302_new_n2822_; 
wire core__abc_21302_new_n2823_; 
wire core__abc_21302_new_n2824_; 
wire core__abc_21302_new_n2825_; 
wire core__abc_21302_new_n2826_; 
wire core__abc_21302_new_n2827_; 
wire core__abc_21302_new_n2828_; 
wire core__abc_21302_new_n2829_; 
wire core__abc_21302_new_n2830_; 
wire core__abc_21302_new_n2831_; 
wire core__abc_21302_new_n2832_; 
wire core__abc_21302_new_n2833_; 
wire core__abc_21302_new_n2834_; 
wire core__abc_21302_new_n2835_; 
wire core__abc_21302_new_n2836_; 
wire core__abc_21302_new_n2837_; 
wire core__abc_21302_new_n2839_; 
wire core__abc_21302_new_n2840_; 
wire core__abc_21302_new_n2841_; 
wire core__abc_21302_new_n2842_; 
wire core__abc_21302_new_n2843_; 
wire core__abc_21302_new_n2844_; 
wire core__abc_21302_new_n2845_; 
wire core__abc_21302_new_n2846_; 
wire core__abc_21302_new_n2847_; 
wire core__abc_21302_new_n2848_; 
wire core__abc_21302_new_n2849_; 
wire core__abc_21302_new_n2850_; 
wire core__abc_21302_new_n2851_; 
wire core__abc_21302_new_n2852_; 
wire core__abc_21302_new_n2853_; 
wire core__abc_21302_new_n2854_; 
wire core__abc_21302_new_n2855_; 
wire core__abc_21302_new_n2856_; 
wire core__abc_21302_new_n2857_; 
wire core__abc_21302_new_n2858_; 
wire core__abc_21302_new_n2859_; 
wire core__abc_21302_new_n2860_; 
wire core__abc_21302_new_n2861_; 
wire core__abc_21302_new_n2862_; 
wire core__abc_21302_new_n2863_; 
wire core__abc_21302_new_n2864_; 
wire core__abc_21302_new_n2865_; 
wire core__abc_21302_new_n2866_; 
wire core__abc_21302_new_n2867_; 
wire core__abc_21302_new_n2868_; 
wire core__abc_21302_new_n2869_; 
wire core__abc_21302_new_n2870_; 
wire core__abc_21302_new_n2871_; 
wire core__abc_21302_new_n2872_; 
wire core__abc_21302_new_n2873_; 
wire core__abc_21302_new_n2874_; 
wire core__abc_21302_new_n2875_; 
wire core__abc_21302_new_n2876_; 
wire core__abc_21302_new_n2877_; 
wire core__abc_21302_new_n2879_; 
wire core__abc_21302_new_n2880_; 
wire core__abc_21302_new_n2881_; 
wire core__abc_21302_new_n2882_; 
wire core__abc_21302_new_n2883_; 
wire core__abc_21302_new_n2884_; 
wire core__abc_21302_new_n2885_; 
wire core__abc_21302_new_n2886_; 
wire core__abc_21302_new_n2887_; 
wire core__abc_21302_new_n2888_; 
wire core__abc_21302_new_n2889_; 
wire core__abc_21302_new_n2890_; 
wire core__abc_21302_new_n2891_; 
wire core__abc_21302_new_n2892_; 
wire core__abc_21302_new_n2893_; 
wire core__abc_21302_new_n2894_; 
wire core__abc_21302_new_n2895_; 
wire core__abc_21302_new_n2896_; 
wire core__abc_21302_new_n2897_; 
wire core__abc_21302_new_n2898_; 
wire core__abc_21302_new_n2899_; 
wire core__abc_21302_new_n2900_; 
wire core__abc_21302_new_n2901_; 
wire core__abc_21302_new_n2902_; 
wire core__abc_21302_new_n2903_; 
wire core__abc_21302_new_n2904_; 
wire core__abc_21302_new_n2905_; 
wire core__abc_21302_new_n2906_; 
wire core__abc_21302_new_n2907_; 
wire core__abc_21302_new_n2908_; 
wire core__abc_21302_new_n2909_; 
wire core__abc_21302_new_n2910_; 
wire core__abc_21302_new_n2911_; 
wire core__abc_21302_new_n2912_; 
wire core__abc_21302_new_n2913_; 
wire core__abc_21302_new_n2915_; 
wire core__abc_21302_new_n2916_; 
wire core__abc_21302_new_n2917_; 
wire core__abc_21302_new_n2918_; 
wire core__abc_21302_new_n2919_; 
wire core__abc_21302_new_n2920_; 
wire core__abc_21302_new_n2921_; 
wire core__abc_21302_new_n2922_; 
wire core__abc_21302_new_n2923_; 
wire core__abc_21302_new_n2924_; 
wire core__abc_21302_new_n2925_; 
wire core__abc_21302_new_n2926_; 
wire core__abc_21302_new_n2927_; 
wire core__abc_21302_new_n2928_; 
wire core__abc_21302_new_n2929_; 
wire core__abc_21302_new_n2930_; 
wire core__abc_21302_new_n2931_; 
wire core__abc_21302_new_n2932_; 
wire core__abc_21302_new_n2933_; 
wire core__abc_21302_new_n2934_; 
wire core__abc_21302_new_n2935_; 
wire core__abc_21302_new_n2936_; 
wire core__abc_21302_new_n2937_; 
wire core__abc_21302_new_n2938_; 
wire core__abc_21302_new_n2939_; 
wire core__abc_21302_new_n2940_; 
wire core__abc_21302_new_n2941_; 
wire core__abc_21302_new_n2942_; 
wire core__abc_21302_new_n2943_; 
wire core__abc_21302_new_n2944_; 
wire core__abc_21302_new_n2945_; 
wire core__abc_21302_new_n2946_; 
wire core__abc_21302_new_n2947_; 
wire core__abc_21302_new_n2948_; 
wire core__abc_21302_new_n2949_; 
wire core__abc_21302_new_n2950_; 
wire core__abc_21302_new_n2951_; 
wire core__abc_21302_new_n2952_; 
wire core__abc_21302_new_n2953_; 
wire core__abc_21302_new_n2954_; 
wire core__abc_21302_new_n2955_; 
wire core__abc_21302_new_n2956_; 
wire core__abc_21302_new_n2957_; 
wire core__abc_21302_new_n2958_; 
wire core__abc_21302_new_n2959_; 
wire core__abc_21302_new_n2960_; 
wire core__abc_21302_new_n2961_; 
wire core__abc_21302_new_n2962_; 
wire core__abc_21302_new_n2964_; 
wire core__abc_21302_new_n2965_; 
wire core__abc_21302_new_n2966_; 
wire core__abc_21302_new_n2967_; 
wire core__abc_21302_new_n2968_; 
wire core__abc_21302_new_n2969_; 
wire core__abc_21302_new_n2970_; 
wire core__abc_21302_new_n2971_; 
wire core__abc_21302_new_n2972_; 
wire core__abc_21302_new_n2973_; 
wire core__abc_21302_new_n2974_; 
wire core__abc_21302_new_n2975_; 
wire core__abc_21302_new_n2976_; 
wire core__abc_21302_new_n2977_; 
wire core__abc_21302_new_n2978_; 
wire core__abc_21302_new_n2979_; 
wire core__abc_21302_new_n2980_; 
wire core__abc_21302_new_n2981_; 
wire core__abc_21302_new_n2982_; 
wire core__abc_21302_new_n2983_; 
wire core__abc_21302_new_n2984_; 
wire core__abc_21302_new_n2985_; 
wire core__abc_21302_new_n2986_; 
wire core__abc_21302_new_n2987_; 
wire core__abc_21302_new_n2988_; 
wire core__abc_21302_new_n2989_; 
wire core__abc_21302_new_n2990_; 
wire core__abc_21302_new_n2991_; 
wire core__abc_21302_new_n2992_; 
wire core__abc_21302_new_n2993_; 
wire core__abc_21302_new_n2994_; 
wire core__abc_21302_new_n2995_; 
wire core__abc_21302_new_n2996_; 
wire core__abc_21302_new_n2997_; 
wire core__abc_21302_new_n2998_; 
wire core__abc_21302_new_n3000_; 
wire core__abc_21302_new_n3001_; 
wire core__abc_21302_new_n3002_; 
wire core__abc_21302_new_n3003_; 
wire core__abc_21302_new_n3004_; 
wire core__abc_21302_new_n3005_; 
wire core__abc_21302_new_n3006_; 
wire core__abc_21302_new_n3007_; 
wire core__abc_21302_new_n3008_; 
wire core__abc_21302_new_n3009_; 
wire core__abc_21302_new_n3010_; 
wire core__abc_21302_new_n3011_; 
wire core__abc_21302_new_n3012_; 
wire core__abc_21302_new_n3013_; 
wire core__abc_21302_new_n3014_; 
wire core__abc_21302_new_n3015_; 
wire core__abc_21302_new_n3016_; 
wire core__abc_21302_new_n3017_; 
wire core__abc_21302_new_n3018_; 
wire core__abc_21302_new_n3019_; 
wire core__abc_21302_new_n3020_; 
wire core__abc_21302_new_n3021_; 
wire core__abc_21302_new_n3022_; 
wire core__abc_21302_new_n3023_; 
wire core__abc_21302_new_n3024_; 
wire core__abc_21302_new_n3025_; 
wire core__abc_21302_new_n3026_; 
wire core__abc_21302_new_n3027_; 
wire core__abc_21302_new_n3028_; 
wire core__abc_21302_new_n3029_; 
wire core__abc_21302_new_n3030_; 
wire core__abc_21302_new_n3031_; 
wire core__abc_21302_new_n3032_; 
wire core__abc_21302_new_n3033_; 
wire core__abc_21302_new_n3034_; 
wire core__abc_21302_new_n3035_; 
wire core__abc_21302_new_n3036_; 
wire core__abc_21302_new_n3037_; 
wire core__abc_21302_new_n3038_; 
wire core__abc_21302_new_n3039_; 
wire core__abc_21302_new_n3040_; 
wire core__abc_21302_new_n3042_; 
wire core__abc_21302_new_n3043_; 
wire core__abc_21302_new_n3044_; 
wire core__abc_21302_new_n3045_; 
wire core__abc_21302_new_n3046_; 
wire core__abc_21302_new_n3047_; 
wire core__abc_21302_new_n3048_; 
wire core__abc_21302_new_n3049_; 
wire core__abc_21302_new_n3050_; 
wire core__abc_21302_new_n3051_; 
wire core__abc_21302_new_n3052_; 
wire core__abc_21302_new_n3053_; 
wire core__abc_21302_new_n3054_; 
wire core__abc_21302_new_n3055_; 
wire core__abc_21302_new_n3056_; 
wire core__abc_21302_new_n3057_; 
wire core__abc_21302_new_n3058_; 
wire core__abc_21302_new_n3059_; 
wire core__abc_21302_new_n3060_; 
wire core__abc_21302_new_n3061_; 
wire core__abc_21302_new_n3062_; 
wire core__abc_21302_new_n3063_; 
wire core__abc_21302_new_n3064_; 
wire core__abc_21302_new_n3065_; 
wire core__abc_21302_new_n3066_; 
wire core__abc_21302_new_n3067_; 
wire core__abc_21302_new_n3068_; 
wire core__abc_21302_new_n3069_; 
wire core__abc_21302_new_n3070_; 
wire core__abc_21302_new_n3071_; 
wire core__abc_21302_new_n3072_; 
wire core__abc_21302_new_n3073_; 
wire core__abc_21302_new_n3074_; 
wire core__abc_21302_new_n3075_; 
wire core__abc_21302_new_n3076_; 
wire core__abc_21302_new_n3077_; 
wire core__abc_21302_new_n3078_; 
wire core__abc_21302_new_n3079_; 
wire core__abc_21302_new_n3080_; 
wire core__abc_21302_new_n3082_; 
wire core__abc_21302_new_n3083_; 
wire core__abc_21302_new_n3084_; 
wire core__abc_21302_new_n3085_; 
wire core__abc_21302_new_n3086_; 
wire core__abc_21302_new_n3087_; 
wire core__abc_21302_new_n3088_; 
wire core__abc_21302_new_n3089_; 
wire core__abc_21302_new_n3090_; 
wire core__abc_21302_new_n3091_; 
wire core__abc_21302_new_n3092_; 
wire core__abc_21302_new_n3093_; 
wire core__abc_21302_new_n3094_; 
wire core__abc_21302_new_n3095_; 
wire core__abc_21302_new_n3096_; 
wire core__abc_21302_new_n3097_; 
wire core__abc_21302_new_n3098_; 
wire core__abc_21302_new_n3099_; 
wire core__abc_21302_new_n3100_; 
wire core__abc_21302_new_n3101_; 
wire core__abc_21302_new_n3102_; 
wire core__abc_21302_new_n3103_; 
wire core__abc_21302_new_n3104_; 
wire core__abc_21302_new_n3105_; 
wire core__abc_21302_new_n3106_; 
wire core__abc_21302_new_n3107_; 
wire core__abc_21302_new_n3108_; 
wire core__abc_21302_new_n3109_; 
wire core__abc_21302_new_n3110_; 
wire core__abc_21302_new_n3111_; 
wire core__abc_21302_new_n3112_; 
wire core__abc_21302_new_n3113_; 
wire core__abc_21302_new_n3114_; 
wire core__abc_21302_new_n3115_; 
wire core__abc_21302_new_n3116_; 
wire core__abc_21302_new_n3117_; 
wire core__abc_21302_new_n3118_; 
wire core__abc_21302_new_n3119_; 
wire core__abc_21302_new_n3120_; 
wire core__abc_21302_new_n3121_; 
wire core__abc_21302_new_n3122_; 
wire core__abc_21302_new_n3123_; 
wire core__abc_21302_new_n3124_; 
wire core__abc_21302_new_n3125_; 
wire core__abc_21302_new_n3126_; 
wire core__abc_21302_new_n3127_; 
wire core__abc_21302_new_n3129_; 
wire core__abc_21302_new_n3130_; 
wire core__abc_21302_new_n3131_; 
wire core__abc_21302_new_n3132_; 
wire core__abc_21302_new_n3133_; 
wire core__abc_21302_new_n3134_; 
wire core__abc_21302_new_n3135_; 
wire core__abc_21302_new_n3136_; 
wire core__abc_21302_new_n3137_; 
wire core__abc_21302_new_n3138_; 
wire core__abc_21302_new_n3139_; 
wire core__abc_21302_new_n3140_; 
wire core__abc_21302_new_n3141_; 
wire core__abc_21302_new_n3142_; 
wire core__abc_21302_new_n3143_; 
wire core__abc_21302_new_n3144_; 
wire core__abc_21302_new_n3145_; 
wire core__abc_21302_new_n3146_; 
wire core__abc_21302_new_n3147_; 
wire core__abc_21302_new_n3148_; 
wire core__abc_21302_new_n3149_; 
wire core__abc_21302_new_n3150_; 
wire core__abc_21302_new_n3151_; 
wire core__abc_21302_new_n3152_; 
wire core__abc_21302_new_n3153_; 
wire core__abc_21302_new_n3154_; 
wire core__abc_21302_new_n3155_; 
wire core__abc_21302_new_n3156_; 
wire core__abc_21302_new_n3157_; 
wire core__abc_21302_new_n3158_; 
wire core__abc_21302_new_n3159_; 
wire core__abc_21302_new_n3160_; 
wire core__abc_21302_new_n3161_; 
wire core__abc_21302_new_n3162_; 
wire core__abc_21302_new_n3163_; 
wire core__abc_21302_new_n3164_; 
wire core__abc_21302_new_n3165_; 
wire core__abc_21302_new_n3166_; 
wire core__abc_21302_new_n3167_; 
wire core__abc_21302_new_n3168_; 
wire core__abc_21302_new_n3169_; 
wire core__abc_21302_new_n3170_; 
wire core__abc_21302_new_n3171_; 
wire core__abc_21302_new_n3172_; 
wire core__abc_21302_new_n3173_; 
wire core__abc_21302_new_n3175_; 
wire core__abc_21302_new_n3176_; 
wire core__abc_21302_new_n3177_; 
wire core__abc_21302_new_n3178_; 
wire core__abc_21302_new_n3179_; 
wire core__abc_21302_new_n3180_; 
wire core__abc_21302_new_n3181_; 
wire core__abc_21302_new_n3182_; 
wire core__abc_21302_new_n3183_; 
wire core__abc_21302_new_n3184_; 
wire core__abc_21302_new_n3185_; 
wire core__abc_21302_new_n3186_; 
wire core__abc_21302_new_n3187_; 
wire core__abc_21302_new_n3188_; 
wire core__abc_21302_new_n3189_; 
wire core__abc_21302_new_n3190_; 
wire core__abc_21302_new_n3191_; 
wire core__abc_21302_new_n3192_; 
wire core__abc_21302_new_n3193_; 
wire core__abc_21302_new_n3194_; 
wire core__abc_21302_new_n3195_; 
wire core__abc_21302_new_n3196_; 
wire core__abc_21302_new_n3197_; 
wire core__abc_21302_new_n3198_; 
wire core__abc_21302_new_n3199_; 
wire core__abc_21302_new_n3200_; 
wire core__abc_21302_new_n3201_; 
wire core__abc_21302_new_n3202_; 
wire core__abc_21302_new_n3203_; 
wire core__abc_21302_new_n3204_; 
wire core__abc_21302_new_n3205_; 
wire core__abc_21302_new_n3206_; 
wire core__abc_21302_new_n3207_; 
wire core__abc_21302_new_n3208_; 
wire core__abc_21302_new_n3209_; 
wire core__abc_21302_new_n3210_; 
wire core__abc_21302_new_n3211_; 
wire core__abc_21302_new_n3212_; 
wire core__abc_21302_new_n3213_; 
wire core__abc_21302_new_n3214_; 
wire core__abc_21302_new_n3215_; 
wire core__abc_21302_new_n3216_; 
wire core__abc_21302_new_n3217_; 
wire core__abc_21302_new_n3218_; 
wire core__abc_21302_new_n3219_; 
wire core__abc_21302_new_n3220_; 
wire core__abc_21302_new_n3221_; 
wire core__abc_21302_new_n3223_; 
wire core__abc_21302_new_n3224_; 
wire core__abc_21302_new_n3225_; 
wire core__abc_21302_new_n3226_; 
wire core__abc_21302_new_n3227_; 
wire core__abc_21302_new_n3228_; 
wire core__abc_21302_new_n3229_; 
wire core__abc_21302_new_n3230_; 
wire core__abc_21302_new_n3231_; 
wire core__abc_21302_new_n3232_; 
wire core__abc_21302_new_n3233_; 
wire core__abc_21302_new_n3234_; 
wire core__abc_21302_new_n3235_; 
wire core__abc_21302_new_n3236_; 
wire core__abc_21302_new_n3237_; 
wire core__abc_21302_new_n3238_; 
wire core__abc_21302_new_n3239_; 
wire core__abc_21302_new_n3240_; 
wire core__abc_21302_new_n3241_; 
wire core__abc_21302_new_n3242_; 
wire core__abc_21302_new_n3243_; 
wire core__abc_21302_new_n3244_; 
wire core__abc_21302_new_n3245_; 
wire core__abc_21302_new_n3246_; 
wire core__abc_21302_new_n3247_; 
wire core__abc_21302_new_n3248_; 
wire core__abc_21302_new_n3249_; 
wire core__abc_21302_new_n3250_; 
wire core__abc_21302_new_n3251_; 
wire core__abc_21302_new_n3252_; 
wire core__abc_21302_new_n3253_; 
wire core__abc_21302_new_n3254_; 
wire core__abc_21302_new_n3255_; 
wire core__abc_21302_new_n3256_; 
wire core__abc_21302_new_n3257_; 
wire core__abc_21302_new_n3258_; 
wire core__abc_21302_new_n3259_; 
wire core__abc_21302_new_n3260_; 
wire core__abc_21302_new_n3261_; 
wire core__abc_21302_new_n3262_; 
wire core__abc_21302_new_n3263_; 
wire core__abc_21302_new_n3265_; 
wire core__abc_21302_new_n3266_; 
wire core__abc_21302_new_n3267_; 
wire core__abc_21302_new_n3268_; 
wire core__abc_21302_new_n3269_; 
wire core__abc_21302_new_n3270_; 
wire core__abc_21302_new_n3271_; 
wire core__abc_21302_new_n3272_; 
wire core__abc_21302_new_n3273_; 
wire core__abc_21302_new_n3274_; 
wire core__abc_21302_new_n3275_; 
wire core__abc_21302_new_n3276_; 
wire core__abc_21302_new_n3277_; 
wire core__abc_21302_new_n3278_; 
wire core__abc_21302_new_n3279_; 
wire core__abc_21302_new_n3280_; 
wire core__abc_21302_new_n3281_; 
wire core__abc_21302_new_n3282_; 
wire core__abc_21302_new_n3283_; 
wire core__abc_21302_new_n3284_; 
wire core__abc_21302_new_n3285_; 
wire core__abc_21302_new_n3286_; 
wire core__abc_21302_new_n3287_; 
wire core__abc_21302_new_n3288_; 
wire core__abc_21302_new_n3289_; 
wire core__abc_21302_new_n3290_; 
wire core__abc_21302_new_n3291_; 
wire core__abc_21302_new_n3292_; 
wire core__abc_21302_new_n3293_; 
wire core__abc_21302_new_n3294_; 
wire core__abc_21302_new_n3295_; 
wire core__abc_21302_new_n3296_; 
wire core__abc_21302_new_n3297_; 
wire core__abc_21302_new_n3298_; 
wire core__abc_21302_new_n3299_; 
wire core__abc_21302_new_n3300_; 
wire core__abc_21302_new_n3301_; 
wire core__abc_21302_new_n3302_; 
wire core__abc_21302_new_n3303_; 
wire core__abc_21302_new_n3304_; 
wire core__abc_21302_new_n3305_; 
wire core__abc_21302_new_n3306_; 
wire core__abc_21302_new_n3307_; 
wire core__abc_21302_new_n3308_; 
wire core__abc_21302_new_n3309_; 
wire core__abc_21302_new_n3310_; 
wire core__abc_21302_new_n3311_; 
wire core__abc_21302_new_n3312_; 
wire core__abc_21302_new_n3313_; 
wire core__abc_21302_new_n3314_; 
wire core__abc_21302_new_n3315_; 
wire core__abc_21302_new_n3316_; 
wire core__abc_21302_new_n3317_; 
wire core__abc_21302_new_n3318_; 
wire core__abc_21302_new_n3319_; 
wire core__abc_21302_new_n3320_; 
wire core__abc_21302_new_n3321_; 
wire core__abc_21302_new_n3322_; 
wire core__abc_21302_new_n3323_; 
wire core__abc_21302_new_n3324_; 
wire core__abc_21302_new_n3325_; 
wire core__abc_21302_new_n3326_; 
wire core__abc_21302_new_n3328_; 
wire core__abc_21302_new_n3329_; 
wire core__abc_21302_new_n3330_; 
wire core__abc_21302_new_n3331_; 
wire core__abc_21302_new_n3332_; 
wire core__abc_21302_new_n3333_; 
wire core__abc_21302_new_n3334_; 
wire core__abc_21302_new_n3335_; 
wire core__abc_21302_new_n3336_; 
wire core__abc_21302_new_n3337_; 
wire core__abc_21302_new_n3338_; 
wire core__abc_21302_new_n3339_; 
wire core__abc_21302_new_n3340_; 
wire core__abc_21302_new_n3341_; 
wire core__abc_21302_new_n3342_; 
wire core__abc_21302_new_n3343_; 
wire core__abc_21302_new_n3344_; 
wire core__abc_21302_new_n3345_; 
wire core__abc_21302_new_n3346_; 
wire core__abc_21302_new_n3347_; 
wire core__abc_21302_new_n3348_; 
wire core__abc_21302_new_n3349_; 
wire core__abc_21302_new_n3350_; 
wire core__abc_21302_new_n3351_; 
wire core__abc_21302_new_n3352_; 
wire core__abc_21302_new_n3353_; 
wire core__abc_21302_new_n3354_; 
wire core__abc_21302_new_n3355_; 
wire core__abc_21302_new_n3356_; 
wire core__abc_21302_new_n3357_; 
wire core__abc_21302_new_n3358_; 
wire core__abc_21302_new_n3359_; 
wire core__abc_21302_new_n3360_; 
wire core__abc_21302_new_n3361_; 
wire core__abc_21302_new_n3362_; 
wire core__abc_21302_new_n3363_; 
wire core__abc_21302_new_n3364_; 
wire core__abc_21302_new_n3365_; 
wire core__abc_21302_new_n3366_; 
wire core__abc_21302_new_n3368_; 
wire core__abc_21302_new_n3369_; 
wire core__abc_21302_new_n3370_; 
wire core__abc_21302_new_n3371_; 
wire core__abc_21302_new_n3372_; 
wire core__abc_21302_new_n3373_; 
wire core__abc_21302_new_n3374_; 
wire core__abc_21302_new_n3375_; 
wire core__abc_21302_new_n3376_; 
wire core__abc_21302_new_n3377_; 
wire core__abc_21302_new_n3378_; 
wire core__abc_21302_new_n3379_; 
wire core__abc_21302_new_n3380_; 
wire core__abc_21302_new_n3381_; 
wire core__abc_21302_new_n3382_; 
wire core__abc_21302_new_n3383_; 
wire core__abc_21302_new_n3384_; 
wire core__abc_21302_new_n3385_; 
wire core__abc_21302_new_n3386_; 
wire core__abc_21302_new_n3387_; 
wire core__abc_21302_new_n3388_; 
wire core__abc_21302_new_n3389_; 
wire core__abc_21302_new_n3390_; 
wire core__abc_21302_new_n3391_; 
wire core__abc_21302_new_n3392_; 
wire core__abc_21302_new_n3393_; 
wire core__abc_21302_new_n3394_; 
wire core__abc_21302_new_n3395_; 
wire core__abc_21302_new_n3396_; 
wire core__abc_21302_new_n3397_; 
wire core__abc_21302_new_n3398_; 
wire core__abc_21302_new_n3399_; 
wire core__abc_21302_new_n3400_; 
wire core__abc_21302_new_n3401_; 
wire core__abc_21302_new_n3402_; 
wire core__abc_21302_new_n3403_; 
wire core__abc_21302_new_n3404_; 
wire core__abc_21302_new_n3405_; 
wire core__abc_21302_new_n3406_; 
wire core__abc_21302_new_n3407_; 
wire core__abc_21302_new_n3408_; 
wire core__abc_21302_new_n3409_; 
wire core__abc_21302_new_n3410_; 
wire core__abc_21302_new_n3411_; 
wire core__abc_21302_new_n3412_; 
wire core__abc_21302_new_n3413_; 
wire core__abc_21302_new_n3415_; 
wire core__abc_21302_new_n3416_; 
wire core__abc_21302_new_n3417_; 
wire core__abc_21302_new_n3418_; 
wire core__abc_21302_new_n3419_; 
wire core__abc_21302_new_n3420_; 
wire core__abc_21302_new_n3421_; 
wire core__abc_21302_new_n3422_; 
wire core__abc_21302_new_n3423_; 
wire core__abc_21302_new_n3424_; 
wire core__abc_21302_new_n3425_; 
wire core__abc_21302_new_n3426_; 
wire core__abc_21302_new_n3427_; 
wire core__abc_21302_new_n3428_; 
wire core__abc_21302_new_n3429_; 
wire core__abc_21302_new_n3430_; 
wire core__abc_21302_new_n3431_; 
wire core__abc_21302_new_n3432_; 
wire core__abc_21302_new_n3433_; 
wire core__abc_21302_new_n3434_; 
wire core__abc_21302_new_n3435_; 
wire core__abc_21302_new_n3436_; 
wire core__abc_21302_new_n3437_; 
wire core__abc_21302_new_n3438_; 
wire core__abc_21302_new_n3439_; 
wire core__abc_21302_new_n3440_; 
wire core__abc_21302_new_n3441_; 
wire core__abc_21302_new_n3442_; 
wire core__abc_21302_new_n3443_; 
wire core__abc_21302_new_n3444_; 
wire core__abc_21302_new_n3445_; 
wire core__abc_21302_new_n3446_; 
wire core__abc_21302_new_n3447_; 
wire core__abc_21302_new_n3448_; 
wire core__abc_21302_new_n3449_; 
wire core__abc_21302_new_n3450_; 
wire core__abc_21302_new_n3451_; 
wire core__abc_21302_new_n3452_; 
wire core__abc_21302_new_n3453_; 
wire core__abc_21302_new_n3454_; 
wire core__abc_21302_new_n3455_; 
wire core__abc_21302_new_n3456_; 
wire core__abc_21302_new_n3458_; 
wire core__abc_21302_new_n3459_; 
wire core__abc_21302_new_n3460_; 
wire core__abc_21302_new_n3461_; 
wire core__abc_21302_new_n3462_; 
wire core__abc_21302_new_n3463_; 
wire core__abc_21302_new_n3464_; 
wire core__abc_21302_new_n3465_; 
wire core__abc_21302_new_n3466_; 
wire core__abc_21302_new_n3467_; 
wire core__abc_21302_new_n3468_; 
wire core__abc_21302_new_n3469_; 
wire core__abc_21302_new_n3470_; 
wire core__abc_21302_new_n3471_; 
wire core__abc_21302_new_n3472_; 
wire core__abc_21302_new_n3473_; 
wire core__abc_21302_new_n3474_; 
wire core__abc_21302_new_n3475_; 
wire core__abc_21302_new_n3476_; 
wire core__abc_21302_new_n3477_; 
wire core__abc_21302_new_n3478_; 
wire core__abc_21302_new_n3479_; 
wire core__abc_21302_new_n3480_; 
wire core__abc_21302_new_n3481_; 
wire core__abc_21302_new_n3482_; 
wire core__abc_21302_new_n3483_; 
wire core__abc_21302_new_n3484_; 
wire core__abc_21302_new_n3485_; 
wire core__abc_21302_new_n3486_; 
wire core__abc_21302_new_n3487_; 
wire core__abc_21302_new_n3488_; 
wire core__abc_21302_new_n3489_; 
wire core__abc_21302_new_n3490_; 
wire core__abc_21302_new_n3491_; 
wire core__abc_21302_new_n3492_; 
wire core__abc_21302_new_n3493_; 
wire core__abc_21302_new_n3494_; 
wire core__abc_21302_new_n3495_; 
wire core__abc_21302_new_n3496_; 
wire core__abc_21302_new_n3497_; 
wire core__abc_21302_new_n3499_; 
wire core__abc_21302_new_n3500_; 
wire core__abc_21302_new_n3501_; 
wire core__abc_21302_new_n3502_; 
wire core__abc_21302_new_n3503_; 
wire core__abc_21302_new_n3504_; 
wire core__abc_21302_new_n3505_; 
wire core__abc_21302_new_n3506_; 
wire core__abc_21302_new_n3507_; 
wire core__abc_21302_new_n3508_; 
wire core__abc_21302_new_n3509_; 
wire core__abc_21302_new_n3510_; 
wire core__abc_21302_new_n3511_; 
wire core__abc_21302_new_n3512_; 
wire core__abc_21302_new_n3513_; 
wire core__abc_21302_new_n3514_; 
wire core__abc_21302_new_n3515_; 
wire core__abc_21302_new_n3516_; 
wire core__abc_21302_new_n3517_; 
wire core__abc_21302_new_n3518_; 
wire core__abc_21302_new_n3519_; 
wire core__abc_21302_new_n3520_; 
wire core__abc_21302_new_n3521_; 
wire core__abc_21302_new_n3522_; 
wire core__abc_21302_new_n3523_; 
wire core__abc_21302_new_n3524_; 
wire core__abc_21302_new_n3525_; 
wire core__abc_21302_new_n3526_; 
wire core__abc_21302_new_n3527_; 
wire core__abc_21302_new_n3528_; 
wire core__abc_21302_new_n3529_; 
wire core__abc_21302_new_n3531_; 
wire core__abc_21302_new_n3532_; 
wire core__abc_21302_new_n3533_; 
wire core__abc_21302_new_n3534_; 
wire core__abc_21302_new_n3535_; 
wire core__abc_21302_new_n3536_; 
wire core__abc_21302_new_n3537_; 
wire core__abc_21302_new_n3538_; 
wire core__abc_21302_new_n3539_; 
wire core__abc_21302_new_n3540_; 
wire core__abc_21302_new_n3541_; 
wire core__abc_21302_new_n3542_; 
wire core__abc_21302_new_n3543_; 
wire core__abc_21302_new_n3544_; 
wire core__abc_21302_new_n3545_; 
wire core__abc_21302_new_n3546_; 
wire core__abc_21302_new_n3547_; 
wire core__abc_21302_new_n3548_; 
wire core__abc_21302_new_n3549_; 
wire core__abc_21302_new_n3550_; 
wire core__abc_21302_new_n3551_; 
wire core__abc_21302_new_n3552_; 
wire core__abc_21302_new_n3553_; 
wire core__abc_21302_new_n3554_; 
wire core__abc_21302_new_n3555_; 
wire core__abc_21302_new_n3556_; 
wire core__abc_21302_new_n3557_; 
wire core__abc_21302_new_n3558_; 
wire core__abc_21302_new_n3559_; 
wire core__abc_21302_new_n3560_; 
wire core__abc_21302_new_n3561_; 
wire core__abc_21302_new_n3562_; 
wire core__abc_21302_new_n3563_; 
wire core__abc_21302_new_n3564_; 
wire core__abc_21302_new_n3565_; 
wire core__abc_21302_new_n3566_; 
wire core__abc_21302_new_n3567_; 
wire core__abc_21302_new_n3568_; 
wire core__abc_21302_new_n3569_; 
wire core__abc_21302_new_n3570_; 
wire core__abc_21302_new_n3571_; 
wire core__abc_21302_new_n3573_; 
wire core__abc_21302_new_n3574_; 
wire core__abc_21302_new_n3575_; 
wire core__abc_21302_new_n3576_; 
wire core__abc_21302_new_n3577_; 
wire core__abc_21302_new_n3578_; 
wire core__abc_21302_new_n3579_; 
wire core__abc_21302_new_n3580_; 
wire core__abc_21302_new_n3581_; 
wire core__abc_21302_new_n3582_; 
wire core__abc_21302_new_n3583_; 
wire core__abc_21302_new_n3584_; 
wire core__abc_21302_new_n3585_; 
wire core__abc_21302_new_n3586_; 
wire core__abc_21302_new_n3587_; 
wire core__abc_21302_new_n3588_; 
wire core__abc_21302_new_n3589_; 
wire core__abc_21302_new_n3590_; 
wire core__abc_21302_new_n3591_; 
wire core__abc_21302_new_n3592_; 
wire core__abc_21302_new_n3593_; 
wire core__abc_21302_new_n3594_; 
wire core__abc_21302_new_n3595_; 
wire core__abc_21302_new_n3596_; 
wire core__abc_21302_new_n3597_; 
wire core__abc_21302_new_n3598_; 
wire core__abc_21302_new_n3599_; 
wire core__abc_21302_new_n3600_; 
wire core__abc_21302_new_n3601_; 
wire core__abc_21302_new_n3602_; 
wire core__abc_21302_new_n3604_; 
wire core__abc_21302_new_n3605_; 
wire core__abc_21302_new_n3606_; 
wire core__abc_21302_new_n3607_; 
wire core__abc_21302_new_n3608_; 
wire core__abc_21302_new_n3609_; 
wire core__abc_21302_new_n3610_; 
wire core__abc_21302_new_n3611_; 
wire core__abc_21302_new_n3612_; 
wire core__abc_21302_new_n3613_; 
wire core__abc_21302_new_n3614_; 
wire core__abc_21302_new_n3615_; 
wire core__abc_21302_new_n3616_; 
wire core__abc_21302_new_n3617_; 
wire core__abc_21302_new_n3618_; 
wire core__abc_21302_new_n3619_; 
wire core__abc_21302_new_n3620_; 
wire core__abc_21302_new_n3621_; 
wire core__abc_21302_new_n3622_; 
wire core__abc_21302_new_n3623_; 
wire core__abc_21302_new_n3624_; 
wire core__abc_21302_new_n3625_; 
wire core__abc_21302_new_n3626_; 
wire core__abc_21302_new_n3627_; 
wire core__abc_21302_new_n3628_; 
wire core__abc_21302_new_n3629_; 
wire core__abc_21302_new_n3630_; 
wire core__abc_21302_new_n3631_; 
wire core__abc_21302_new_n3632_; 
wire core__abc_21302_new_n3633_; 
wire core__abc_21302_new_n3634_; 
wire core__abc_21302_new_n3635_; 
wire core__abc_21302_new_n3636_; 
wire core__abc_21302_new_n3637_; 
wire core__abc_21302_new_n3638_; 
wire core__abc_21302_new_n3639_; 
wire core__abc_21302_new_n3640_; 
wire core__abc_21302_new_n3641_; 
wire core__abc_21302_new_n3642_; 
wire core__abc_21302_new_n3643_; 
wire core__abc_21302_new_n3644_; 
wire core__abc_21302_new_n3645_; 
wire core__abc_21302_new_n3646_; 
wire core__abc_21302_new_n3647_; 
wire core__abc_21302_new_n3648_; 
wire core__abc_21302_new_n3649_; 
wire core__abc_21302_new_n3650_; 
wire core__abc_21302_new_n3651_; 
wire core__abc_21302_new_n3652_; 
wire core__abc_21302_new_n3653_; 
wire core__abc_21302_new_n3655_; 
wire core__abc_21302_new_n3656_; 
wire core__abc_21302_new_n3657_; 
wire core__abc_21302_new_n3658_; 
wire core__abc_21302_new_n3659_; 
wire core__abc_21302_new_n3660_; 
wire core__abc_21302_new_n3661_; 
wire core__abc_21302_new_n3662_; 
wire core__abc_21302_new_n3663_; 
wire core__abc_21302_new_n3664_; 
wire core__abc_21302_new_n3665_; 
wire core__abc_21302_new_n3666_; 
wire core__abc_21302_new_n3667_; 
wire core__abc_21302_new_n3668_; 
wire core__abc_21302_new_n3669_; 
wire core__abc_21302_new_n3670_; 
wire core__abc_21302_new_n3671_; 
wire core__abc_21302_new_n3672_; 
wire core__abc_21302_new_n3673_; 
wire core__abc_21302_new_n3674_; 
wire core__abc_21302_new_n3675_; 
wire core__abc_21302_new_n3676_; 
wire core__abc_21302_new_n3677_; 
wire core__abc_21302_new_n3678_; 
wire core__abc_21302_new_n3679_; 
wire core__abc_21302_new_n3680_; 
wire core__abc_21302_new_n3681_; 
wire core__abc_21302_new_n3682_; 
wire core__abc_21302_new_n3683_; 
wire core__abc_21302_new_n3684_; 
wire core__abc_21302_new_n3685_; 
wire core__abc_21302_new_n3687_; 
wire core__abc_21302_new_n3688_; 
wire core__abc_21302_new_n3689_; 
wire core__abc_21302_new_n3690_; 
wire core__abc_21302_new_n3691_; 
wire core__abc_21302_new_n3692_; 
wire core__abc_21302_new_n3693_; 
wire core__abc_21302_new_n3694_; 
wire core__abc_21302_new_n3695_; 
wire core__abc_21302_new_n3696_; 
wire core__abc_21302_new_n3697_; 
wire core__abc_21302_new_n3698_; 
wire core__abc_21302_new_n3699_; 
wire core__abc_21302_new_n3700_; 
wire core__abc_21302_new_n3701_; 
wire core__abc_21302_new_n3702_; 
wire core__abc_21302_new_n3703_; 
wire core__abc_21302_new_n3704_; 
wire core__abc_21302_new_n3705_; 
wire core__abc_21302_new_n3706_; 
wire core__abc_21302_new_n3707_; 
wire core__abc_21302_new_n3708_; 
wire core__abc_21302_new_n3709_; 
wire core__abc_21302_new_n3710_; 
wire core__abc_21302_new_n3711_; 
wire core__abc_21302_new_n3712_; 
wire core__abc_21302_new_n3713_; 
wire core__abc_21302_new_n3714_; 
wire core__abc_21302_new_n3715_; 
wire core__abc_21302_new_n3716_; 
wire core__abc_21302_new_n3717_; 
wire core__abc_21302_new_n3718_; 
wire core__abc_21302_new_n3719_; 
wire core__abc_21302_new_n3720_; 
wire core__abc_21302_new_n3721_; 
wire core__abc_21302_new_n3722_; 
wire core__abc_21302_new_n3723_; 
wire core__abc_21302_new_n3725_; 
wire core__abc_21302_new_n3726_; 
wire core__abc_21302_new_n3727_; 
wire core__abc_21302_new_n3728_; 
wire core__abc_21302_new_n3729_; 
wire core__abc_21302_new_n3730_; 
wire core__abc_21302_new_n3731_; 
wire core__abc_21302_new_n3732_; 
wire core__abc_21302_new_n3733_; 
wire core__abc_21302_new_n3734_; 
wire core__abc_21302_new_n3735_; 
wire core__abc_21302_new_n3736_; 
wire core__abc_21302_new_n3737_; 
wire core__abc_21302_new_n3738_; 
wire core__abc_21302_new_n3739_; 
wire core__abc_21302_new_n3740_; 
wire core__abc_21302_new_n3741_; 
wire core__abc_21302_new_n3742_; 
wire core__abc_21302_new_n3743_; 
wire core__abc_21302_new_n3744_; 
wire core__abc_21302_new_n3745_; 
wire core__abc_21302_new_n3746_; 
wire core__abc_21302_new_n3747_; 
wire core__abc_21302_new_n3748_; 
wire core__abc_21302_new_n3749_; 
wire core__abc_21302_new_n3750_; 
wire core__abc_21302_new_n3751_; 
wire core__abc_21302_new_n3752_; 
wire core__abc_21302_new_n3753_; 
wire core__abc_21302_new_n3754_; 
wire core__abc_21302_new_n3755_; 
wire core__abc_21302_new_n3756_; 
wire core__abc_21302_new_n3757_; 
wire core__abc_21302_new_n3759_; 
wire core__abc_21302_new_n3760_; 
wire core__abc_21302_new_n3761_; 
wire core__abc_21302_new_n3762_; 
wire core__abc_21302_new_n3763_; 
wire core__abc_21302_new_n3764_; 
wire core__abc_21302_new_n3765_; 
wire core__abc_21302_new_n3766_; 
wire core__abc_21302_new_n3767_; 
wire core__abc_21302_new_n3768_; 
wire core__abc_21302_new_n3769_; 
wire core__abc_21302_new_n3770_; 
wire core__abc_21302_new_n3771_; 
wire core__abc_21302_new_n3772_; 
wire core__abc_21302_new_n3773_; 
wire core__abc_21302_new_n3774_; 
wire core__abc_21302_new_n3775_; 
wire core__abc_21302_new_n3776_; 
wire core__abc_21302_new_n3777_; 
wire core__abc_21302_new_n3778_; 
wire core__abc_21302_new_n3779_; 
wire core__abc_21302_new_n3780_; 
wire core__abc_21302_new_n3781_; 
wire core__abc_21302_new_n3782_; 
wire core__abc_21302_new_n3783_; 
wire core__abc_21302_new_n3784_; 
wire core__abc_21302_new_n3785_; 
wire core__abc_21302_new_n3786_; 
wire core__abc_21302_new_n3787_; 
wire core__abc_21302_new_n3788_; 
wire core__abc_21302_new_n3790_; 
wire core__abc_21302_new_n3791_; 
wire core__abc_21302_new_n3792_; 
wire core__abc_21302_new_n3793_; 
wire core__abc_21302_new_n3794_; 
wire core__abc_21302_new_n3795_; 
wire core__abc_21302_new_n3796_; 
wire core__abc_21302_new_n3797_; 
wire core__abc_21302_new_n3798_; 
wire core__abc_21302_new_n3799_; 
wire core__abc_21302_new_n3800_; 
wire core__abc_21302_new_n3801_; 
wire core__abc_21302_new_n3802_; 
wire core__abc_21302_new_n3803_; 
wire core__abc_21302_new_n3804_; 
wire core__abc_21302_new_n3805_; 
wire core__abc_21302_new_n3806_; 
wire core__abc_21302_new_n3807_; 
wire core__abc_21302_new_n3808_; 
wire core__abc_21302_new_n3809_; 
wire core__abc_21302_new_n3810_; 
wire core__abc_21302_new_n3811_; 
wire core__abc_21302_new_n3812_; 
wire core__abc_21302_new_n3813_; 
wire core__abc_21302_new_n3814_; 
wire core__abc_21302_new_n3815_; 
wire core__abc_21302_new_n3816_; 
wire core__abc_21302_new_n3817_; 
wire core__abc_21302_new_n3818_; 
wire core__abc_21302_new_n3819_; 
wire core__abc_21302_new_n3820_; 
wire core__abc_21302_new_n3821_; 
wire core__abc_21302_new_n3822_; 
wire core__abc_21302_new_n3823_; 
wire core__abc_21302_new_n3824_; 
wire core__abc_21302_new_n3825_; 
wire core__abc_21302_new_n3826_; 
wire core__abc_21302_new_n3827_; 
wire core__abc_21302_new_n3828_; 
wire core__abc_21302_new_n3830_; 
wire core__abc_21302_new_n3831_; 
wire core__abc_21302_new_n3832_; 
wire core__abc_21302_new_n3833_; 
wire core__abc_21302_new_n3834_; 
wire core__abc_21302_new_n3835_; 
wire core__abc_21302_new_n3836_; 
wire core__abc_21302_new_n3837_; 
wire core__abc_21302_new_n3838_; 
wire core__abc_21302_new_n3839_; 
wire core__abc_21302_new_n3840_; 
wire core__abc_21302_new_n3841_; 
wire core__abc_21302_new_n3842_; 
wire core__abc_21302_new_n3843_; 
wire core__abc_21302_new_n3844_; 
wire core__abc_21302_new_n3845_; 
wire core__abc_21302_new_n3846_; 
wire core__abc_21302_new_n3847_; 
wire core__abc_21302_new_n3848_; 
wire core__abc_21302_new_n3849_; 
wire core__abc_21302_new_n3850_; 
wire core__abc_21302_new_n3851_; 
wire core__abc_21302_new_n3852_; 
wire core__abc_21302_new_n3853_; 
wire core__abc_21302_new_n3854_; 
wire core__abc_21302_new_n3855_; 
wire core__abc_21302_new_n3856_; 
wire core__abc_21302_new_n3857_; 
wire core__abc_21302_new_n3858_; 
wire core__abc_21302_new_n3859_; 
wire core__abc_21302_new_n3860_; 
wire core__abc_21302_new_n3861_; 
wire core__abc_21302_new_n3862_; 
wire core__abc_21302_new_n3863_; 
wire core__abc_21302_new_n3864_; 
wire core__abc_21302_new_n3865_; 
wire core__abc_21302_new_n3866_; 
wire core__abc_21302_new_n3867_; 
wire core__abc_21302_new_n3868_; 
wire core__abc_21302_new_n3869_; 
wire core__abc_21302_new_n3870_; 
wire core__abc_21302_new_n3871_; 
wire core__abc_21302_new_n3872_; 
wire core__abc_21302_new_n3873_; 
wire core__abc_21302_new_n3874_; 
wire core__abc_21302_new_n3875_; 
wire core__abc_21302_new_n3877_; 
wire core__abc_21302_new_n3878_; 
wire core__abc_21302_new_n3879_; 
wire core__abc_21302_new_n3880_; 
wire core__abc_21302_new_n3881_; 
wire core__abc_21302_new_n3882_; 
wire core__abc_21302_new_n3883_; 
wire core__abc_21302_new_n3884_; 
wire core__abc_21302_new_n3885_; 
wire core__abc_21302_new_n3886_; 
wire core__abc_21302_new_n3887_; 
wire core__abc_21302_new_n3888_; 
wire core__abc_21302_new_n3889_; 
wire core__abc_21302_new_n3890_; 
wire core__abc_21302_new_n3891_; 
wire core__abc_21302_new_n3892_; 
wire core__abc_21302_new_n3893_; 
wire core__abc_21302_new_n3894_; 
wire core__abc_21302_new_n3895_; 
wire core__abc_21302_new_n3896_; 
wire core__abc_21302_new_n3897_; 
wire core__abc_21302_new_n3898_; 
wire core__abc_21302_new_n3899_; 
wire core__abc_21302_new_n3900_; 
wire core__abc_21302_new_n3901_; 
wire core__abc_21302_new_n3902_; 
wire core__abc_21302_new_n3903_; 
wire core__abc_21302_new_n3904_; 
wire core__abc_21302_new_n3905_; 
wire core__abc_21302_new_n3906_; 
wire core__abc_21302_new_n3908_; 
wire core__abc_21302_new_n3909_; 
wire core__abc_21302_new_n3910_; 
wire core__abc_21302_new_n3911_; 
wire core__abc_21302_new_n3912_; 
wire core__abc_21302_new_n3913_; 
wire core__abc_21302_new_n3914_; 
wire core__abc_21302_new_n3915_; 
wire core__abc_21302_new_n3916_; 
wire core__abc_21302_new_n3917_; 
wire core__abc_21302_new_n3918_; 
wire core__abc_21302_new_n3919_; 
wire core__abc_21302_new_n3920_; 
wire core__abc_21302_new_n3921_; 
wire core__abc_21302_new_n3922_; 
wire core__abc_21302_new_n3923_; 
wire core__abc_21302_new_n3924_; 
wire core__abc_21302_new_n3925_; 
wire core__abc_21302_new_n3926_; 
wire core__abc_21302_new_n3927_; 
wire core__abc_21302_new_n3928_; 
wire core__abc_21302_new_n3929_; 
wire core__abc_21302_new_n3930_; 
wire core__abc_21302_new_n3931_; 
wire core__abc_21302_new_n3932_; 
wire core__abc_21302_new_n3933_; 
wire core__abc_21302_new_n3934_; 
wire core__abc_21302_new_n3935_; 
wire core__abc_21302_new_n3936_; 
wire core__abc_21302_new_n3937_; 
wire core__abc_21302_new_n3938_; 
wire core__abc_21302_new_n3939_; 
wire core__abc_21302_new_n3940_; 
wire core__abc_21302_new_n3942_; 
wire core__abc_21302_new_n3943_; 
wire core__abc_21302_new_n3944_; 
wire core__abc_21302_new_n3945_; 
wire core__abc_21302_new_n3946_; 
wire core__abc_21302_new_n3947_; 
wire core__abc_21302_new_n3948_; 
wire core__abc_21302_new_n3949_; 
wire core__abc_21302_new_n3950_; 
wire core__abc_21302_new_n3951_; 
wire core__abc_21302_new_n3952_; 
wire core__abc_21302_new_n3953_; 
wire core__abc_21302_new_n3954_; 
wire core__abc_21302_new_n3955_; 
wire core__abc_21302_new_n3956_; 
wire core__abc_21302_new_n3957_; 
wire core__abc_21302_new_n3958_; 
wire core__abc_21302_new_n3959_; 
wire core__abc_21302_new_n3960_; 
wire core__abc_21302_new_n3961_; 
wire core__abc_21302_new_n3962_; 
wire core__abc_21302_new_n3963_; 
wire core__abc_21302_new_n3964_; 
wire core__abc_21302_new_n3965_; 
wire core__abc_21302_new_n3966_; 
wire core__abc_21302_new_n3967_; 
wire core__abc_21302_new_n3969_; 
wire core__abc_21302_new_n3970_; 
wire core__abc_21302_new_n3971_; 
wire core__abc_21302_new_n3972_; 
wire core__abc_21302_new_n3973_; 
wire core__abc_21302_new_n3974_; 
wire core__abc_21302_new_n3975_; 
wire core__abc_21302_new_n3976_; 
wire core__abc_21302_new_n3977_; 
wire core__abc_21302_new_n3978_; 
wire core__abc_21302_new_n3979_; 
wire core__abc_21302_new_n3980_; 
wire core__abc_21302_new_n3981_; 
wire core__abc_21302_new_n3982_; 
wire core__abc_21302_new_n3983_; 
wire core__abc_21302_new_n3984_; 
wire core__abc_21302_new_n3985_; 
wire core__abc_21302_new_n3986_; 
wire core__abc_21302_new_n3987_; 
wire core__abc_21302_new_n3988_; 
wire core__abc_21302_new_n3989_; 
wire core__abc_21302_new_n3990_; 
wire core__abc_21302_new_n3991_; 
wire core__abc_21302_new_n3992_; 
wire core__abc_21302_new_n3993_; 
wire core__abc_21302_new_n3994_; 
wire core__abc_21302_new_n3995_; 
wire core__abc_21302_new_n3996_; 
wire core__abc_21302_new_n3997_; 
wire core__abc_21302_new_n3998_; 
wire core__abc_21302_new_n3999_; 
wire core__abc_21302_new_n4001_; 
wire core__abc_21302_new_n4002_; 
wire core__abc_21302_new_n4003_; 
wire core__abc_21302_new_n4004_; 
wire core__abc_21302_new_n4005_; 
wire core__abc_21302_new_n4006_; 
wire core__abc_21302_new_n4007_; 
wire core__abc_21302_new_n4008_; 
wire core__abc_21302_new_n4009_; 
wire core__abc_21302_new_n4010_; 
wire core__abc_21302_new_n4011_; 
wire core__abc_21302_new_n4012_; 
wire core__abc_21302_new_n4013_; 
wire core__abc_21302_new_n4014_; 
wire core__abc_21302_new_n4015_; 
wire core__abc_21302_new_n4016_; 
wire core__abc_21302_new_n4017_; 
wire core__abc_21302_new_n4018_; 
wire core__abc_21302_new_n4019_; 
wire core__abc_21302_new_n4020_; 
wire core__abc_21302_new_n4021_; 
wire core__abc_21302_new_n4022_; 
wire core__abc_21302_new_n4023_; 
wire core__abc_21302_new_n4024_; 
wire core__abc_21302_new_n4025_; 
wire core__abc_21302_new_n4026_; 
wire core__abc_21302_new_n4027_; 
wire core__abc_21302_new_n4028_; 
wire core__abc_21302_new_n4030_; 
wire core__abc_21302_new_n4031_; 
wire core__abc_21302_new_n4032_; 
wire core__abc_21302_new_n4033_; 
wire core__abc_21302_new_n4034_; 
wire core__abc_21302_new_n4035_; 
wire core__abc_21302_new_n4036_; 
wire core__abc_21302_new_n4037_; 
wire core__abc_21302_new_n4038_; 
wire core__abc_21302_new_n4039_; 
wire core__abc_21302_new_n4040_; 
wire core__abc_21302_new_n4041_; 
wire core__abc_21302_new_n4042_; 
wire core__abc_21302_new_n4043_; 
wire core__abc_21302_new_n4044_; 
wire core__abc_21302_new_n4045_; 
wire core__abc_21302_new_n4046_; 
wire core__abc_21302_new_n4047_; 
wire core__abc_21302_new_n4048_; 
wire core__abc_21302_new_n4049_; 
wire core__abc_21302_new_n4050_; 
wire core__abc_21302_new_n4051_; 
wire core__abc_21302_new_n4052_; 
wire core__abc_21302_new_n4053_; 
wire core__abc_21302_new_n4054_; 
wire core__abc_21302_new_n4055_; 
wire core__abc_21302_new_n4056_; 
wire core__abc_21302_new_n4057_; 
wire core__abc_21302_new_n4058_; 
wire core__abc_21302_new_n4059_; 
wire core__abc_21302_new_n4060_; 
wire core__abc_21302_new_n4062_; 
wire core__abc_21302_new_n4063_; 
wire core__abc_21302_new_n4064_; 
wire core__abc_21302_new_n4065_; 
wire core__abc_21302_new_n4066_; 
wire core__abc_21302_new_n4067_; 
wire core__abc_21302_new_n4068_; 
wire core__abc_21302_new_n4069_; 
wire core__abc_21302_new_n4070_; 
wire core__abc_21302_new_n4071_; 
wire core__abc_21302_new_n4072_; 
wire core__abc_21302_new_n4073_; 
wire core__abc_21302_new_n4074_; 
wire core__abc_21302_new_n4075_; 
wire core__abc_21302_new_n4076_; 
wire core__abc_21302_new_n4077_; 
wire core__abc_21302_new_n4078_; 
wire core__abc_21302_new_n4079_; 
wire core__abc_21302_new_n4080_; 
wire core__abc_21302_new_n4081_; 
wire core__abc_21302_new_n4082_; 
wire core__abc_21302_new_n4083_; 
wire core__abc_21302_new_n4084_; 
wire core__abc_21302_new_n4085_; 
wire core__abc_21302_new_n4086_; 
wire core__abc_21302_new_n4087_; 
wire core__abc_21302_new_n4088_; 
wire core__abc_21302_new_n4090_; 
wire core__abc_21302_new_n4091_; 
wire core__abc_21302_new_n4092_; 
wire core__abc_21302_new_n4093_; 
wire core__abc_21302_new_n4094_; 
wire core__abc_21302_new_n4095_; 
wire core__abc_21302_new_n4096_; 
wire core__abc_21302_new_n4097_; 
wire core__abc_21302_new_n4098_; 
wire core__abc_21302_new_n4099_; 
wire core__abc_21302_new_n4100_; 
wire core__abc_21302_new_n4101_; 
wire core__abc_21302_new_n4102_; 
wire core__abc_21302_new_n4103_; 
wire core__abc_21302_new_n4104_; 
wire core__abc_21302_new_n4105_; 
wire core__abc_21302_new_n4106_; 
wire core__abc_21302_new_n4107_; 
wire core__abc_21302_new_n4108_; 
wire core__abc_21302_new_n4109_; 
wire core__abc_21302_new_n4110_; 
wire core__abc_21302_new_n4111_; 
wire core__abc_21302_new_n4112_; 
wire core__abc_21302_new_n4113_; 
wire core__abc_21302_new_n4114_; 
wire core__abc_21302_new_n4115_; 
wire core__abc_21302_new_n4116_; 
wire core__abc_21302_new_n4117_; 
wire core__abc_21302_new_n4118_; 
wire core__abc_21302_new_n4119_; 
wire core__abc_21302_new_n4120_; 
wire core__abc_21302_new_n4121_; 
wire core__abc_21302_new_n4122_; 
wire core__abc_21302_new_n4123_; 
wire core__abc_21302_new_n4125_; 
wire core__abc_21302_new_n4126_; 
wire core__abc_21302_new_n4127_; 
wire core__abc_21302_new_n4128_; 
wire core__abc_21302_new_n4129_; 
wire core__abc_21302_new_n4130_; 
wire core__abc_21302_new_n4131_; 
wire core__abc_21302_new_n4132_; 
wire core__abc_21302_new_n4133_; 
wire core__abc_21302_new_n4134_; 
wire core__abc_21302_new_n4135_; 
wire core__abc_21302_new_n4136_; 
wire core__abc_21302_new_n4137_; 
wire core__abc_21302_new_n4138_; 
wire core__abc_21302_new_n4139_; 
wire core__abc_21302_new_n4140_; 
wire core__abc_21302_new_n4141_; 
wire core__abc_21302_new_n4142_; 
wire core__abc_21302_new_n4143_; 
wire core__abc_21302_new_n4144_; 
wire core__abc_21302_new_n4145_; 
wire core__abc_21302_new_n4146_; 
wire core__abc_21302_new_n4147_; 
wire core__abc_21302_new_n4148_; 
wire core__abc_21302_new_n4149_; 
wire core__abc_21302_new_n4150_; 
wire core__abc_21302_new_n4151_; 
wire core__abc_21302_new_n4153_; 
wire core__abc_21302_new_n4154_; 
wire core__abc_21302_new_n4155_; 
wire core__abc_21302_new_n4156_; 
wire core__abc_21302_new_n4157_; 
wire core__abc_21302_new_n4158_; 
wire core__abc_21302_new_n4159_; 
wire core__abc_21302_new_n4160_; 
wire core__abc_21302_new_n4161_; 
wire core__abc_21302_new_n4162_; 
wire core__abc_21302_new_n4163_; 
wire core__abc_21302_new_n4164_; 
wire core__abc_21302_new_n4165_; 
wire core__abc_21302_new_n4166_; 
wire core__abc_21302_new_n4167_; 
wire core__abc_21302_new_n4168_; 
wire core__abc_21302_new_n4169_; 
wire core__abc_21302_new_n4170_; 
wire core__abc_21302_new_n4171_; 
wire core__abc_21302_new_n4172_; 
wire core__abc_21302_new_n4173_; 
wire core__abc_21302_new_n4174_; 
wire core__abc_21302_new_n4175_; 
wire core__abc_21302_new_n4176_; 
wire core__abc_21302_new_n4177_; 
wire core__abc_21302_new_n4178_; 
wire core__abc_21302_new_n4179_; 
wire core__abc_21302_new_n4180_; 
wire core__abc_21302_new_n4181_; 
wire core__abc_21302_new_n4182_; 
wire core__abc_21302_new_n4183_; 
wire core__abc_21302_new_n4184_; 
wire core__abc_21302_new_n4185_; 
wire core__abc_21302_new_n4186_; 
wire core__abc_21302_new_n4187_; 
wire core__abc_21302_new_n4188_; 
wire core__abc_21302_new_n4190_; 
wire core__abc_21302_new_n4191_; 
wire core__abc_21302_new_n4192_; 
wire core__abc_21302_new_n4193_; 
wire core__abc_21302_new_n4194_; 
wire core__abc_21302_new_n4195_; 
wire core__abc_21302_new_n4196_; 
wire core__abc_21302_new_n4197_; 
wire core__abc_21302_new_n4198_; 
wire core__abc_21302_new_n4199_; 
wire core__abc_21302_new_n4200_; 
wire core__abc_21302_new_n4201_; 
wire core__abc_21302_new_n4202_; 
wire core__abc_21302_new_n4203_; 
wire core__abc_21302_new_n4204_; 
wire core__abc_21302_new_n4205_; 
wire core__abc_21302_new_n4206_; 
wire core__abc_21302_new_n4207_; 
wire core__abc_21302_new_n4208_; 
wire core__abc_21302_new_n4209_; 
wire core__abc_21302_new_n4210_; 
wire core__abc_21302_new_n4211_; 
wire core__abc_21302_new_n4212_; 
wire core__abc_21302_new_n4213_; 
wire core__abc_21302_new_n4214_; 
wire core__abc_21302_new_n4215_; 
wire core__abc_21302_new_n4217_; 
wire core__abc_21302_new_n4218_; 
wire core__abc_21302_new_n4219_; 
wire core__abc_21302_new_n4220_; 
wire core__abc_21302_new_n4221_; 
wire core__abc_21302_new_n4222_; 
wire core__abc_21302_new_n4223_; 
wire core__abc_21302_new_n4224_; 
wire core__abc_21302_new_n4225_; 
wire core__abc_21302_new_n4226_; 
wire core__abc_21302_new_n4227_; 
wire core__abc_21302_new_n4228_; 
wire core__abc_21302_new_n4229_; 
wire core__abc_21302_new_n4230_; 
wire core__abc_21302_new_n4231_; 
wire core__abc_21302_new_n4232_; 
wire core__abc_21302_new_n4233_; 
wire core__abc_21302_new_n4234_; 
wire core__abc_21302_new_n4235_; 
wire core__abc_21302_new_n4236_; 
wire core__abc_21302_new_n4237_; 
wire core__abc_21302_new_n4238_; 
wire core__abc_21302_new_n4239_; 
wire core__abc_21302_new_n4240_; 
wire core__abc_21302_new_n4241_; 
wire core__abc_21302_new_n4242_; 
wire core__abc_21302_new_n4243_; 
wire core__abc_21302_new_n4244_; 
wire core__abc_21302_new_n4245_; 
wire core__abc_21302_new_n4246_; 
wire core__abc_21302_new_n4248_; 
wire core__abc_21302_new_n4249_; 
wire core__abc_21302_new_n4250_; 
wire core__abc_21302_new_n4251_; 
wire core__abc_21302_new_n4252_; 
wire core__abc_21302_new_n4253_; 
wire core__abc_21302_new_n4254_; 
wire core__abc_21302_new_n4255_; 
wire core__abc_21302_new_n4256_; 
wire core__abc_21302_new_n4257_; 
wire core__abc_21302_new_n4258_; 
wire core__abc_21302_new_n4259_; 
wire core__abc_21302_new_n4260_; 
wire core__abc_21302_new_n4261_; 
wire core__abc_21302_new_n4262_; 
wire core__abc_21302_new_n4263_; 
wire core__abc_21302_new_n4264_; 
wire core__abc_21302_new_n4265_; 
wire core__abc_21302_new_n4266_; 
wire core__abc_21302_new_n4267_; 
wire core__abc_21302_new_n4268_; 
wire core__abc_21302_new_n4269_; 
wire core__abc_21302_new_n4270_; 
wire core__abc_21302_new_n4271_; 
wire core__abc_21302_new_n4273_; 
wire core__abc_21302_new_n4274_; 
wire core__abc_21302_new_n4275_; 
wire core__abc_21302_new_n4276_; 
wire core__abc_21302_new_n4277_; 
wire core__abc_21302_new_n4278_; 
wire core__abc_21302_new_n4279_; 
wire core__abc_21302_new_n4280_; 
wire core__abc_21302_new_n4281_; 
wire core__abc_21302_new_n4282_; 
wire core__abc_21302_new_n4283_; 
wire core__abc_21302_new_n4284_; 
wire core__abc_21302_new_n4285_; 
wire core__abc_21302_new_n4286_; 
wire core__abc_21302_new_n4287_; 
wire core__abc_21302_new_n4288_; 
wire core__abc_21302_new_n4289_; 
wire core__abc_21302_new_n4290_; 
wire core__abc_21302_new_n4291_; 
wire core__abc_21302_new_n4292_; 
wire core__abc_21302_new_n4293_; 
wire core__abc_21302_new_n4294_; 
wire core__abc_21302_new_n4295_; 
wire core__abc_21302_new_n4296_; 
wire core__abc_21302_new_n4297_; 
wire core__abc_21302_new_n4299_; 
wire core__abc_21302_new_n4300_; 
wire core__abc_21302_new_n4301_; 
wire core__abc_21302_new_n4302_; 
wire core__abc_21302_new_n4303_; 
wire core__abc_21302_new_n4304_; 
wire core__abc_21302_new_n4305_; 
wire core__abc_21302_new_n4306_; 
wire core__abc_21302_new_n4307_; 
wire core__abc_21302_new_n4308_; 
wire core__abc_21302_new_n4309_; 
wire core__abc_21302_new_n4310_; 
wire core__abc_21302_new_n4311_; 
wire core__abc_21302_new_n4312_; 
wire core__abc_21302_new_n4313_; 
wire core__abc_21302_new_n4314_; 
wire core__abc_21302_new_n4315_; 
wire core__abc_21302_new_n4316_; 
wire core__abc_21302_new_n4317_; 
wire core__abc_21302_new_n4318_; 
wire core__abc_21302_new_n4319_; 
wire core__abc_21302_new_n4320_; 
wire core__abc_21302_new_n4322_; 
wire core__abc_21302_new_n4323_; 
wire core__abc_21302_new_n4324_; 
wire core__abc_21302_new_n4325_; 
wire core__abc_21302_new_n4326_; 
wire core__abc_21302_new_n4327_; 
wire core__abc_21302_new_n4328_; 
wire core__abc_21302_new_n4329_; 
wire core__abc_21302_new_n4330_; 
wire core__abc_21302_new_n4331_; 
wire core__abc_21302_new_n4332_; 
wire core__abc_21302_new_n4333_; 
wire core__abc_21302_new_n4334_; 
wire core__abc_21302_new_n4335_; 
wire core__abc_21302_new_n4336_; 
wire core__abc_21302_new_n4337_; 
wire core__abc_21302_new_n4338_; 
wire core__abc_21302_new_n4339_; 
wire core__abc_21302_new_n4340_; 
wire core__abc_21302_new_n4341_; 
wire core__abc_21302_new_n4342_; 
wire core__abc_21302_new_n4343_; 
wire core__abc_21302_new_n4344_; 
wire core__abc_21302_new_n4345_; 
wire core__abc_21302_new_n4346_; 
wire core__abc_21302_new_n4347_; 
wire core__abc_21302_new_n4348_; 
wire core__abc_21302_new_n4349_; 
wire core__abc_21302_new_n4350_; 
wire core__abc_21302_new_n4351_; 
wire core__abc_21302_new_n4352_; 
wire core__abc_21302_new_n4353_; 
wire core__abc_21302_new_n4354_; 
wire core__abc_21302_new_n4355_; 
wire core__abc_21302_new_n4357_; 
wire core__abc_21302_new_n4358_; 
wire core__abc_21302_new_n4359_; 
wire core__abc_21302_new_n4360_; 
wire core__abc_21302_new_n4361_; 
wire core__abc_21302_new_n4362_; 
wire core__abc_21302_new_n4363_; 
wire core__abc_21302_new_n4364_; 
wire core__abc_21302_new_n4365_; 
wire core__abc_21302_new_n4366_; 
wire core__abc_21302_new_n4367_; 
wire core__abc_21302_new_n4368_; 
wire core__abc_21302_new_n4369_; 
wire core__abc_21302_new_n4370_; 
wire core__abc_21302_new_n4371_; 
wire core__abc_21302_new_n4372_; 
wire core__abc_21302_new_n4373_; 
wire core__abc_21302_new_n4374_; 
wire core__abc_21302_new_n4375_; 
wire core__abc_21302_new_n4376_; 
wire core__abc_21302_new_n4377_; 
wire core__abc_21302_new_n4378_; 
wire core__abc_21302_new_n4379_; 
wire core__abc_21302_new_n4380_; 
wire core__abc_21302_new_n4381_; 
wire core__abc_21302_new_n4382_; 
wire core__abc_21302_new_n4384_; 
wire core__abc_21302_new_n4385_; 
wire core__abc_21302_new_n4386_; 
wire core__abc_21302_new_n4387_; 
wire core__abc_21302_new_n4388_; 
wire core__abc_21302_new_n4389_; 
wire core__abc_21302_new_n4390_; 
wire core__abc_21302_new_n4391_; 
wire core__abc_21302_new_n4392_; 
wire core__abc_21302_new_n4393_; 
wire core__abc_21302_new_n4394_; 
wire core__abc_21302_new_n4395_; 
wire core__abc_21302_new_n4396_; 
wire core__abc_21302_new_n4397_; 
wire core__abc_21302_new_n4398_; 
wire core__abc_21302_new_n4399_; 
wire core__abc_21302_new_n4400_; 
wire core__abc_21302_new_n4401_; 
wire core__abc_21302_new_n4402_; 
wire core__abc_21302_new_n4403_; 
wire core__abc_21302_new_n4404_; 
wire core__abc_21302_new_n4405_; 
wire core__abc_21302_new_n4406_; 
wire core__abc_21302_new_n4407_; 
wire core__abc_21302_new_n4408_; 
wire core__abc_21302_new_n4410_; 
wire core__abc_21302_new_n4411_; 
wire core__abc_21302_new_n4412_; 
wire core__abc_21302_new_n4413_; 
wire core__abc_21302_new_n4414_; 
wire core__abc_21302_new_n4415_; 
wire core__abc_21302_new_n4416_; 
wire core__abc_21302_new_n4417_; 
wire core__abc_21302_new_n4418_; 
wire core__abc_21302_new_n4419_; 
wire core__abc_21302_new_n4420_; 
wire core__abc_21302_new_n4421_; 
wire core__abc_21302_new_n4422_; 
wire core__abc_21302_new_n4423_; 
wire core__abc_21302_new_n4424_; 
wire core__abc_21302_new_n4425_; 
wire core__abc_21302_new_n4426_; 
wire core__abc_21302_new_n4427_; 
wire core__abc_21302_new_n4428_; 
wire core__abc_21302_new_n4429_; 
wire core__abc_21302_new_n4430_; 
wire core__abc_21302_new_n4431_; 
wire core__abc_21302_new_n4432_; 
wire core__abc_21302_new_n4433_; 
wire core__abc_21302_new_n4434_; 
wire core__abc_21302_new_n4435_; 
wire core__abc_21302_new_n4436_; 
wire core__abc_21302_new_n4437_; 
wire core__abc_21302_new_n4438_; 
wire core__abc_21302_new_n4439_; 
wire core__abc_21302_new_n4440_; 
wire core__abc_21302_new_n4442_; 
wire core__abc_21302_new_n4443_; 
wire core__abc_21302_new_n4444_; 
wire core__abc_21302_new_n4445_; 
wire core__abc_21302_new_n4446_; 
wire core__abc_21302_new_n4447_; 
wire core__abc_21302_new_n4448_; 
wire core__abc_21302_new_n4449_; 
wire core__abc_21302_new_n4450_; 
wire core__abc_21302_new_n4451_; 
wire core__abc_21302_new_n4452_; 
wire core__abc_21302_new_n4453_; 
wire core__abc_21302_new_n4454_; 
wire core__abc_21302_new_n4455_; 
wire core__abc_21302_new_n4456_; 
wire core__abc_21302_new_n4457_; 
wire core__abc_21302_new_n4458_; 
wire core__abc_21302_new_n4459_; 
wire core__abc_21302_new_n4460_; 
wire core__abc_21302_new_n4461_; 
wire core__abc_21302_new_n4462_; 
wire core__abc_21302_new_n4463_; 
wire core__abc_21302_new_n4464_; 
wire core__abc_21302_new_n4465_; 
wire core__abc_21302_new_n4466_; 
wire core__abc_21302_new_n4467_; 
wire core__abc_21302_new_n4469_; 
wire core__abc_21302_new_n4470_; 
wire core__abc_21302_new_n4471_; 
wire core__abc_21302_new_n4472_; 
wire core__abc_21302_new_n4473_; 
wire core__abc_21302_new_n4474_; 
wire core__abc_21302_new_n4475_; 
wire core__abc_21302_new_n4476_; 
wire core__abc_21302_new_n4477_; 
wire core__abc_21302_new_n4478_; 
wire core__abc_21302_new_n4479_; 
wire core__abc_21302_new_n4480_; 
wire core__abc_21302_new_n4481_; 
wire core__abc_21302_new_n4482_; 
wire core__abc_21302_new_n4483_; 
wire core__abc_21302_new_n4484_; 
wire core__abc_21302_new_n4485_; 
wire core__abc_21302_new_n4486_; 
wire core__abc_21302_new_n4487_; 
wire core__abc_21302_new_n4488_; 
wire core__abc_21302_new_n4489_; 
wire core__abc_21302_new_n4491_; 
wire core__abc_21302_new_n4492_; 
wire core__abc_21302_new_n4493_; 
wire core__abc_21302_new_n4494_; 
wire core__abc_21302_new_n4495_; 
wire core__abc_21302_new_n4496_; 
wire core__abc_21302_new_n4497_; 
wire core__abc_21302_new_n4498_; 
wire core__abc_21302_new_n4499_; 
wire core__abc_21302_new_n4500_; 
wire core__abc_21302_new_n4501_; 
wire core__abc_21302_new_n4502_; 
wire core__abc_21302_new_n4503_; 
wire core__abc_21302_new_n4504_; 
wire core__abc_21302_new_n4505_; 
wire core__abc_21302_new_n4506_; 
wire core__abc_21302_new_n4507_; 
wire core__abc_21302_new_n4508_; 
wire core__abc_21302_new_n4509_; 
wire core__abc_21302_new_n4510_; 
wire core__abc_21302_new_n4511_; 
wire core__abc_21302_new_n4512_; 
wire core__abc_21302_new_n4514_; 
wire core__abc_21302_new_n4515_; 
wire core__abc_21302_new_n4516_; 
wire core__abc_21302_new_n4517_; 
wire core__abc_21302_new_n4518_; 
wire core__abc_21302_new_n4519_; 
wire core__abc_21302_new_n4520_; 
wire core__abc_21302_new_n4521_; 
wire core__abc_21302_new_n4522_; 
wire core__abc_21302_new_n4523_; 
wire core__abc_21302_new_n4524_; 
wire core__abc_21302_new_n4525_; 
wire core__abc_21302_new_n4526_; 
wire core__abc_21302_new_n4527_; 
wire core__abc_21302_new_n4528_; 
wire core__abc_21302_new_n4529_; 
wire core__abc_21302_new_n4530_; 
wire core__abc_21302_new_n4531_; 
wire core__abc_21302_new_n4532_; 
wire core__abc_21302_new_n4533_; 
wire core__abc_21302_new_n4534_; 
wire core__abc_21302_new_n4535_; 
wire core__abc_21302_new_n4536_; 
wire core__abc_21302_new_n4538_; 
wire core__abc_21302_new_n4539_; 
wire core__abc_21302_new_n4540_; 
wire core__abc_21302_new_n4541_; 
wire core__abc_21302_new_n4542_; 
wire core__abc_21302_new_n4543_; 
wire core__abc_21302_new_n4544_; 
wire core__abc_21302_new_n4545_; 
wire core__abc_21302_new_n4546_; 
wire core__abc_21302_new_n4547_; 
wire core__abc_21302_new_n4548_; 
wire core__abc_21302_new_n4549_; 
wire core__abc_21302_new_n4550_; 
wire core__abc_21302_new_n4551_; 
wire core__abc_21302_new_n4552_; 
wire core__abc_21302_new_n4553_; 
wire core__abc_21302_new_n4554_; 
wire core__abc_21302_new_n4555_; 
wire core__abc_21302_new_n4556_; 
wire core__abc_21302_new_n4557_; 
wire core__abc_21302_new_n4558_; 
wire core__abc_21302_new_n4559_; 
wire core__abc_21302_new_n4560_; 
wire core__abc_21302_new_n4561_; 
wire core__abc_21302_new_n4563_; 
wire core__abc_21302_new_n4564_; 
wire core__abc_21302_new_n4565_; 
wire core__abc_21302_new_n4566_; 
wire core__abc_21302_new_n4567_; 
wire core__abc_21302_new_n4568_; 
wire core__abc_21302_new_n4569_; 
wire core__abc_21302_new_n4570_; 
wire core__abc_21302_new_n4571_; 
wire core__abc_21302_new_n4572_; 
wire core__abc_21302_new_n4573_; 
wire core__abc_21302_new_n4574_; 
wire core__abc_21302_new_n4575_; 
wire core__abc_21302_new_n4576_; 
wire core__abc_21302_new_n4577_; 
wire core__abc_21302_new_n4578_; 
wire core__abc_21302_new_n4579_; 
wire core__abc_21302_new_n4580_; 
wire core__abc_21302_new_n4581_; 
wire core__abc_21302_new_n4582_; 
wire core__abc_21302_new_n4583_; 
wire core__abc_21302_new_n4584_; 
wire core__abc_21302_new_n4585_; 
wire core__abc_21302_new_n4586_; 
wire core__abc_21302_new_n4587_; 
wire core__abc_21302_new_n4588_; 
wire core__abc_21302_new_n4589_; 
wire core__abc_21302_new_n4590_; 
wire core__abc_21302_new_n4592_; 
wire core__abc_21302_new_n4593_; 
wire core__abc_21302_new_n4594_; 
wire core__abc_21302_new_n4595_; 
wire core__abc_21302_new_n4596_; 
wire core__abc_21302_new_n4597_; 
wire core__abc_21302_new_n4598_; 
wire core__abc_21302_new_n4599_; 
wire core__abc_21302_new_n4600_; 
wire core__abc_21302_new_n4601_; 
wire core__abc_21302_new_n4602_; 
wire core__abc_21302_new_n4603_; 
wire core__abc_21302_new_n4604_; 
wire core__abc_21302_new_n4605_; 
wire core__abc_21302_new_n4606_; 
wire core__abc_21302_new_n4607_; 
wire core__abc_21302_new_n4608_; 
wire core__abc_21302_new_n4609_; 
wire core__abc_21302_new_n4610_; 
wire core__abc_21302_new_n4611_; 
wire core__abc_21302_new_n4612_; 
wire core__abc_21302_new_n4613_; 
wire core__abc_21302_new_n4614_; 
wire core__abc_21302_new_n4616_; 
wire core__abc_21302_new_n4617_; 
wire core__abc_21302_new_n4618_; 
wire core__abc_21302_new_n4619_; 
wire core__abc_21302_new_n4620_; 
wire core__abc_21302_new_n4621_; 
wire core__abc_21302_new_n4622_; 
wire core__abc_21302_new_n4623_; 
wire core__abc_21302_new_n4624_; 
wire core__abc_21302_new_n4625_; 
wire core__abc_21302_new_n4626_; 
wire core__abc_21302_new_n4627_; 
wire core__abc_21302_new_n4628_; 
wire core__abc_21302_new_n4629_; 
wire core__abc_21302_new_n4630_; 
wire core__abc_21302_new_n4631_; 
wire core__abc_21302_new_n4632_; 
wire core__abc_21302_new_n4633_; 
wire core__abc_21302_new_n4634_; 
wire core__abc_21302_new_n4635_; 
wire core__abc_21302_new_n4636_; 
wire core__abc_21302_new_n4637_; 
wire core__abc_21302_new_n4638_; 
wire core__abc_21302_new_n4639_; 
wire core__abc_21302_new_n4641_; 
wire core__abc_21302_new_n4642_; 
wire core__abc_21302_new_n4643_; 
wire core__abc_21302_new_n4644_; 
wire core__abc_21302_new_n4645_; 
wire core__abc_21302_new_n4646_; 
wire core__abc_21302_new_n4647_; 
wire core__abc_21302_new_n4648_; 
wire core__abc_21302_new_n4649_; 
wire core__abc_21302_new_n4650_; 
wire core__abc_21302_new_n4651_; 
wire core__abc_21302_new_n4652_; 
wire core__abc_21302_new_n4653_; 
wire core__abc_21302_new_n4654_; 
wire core__abc_21302_new_n4655_; 
wire core__abc_21302_new_n4656_; 
wire core__abc_21302_new_n4657_; 
wire core__abc_21302_new_n4658_; 
wire core__abc_21302_new_n4659_; 
wire core__abc_21302_new_n4660_; 
wire core__abc_21302_new_n4661_; 
wire core__abc_21302_new_n4662_; 
wire core__abc_21302_new_n4663_; 
wire core__abc_21302_new_n4664_; 
wire core__abc_21302_new_n4665_; 
wire core__abc_21302_new_n4666_; 
wire core__abc_21302_new_n4667_; 
wire core__abc_21302_new_n4668_; 
wire core__abc_21302_new_n4669_; 
wire core__abc_21302_new_n4671_; 
wire core__abc_21302_new_n4672_; 
wire core__abc_21302_new_n4673_; 
wire core__abc_21302_new_n4674_; 
wire core__abc_21302_new_n4675_; 
wire core__abc_21302_new_n4676_; 
wire core__abc_21302_new_n4677_; 
wire core__abc_21302_new_n4678_; 
wire core__abc_21302_new_n4679_; 
wire core__abc_21302_new_n4680_; 
wire core__abc_21302_new_n4681_; 
wire core__abc_21302_new_n4682_; 
wire core__abc_21302_new_n4683_; 
wire core__abc_21302_new_n4684_; 
wire core__abc_21302_new_n4685_; 
wire core__abc_21302_new_n4686_; 
wire core__abc_21302_new_n4687_; 
wire core__abc_21302_new_n4688_; 
wire core__abc_21302_new_n4689_; 
wire core__abc_21302_new_n4690_; 
wire core__abc_21302_new_n4691_; 
wire core__abc_21302_new_n4692_; 
wire core__abc_21302_new_n4693_; 
wire core__abc_21302_new_n4694_; 
wire core__abc_21302_new_n4695_; 
wire core__abc_21302_new_n4697_; 
wire core__abc_21302_new_n4698_; 
wire core__abc_21302_new_n4699_; 
wire core__abc_21302_new_n4700_; 
wire core__abc_21302_new_n4701_; 
wire core__abc_21302_new_n4702_; 
wire core__abc_21302_new_n4703_; 
wire core__abc_21302_new_n4704_; 
wire core__abc_21302_new_n4705_; 
wire core__abc_21302_new_n4706_; 
wire core__abc_21302_new_n4707_; 
wire core__abc_21302_new_n4708_; 
wire core__abc_21302_new_n4709_; 
wire core__abc_21302_new_n4710_; 
wire core__abc_21302_new_n4711_; 
wire core__abc_21302_new_n4712_; 
wire core__abc_21302_new_n4713_; 
wire core__abc_21302_new_n4714_; 
wire core__abc_21302_new_n4715_; 
wire core__abc_21302_new_n4716_; 
wire core__abc_21302_new_n4717_; 
wire core__abc_21302_new_n4718_; 
wire core__abc_21302_new_n4719_; 
wire core__abc_21302_new_n4720_; 
wire core__abc_21302_new_n4721_; 
wire core__abc_21302_new_n4722_; 
wire core__abc_21302_new_n4723_; 
wire core__abc_21302_new_n4724_; 
wire core__abc_21302_new_n4725_; 
wire core__abc_21302_new_n4726_; 
wire core__abc_21302_new_n4727_; 
wire core__abc_21302_new_n4728_; 
wire core__abc_21302_new_n4730_; 
wire core__abc_21302_new_n4731_; 
wire core__abc_21302_new_n4732_; 
wire core__abc_21302_new_n4733_; 
wire core__abc_21302_new_n4734_; 
wire core__abc_21302_new_n4735_; 
wire core__abc_21302_new_n4736_; 
wire core__abc_21302_new_n4737_; 
wire core__abc_21302_new_n4738_; 
wire core__abc_21302_new_n4739_; 
wire core__abc_21302_new_n4740_; 
wire core__abc_21302_new_n4741_; 
wire core__abc_21302_new_n4742_; 
wire core__abc_21302_new_n4743_; 
wire core__abc_21302_new_n4744_; 
wire core__abc_21302_new_n4745_; 
wire core__abc_21302_new_n4746_; 
wire core__abc_21302_new_n4747_; 
wire core__abc_21302_new_n4748_; 
wire core__abc_21302_new_n4749_; 
wire core__abc_21302_new_n4750_; 
wire core__abc_21302_new_n4751_; 
wire core__abc_21302_new_n4752_; 
wire core__abc_21302_new_n4753_; 
wire core__abc_21302_new_n4754_; 
wire core__abc_21302_new_n4755_; 
wire core__abc_21302_new_n4756_; 
wire core__abc_21302_new_n4757_; 
wire core__abc_21302_new_n4758_; 
wire core__abc_21302_new_n4759_; 
wire core__abc_21302_new_n4760_; 
wire core__abc_21302_new_n4762_; 
wire core__abc_21302_new_n4763_; 
wire core__abc_21302_new_n4764_; 
wire core__abc_21302_new_n4765_; 
wire core__abc_21302_new_n4766_; 
wire core__abc_21302_new_n4767_; 
wire core__abc_21302_new_n4768_; 
wire core__abc_21302_new_n4769_; 
wire core__abc_21302_new_n4770_; 
wire core__abc_21302_new_n4771_; 
wire core__abc_21302_new_n4772_; 
wire core__abc_21302_new_n4773_; 
wire core__abc_21302_new_n4774_; 
wire core__abc_21302_new_n4775_; 
wire core__abc_21302_new_n4776_; 
wire core__abc_21302_new_n4777_; 
wire core__abc_21302_new_n4778_; 
wire core__abc_21302_new_n4779_; 
wire core__abc_21302_new_n4780_; 
wire core__abc_21302_new_n4781_; 
wire core__abc_21302_new_n4782_; 
wire core__abc_21302_new_n4783_; 
wire core__abc_21302_new_n4784_; 
wire core__abc_21302_new_n4785_; 
wire core__abc_21302_new_n4786_; 
wire core__abc_21302_new_n4787_; 
wire core__abc_21302_new_n4788_; 
wire core__abc_21302_new_n4789_; 
wire core__abc_21302_new_n4790_; 
wire core__abc_21302_new_n4791_; 
wire core__abc_21302_new_n4792_; 
wire core__abc_21302_new_n4793_; 
wire core__abc_21302_new_n4795_; 
wire core__abc_21302_new_n4796_; 
wire core__abc_21302_new_n4797_; 
wire core__abc_21302_new_n4798_; 
wire core__abc_21302_new_n4799_; 
wire core__abc_21302_new_n4800_; 
wire core__abc_21302_new_n4801_; 
wire core__abc_21302_new_n4802_; 
wire core__abc_21302_new_n4803_; 
wire core__abc_21302_new_n4804_; 
wire core__abc_21302_new_n4805_; 
wire core__abc_21302_new_n4806_; 
wire core__abc_21302_new_n4807_; 
wire core__abc_21302_new_n4808_; 
wire core__abc_21302_new_n4809_; 
wire core__abc_21302_new_n4810_; 
wire core__abc_21302_new_n4811_; 
wire core__abc_21302_new_n4812_; 
wire core__abc_21302_new_n4813_; 
wire core__abc_21302_new_n4814_; 
wire core__abc_21302_new_n4815_; 
wire core__abc_21302_new_n4816_; 
wire core__abc_21302_new_n4817_; 
wire core__abc_21302_new_n4818_; 
wire core__abc_21302_new_n4819_; 
wire core__abc_21302_new_n4820_; 
wire core__abc_21302_new_n4822_; 
wire core__abc_21302_new_n4823_; 
wire core__abc_21302_new_n4824_; 
wire core__abc_21302_new_n4825_; 
wire core__abc_21302_new_n4826_; 
wire core__abc_21302_new_n4827_; 
wire core__abc_21302_new_n4828_; 
wire core__abc_21302_new_n4829_; 
wire core__abc_21302_new_n4830_; 
wire core__abc_21302_new_n4831_; 
wire core__abc_21302_new_n4832_; 
wire core__abc_21302_new_n4833_; 
wire core__abc_21302_new_n4834_; 
wire core__abc_21302_new_n4835_; 
wire core__abc_21302_new_n4836_; 
wire core__abc_21302_new_n4837_; 
wire core__abc_21302_new_n4838_; 
wire core__abc_21302_new_n4839_; 
wire core__abc_21302_new_n4840_; 
wire core__abc_21302_new_n4841_; 
wire core__abc_21302_new_n4842_; 
wire core__abc_21302_new_n4843_; 
wire core__abc_21302_new_n4844_; 
wire core__abc_21302_new_n4845_; 
wire core__abc_21302_new_n4846_; 
wire core__abc_21302_new_n4847_; 
wire core__abc_21302_new_n4848_; 
wire core__abc_21302_new_n4849_; 
wire core__abc_21302_new_n4850_; 
wire core__abc_21302_new_n4851_; 
wire core__abc_21302_new_n4852_; 
wire core__abc_21302_new_n4853_; 
wire core__abc_21302_new_n4854_; 
wire core__abc_21302_new_n4855_; 
wire core__abc_21302_new_n4856_; 
wire core__abc_21302_new_n4857_; 
wire core__abc_21302_new_n4858_; 
wire core__abc_21302_new_n4859_; 
wire core__abc_21302_new_n4860_; 
wire core__abc_21302_new_n4861_; 
wire core__abc_21302_new_n4862_; 
wire core__abc_21302_new_n4863_; 
wire core__abc_21302_new_n4864_; 
wire core__abc_21302_new_n4865_; 
wire core__abc_21302_new_n4866_; 
wire core__abc_21302_new_n4867_; 
wire core__abc_21302_new_n4868_; 
wire core__abc_21302_new_n4869_; 
wire core__abc_21302_new_n4870_; 
wire core__abc_21302_new_n4871_; 
wire core__abc_21302_new_n4872_; 
wire core__abc_21302_new_n4873_; 
wire core__abc_21302_new_n4874_; 
wire core__abc_21302_new_n4875_; 
wire core__abc_21302_new_n4876_; 
wire core__abc_21302_new_n4877_; 
wire core__abc_21302_new_n4878_; 
wire core__abc_21302_new_n4879_; 
wire core__abc_21302_new_n4880_; 
wire core__abc_21302_new_n4881_; 
wire core__abc_21302_new_n4882_; 
wire core__abc_21302_new_n4883_; 
wire core__abc_21302_new_n4884_; 
wire core__abc_21302_new_n4885_; 
wire core__abc_21302_new_n4886_; 
wire core__abc_21302_new_n4887_; 
wire core__abc_21302_new_n4888_; 
wire core__abc_21302_new_n4889_; 
wire core__abc_21302_new_n4890_; 
wire core__abc_21302_new_n4891_; 
wire core__abc_21302_new_n4892_; 
wire core__abc_21302_new_n4893_; 
wire core__abc_21302_new_n4894_; 
wire core__abc_21302_new_n4895_; 
wire core__abc_21302_new_n4896_; 
wire core__abc_21302_new_n4897_; 
wire core__abc_21302_new_n4898_; 
wire core__abc_21302_new_n4899_; 
wire core__abc_21302_new_n4900_; 
wire core__abc_21302_new_n4901_; 
wire core__abc_21302_new_n4902_; 
wire core__abc_21302_new_n4903_; 
wire core__abc_21302_new_n4904_; 
wire core__abc_21302_new_n4905_; 
wire core__abc_21302_new_n4906_; 
wire core__abc_21302_new_n4907_; 
wire core__abc_21302_new_n4908_; 
wire core__abc_21302_new_n4909_; 
wire core__abc_21302_new_n4910_; 
wire core__abc_21302_new_n4911_; 
wire core__abc_21302_new_n4912_; 
wire core__abc_21302_new_n4913_; 
wire core__abc_21302_new_n4914_; 
wire core__abc_21302_new_n4915_; 
wire core__abc_21302_new_n4916_; 
wire core__abc_21302_new_n4917_; 
wire core__abc_21302_new_n4918_; 
wire core__abc_21302_new_n4919_; 
wire core__abc_21302_new_n4920_; 
wire core__abc_21302_new_n4921_; 
wire core__abc_21302_new_n4922_; 
wire core__abc_21302_new_n4923_; 
wire core__abc_21302_new_n4924_; 
wire core__abc_21302_new_n4925_; 
wire core__abc_21302_new_n4926_; 
wire core__abc_21302_new_n4927_; 
wire core__abc_21302_new_n4928_; 
wire core__abc_21302_new_n4929_; 
wire core__abc_21302_new_n4930_; 
wire core__abc_21302_new_n4931_; 
wire core__abc_21302_new_n4932_; 
wire core__abc_21302_new_n4933_; 
wire core__abc_21302_new_n4934_; 
wire core__abc_21302_new_n4935_; 
wire core__abc_21302_new_n4936_; 
wire core__abc_21302_new_n4937_; 
wire core__abc_21302_new_n4938_; 
wire core__abc_21302_new_n4939_; 
wire core__abc_21302_new_n4940_; 
wire core__abc_21302_new_n4941_; 
wire core__abc_21302_new_n4942_; 
wire core__abc_21302_new_n4943_; 
wire core__abc_21302_new_n4944_; 
wire core__abc_21302_new_n4945_; 
wire core__abc_21302_new_n4946_; 
wire core__abc_21302_new_n4947_; 
wire core__abc_21302_new_n4948_; 
wire core__abc_21302_new_n4949_; 
wire core__abc_21302_new_n4950_; 
wire core__abc_21302_new_n4951_; 
wire core__abc_21302_new_n4952_; 
wire core__abc_21302_new_n4953_; 
wire core__abc_21302_new_n4954_; 
wire core__abc_21302_new_n4955_; 
wire core__abc_21302_new_n4956_; 
wire core__abc_21302_new_n4957_; 
wire core__abc_21302_new_n4958_; 
wire core__abc_21302_new_n4959_; 
wire core__abc_21302_new_n4960_; 
wire core__abc_21302_new_n4961_; 
wire core__abc_21302_new_n4962_; 
wire core__abc_21302_new_n4963_; 
wire core__abc_21302_new_n4964_; 
wire core__abc_21302_new_n4965_; 
wire core__abc_21302_new_n4966_; 
wire core__abc_21302_new_n4967_; 
wire core__abc_21302_new_n4968_; 
wire core__abc_21302_new_n4969_; 
wire core__abc_21302_new_n4970_; 
wire core__abc_21302_new_n4971_; 
wire core__abc_21302_new_n4972_; 
wire core__abc_21302_new_n4973_; 
wire core__abc_21302_new_n4974_; 
wire core__abc_21302_new_n4975_; 
wire core__abc_21302_new_n4976_; 
wire core__abc_21302_new_n4977_; 
wire core__abc_21302_new_n4978_; 
wire core__abc_21302_new_n4979_; 
wire core__abc_21302_new_n4980_; 
wire core__abc_21302_new_n4981_; 
wire core__abc_21302_new_n4982_; 
wire core__abc_21302_new_n4983_; 
wire core__abc_21302_new_n4984_; 
wire core__abc_21302_new_n4985_; 
wire core__abc_21302_new_n4986_; 
wire core__abc_21302_new_n4987_; 
wire core__abc_21302_new_n4988_; 
wire core__abc_21302_new_n4989_; 
wire core__abc_21302_new_n4990_; 
wire core__abc_21302_new_n4991_; 
wire core__abc_21302_new_n4992_; 
wire core__abc_21302_new_n4993_; 
wire core__abc_21302_new_n4994_; 
wire core__abc_21302_new_n4995_; 
wire core__abc_21302_new_n4996_; 
wire core__abc_21302_new_n4997_; 
wire core__abc_21302_new_n4998_; 
wire core__abc_21302_new_n4999_; 
wire core__abc_21302_new_n5000_; 
wire core__abc_21302_new_n5001_; 
wire core__abc_21302_new_n5002_; 
wire core__abc_21302_new_n5003_; 
wire core__abc_21302_new_n5004_; 
wire core__abc_21302_new_n5005_; 
wire core__abc_21302_new_n5006_; 
wire core__abc_21302_new_n5007_; 
wire core__abc_21302_new_n5008_; 
wire core__abc_21302_new_n5009_; 
wire core__abc_21302_new_n5010_; 
wire core__abc_21302_new_n5011_; 
wire core__abc_21302_new_n5012_; 
wire core__abc_21302_new_n5013_; 
wire core__abc_21302_new_n5014_; 
wire core__abc_21302_new_n5015_; 
wire core__abc_21302_new_n5016_; 
wire core__abc_21302_new_n5017_; 
wire core__abc_21302_new_n5018_; 
wire core__abc_21302_new_n5019_; 
wire core__abc_21302_new_n5020_; 
wire core__abc_21302_new_n5021_; 
wire core__abc_21302_new_n5022_; 
wire core__abc_21302_new_n5023_; 
wire core__abc_21302_new_n5024_; 
wire core__abc_21302_new_n5025_; 
wire core__abc_21302_new_n5026_; 
wire core__abc_21302_new_n5027_; 
wire core__abc_21302_new_n5028_; 
wire core__abc_21302_new_n5029_; 
wire core__abc_21302_new_n5030_; 
wire core__abc_21302_new_n5031_; 
wire core__abc_21302_new_n5032_; 
wire core__abc_21302_new_n5033_; 
wire core__abc_21302_new_n5034_; 
wire core__abc_21302_new_n5035_; 
wire core__abc_21302_new_n5036_; 
wire core__abc_21302_new_n5037_; 
wire core__abc_21302_new_n5038_; 
wire core__abc_21302_new_n5039_; 
wire core__abc_21302_new_n5040_; 
wire core__abc_21302_new_n5041_; 
wire core__abc_21302_new_n5042_; 
wire core__abc_21302_new_n5043_; 
wire core__abc_21302_new_n5044_; 
wire core__abc_21302_new_n5045_; 
wire core__abc_21302_new_n5046_; 
wire core__abc_21302_new_n5047_; 
wire core__abc_21302_new_n5048_; 
wire core__abc_21302_new_n5049_; 
wire core__abc_21302_new_n5050_; 
wire core__abc_21302_new_n5051_; 
wire core__abc_21302_new_n5052_; 
wire core__abc_21302_new_n5053_; 
wire core__abc_21302_new_n5054_; 
wire core__abc_21302_new_n5055_; 
wire core__abc_21302_new_n5056_; 
wire core__abc_21302_new_n5057_; 
wire core__abc_21302_new_n5058_; 
wire core__abc_21302_new_n5059_; 
wire core__abc_21302_new_n5060_; 
wire core__abc_21302_new_n5061_; 
wire core__abc_21302_new_n5062_; 
wire core__abc_21302_new_n5063_; 
wire core__abc_21302_new_n5064_; 
wire core__abc_21302_new_n5065_; 
wire core__abc_21302_new_n5066_; 
wire core__abc_21302_new_n5067_; 
wire core__abc_21302_new_n5068_; 
wire core__abc_21302_new_n5069_; 
wire core__abc_21302_new_n5070_; 
wire core__abc_21302_new_n5071_; 
wire core__abc_21302_new_n5072_; 
wire core__abc_21302_new_n5073_; 
wire core__abc_21302_new_n5074_; 
wire core__abc_21302_new_n5075_; 
wire core__abc_21302_new_n5076_; 
wire core__abc_21302_new_n5077_; 
wire core__abc_21302_new_n5078_; 
wire core__abc_21302_new_n5079_; 
wire core__abc_21302_new_n5080_; 
wire core__abc_21302_new_n5081_; 
wire core__abc_21302_new_n5082_; 
wire core__abc_21302_new_n5083_; 
wire core__abc_21302_new_n5084_; 
wire core__abc_21302_new_n5085_; 
wire core__abc_21302_new_n5085__bF_buf0; 
wire core__abc_21302_new_n5085__bF_buf1; 
wire core__abc_21302_new_n5085__bF_buf2; 
wire core__abc_21302_new_n5085__bF_buf3; 
wire core__abc_21302_new_n5085__bF_buf4; 
wire core__abc_21302_new_n5085__bF_buf5; 
wire core__abc_21302_new_n5086_; 
wire core__abc_21302_new_n5088_; 
wire core__abc_21302_new_n5089_; 
wire core__abc_21302_new_n5090_; 
wire core__abc_21302_new_n5091_; 
wire core__abc_21302_new_n5092_; 
wire core__abc_21302_new_n5093_; 
wire core__abc_21302_new_n5094_; 
wire core__abc_21302_new_n5095_; 
wire core__abc_21302_new_n5096_; 
wire core__abc_21302_new_n5097_; 
wire core__abc_21302_new_n5098_; 
wire core__abc_21302_new_n5099_; 
wire core__abc_21302_new_n5100_; 
wire core__abc_21302_new_n5101_; 
wire core__abc_21302_new_n5102_; 
wire core__abc_21302_new_n5104_; 
wire core__abc_21302_new_n5104__bF_buf0; 
wire core__abc_21302_new_n5104__bF_buf1; 
wire core__abc_21302_new_n5104__bF_buf2; 
wire core__abc_21302_new_n5104__bF_buf3; 
wire core__abc_21302_new_n5104__bF_buf4; 
wire core__abc_21302_new_n5104__bF_buf5; 
wire core__abc_21302_new_n5104__bF_buf6; 
wire core__abc_21302_new_n5104__bF_buf7; 
wire core__abc_21302_new_n5105_; 
wire core__abc_21302_new_n5106_; 
wire core__abc_21302_new_n5107_; 
wire core__abc_21302_new_n5108_; 
wire core__abc_21302_new_n5109_; 
wire core__abc_21302_new_n5110_; 
wire core__abc_21302_new_n5111_; 
wire core__abc_21302_new_n5112_; 
wire core__abc_21302_new_n5113_; 
wire core__abc_21302_new_n5114_; 
wire core__abc_21302_new_n5115_; 
wire core__abc_21302_new_n5116_; 
wire core__abc_21302_new_n5117_; 
wire core__abc_21302_new_n5118_; 
wire core__abc_21302_new_n5119_; 
wire core__abc_21302_new_n5120_; 
wire core__abc_21302_new_n5121_; 
wire core__abc_21302_new_n5122_; 
wire core__abc_21302_new_n5123_; 
wire core__abc_21302_new_n5124_; 
wire core__abc_21302_new_n5125_; 
wire core__abc_21302_new_n5126_; 
wire core__abc_21302_new_n5127_; 
wire core__abc_21302_new_n5128_; 
wire core__abc_21302_new_n5129_; 
wire core__abc_21302_new_n5131_; 
wire core__abc_21302_new_n5132_; 
wire core__abc_21302_new_n5133_; 
wire core__abc_21302_new_n5134_; 
wire core__abc_21302_new_n5135_; 
wire core__abc_21302_new_n5136_; 
wire core__abc_21302_new_n5137_; 
wire core__abc_21302_new_n5138_; 
wire core__abc_21302_new_n5139_; 
wire core__abc_21302_new_n5140_; 
wire core__abc_21302_new_n5141_; 
wire core__abc_21302_new_n5142_; 
wire core__abc_21302_new_n5143_; 
wire core__abc_21302_new_n5144_; 
wire core__abc_21302_new_n5145_; 
wire core__abc_21302_new_n5146_; 
wire core__abc_21302_new_n5147_; 
wire core__abc_21302_new_n5148_; 
wire core__abc_21302_new_n5149_; 
wire core__abc_21302_new_n5151_; 
wire core__abc_21302_new_n5152_; 
wire core__abc_21302_new_n5153_; 
wire core__abc_21302_new_n5154_; 
wire core__abc_21302_new_n5155_; 
wire core__abc_21302_new_n5156_; 
wire core__abc_21302_new_n5157_; 
wire core__abc_21302_new_n5158_; 
wire core__abc_21302_new_n5159_; 
wire core__abc_21302_new_n5160_; 
wire core__abc_21302_new_n5161_; 
wire core__abc_21302_new_n5162_; 
wire core__abc_21302_new_n5163_; 
wire core__abc_21302_new_n5164_; 
wire core__abc_21302_new_n5165_; 
wire core__abc_21302_new_n5166_; 
wire core__abc_21302_new_n5167_; 
wire core__abc_21302_new_n5168_; 
wire core__abc_21302_new_n5169_; 
wire core__abc_21302_new_n5170_; 
wire core__abc_21302_new_n5171_; 
wire core__abc_21302_new_n5172_; 
wire core__abc_21302_new_n5174_; 
wire core__abc_21302_new_n5175_; 
wire core__abc_21302_new_n5176_; 
wire core__abc_21302_new_n5177_; 
wire core__abc_21302_new_n5178_; 
wire core__abc_21302_new_n5179_; 
wire core__abc_21302_new_n5180_; 
wire core__abc_21302_new_n5181_; 
wire core__abc_21302_new_n5182_; 
wire core__abc_21302_new_n5183_; 
wire core__abc_21302_new_n5184_; 
wire core__abc_21302_new_n5185_; 
wire core__abc_21302_new_n5187_; 
wire core__abc_21302_new_n5188_; 
wire core__abc_21302_new_n5189_; 
wire core__abc_21302_new_n5190_; 
wire core__abc_21302_new_n5191_; 
wire core__abc_21302_new_n5192_; 
wire core__abc_21302_new_n5193_; 
wire core__abc_21302_new_n5194_; 
wire core__abc_21302_new_n5195_; 
wire core__abc_21302_new_n5196_; 
wire core__abc_21302_new_n5197_; 
wire core__abc_21302_new_n5198_; 
wire core__abc_21302_new_n5199_; 
wire core__abc_21302_new_n5200_; 
wire core__abc_21302_new_n5201_; 
wire core__abc_21302_new_n5202_; 
wire core__abc_21302_new_n5203_; 
wire core__abc_21302_new_n5205_; 
wire core__abc_21302_new_n5206_; 
wire core__abc_21302_new_n5207_; 
wire core__abc_21302_new_n5208_; 
wire core__abc_21302_new_n5209_; 
wire core__abc_21302_new_n5210_; 
wire core__abc_21302_new_n5211_; 
wire core__abc_21302_new_n5212_; 
wire core__abc_21302_new_n5213_; 
wire core__abc_21302_new_n5214_; 
wire core__abc_21302_new_n5215_; 
wire core__abc_21302_new_n5216_; 
wire core__abc_21302_new_n5217_; 
wire core__abc_21302_new_n5218_; 
wire core__abc_21302_new_n5219_; 
wire core__abc_21302_new_n5220_; 
wire core__abc_21302_new_n5221_; 
wire core__abc_21302_new_n5222_; 
wire core__abc_21302_new_n5223_; 
wire core__abc_21302_new_n5224_; 
wire core__abc_21302_new_n5226_; 
wire core__abc_21302_new_n5227_; 
wire core__abc_21302_new_n5228_; 
wire core__abc_21302_new_n5229_; 
wire core__abc_21302_new_n5230_; 
wire core__abc_21302_new_n5231_; 
wire core__abc_21302_new_n5232_; 
wire core__abc_21302_new_n5233_; 
wire core__abc_21302_new_n5234_; 
wire core__abc_21302_new_n5235_; 
wire core__abc_21302_new_n5236_; 
wire core__abc_21302_new_n5237_; 
wire core__abc_21302_new_n5238_; 
wire core__abc_21302_new_n5239_; 
wire core__abc_21302_new_n5240_; 
wire core__abc_21302_new_n5241_; 
wire core__abc_21302_new_n5242_; 
wire core__abc_21302_new_n5243_; 
wire core__abc_21302_new_n5244_; 
wire core__abc_21302_new_n5245_; 
wire core__abc_21302_new_n5246_; 
wire core__abc_21302_new_n5248_; 
wire core__abc_21302_new_n5249_; 
wire core__abc_21302_new_n5250_; 
wire core__abc_21302_new_n5251_; 
wire core__abc_21302_new_n5252_; 
wire core__abc_21302_new_n5253_; 
wire core__abc_21302_new_n5254_; 
wire core__abc_21302_new_n5255_; 
wire core__abc_21302_new_n5256_; 
wire core__abc_21302_new_n5257_; 
wire core__abc_21302_new_n5258_; 
wire core__abc_21302_new_n5259_; 
wire core__abc_21302_new_n5260_; 
wire core__abc_21302_new_n5262_; 
wire core__abc_21302_new_n5263_; 
wire core__abc_21302_new_n5264_; 
wire core__abc_21302_new_n5265_; 
wire core__abc_21302_new_n5266_; 
wire core__abc_21302_new_n5267_; 
wire core__abc_21302_new_n5268_; 
wire core__abc_21302_new_n5269_; 
wire core__abc_21302_new_n5270_; 
wire core__abc_21302_new_n5271_; 
wire core__abc_21302_new_n5272_; 
wire core__abc_21302_new_n5273_; 
wire core__abc_21302_new_n5274_; 
wire core__abc_21302_new_n5275_; 
wire core__abc_21302_new_n5276_; 
wire core__abc_21302_new_n5277_; 
wire core__abc_21302_new_n5278_; 
wire core__abc_21302_new_n5279_; 
wire core__abc_21302_new_n5280_; 
wire core__abc_21302_new_n5281_; 
wire core__abc_21302_new_n5282_; 
wire core__abc_21302_new_n5283_; 
wire core__abc_21302_new_n5285_; 
wire core__abc_21302_new_n5286_; 
wire core__abc_21302_new_n5287_; 
wire core__abc_21302_new_n5288_; 
wire core__abc_21302_new_n5289_; 
wire core__abc_21302_new_n5290_; 
wire core__abc_21302_new_n5291_; 
wire core__abc_21302_new_n5292_; 
wire core__abc_21302_new_n5293_; 
wire core__abc_21302_new_n5294_; 
wire core__abc_21302_new_n5295_; 
wire core__abc_21302_new_n5296_; 
wire core__abc_21302_new_n5297_; 
wire core__abc_21302_new_n5298_; 
wire core__abc_21302_new_n5299_; 
wire core__abc_21302_new_n5300_; 
wire core__abc_21302_new_n5301_; 
wire core__abc_21302_new_n5303_; 
wire core__abc_21302_new_n5304_; 
wire core__abc_21302_new_n5305_; 
wire core__abc_21302_new_n5306_; 
wire core__abc_21302_new_n5307_; 
wire core__abc_21302_new_n5308_; 
wire core__abc_21302_new_n5309_; 
wire core__abc_21302_new_n5310_; 
wire core__abc_21302_new_n5311_; 
wire core__abc_21302_new_n5312_; 
wire core__abc_21302_new_n5313_; 
wire core__abc_21302_new_n5314_; 
wire core__abc_21302_new_n5315_; 
wire core__abc_21302_new_n5316_; 
wire core__abc_21302_new_n5317_; 
wire core__abc_21302_new_n5318_; 
wire core__abc_21302_new_n5319_; 
wire core__abc_21302_new_n5320_; 
wire core__abc_21302_new_n5322_; 
wire core__abc_21302_new_n5323_; 
wire core__abc_21302_new_n5324_; 
wire core__abc_21302_new_n5325_; 
wire core__abc_21302_new_n5326_; 
wire core__abc_21302_new_n5327_; 
wire core__abc_21302_new_n5328_; 
wire core__abc_21302_new_n5329_; 
wire core__abc_21302_new_n5330_; 
wire core__abc_21302_new_n5331_; 
wire core__abc_21302_new_n5332_; 
wire core__abc_21302_new_n5333_; 
wire core__abc_21302_new_n5334_; 
wire core__abc_21302_new_n5335_; 
wire core__abc_21302_new_n5336_; 
wire core__abc_21302_new_n5337_; 
wire core__abc_21302_new_n5338_; 
wire core__abc_21302_new_n5339_; 
wire core__abc_21302_new_n5340_; 
wire core__abc_21302_new_n5342_; 
wire core__abc_21302_new_n5343_; 
wire core__abc_21302_new_n5344_; 
wire core__abc_21302_new_n5345_; 
wire core__abc_21302_new_n5346_; 
wire core__abc_21302_new_n5347_; 
wire core__abc_21302_new_n5348_; 
wire core__abc_21302_new_n5349_; 
wire core__abc_21302_new_n5350_; 
wire core__abc_21302_new_n5351_; 
wire core__abc_21302_new_n5352_; 
wire core__abc_21302_new_n5353_; 
wire core__abc_21302_new_n5354_; 
wire core__abc_21302_new_n5355_; 
wire core__abc_21302_new_n5356_; 
wire core__abc_21302_new_n5357_; 
wire core__abc_21302_new_n5358_; 
wire core__abc_21302_new_n5359_; 
wire core__abc_21302_new_n5360_; 
wire core__abc_21302_new_n5361_; 
wire core__abc_21302_new_n5362_; 
wire core__abc_21302_new_n5363_; 
wire core__abc_21302_new_n5364_; 
wire core__abc_21302_new_n5365_; 
wire core__abc_21302_new_n5366_; 
wire core__abc_21302_new_n5368_; 
wire core__abc_21302_new_n5369_; 
wire core__abc_21302_new_n5370_; 
wire core__abc_21302_new_n5371_; 
wire core__abc_21302_new_n5372_; 
wire core__abc_21302_new_n5373_; 
wire core__abc_21302_new_n5374_; 
wire core__abc_21302_new_n5375_; 
wire core__abc_21302_new_n5376_; 
wire core__abc_21302_new_n5377_; 
wire core__abc_21302_new_n5378_; 
wire core__abc_21302_new_n5379_; 
wire core__abc_21302_new_n5380_; 
wire core__abc_21302_new_n5381_; 
wire core__abc_21302_new_n5382_; 
wire core__abc_21302_new_n5383_; 
wire core__abc_21302_new_n5384_; 
wire core__abc_21302_new_n5385_; 
wire core__abc_21302_new_n5386_; 
wire core__abc_21302_new_n5388_; 
wire core__abc_21302_new_n5389_; 
wire core__abc_21302_new_n5390_; 
wire core__abc_21302_new_n5391_; 
wire core__abc_21302_new_n5392_; 
wire core__abc_21302_new_n5393_; 
wire core__abc_21302_new_n5394_; 
wire core__abc_21302_new_n5395_; 
wire core__abc_21302_new_n5396_; 
wire core__abc_21302_new_n5397_; 
wire core__abc_21302_new_n5398_; 
wire core__abc_21302_new_n5399_; 
wire core__abc_21302_new_n5400_; 
wire core__abc_21302_new_n5401_; 
wire core__abc_21302_new_n5402_; 
wire core__abc_21302_new_n5403_; 
wire core__abc_21302_new_n5404_; 
wire core__abc_21302_new_n5405_; 
wire core__abc_21302_new_n5406_; 
wire core__abc_21302_new_n5407_; 
wire core__abc_21302_new_n5408_; 
wire core__abc_21302_new_n5409_; 
wire core__abc_21302_new_n5410_; 
wire core__abc_21302_new_n5411_; 
wire core__abc_21302_new_n5412_; 
wire core__abc_21302_new_n5413_; 
wire core__abc_21302_new_n5415_; 
wire core__abc_21302_new_n5416_; 
wire core__abc_21302_new_n5417_; 
wire core__abc_21302_new_n5418_; 
wire core__abc_21302_new_n5419_; 
wire core__abc_21302_new_n5420_; 
wire core__abc_21302_new_n5421_; 
wire core__abc_21302_new_n5422_; 
wire core__abc_21302_new_n5423_; 
wire core__abc_21302_new_n5424_; 
wire core__abc_21302_new_n5425_; 
wire core__abc_21302_new_n5426_; 
wire core__abc_21302_new_n5427_; 
wire core__abc_21302_new_n5428_; 
wire core__abc_21302_new_n5429_; 
wire core__abc_21302_new_n5430_; 
wire core__abc_21302_new_n5431_; 
wire core__abc_21302_new_n5432_; 
wire core__abc_21302_new_n5434_; 
wire core__abc_21302_new_n5435_; 
wire core__abc_21302_new_n5436_; 
wire core__abc_21302_new_n5437_; 
wire core__abc_21302_new_n5438_; 
wire core__abc_21302_new_n5439_; 
wire core__abc_21302_new_n5440_; 
wire core__abc_21302_new_n5441_; 
wire core__abc_21302_new_n5442_; 
wire core__abc_21302_new_n5443_; 
wire core__abc_21302_new_n5444_; 
wire core__abc_21302_new_n5445_; 
wire core__abc_21302_new_n5446_; 
wire core__abc_21302_new_n5447_; 
wire core__abc_21302_new_n5448_; 
wire core__abc_21302_new_n5449_; 
wire core__abc_21302_new_n5450_; 
wire core__abc_21302_new_n5451_; 
wire core__abc_21302_new_n5452_; 
wire core__abc_21302_new_n5454_; 
wire core__abc_21302_new_n5455_; 
wire core__abc_21302_new_n5456_; 
wire core__abc_21302_new_n5457_; 
wire core__abc_21302_new_n5458_; 
wire core__abc_21302_new_n5459_; 
wire core__abc_21302_new_n5460_; 
wire core__abc_21302_new_n5461_; 
wire core__abc_21302_new_n5462_; 
wire core__abc_21302_new_n5463_; 
wire core__abc_21302_new_n5464_; 
wire core__abc_21302_new_n5466_; 
wire core__abc_21302_new_n5467_; 
wire core__abc_21302_new_n5468_; 
wire core__abc_21302_new_n5469_; 
wire core__abc_21302_new_n5470_; 
wire core__abc_21302_new_n5471_; 
wire core__abc_21302_new_n5472_; 
wire core__abc_21302_new_n5473_; 
wire core__abc_21302_new_n5474_; 
wire core__abc_21302_new_n5475_; 
wire core__abc_21302_new_n5476_; 
wire core__abc_21302_new_n5477_; 
wire core__abc_21302_new_n5478_; 
wire core__abc_21302_new_n5479_; 
wire core__abc_21302_new_n5480_; 
wire core__abc_21302_new_n5481_; 
wire core__abc_21302_new_n5482_; 
wire core__abc_21302_new_n5483_; 
wire core__abc_21302_new_n5484_; 
wire core__abc_21302_new_n5485_; 
wire core__abc_21302_new_n5486_; 
wire core__abc_21302_new_n5487_; 
wire core__abc_21302_new_n5488_; 
wire core__abc_21302_new_n5489_; 
wire core__abc_21302_new_n5490_; 
wire core__abc_21302_new_n5492_; 
wire core__abc_21302_new_n5493_; 
wire core__abc_21302_new_n5494_; 
wire core__abc_21302_new_n5495_; 
wire core__abc_21302_new_n5496_; 
wire core__abc_21302_new_n5497_; 
wire core__abc_21302_new_n5498_; 
wire core__abc_21302_new_n5499_; 
wire core__abc_21302_new_n5500_; 
wire core__abc_21302_new_n5501_; 
wire core__abc_21302_new_n5502_; 
wire core__abc_21302_new_n5503_; 
wire core__abc_21302_new_n5504_; 
wire core__abc_21302_new_n5505_; 
wire core__abc_21302_new_n5507_; 
wire core__abc_21302_new_n5508_; 
wire core__abc_21302_new_n5509_; 
wire core__abc_21302_new_n5510_; 
wire core__abc_21302_new_n5511_; 
wire core__abc_21302_new_n5512_; 
wire core__abc_21302_new_n5513_; 
wire core__abc_21302_new_n5514_; 
wire core__abc_21302_new_n5515_; 
wire core__abc_21302_new_n5516_; 
wire core__abc_21302_new_n5517_; 
wire core__abc_21302_new_n5518_; 
wire core__abc_21302_new_n5519_; 
wire core__abc_21302_new_n5520_; 
wire core__abc_21302_new_n5521_; 
wire core__abc_21302_new_n5522_; 
wire core__abc_21302_new_n5523_; 
wire core__abc_21302_new_n5524_; 
wire core__abc_21302_new_n5525_; 
wire core__abc_21302_new_n5526_; 
wire core__abc_21302_new_n5528_; 
wire core__abc_21302_new_n5529_; 
wire core__abc_21302_new_n5530_; 
wire core__abc_21302_new_n5531_; 
wire core__abc_21302_new_n5532_; 
wire core__abc_21302_new_n5533_; 
wire core__abc_21302_new_n5534_; 
wire core__abc_21302_new_n5535_; 
wire core__abc_21302_new_n5536_; 
wire core__abc_21302_new_n5537_; 
wire core__abc_21302_new_n5538_; 
wire core__abc_21302_new_n5539_; 
wire core__abc_21302_new_n5540_; 
wire core__abc_21302_new_n5541_; 
wire core__abc_21302_new_n5542_; 
wire core__abc_21302_new_n5543_; 
wire core__abc_21302_new_n5545_; 
wire core__abc_21302_new_n5546_; 
wire core__abc_21302_new_n5547_; 
wire core__abc_21302_new_n5548_; 
wire core__abc_21302_new_n5549_; 
wire core__abc_21302_new_n5550_; 
wire core__abc_21302_new_n5551_; 
wire core__abc_21302_new_n5552_; 
wire core__abc_21302_new_n5553_; 
wire core__abc_21302_new_n5554_; 
wire core__abc_21302_new_n5555_; 
wire core__abc_21302_new_n5556_; 
wire core__abc_21302_new_n5557_; 
wire core__abc_21302_new_n5558_; 
wire core__abc_21302_new_n5559_; 
wire core__abc_21302_new_n5560_; 
wire core__abc_21302_new_n5561_; 
wire core__abc_21302_new_n5562_; 
wire core__abc_21302_new_n5563_; 
wire core__abc_21302_new_n5564_; 
wire core__abc_21302_new_n5565_; 
wire core__abc_21302_new_n5566_; 
wire core__abc_21302_new_n5567_; 
wire core__abc_21302_new_n5568_; 
wire core__abc_21302_new_n5570_; 
wire core__abc_21302_new_n5571_; 
wire core__abc_21302_new_n5572_; 
wire core__abc_21302_new_n5573_; 
wire core__abc_21302_new_n5574_; 
wire core__abc_21302_new_n5575_; 
wire core__abc_21302_new_n5576_; 
wire core__abc_21302_new_n5577_; 
wire core__abc_21302_new_n5578_; 
wire core__abc_21302_new_n5579_; 
wire core__abc_21302_new_n5580_; 
wire core__abc_21302_new_n5581_; 
wire core__abc_21302_new_n5583_; 
wire core__abc_21302_new_n5584_; 
wire core__abc_21302_new_n5585_; 
wire core__abc_21302_new_n5586_; 
wire core__abc_21302_new_n5587_; 
wire core__abc_21302_new_n5588_; 
wire core__abc_21302_new_n5589_; 
wire core__abc_21302_new_n5590_; 
wire core__abc_21302_new_n5591_; 
wire core__abc_21302_new_n5592_; 
wire core__abc_21302_new_n5593_; 
wire core__abc_21302_new_n5594_; 
wire core__abc_21302_new_n5595_; 
wire core__abc_21302_new_n5596_; 
wire core__abc_21302_new_n5597_; 
wire core__abc_21302_new_n5598_; 
wire core__abc_21302_new_n5599_; 
wire core__abc_21302_new_n5601_; 
wire core__abc_21302_new_n5602_; 
wire core__abc_21302_new_n5603_; 
wire core__abc_21302_new_n5604_; 
wire core__abc_21302_new_n5605_; 
wire core__abc_21302_new_n5606_; 
wire core__abc_21302_new_n5607_; 
wire core__abc_21302_new_n5608_; 
wire core__abc_21302_new_n5609_; 
wire core__abc_21302_new_n5610_; 
wire core__abc_21302_new_n5611_; 
wire core__abc_21302_new_n5612_; 
wire core__abc_21302_new_n5613_; 
wire core__abc_21302_new_n5614_; 
wire core__abc_21302_new_n5615_; 
wire core__abc_21302_new_n5617_; 
wire core__abc_21302_new_n5618_; 
wire core__abc_21302_new_n5619_; 
wire core__abc_21302_new_n5620_; 
wire core__abc_21302_new_n5621_; 
wire core__abc_21302_new_n5622_; 
wire core__abc_21302_new_n5623_; 
wire core__abc_21302_new_n5624_; 
wire core__abc_21302_new_n5625_; 
wire core__abc_21302_new_n5626_; 
wire core__abc_21302_new_n5627_; 
wire core__abc_21302_new_n5628_; 
wire core__abc_21302_new_n5629_; 
wire core__abc_21302_new_n5630_; 
wire core__abc_21302_new_n5631_; 
wire core__abc_21302_new_n5632_; 
wire core__abc_21302_new_n5633_; 
wire core__abc_21302_new_n5634_; 
wire core__abc_21302_new_n5635_; 
wire core__abc_21302_new_n5636_; 
wire core__abc_21302_new_n5637_; 
wire core__abc_21302_new_n5638_; 
wire core__abc_21302_new_n5639_; 
wire core__abc_21302_new_n5640_; 
wire core__abc_21302_new_n5641_; 
wire core__abc_21302_new_n5642_; 
wire core__abc_21302_new_n5643_; 
wire core__abc_21302_new_n5645_; 
wire core__abc_21302_new_n5646_; 
wire core__abc_21302_new_n5647_; 
wire core__abc_21302_new_n5648_; 
wire core__abc_21302_new_n5649_; 
wire core__abc_21302_new_n5650_; 
wire core__abc_21302_new_n5651_; 
wire core__abc_21302_new_n5652_; 
wire core__abc_21302_new_n5653_; 
wire core__abc_21302_new_n5654_; 
wire core__abc_21302_new_n5655_; 
wire core__abc_21302_new_n5656_; 
wire core__abc_21302_new_n5657_; 
wire core__abc_21302_new_n5658_; 
wire core__abc_21302_new_n5659_; 
wire core__abc_21302_new_n5660_; 
wire core__abc_21302_new_n5661_; 
wire core__abc_21302_new_n5663_; 
wire core__abc_21302_new_n5664_; 
wire core__abc_21302_new_n5665_; 
wire core__abc_21302_new_n5666_; 
wire core__abc_21302_new_n5667_; 
wire core__abc_21302_new_n5668_; 
wire core__abc_21302_new_n5669_; 
wire core__abc_21302_new_n5670_; 
wire core__abc_21302_new_n5671_; 
wire core__abc_21302_new_n5672_; 
wire core__abc_21302_new_n5673_; 
wire core__abc_21302_new_n5674_; 
wire core__abc_21302_new_n5675_; 
wire core__abc_21302_new_n5676_; 
wire core__abc_21302_new_n5677_; 
wire core__abc_21302_new_n5678_; 
wire core__abc_21302_new_n5679_; 
wire core__abc_21302_new_n5680_; 
wire core__abc_21302_new_n5681_; 
wire core__abc_21302_new_n5683_; 
wire core__abc_21302_new_n5684_; 
wire core__abc_21302_new_n5685_; 
wire core__abc_21302_new_n5686_; 
wire core__abc_21302_new_n5687_; 
wire core__abc_21302_new_n5688_; 
wire core__abc_21302_new_n5689_; 
wire core__abc_21302_new_n5690_; 
wire core__abc_21302_new_n5691_; 
wire core__abc_21302_new_n5692_; 
wire core__abc_21302_new_n5693_; 
wire core__abc_21302_new_n5694_; 
wire core__abc_21302_new_n5695_; 
wire core__abc_21302_new_n5696_; 
wire core__abc_21302_new_n5697_; 
wire core__abc_21302_new_n5699_; 
wire core__abc_21302_new_n5700_; 
wire core__abc_21302_new_n5701_; 
wire core__abc_21302_new_n5702_; 
wire core__abc_21302_new_n5703_; 
wire core__abc_21302_new_n5704_; 
wire core__abc_21302_new_n5706_; 
wire core__abc_21302_new_n5707_; 
wire core__abc_21302_new_n5708_; 
wire core__abc_21302_new_n5709_; 
wire core__abc_21302_new_n5710_; 
wire core__abc_21302_new_n5711_; 
wire core__abc_21302_new_n5712_; 
wire core__abc_21302_new_n5714_; 
wire core__abc_21302_new_n5715_; 
wire core__abc_21302_new_n5716_; 
wire core__abc_21302_new_n5717_; 
wire core__abc_21302_new_n5718_; 
wire core__abc_21302_new_n5720_; 
wire core__abc_21302_new_n5721_; 
wire core__abc_21302_new_n5722_; 
wire core__abc_21302_new_n5723_; 
wire core__abc_21302_new_n5724_; 
wire core__abc_21302_new_n5725_; 
wire core__abc_21302_new_n5726_; 
wire core__abc_21302_new_n5728_; 
wire core__abc_21302_new_n5729_; 
wire core__abc_21302_new_n5730_; 
wire core__abc_21302_new_n5731_; 
wire core__abc_21302_new_n5732_; 
wire core__abc_21302_new_n5733_; 
wire core__abc_21302_new_n5734_; 
wire core__abc_21302_new_n5735_; 
wire core__abc_21302_new_n5737_; 
wire core__abc_21302_new_n5738_; 
wire core__abc_21302_new_n5739_; 
wire core__abc_21302_new_n5740_; 
wire core__abc_21302_new_n5741_; 
wire core__abc_21302_new_n5742_; 
wire core__abc_21302_new_n5743_; 
wire core__abc_21302_new_n5745_; 
wire core__abc_21302_new_n5746_; 
wire core__abc_21302_new_n5747_; 
wire core__abc_21302_new_n5748_; 
wire core__abc_21302_new_n5749_; 
wire core__abc_21302_new_n5750_; 
wire core__abc_21302_new_n5752_; 
wire core__abc_21302_new_n5753_; 
wire core__abc_21302_new_n5754_; 
wire core__abc_21302_new_n5755_; 
wire core__abc_21302_new_n5756_; 
wire core__abc_21302_new_n5757_; 
wire core__abc_21302_new_n5758_; 
wire core__abc_21302_new_n5759_; 
wire core__abc_21302_new_n5760_; 
wire core__abc_21302_new_n5761_; 
wire core__abc_21302_new_n5762_; 
wire core__abc_21302_new_n5764_; 
wire core__abc_21302_new_n5765_; 
wire core__abc_21302_new_n5766_; 
wire core__abc_21302_new_n5767_; 
wire core__abc_21302_new_n5768_; 
wire core__abc_21302_new_n5769_; 
wire core__abc_21302_new_n5770_; 
wire core__abc_21302_new_n5772_; 
wire core__abc_21302_new_n5773_; 
wire core__abc_21302_new_n5774_; 
wire core__abc_21302_new_n5775_; 
wire core__abc_21302_new_n5776_; 
wire core__abc_21302_new_n5777_; 
wire core__abc_21302_new_n5778_; 
wire core__abc_21302_new_n5779_; 
wire core__abc_21302_new_n5780_; 
wire core__abc_21302_new_n5782_; 
wire core__abc_21302_new_n5783_; 
wire core__abc_21302_new_n5784_; 
wire core__abc_21302_new_n5785_; 
wire core__abc_21302_new_n5786_; 
wire core__abc_21302_new_n5787_; 
wire core__abc_21302_new_n5788_; 
wire core__abc_21302_new_n5790_; 
wire core__abc_21302_new_n5791_; 
wire core__abc_21302_new_n5792_; 
wire core__abc_21302_new_n5793_; 
wire core__abc_21302_new_n5794_; 
wire core__abc_21302_new_n5795_; 
wire core__abc_21302_new_n5797_; 
wire core__abc_21302_new_n5798_; 
wire core__abc_21302_new_n5799_; 
wire core__abc_21302_new_n5800_; 
wire core__abc_21302_new_n5801_; 
wire core__abc_21302_new_n5802_; 
wire core__abc_21302_new_n5803_; 
wire core__abc_21302_new_n5804_; 
wire core__abc_21302_new_n5805_; 
wire core__abc_21302_new_n5806_; 
wire core__abc_21302_new_n5807_; 
wire core__abc_21302_new_n5808_; 
wire core__abc_21302_new_n5809_; 
wire core__abc_21302_new_n5811_; 
wire core__abc_21302_new_n5812_; 
wire core__abc_21302_new_n5813_; 
wire core__abc_21302_new_n5814_; 
wire core__abc_21302_new_n5815_; 
wire core__abc_21302_new_n5816_; 
wire core__abc_21302_new_n5817_; 
wire core__abc_21302_new_n5819_; 
wire core__abc_21302_new_n5820_; 
wire core__abc_21302_new_n5821_; 
wire core__abc_21302_new_n5822_; 
wire core__abc_21302_new_n5823_; 
wire core__abc_21302_new_n5824_; 
wire core__abc_21302_new_n5825_; 
wire core__abc_21302_new_n5827_; 
wire core__abc_21302_new_n5828_; 
wire core__abc_21302_new_n5829_; 
wire core__abc_21302_new_n5830_; 
wire core__abc_21302_new_n5831_; 
wire core__abc_21302_new_n5832_; 
wire core__abc_21302_new_n5833_; 
wire core__abc_21302_new_n5834_; 
wire core__abc_21302_new_n5835_; 
wire core__abc_21302_new_n5836_; 
wire core__abc_21302_new_n5838_; 
wire core__abc_21302_new_n5839_; 
wire core__abc_21302_new_n5840_; 
wire core__abc_21302_new_n5841_; 
wire core__abc_21302_new_n5842_; 
wire core__abc_21302_new_n5843_; 
wire core__abc_21302_new_n5844_; 
wire core__abc_21302_new_n5845_; 
wire core__abc_21302_new_n5846_; 
wire core__abc_21302_new_n5847_; 
wire core__abc_21302_new_n5849_; 
wire core__abc_21302_new_n5850_; 
wire core__abc_21302_new_n5851_; 
wire core__abc_21302_new_n5852_; 
wire core__abc_21302_new_n5853_; 
wire core__abc_21302_new_n5854_; 
wire core__abc_21302_new_n5855_; 
wire core__abc_21302_new_n5856_; 
wire core__abc_21302_new_n5858_; 
wire core__abc_21302_new_n5859_; 
wire core__abc_21302_new_n5860_; 
wire core__abc_21302_new_n5861_; 
wire core__abc_21302_new_n5862_; 
wire core__abc_21302_new_n5863_; 
wire core__abc_21302_new_n5864_; 
wire core__abc_21302_new_n5865_; 
wire core__abc_21302_new_n5866_; 
wire core__abc_21302_new_n5867_; 
wire core__abc_21302_new_n5868_; 
wire core__abc_21302_new_n5869_; 
wire core__abc_21302_new_n5871_; 
wire core__abc_21302_new_n5872_; 
wire core__abc_21302_new_n5873_; 
wire core__abc_21302_new_n5874_; 
wire core__abc_21302_new_n5875_; 
wire core__abc_21302_new_n5876_; 
wire core__abc_21302_new_n5878_; 
wire core__abc_21302_new_n5879_; 
wire core__abc_21302_new_n5880_; 
wire core__abc_21302_new_n5881_; 
wire core__abc_21302_new_n5882_; 
wire core__abc_21302_new_n5883_; 
wire core__abc_21302_new_n5884_; 
wire core__abc_21302_new_n5885_; 
wire core__abc_21302_new_n5886_; 
wire core__abc_21302_new_n5887_; 
wire core__abc_21302_new_n5889_; 
wire core__abc_21302_new_n5890_; 
wire core__abc_21302_new_n5891_; 
wire core__abc_21302_new_n5892_; 
wire core__abc_21302_new_n5893_; 
wire core__abc_21302_new_n5894_; 
wire core__abc_21302_new_n5895_; 
wire core__abc_21302_new_n5896_; 
wire core__abc_21302_new_n5897_; 
wire core__abc_21302_new_n5899_; 
wire core__abc_21302_new_n5900_; 
wire core__abc_21302_new_n5901_; 
wire core__abc_21302_new_n5902_; 
wire core__abc_21302_new_n5903_; 
wire core__abc_21302_new_n5904_; 
wire core__abc_21302_new_n5905_; 
wire core__abc_21302_new_n5906_; 
wire core__abc_21302_new_n5907_; 
wire core__abc_21302_new_n5909_; 
wire core__abc_21302_new_n5910_; 
wire core__abc_21302_new_n5911_; 
wire core__abc_21302_new_n5912_; 
wire core__abc_21302_new_n5913_; 
wire core__abc_21302_new_n5914_; 
wire core__abc_21302_new_n5915_; 
wire core__abc_21302_new_n5916_; 
wire core__abc_21302_new_n5917_; 
wire core__abc_21302_new_n5918_; 
wire core__abc_21302_new_n5919_; 
wire core__abc_21302_new_n5921_; 
wire core__abc_21302_new_n5922_; 
wire core__abc_21302_new_n5923_; 
wire core__abc_21302_new_n5924_; 
wire core__abc_21302_new_n5925_; 
wire core__abc_21302_new_n5926_; 
wire core__abc_21302_new_n5927_; 
wire core__abc_21302_new_n5928_; 
wire core__abc_21302_new_n5930_; 
wire core__abc_21302_new_n5931_; 
wire core__abc_21302_new_n5932_; 
wire core__abc_21302_new_n5933_; 
wire core__abc_21302_new_n5934_; 
wire core__abc_21302_new_n5935_; 
wire core__abc_21302_new_n5937_; 
wire core__abc_21302_new_n5938_; 
wire core__abc_21302_new_n5939_; 
wire core__abc_21302_new_n5940_; 
wire core__abc_21302_new_n5941_; 
wire core__abc_21302_new_n5942_; 
wire core__abc_21302_new_n5944_; 
wire core__abc_21302_new_n5945_; 
wire core__abc_21302_new_n5946_; 
wire core__abc_21302_new_n5947_; 
wire core__abc_21302_new_n5948_; 
wire core__abc_21302_new_n5949_; 
wire core__abc_21302_new_n5950_; 
wire core__abc_21302_new_n5951_; 
wire core__abc_21302_new_n5953_; 
wire core__abc_21302_new_n5954_; 
wire core__abc_21302_new_n5955_; 
wire core__abc_21302_new_n5956_; 
wire core__abc_21302_new_n5957_; 
wire core__abc_21302_new_n5958_; 
wire core__abc_21302_new_n5959_; 
wire core__abc_21302_new_n5960_; 
wire core__abc_21302_new_n5961_; 
wire core__abc_21302_new_n5962_; 
wire core__abc_21302_new_n5963_; 
wire core__abc_21302_new_n5965_; 
wire core__abc_21302_new_n5966_; 
wire core__abc_21302_new_n5967_; 
wire core__abc_21302_new_n5968_; 
wire core__abc_21302_new_n5969_; 
wire core__abc_21302_new_n5970_; 
wire core__abc_21302_new_n5971_; 
wire core__abc_21302_new_n5972_; 
wire core__abc_21302_new_n5973_; 
wire core__abc_21302_new_n5974_; 
wire core__abc_21302_new_n5976_; 
wire core__abc_21302_new_n5977_; 
wire core__abc_21302_new_n5978_; 
wire core__abc_21302_new_n5979_; 
wire core__abc_21302_new_n5980_; 
wire core__abc_21302_new_n5981_; 
wire core__abc_21302_new_n5982_; 
wire core__abc_21302_new_n5983_; 
wire core__abc_21302_new_n5985_; 
wire core__abc_21302_new_n5986_; 
wire core__abc_21302_new_n5987_; 
wire core__abc_21302_new_n5988_; 
wire core__abc_21302_new_n5989_; 
wire core__abc_21302_new_n5990_; 
wire core__abc_21302_new_n5991_; 
wire core__abc_21302_new_n5992_; 
wire core__abc_21302_new_n5993_; 
wire core__abc_21302_new_n5995_; 
wire core__abc_21302_new_n5996_; 
wire core__abc_21302_new_n5997_; 
wire core__abc_21302_new_n5998_; 
wire core__abc_21302_new_n5998__bF_buf0; 
wire core__abc_21302_new_n5998__bF_buf1; 
wire core__abc_21302_new_n5998__bF_buf2; 
wire core__abc_21302_new_n5998__bF_buf3; 
wire core__abc_21302_new_n5999_; 
wire core__abc_21302_new_n5999__bF_buf0; 
wire core__abc_21302_new_n5999__bF_buf1; 
wire core__abc_21302_new_n5999__bF_buf2; 
wire core__abc_21302_new_n5999__bF_buf3; 
wire core__abc_21302_new_n5999__bF_buf4; 
wire core__abc_21302_new_n5999__bF_buf5; 
wire core__abc_21302_new_n6000_; 
wire core__abc_21302_new_n6001_; 
wire core__abc_21302_new_n6002_; 
wire core__abc_21302_new_n6003_; 
wire core__abc_21302_new_n6004_; 
wire core__abc_21302_new_n6006_; 
wire core__abc_21302_new_n6007_; 
wire core__abc_21302_new_n6008_; 
wire core__abc_21302_new_n6009_; 
wire core__abc_21302_new_n6009__bF_buf0; 
wire core__abc_21302_new_n6009__bF_buf1; 
wire core__abc_21302_new_n6009__bF_buf2; 
wire core__abc_21302_new_n6009__bF_buf3; 
wire core__abc_21302_new_n6009__bF_buf4; 
wire core__abc_21302_new_n6009__bF_buf5; 
wire core__abc_21302_new_n6009__bF_buf6; 
wire core__abc_21302_new_n6009__bF_buf7; 
wire core__abc_21302_new_n6009__bF_buf8; 
wire core__abc_21302_new_n6009__bF_buf9; 
wire core__abc_21302_new_n6010_; 
wire core__abc_21302_new_n6011_; 
wire core__abc_21302_new_n6012_; 
wire core__abc_21302_new_n6014_; 
wire core__abc_21302_new_n6015_; 
wire core__abc_21302_new_n6016_; 
wire core__abc_21302_new_n6017_; 
wire core__abc_21302_new_n6018_; 
wire core__abc_21302_new_n6019_; 
wire core__abc_21302_new_n6020_; 
wire core__abc_21302_new_n6022_; 
wire core__abc_21302_new_n6023_; 
wire core__abc_21302_new_n6024_; 
wire core__abc_21302_new_n6025_; 
wire core__abc_21302_new_n6026_; 
wire core__abc_21302_new_n6027_; 
wire core__abc_21302_new_n6028_; 
wire core__abc_21302_new_n6030_; 
wire core__abc_21302_new_n6031_; 
wire core__abc_21302_new_n6032_; 
wire core__abc_21302_new_n6033_; 
wire core__abc_21302_new_n6034_; 
wire core__abc_21302_new_n6035_; 
wire core__abc_21302_new_n6036_; 
wire core__abc_21302_new_n6038_; 
wire core__abc_21302_new_n6039_; 
wire core__abc_21302_new_n6040_; 
wire core__abc_21302_new_n6041_; 
wire core__abc_21302_new_n6042_; 
wire core__abc_21302_new_n6043_; 
wire core__abc_21302_new_n6044_; 
wire core__abc_21302_new_n6046_; 
wire core__abc_21302_new_n6047_; 
wire core__abc_21302_new_n6048_; 
wire core__abc_21302_new_n6049_; 
wire core__abc_21302_new_n6050_; 
wire core__abc_21302_new_n6051_; 
wire core__abc_21302_new_n6053_; 
wire core__abc_21302_new_n6054_; 
wire core__abc_21302_new_n6055_; 
wire core__abc_21302_new_n6056_; 
wire core__abc_21302_new_n6057_; 
wire core__abc_21302_new_n6058_; 
wire core__abc_21302_new_n6059_; 
wire core__abc_21302_new_n6061_; 
wire core__abc_21302_new_n6062_; 
wire core__abc_21302_new_n6063_; 
wire core__abc_21302_new_n6064_; 
wire core__abc_21302_new_n6065_; 
wire core__abc_21302_new_n6066_; 
wire core__abc_21302_new_n6068_; 
wire core__abc_21302_new_n6069_; 
wire core__abc_21302_new_n6070_; 
wire core__abc_21302_new_n6071_; 
wire core__abc_21302_new_n6072_; 
wire core__abc_21302_new_n6073_; 
wire core__abc_21302_new_n6075_; 
wire core__abc_21302_new_n6076_; 
wire core__abc_21302_new_n6077_; 
wire core__abc_21302_new_n6078_; 
wire core__abc_21302_new_n6079_; 
wire core__abc_21302_new_n6081_; 
wire core__abc_21302_new_n6082_; 
wire core__abc_21302_new_n6083_; 
wire core__abc_21302_new_n6084_; 
wire core__abc_21302_new_n6085_; 
wire core__abc_21302_new_n6086_; 
wire core__abc_21302_new_n6088_; 
wire core__abc_21302_new_n6089_; 
wire core__abc_21302_new_n6090_; 
wire core__abc_21302_new_n6091_; 
wire core__abc_21302_new_n6092_; 
wire core__abc_21302_new_n6094_; 
wire core__abc_21302_new_n6095_; 
wire core__abc_21302_new_n6096_; 
wire core__abc_21302_new_n6097_; 
wire core__abc_21302_new_n6098_; 
wire core__abc_21302_new_n6100_; 
wire core__abc_21302_new_n6101_; 
wire core__abc_21302_new_n6102_; 
wire core__abc_21302_new_n6103_; 
wire core__abc_21302_new_n6104_; 
wire core__abc_21302_new_n6105_; 
wire core__abc_21302_new_n6107_; 
wire core__abc_21302_new_n6108_; 
wire core__abc_21302_new_n6109_; 
wire core__abc_21302_new_n6110_; 
wire core__abc_21302_new_n6111_; 
wire core__abc_21302_new_n6113_; 
wire core__abc_21302_new_n6114_; 
wire core__abc_21302_new_n6115_; 
wire core__abc_21302_new_n6116_; 
wire core__abc_21302_new_n6117_; 
wire core__abc_21302_new_n6119_; 
wire core__abc_21302_new_n6120_; 
wire core__abc_21302_new_n6121_; 
wire core__abc_21302_new_n6122_; 
wire core__abc_21302_new_n6123_; 
wire core__abc_21302_new_n6125_; 
wire core__abc_21302_new_n6126_; 
wire core__abc_21302_new_n6127_; 
wire core__abc_21302_new_n6128_; 
wire core__abc_21302_new_n6129_; 
wire core__abc_21302_new_n6130_; 
wire core__abc_21302_new_n6132_; 
wire core__abc_21302_new_n6133_; 
wire core__abc_21302_new_n6134_; 
wire core__abc_21302_new_n6135_; 
wire core__abc_21302_new_n6136_; 
wire core__abc_21302_new_n6137_; 
wire core__abc_21302_new_n6139_; 
wire core__abc_21302_new_n6140_; 
wire core__abc_21302_new_n6141_; 
wire core__abc_21302_new_n6142_; 
wire core__abc_21302_new_n6143_; 
wire core__abc_21302_new_n6144_; 
wire core__abc_21302_new_n6145_; 
wire core__abc_21302_new_n6147_; 
wire core__abc_21302_new_n6148_; 
wire core__abc_21302_new_n6149_; 
wire core__abc_21302_new_n6150_; 
wire core__abc_21302_new_n6151_; 
wire core__abc_21302_new_n6153_; 
wire core__abc_21302_new_n6154_; 
wire core__abc_21302_new_n6155_; 
wire core__abc_21302_new_n6156_; 
wire core__abc_21302_new_n6157_; 
wire core__abc_21302_new_n6158_; 
wire core__abc_21302_new_n6160_; 
wire core__abc_21302_new_n6161_; 
wire core__abc_21302_new_n6162_; 
wire core__abc_21302_new_n6163_; 
wire core__abc_21302_new_n6164_; 
wire core__abc_21302_new_n6165_; 
wire core__abc_21302_new_n6167_; 
wire core__abc_21302_new_n6168_; 
wire core__abc_21302_new_n6169_; 
wire core__abc_21302_new_n6170_; 
wire core__abc_21302_new_n6171_; 
wire core__abc_21302_new_n6172_; 
wire core__abc_21302_new_n6174_; 
wire core__abc_21302_new_n6175_; 
wire core__abc_21302_new_n6176_; 
wire core__abc_21302_new_n6177_; 
wire core__abc_21302_new_n6178_; 
wire core__abc_21302_new_n6179_; 
wire core__abc_21302_new_n6181_; 
wire core__abc_21302_new_n6182_; 
wire core__abc_21302_new_n6183_; 
wire core__abc_21302_new_n6184_; 
wire core__abc_21302_new_n6185_; 
wire core__abc_21302_new_n6186_; 
wire core__abc_21302_new_n6188_; 
wire core__abc_21302_new_n6189_; 
wire core__abc_21302_new_n6190_; 
wire core__abc_21302_new_n6191_; 
wire core__abc_21302_new_n6192_; 
wire core__abc_21302_new_n6194_; 
wire core__abc_21302_new_n6195_; 
wire core__abc_21302_new_n6196_; 
wire core__abc_21302_new_n6197_; 
wire core__abc_21302_new_n6198_; 
wire core__abc_21302_new_n6199_; 
wire core__abc_21302_new_n6201_; 
wire core__abc_21302_new_n6202_; 
wire core__abc_21302_new_n6203_; 
wire core__abc_21302_new_n6204_; 
wire core__abc_21302_new_n6205_; 
wire core__abc_21302_new_n6207_; 
wire core__abc_21302_new_n6208_; 
wire core__abc_21302_new_n6209_; 
wire core__abc_21302_new_n6210_; 
wire core__abc_21302_new_n6211_; 
wire core__abc_21302_new_n6212_; 
wire core__abc_21302_new_n6214_; 
wire core__abc_21302_new_n6215_; 
wire core__abc_21302_new_n6216_; 
wire core__abc_21302_new_n6217_; 
wire core__abc_21302_new_n6218_; 
wire core__abc_21302_new_n6220_; 
wire core__abc_21302_new_n6221_; 
wire core__abc_21302_new_n6222_; 
wire core__abc_21302_new_n6223_; 
wire core__abc_21302_new_n6224_; 
wire core__abc_21302_new_n6225_; 
wire core__abc_21302_new_n6227_; 
wire core__abc_21302_new_n6228_; 
wire core__abc_21302_new_n6229_; 
wire core__abc_21302_new_n6230_; 
wire core__abc_21302_new_n6231_; 
wire core__abc_21302_new_n6233_; 
wire core__abc_21302_new_n6234_; 
wire core__abc_21302_new_n6235_; 
wire core__abc_21302_new_n6236_; 
wire core__abc_21302_new_n6237_; 
wire core__abc_21302_new_n6239_; 
wire core__abc_21302_new_n6240_; 
wire core__abc_21302_new_n6241_; 
wire core__abc_21302_new_n6242_; 
wire core__abc_21302_new_n6243_; 
wire core__abc_21302_new_n6245_; 
wire core__abc_21302_new_n6246_; 
wire core__abc_21302_new_n6247_; 
wire core__abc_21302_new_n6248_; 
wire core__abc_21302_new_n6249_; 
wire core__abc_21302_new_n6250_; 
wire core__abc_21302_new_n6252_; 
wire core__abc_21302_new_n6253_; 
wire core__abc_21302_new_n6254_; 
wire core__abc_21302_new_n6255_; 
wire core__abc_21302_new_n6256_; 
wire core__abc_21302_new_n6258_; 
wire core__abc_21302_new_n6259_; 
wire core__abc_21302_new_n6260_; 
wire core__abc_21302_new_n6261_; 
wire core__abc_21302_new_n6262_; 
wire core__abc_21302_new_n6263_; 
wire core__abc_21302_new_n6265_; 
wire core__abc_21302_new_n6266_; 
wire core__abc_21302_new_n6267_; 
wire core__abc_21302_new_n6268_; 
wire core__abc_21302_new_n6269_; 
wire core__abc_21302_new_n6270_; 
wire core__abc_21302_new_n6271_; 
wire core__abc_21302_new_n6272_; 
wire core__abc_21302_new_n6274_; 
wire core__abc_21302_new_n6275_; 
wire core__abc_21302_new_n6276_; 
wire core__abc_21302_new_n6277_; 
wire core__abc_21302_new_n6278_; 
wire core__abc_21302_new_n6279_; 
wire core__abc_21302_new_n6280_; 
wire core__abc_21302_new_n6282_; 
wire core__abc_21302_new_n6283_; 
wire core__abc_21302_new_n6284_; 
wire core__abc_21302_new_n6285_; 
wire core__abc_21302_new_n6286_; 
wire core__abc_21302_new_n6287_; 
wire core__abc_21302_new_n6289_; 
wire core__abc_21302_new_n6290_; 
wire core__abc_21302_new_n6291_; 
wire core__abc_21302_new_n6292_; 
wire core__abc_21302_new_n6293_; 
wire core__abc_21302_new_n6295_; 
wire core__abc_21302_new_n6296_; 
wire core__abc_21302_new_n6297_; 
wire core__abc_21302_new_n6298_; 
wire core__abc_21302_new_n6299_; 
wire core__abc_21302_new_n6301_; 
wire core__abc_21302_new_n6302_; 
wire core__abc_21302_new_n6303_; 
wire core__abc_21302_new_n6304_; 
wire core__abc_21302_new_n6305_; 
wire core__abc_21302_new_n6306_; 
wire core__abc_21302_new_n6307_; 
wire core__abc_21302_new_n6309_; 
wire core__abc_21302_new_n6310_; 
wire core__abc_21302_new_n6311_; 
wire core__abc_21302_new_n6312_; 
wire core__abc_21302_new_n6313_; 
wire core__abc_21302_new_n6314_; 
wire core__abc_21302_new_n6316_; 
wire core__abc_21302_new_n6317_; 
wire core__abc_21302_new_n6318_; 
wire core__abc_21302_new_n6319_; 
wire core__abc_21302_new_n6320_; 
wire core__abc_21302_new_n6321_; 
wire core__abc_21302_new_n6322_; 
wire core__abc_21302_new_n6324_; 
wire core__abc_21302_new_n6325_; 
wire core__abc_21302_new_n6326_; 
wire core__abc_21302_new_n6327_; 
wire core__abc_21302_new_n6328_; 
wire core__abc_21302_new_n6330_; 
wire core__abc_21302_new_n6331_; 
wire core__abc_21302_new_n6332_; 
wire core__abc_21302_new_n6333_; 
wire core__abc_21302_new_n6334_; 
wire core__abc_21302_new_n6335_; 
wire core__abc_21302_new_n6337_; 
wire core__abc_21302_new_n6338_; 
wire core__abc_21302_new_n6339_; 
wire core__abc_21302_new_n6340_; 
wire core__abc_21302_new_n6341_; 
wire core__abc_21302_new_n6342_; 
wire core__abc_21302_new_n6344_; 
wire core__abc_21302_new_n6345_; 
wire core__abc_21302_new_n6346_; 
wire core__abc_21302_new_n6347_; 
wire core__abc_21302_new_n6348_; 
wire core__abc_21302_new_n6349_; 
wire core__abc_21302_new_n6350_; 
wire core__abc_21302_new_n6352_; 
wire core__abc_21302_new_n6353_; 
wire core__abc_21302_new_n6354_; 
wire core__abc_21302_new_n6355_; 
wire core__abc_21302_new_n6356_; 
wire core__abc_21302_new_n6357_; 
wire core__abc_21302_new_n6359_; 
wire core__abc_21302_new_n6360_; 
wire core__abc_21302_new_n6361_; 
wire core__abc_21302_new_n6362_; 
wire core__abc_21302_new_n6363_; 
wire core__abc_21302_new_n6364_; 
wire core__abc_21302_new_n6366_; 
wire core__abc_21302_new_n6367_; 
wire core__abc_21302_new_n6368_; 
wire core__abc_21302_new_n6369_; 
wire core__abc_21302_new_n6370_; 
wire core__abc_21302_new_n6372_; 
wire core__abc_21302_new_n6373_; 
wire core__abc_21302_new_n6374_; 
wire core__abc_21302_new_n6375_; 
wire core__abc_21302_new_n6376_; 
wire core__abc_21302_new_n6378_; 
wire core__abc_21302_new_n6379_; 
wire core__abc_21302_new_n6380_; 
wire core__abc_21302_new_n6381_; 
wire core__abc_21302_new_n6382_; 
wire core__abc_21302_new_n6383_; 
wire core__abc_21302_new_n6384_; 
wire core__abc_21302_new_n6385_; 
wire core__abc_21302_new_n6387_; 
wire core__abc_21302_new_n6388_; 
wire core__abc_21302_new_n6389_; 
wire core__abc_21302_new_n6390_; 
wire core__abc_21302_new_n6391_; 
wire core__abc_21302_new_n6393_; 
wire core__abc_21302_new_n6394_; 
wire core__abc_21302_new_n6395_; 
wire core__abc_21302_new_n6396_; 
wire core__abc_21302_new_n6397_; 
wire core__abc_21302_new_n6398_; 
wire core__abc_21302_new_n6399_; 
wire core__abc_21302_new_n6400_; 
wire core__abc_21302_new_n6402_; 
wire core__abc_21302_new_n6403_; 
wire core__abc_21302_new_n6404_; 
wire core__abc_21302_new_n6405_; 
wire core__abc_21302_new_n6406_; 
wire core__abc_21302_new_n6408_; 
wire core__abc_21302_new_n6409_; 
wire core__abc_21302_new_n6410_; 
wire core__abc_21302_new_n6411_; 
wire core__abc_21302_new_n6412_; 
wire core__abc_21302_new_n6413_; 
wire core__abc_21302_new_n6414_; 
wire core__abc_21302_new_n6415_; 
wire core__abc_21302_new_n6416_; 
wire core__abc_21302_new_n6418_; 
wire core__abc_21302_new_n6419_; 
wire core__abc_21302_new_n6420_; 
wire core__abc_21302_new_n6421_; 
wire core__abc_21302_new_n6422_; 
wire core__abc_21302_new_n6423_; 
wire core__abc_21302_new_n6424_; 
wire core__abc_21302_new_n6425_; 
wire core__abc_21302_new_n6427_; 
wire core__abc_21302_new_n6428_; 
wire core__abc_21302_new_n6429_; 
wire core__abc_21302_new_n6430_; 
wire core__abc_21302_new_n6431_; 
wire core__abc_21302_new_n6433_; 
wire core__abc_21302_new_n6434_; 
wire core__abc_21302_new_n6435_; 
wire core__abc_21302_new_n6436_; 
wire core__abc_21302_new_n6437_; 
wire core__abc_21302_new_n6439_; 
wire core__abc_21302_new_n6440_; 
wire core__abc_21302_new_n6441_; 
wire core__abc_21302_new_n6442_; 
wire core__abc_21302_new_n6443_; 
wire core__abc_21302_new_n6444_; 
wire core__abc_21302_new_n6445_; 
wire core__abc_21302_new_n6446_; 
wire core__abc_21302_new_n6448_; 
wire core__abc_21302_new_n6449_; 
wire core__abc_21302_new_n6449__bF_buf0; 
wire core__abc_21302_new_n6449__bF_buf1; 
wire core__abc_21302_new_n6449__bF_buf2; 
wire core__abc_21302_new_n6449__bF_buf3; 
wire core__abc_21302_new_n6449__bF_buf4; 
wire core__abc_21302_new_n6449__bF_buf5; 
wire core__abc_21302_new_n6449__bF_buf6; 
wire core__abc_21302_new_n6449__bF_buf7; 
wire core__abc_21302_new_n6450_; 
wire core__abc_21302_new_n6450__bF_buf0; 
wire core__abc_21302_new_n6450__bF_buf1; 
wire core__abc_21302_new_n6450__bF_buf2; 
wire core__abc_21302_new_n6450__bF_buf3; 
wire core__abc_21302_new_n6450__bF_buf4; 
wire core__abc_21302_new_n6450__bF_buf5; 
wire core__abc_21302_new_n6450__bF_buf6; 
wire core__abc_21302_new_n6450__bF_buf7; 
wire core__abc_21302_new_n6451_; 
wire core__abc_21302_new_n6452_; 
wire core__abc_21302_new_n6453_; 
wire core__abc_21302_new_n6454_; 
wire core__abc_21302_new_n6455_; 
wire core__abc_21302_new_n6457_; 
wire core__abc_21302_new_n6458_; 
wire core__abc_21302_new_n6459_; 
wire core__abc_21302_new_n6460_; 
wire core__abc_21302_new_n6461_; 
wire core__abc_21302_new_n6462_; 
wire core__abc_21302_new_n6464_; 
wire core__abc_21302_new_n6465_; 
wire core__abc_21302_new_n6466_; 
wire core__abc_21302_new_n6467_; 
wire core__abc_21302_new_n6468_; 
wire core__abc_21302_new_n6469_; 
wire core__abc_21302_new_n6470_; 
wire core__abc_21302_new_n6472_; 
wire core__abc_21302_new_n6473_; 
wire core__abc_21302_new_n6474_; 
wire core__abc_21302_new_n6475_; 
wire core__abc_21302_new_n6476_; 
wire core__abc_21302_new_n6478_; 
wire core__abc_21302_new_n6479_; 
wire core__abc_21302_new_n6480_; 
wire core__abc_21302_new_n6481_; 
wire core__abc_21302_new_n6482_; 
wire core__abc_21302_new_n6483_; 
wire core__abc_21302_new_n6485_; 
wire core__abc_21302_new_n6486_; 
wire core__abc_21302_new_n6487_; 
wire core__abc_21302_new_n6488_; 
wire core__abc_21302_new_n6489_; 
wire core__abc_21302_new_n6490_; 
wire core__abc_21302_new_n6492_; 
wire core__abc_21302_new_n6493_; 
wire core__abc_21302_new_n6494_; 
wire core__abc_21302_new_n6495_; 
wire core__abc_21302_new_n6496_; 
wire core__abc_21302_new_n6497_; 
wire core__abc_21302_new_n6499_; 
wire core__abc_21302_new_n6500_; 
wire core__abc_21302_new_n6501_; 
wire core__abc_21302_new_n6502_; 
wire core__abc_21302_new_n6503_; 
wire core__abc_21302_new_n6504_; 
wire core__abc_21302_new_n6506_; 
wire core__abc_21302_new_n6507_; 
wire core__abc_21302_new_n6508_; 
wire core__abc_21302_new_n6509_; 
wire core__abc_21302_new_n6510_; 
wire core__abc_21302_new_n6511_; 
wire core__abc_21302_new_n6513_; 
wire core__abc_21302_new_n6514_; 
wire core__abc_21302_new_n6515_; 
wire core__abc_21302_new_n6516_; 
wire core__abc_21302_new_n6517_; 
wire core__abc_21302_new_n6518_; 
wire core__abc_21302_new_n6519_; 
wire core__abc_21302_new_n6521_; 
wire core__abc_21302_new_n6522_; 
wire core__abc_21302_new_n6523_; 
wire core__abc_21302_new_n6524_; 
wire core__abc_21302_new_n6525_; 
wire core__abc_21302_new_n6526_; 
wire core__abc_21302_new_n6528_; 
wire core__abc_21302_new_n6529_; 
wire core__abc_21302_new_n6530_; 
wire core__abc_21302_new_n6531_; 
wire core__abc_21302_new_n6532_; 
wire core__abc_21302_new_n6533_; 
wire core__abc_21302_new_n6535_; 
wire core__abc_21302_new_n6536_; 
wire core__abc_21302_new_n6537_; 
wire core__abc_21302_new_n6538_; 
wire core__abc_21302_new_n6539_; 
wire core__abc_21302_new_n6540_; 
wire core__abc_21302_new_n6541_; 
wire core__abc_21302_new_n6543_; 
wire core__abc_21302_new_n6544_; 
wire core__abc_21302_new_n6545_; 
wire core__abc_21302_new_n6546_; 
wire core__abc_21302_new_n6547_; 
wire core__abc_21302_new_n6548_; 
wire core__abc_21302_new_n6550_; 
wire core__abc_21302_new_n6551_; 
wire core__abc_21302_new_n6552_; 
wire core__abc_21302_new_n6553_; 
wire core__abc_21302_new_n6554_; 
wire core__abc_21302_new_n6555_; 
wire core__abc_21302_new_n6557_; 
wire core__abc_21302_new_n6558_; 
wire core__abc_21302_new_n6559_; 
wire core__abc_21302_new_n6560_; 
wire core__abc_21302_new_n6561_; 
wire core__abc_21302_new_n6562_; 
wire core__abc_21302_new_n6564_; 
wire core__abc_21302_new_n6565_; 
wire core__abc_21302_new_n6566_; 
wire core__abc_21302_new_n6567_; 
wire core__abc_21302_new_n6568_; 
wire core__abc_21302_new_n6569_; 
wire core__abc_21302_new_n6571_; 
wire core__abc_21302_new_n6572_; 
wire core__abc_21302_new_n6573_; 
wire core__abc_21302_new_n6574_; 
wire core__abc_21302_new_n6575_; 
wire core__abc_21302_new_n6576_; 
wire core__abc_21302_new_n6578_; 
wire core__abc_21302_new_n6579_; 
wire core__abc_21302_new_n6580_; 
wire core__abc_21302_new_n6581_; 
wire core__abc_21302_new_n6582_; 
wire core__abc_21302_new_n6583_; 
wire core__abc_21302_new_n6584_; 
wire core__abc_21302_new_n6586_; 
wire core__abc_21302_new_n6587_; 
wire core__abc_21302_new_n6588_; 
wire core__abc_21302_new_n6589_; 
wire core__abc_21302_new_n6590_; 
wire core__abc_21302_new_n6591_; 
wire core__abc_21302_new_n6593_; 
wire core__abc_21302_new_n6594_; 
wire core__abc_21302_new_n6595_; 
wire core__abc_21302_new_n6596_; 
wire core__abc_21302_new_n6597_; 
wire core__abc_21302_new_n6598_; 
wire core__abc_21302_new_n6600_; 
wire core__abc_21302_new_n6601_; 
wire core__abc_21302_new_n6602_; 
wire core__abc_21302_new_n6603_; 
wire core__abc_21302_new_n6604_; 
wire core__abc_21302_new_n6605_; 
wire core__abc_21302_new_n6607_; 
wire core__abc_21302_new_n6608_; 
wire core__abc_21302_new_n6609_; 
wire core__abc_21302_new_n6610_; 
wire core__abc_21302_new_n6611_; 
wire core__abc_21302_new_n6612_; 
wire core__abc_21302_new_n6614_; 
wire core__abc_21302_new_n6615_; 
wire core__abc_21302_new_n6616_; 
wire core__abc_21302_new_n6617_; 
wire core__abc_21302_new_n6618_; 
wire core__abc_21302_new_n6619_; 
wire core__abc_21302_new_n6621_; 
wire core__abc_21302_new_n6622_; 
wire core__abc_21302_new_n6623_; 
wire core__abc_21302_new_n6624_; 
wire core__abc_21302_new_n6625_; 
wire core__abc_21302_new_n6626_; 
wire core__abc_21302_new_n6628_; 
wire core__abc_21302_new_n6629_; 
wire core__abc_21302_new_n6630_; 
wire core__abc_21302_new_n6631_; 
wire core__abc_21302_new_n6632_; 
wire core__abc_21302_new_n6633_; 
wire core__abc_21302_new_n6634_; 
wire core__abc_21302_new_n6636_; 
wire core__abc_21302_new_n6637_; 
wire core__abc_21302_new_n6638_; 
wire core__abc_21302_new_n6639_; 
wire core__abc_21302_new_n6640_; 
wire core__abc_21302_new_n6641_; 
wire core__abc_21302_new_n6642_; 
wire core__abc_21302_new_n6644_; 
wire core__abc_21302_new_n6645_; 
wire core__abc_21302_new_n6646_; 
wire core__abc_21302_new_n6647_; 
wire core__abc_21302_new_n6648_; 
wire core__abc_21302_new_n6649_; 
wire core__abc_21302_new_n6650_; 
wire core__abc_21302_new_n6652_; 
wire core__abc_21302_new_n6653_; 
wire core__abc_21302_new_n6654_; 
wire core__abc_21302_new_n6655_; 
wire core__abc_21302_new_n6656_; 
wire core__abc_21302_new_n6657_; 
wire core__abc_21302_new_n6659_; 
wire core__abc_21302_new_n6660_; 
wire core__abc_21302_new_n6661_; 
wire core__abc_21302_new_n6662_; 
wire core__abc_21302_new_n6663_; 
wire core__abc_21302_new_n6664_; 
wire core__abc_21302_new_n6666_; 
wire core__abc_21302_new_n6667_; 
wire core__abc_21302_new_n6668_; 
wire core__abc_21302_new_n6669_; 
wire core__abc_21302_new_n6670_; 
wire core__abc_21302_new_n6671_; 
wire core__abc_21302_new_n6673_; 
wire core__abc_21302_new_n6674_; 
wire core__abc_21302_new_n6675_; 
wire core__abc_21302_new_n6676_; 
wire core__abc_21302_new_n6677_; 
wire core__abc_21302_new_n6678_; 
wire core__abc_21302_new_n6680_; 
wire core__abc_21302_new_n6681_; 
wire core__abc_21302_new_n6682_; 
wire core__abc_21302_new_n6683_; 
wire core__abc_21302_new_n6684_; 
wire core__abc_21302_new_n6686_; 
wire core__abc_21302_new_n6687_; 
wire core__abc_21302_new_n6688_; 
wire core__abc_21302_new_n6689_; 
wire core__abc_21302_new_n6690_; 
wire core__abc_21302_new_n6692_; 
wire core__abc_21302_new_n6693_; 
wire core__abc_21302_new_n6694_; 
wire core__abc_21302_new_n6695_; 
wire core__abc_21302_new_n6696_; 
wire core__abc_21302_new_n6697_; 
wire core__abc_21302_new_n6699_; 
wire core__abc_21302_new_n6700_; 
wire core__abc_21302_new_n6701_; 
wire core__abc_21302_new_n6702_; 
wire core__abc_21302_new_n6703_; 
wire core__abc_21302_new_n6704_; 
wire core__abc_21302_new_n6706_; 
wire core__abc_21302_new_n6707_; 
wire core__abc_21302_new_n6708_; 
wire core__abc_21302_new_n6709_; 
wire core__abc_21302_new_n6710_; 
wire core__abc_21302_new_n6711_; 
wire core__abc_21302_new_n6713_; 
wire core__abc_21302_new_n6714_; 
wire core__abc_21302_new_n6715_; 
wire core__abc_21302_new_n6716_; 
wire core__abc_21302_new_n6717_; 
wire core__abc_21302_new_n6719_; 
wire core__abc_21302_new_n6720_; 
wire core__abc_21302_new_n6721_; 
wire core__abc_21302_new_n6722_; 
wire core__abc_21302_new_n6723_; 
wire core__abc_21302_new_n6724_; 
wire core__abc_21302_new_n6726_; 
wire core__abc_21302_new_n6727_; 
wire core__abc_21302_new_n6728_; 
wire core__abc_21302_new_n6729_; 
wire core__abc_21302_new_n6730_; 
wire core__abc_21302_new_n6731_; 
wire core__abc_21302_new_n6733_; 
wire core__abc_21302_new_n6734_; 
wire core__abc_21302_new_n6735_; 
wire core__abc_21302_new_n6736_; 
wire core__abc_21302_new_n6737_; 
wire core__abc_21302_new_n6739_; 
wire core__abc_21302_new_n6740_; 
wire core__abc_21302_new_n6741_; 
wire core__abc_21302_new_n6742_; 
wire core__abc_21302_new_n6743_; 
wire core__abc_21302_new_n6744_; 
wire core__abc_21302_new_n6745_; 
wire core__abc_21302_new_n6747_; 
wire core__abc_21302_new_n6748_; 
wire core__abc_21302_new_n6749_; 
wire core__abc_21302_new_n6750_; 
wire core__abc_21302_new_n6751_; 
wire core__abc_21302_new_n6752_; 
wire core__abc_21302_new_n6754_; 
wire core__abc_21302_new_n6755_; 
wire core__abc_21302_new_n6756_; 
wire core__abc_21302_new_n6757_; 
wire core__abc_21302_new_n6758_; 
wire core__abc_21302_new_n6759_; 
wire core__abc_21302_new_n6761_; 
wire core__abc_21302_new_n6762_; 
wire core__abc_21302_new_n6763_; 
wire core__abc_21302_new_n6764_; 
wire core__abc_21302_new_n6765_; 
wire core__abc_21302_new_n6766_; 
wire core__abc_21302_new_n6768_; 
wire core__abc_21302_new_n6769_; 
wire core__abc_21302_new_n6770_; 
wire core__abc_21302_new_n6771_; 
wire core__abc_21302_new_n6772_; 
wire core__abc_21302_new_n6773_; 
wire core__abc_21302_new_n6775_; 
wire core__abc_21302_new_n6776_; 
wire core__abc_21302_new_n6777_; 
wire core__abc_21302_new_n6778_; 
wire core__abc_21302_new_n6779_; 
wire core__abc_21302_new_n6780_; 
wire core__abc_21302_new_n6782_; 
wire core__abc_21302_new_n6783_; 
wire core__abc_21302_new_n6784_; 
wire core__abc_21302_new_n6785_; 
wire core__abc_21302_new_n6786_; 
wire core__abc_21302_new_n6787_; 
wire core__abc_21302_new_n6789_; 
wire core__abc_21302_new_n6790_; 
wire core__abc_21302_new_n6791_; 
wire core__abc_21302_new_n6792_; 
wire core__abc_21302_new_n6793_; 
wire core__abc_21302_new_n6795_; 
wire core__abc_21302_new_n6796_; 
wire core__abc_21302_new_n6797_; 
wire core__abc_21302_new_n6798_; 
wire core__abc_21302_new_n6799_; 
wire core__abc_21302_new_n6800_; 
wire core__abc_21302_new_n6802_; 
wire core__abc_21302_new_n6803_; 
wire core__abc_21302_new_n6804_; 
wire core__abc_21302_new_n6805_; 
wire core__abc_21302_new_n6806_; 
wire core__abc_21302_new_n6807_; 
wire core__abc_21302_new_n6809_; 
wire core__abc_21302_new_n6810_; 
wire core__abc_21302_new_n6811_; 
wire core__abc_21302_new_n6812_; 
wire core__abc_21302_new_n6813_; 
wire core__abc_21302_new_n6814_; 
wire core__abc_21302_new_n6816_; 
wire core__abc_21302_new_n6817_; 
wire core__abc_21302_new_n6818_; 
wire core__abc_21302_new_n6819_; 
wire core__abc_21302_new_n6820_; 
wire core__abc_21302_new_n6821_; 
wire core__abc_21302_new_n6822_; 
wire core__abc_21302_new_n6824_; 
wire core__abc_21302_new_n6825_; 
wire core__abc_21302_new_n6826_; 
wire core__abc_21302_new_n6827_; 
wire core__abc_21302_new_n6828_; 
wire core__abc_21302_new_n6829_; 
wire core__abc_21302_new_n6831_; 
wire core__abc_21302_new_n6832_; 
wire core__abc_21302_new_n6833_; 
wire core__abc_21302_new_n6834_; 
wire core__abc_21302_new_n6835_; 
wire core__abc_21302_new_n6836_; 
wire core__abc_21302_new_n6838_; 
wire core__abc_21302_new_n6839_; 
wire core__abc_21302_new_n6840_; 
wire core__abc_21302_new_n6841_; 
wire core__abc_21302_new_n6842_; 
wire core__abc_21302_new_n6843_; 
wire core__abc_21302_new_n6845_; 
wire core__abc_21302_new_n6846_; 
wire core__abc_21302_new_n6847_; 
wire core__abc_21302_new_n6848_; 
wire core__abc_21302_new_n6849_; 
wire core__abc_21302_new_n6850_; 
wire core__abc_21302_new_n6852_; 
wire core__abc_21302_new_n6853_; 
wire core__abc_21302_new_n6854_; 
wire core__abc_21302_new_n6855_; 
wire core__abc_21302_new_n6856_; 
wire core__abc_21302_new_n6857_; 
wire core__abc_21302_new_n6858_; 
wire core__abc_21302_new_n6860_; 
wire core__abc_21302_new_n6861_; 
wire core__abc_21302_new_n6862_; 
wire core__abc_21302_new_n6863_; 
wire core__abc_21302_new_n6864_; 
wire core__abc_21302_new_n6865_; 
wire core__abc_21302_new_n6866_; 
wire core__abc_21302_new_n6868_; 
wire core__abc_21302_new_n6869_; 
wire core__abc_21302_new_n6870_; 
wire core__abc_21302_new_n6871_; 
wire core__abc_21302_new_n6872_; 
wire core__abc_21302_new_n6873_; 
wire core__abc_21302_new_n6874_; 
wire core__abc_21302_new_n6876_; 
wire core__abc_21302_new_n6877_; 
wire core__abc_21302_new_n6878_; 
wire core__abc_21302_new_n6879_; 
wire core__abc_21302_new_n6880_; 
wire core__abc_21302_new_n6881_; 
wire core__abc_21302_new_n6883_; 
wire core__abc_21302_new_n6884_; 
wire core__abc_21302_new_n6885_; 
wire core__abc_21302_new_n6886_; 
wire core__abc_21302_new_n6887_; 
wire core__abc_21302_new_n6888_; 
wire core__abc_21302_new_n6890_; 
wire core__abc_21302_new_n6891_; 
wire core__abc_21302_new_n6892_; 
wire core__abc_21302_new_n6893_; 
wire core__abc_21302_new_n6894_; 
wire core__abc_21302_new_n6895_; 
wire core__abc_21302_new_n6896_; 
wire core__abc_21302_new_n6898_; 
wire core__abc_21302_new_n6899_; 
wire core__abc_21302_new_n6900_; 
wire core__abc_21302_new_n6901_; 
wire core__abc_21302_new_n6902_; 
wire core__abc_21302_new_n6903_; 
wire core__abc_21302_new_n6906_; 
wire core__abc_21302_new_n6907_; 
wire core__abc_21302_new_n6909_; 
wire core__abc_21302_new_n6912_; 
wire core_compress; 
wire core_compression_rounds_0_; 
wire core_compression_rounds_1_; 
wire core_compression_rounds_2_; 
wire core_compression_rounds_3_; 
wire core_final_rounds_0_; 
wire core_final_rounds_1_; 
wire core_final_rounds_2_; 
wire core_final_rounds_3_; 
wire core_finalize; 
wire core_initalize; 
wire core_key_0_; 
wire core_key_100_; 
wire core_key_101_; 
wire core_key_102_; 
wire core_key_103_; 
wire core_key_104_; 
wire core_key_105_; 
wire core_key_106_; 
wire core_key_107_; 
wire core_key_108_; 
wire core_key_109_; 
wire core_key_10_; 
wire core_key_110_; 
wire core_key_111_; 
wire core_key_112_; 
wire core_key_113_; 
wire core_key_114_; 
wire core_key_115_; 
wire core_key_116_; 
wire core_key_117_; 
wire core_key_118_; 
wire core_key_119_; 
wire core_key_11_; 
wire core_key_120_; 
wire core_key_121_; 
wire core_key_122_; 
wire core_key_123_; 
wire core_key_124_; 
wire core_key_125_; 
wire core_key_126_; 
wire core_key_127_; 
wire core_key_12_; 
wire core_key_13_; 
wire core_key_14_; 
wire core_key_15_; 
wire core_key_16_; 
wire core_key_17_; 
wire core_key_18_; 
wire core_key_19_; 
wire core_key_1_; 
wire core_key_20_; 
wire core_key_21_; 
wire core_key_22_; 
wire core_key_23_; 
wire core_key_24_; 
wire core_key_25_; 
wire core_key_26_; 
wire core_key_27_; 
wire core_key_28_; 
wire core_key_29_; 
wire core_key_2_; 
wire core_key_30_; 
wire core_key_31_; 
wire core_key_32_; 
wire core_key_33_; 
wire core_key_34_; 
wire core_key_35_; 
wire core_key_36_; 
wire core_key_37_; 
wire core_key_38_; 
wire core_key_39_; 
wire core_key_3_; 
wire core_key_40_; 
wire core_key_41_; 
wire core_key_42_; 
wire core_key_43_; 
wire core_key_44_; 
wire core_key_45_; 
wire core_key_46_; 
wire core_key_47_; 
wire core_key_48_; 
wire core_key_49_; 
wire core_key_4_; 
wire core_key_50_; 
wire core_key_51_; 
wire core_key_52_; 
wire core_key_53_; 
wire core_key_54_; 
wire core_key_55_; 
wire core_key_56_; 
wire core_key_57_; 
wire core_key_58_; 
wire core_key_59_; 
wire core_key_5_; 
wire core_key_60_; 
wire core_key_61_; 
wire core_key_62_; 
wire core_key_63_; 
wire core_key_64_; 
wire core_key_65_; 
wire core_key_66_; 
wire core_key_67_; 
wire core_key_68_; 
wire core_key_69_; 
wire core_key_6_; 
wire core_key_70_; 
wire core_key_71_; 
wire core_key_72_; 
wire core_key_73_; 
wire core_key_74_; 
wire core_key_75_; 
wire core_key_76_; 
wire core_key_77_; 
wire core_key_78_; 
wire core_key_79_; 
wire core_key_7_; 
wire core_key_80_; 
wire core_key_81_; 
wire core_key_82_; 
wire core_key_83_; 
wire core_key_84_; 
wire core_key_85_; 
wire core_key_86_; 
wire core_key_87_; 
wire core_key_88_; 
wire core_key_89_; 
wire core_key_8_; 
wire core_key_90_; 
wire core_key_91_; 
wire core_key_92_; 
wire core_key_93_; 
wire core_key_94_; 
wire core_key_95_; 
wire core_key_96_; 
wire core_key_97_; 
wire core_key_98_; 
wire core_key_99_; 
wire core_key_9_; 
wire core_long; 
wire core_loop_ctr_reg_0_; 
wire core_loop_ctr_reg_1_; 
wire core_loop_ctr_reg_2_; 
wire core_loop_ctr_reg_3_; 
wire core_mi_0_; 
wire core_mi_10_; 
wire core_mi_11_; 
wire core_mi_12_; 
wire core_mi_13_; 
wire core_mi_14_; 
wire core_mi_15_; 
wire core_mi_16_; 
wire core_mi_17_; 
wire core_mi_18_; 
wire core_mi_19_; 
wire core_mi_1_; 
wire core_mi_20_; 
wire core_mi_21_; 
wire core_mi_22_; 
wire core_mi_23_; 
wire core_mi_24_; 
wire core_mi_25_; 
wire core_mi_26_; 
wire core_mi_27_; 
wire core_mi_28_; 
wire core_mi_29_; 
wire core_mi_2_; 
wire core_mi_30_; 
wire core_mi_31_; 
wire core_mi_32_; 
wire core_mi_33_; 
wire core_mi_34_; 
wire core_mi_35_; 
wire core_mi_36_; 
wire core_mi_37_; 
wire core_mi_38_; 
wire core_mi_39_; 
wire core_mi_3_; 
wire core_mi_40_; 
wire core_mi_41_; 
wire core_mi_42_; 
wire core_mi_43_; 
wire core_mi_44_; 
wire core_mi_45_; 
wire core_mi_46_; 
wire core_mi_47_; 
wire core_mi_48_; 
wire core_mi_49_; 
wire core_mi_4_; 
wire core_mi_50_; 
wire core_mi_51_; 
wire core_mi_52_; 
wire core_mi_53_; 
wire core_mi_54_; 
wire core_mi_55_; 
wire core_mi_56_; 
wire core_mi_57_; 
wire core_mi_58_; 
wire core_mi_59_; 
wire core_mi_5_; 
wire core_mi_60_; 
wire core_mi_61_; 
wire core_mi_62_; 
wire core_mi_63_; 
wire core_mi_6_; 
wire core_mi_7_; 
wire core_mi_8_; 
wire core_mi_9_; 
wire core_mi_reg_0_; 
wire core_mi_reg_10_; 
wire core_mi_reg_11_; 
wire core_mi_reg_12_; 
wire core_mi_reg_13_; 
wire core_mi_reg_14_; 
wire core_mi_reg_15_; 
wire core_mi_reg_16_; 
wire core_mi_reg_17_; 
wire core_mi_reg_18_; 
wire core_mi_reg_19_; 
wire core_mi_reg_1_; 
wire core_mi_reg_20_; 
wire core_mi_reg_21_; 
wire core_mi_reg_22_; 
wire core_mi_reg_23_; 
wire core_mi_reg_24_; 
wire core_mi_reg_25_; 
wire core_mi_reg_26_; 
wire core_mi_reg_27_; 
wire core_mi_reg_28_; 
wire core_mi_reg_29_; 
wire core_mi_reg_2_; 
wire core_mi_reg_30_; 
wire core_mi_reg_31_; 
wire core_mi_reg_32_; 
wire core_mi_reg_33_; 
wire core_mi_reg_34_; 
wire core_mi_reg_35_; 
wire core_mi_reg_36_; 
wire core_mi_reg_37_; 
wire core_mi_reg_38_; 
wire core_mi_reg_39_; 
wire core_mi_reg_3_; 
wire core_mi_reg_40_; 
wire core_mi_reg_41_; 
wire core_mi_reg_42_; 
wire core_mi_reg_43_; 
wire core_mi_reg_44_; 
wire core_mi_reg_45_; 
wire core_mi_reg_46_; 
wire core_mi_reg_47_; 
wire core_mi_reg_48_; 
wire core_mi_reg_49_; 
wire core_mi_reg_4_; 
wire core_mi_reg_50_; 
wire core_mi_reg_51_; 
wire core_mi_reg_52_; 
wire core_mi_reg_53_; 
wire core_mi_reg_54_; 
wire core_mi_reg_55_; 
wire core_mi_reg_56_; 
wire core_mi_reg_57_; 
wire core_mi_reg_58_; 
wire core_mi_reg_59_; 
wire core_mi_reg_5_; 
wire core_mi_reg_60_; 
wire core_mi_reg_61_; 
wire core_mi_reg_62_; 
wire core_mi_reg_63_; 
wire core_mi_reg_6_; 
wire core_mi_reg_7_; 
wire core_mi_reg_8_; 
wire core_mi_reg_9_; 
wire core_ready; 
wire core_siphash_ctrl_reg_0_; 
wire core_siphash_ctrl_reg_1_; 
wire core_siphash_ctrl_reg_2_; 
wire core_siphash_ctrl_reg_3_; 
wire core_siphash_ctrl_reg_4_; 
wire core_siphash_ctrl_reg_5_; 
wire core_siphash_ctrl_reg_6_; 
wire core_siphash_valid_reg; 
wire core_siphash_word1_we; 
wire core_siphash_word1_we_bF_buf0; 
wire core_siphash_word1_we_bF_buf1; 
wire core_siphash_word1_we_bF_buf10; 
wire core_siphash_word1_we_bF_buf2; 
wire core_siphash_word1_we_bF_buf3; 
wire core_siphash_word1_we_bF_buf4; 
wire core_siphash_word1_we_bF_buf5; 
wire core_siphash_word1_we_bF_buf6; 
wire core_siphash_word1_we_bF_buf7; 
wire core_siphash_word1_we_bF_buf8; 
wire core_siphash_word1_we_bF_buf9; 
wire core_siphash_word_0_; 
wire core_siphash_word_100_; 
wire core_siphash_word_101_; 
wire core_siphash_word_102_; 
wire core_siphash_word_103_; 
wire core_siphash_word_104_; 
wire core_siphash_word_105_; 
wire core_siphash_word_106_; 
wire core_siphash_word_107_; 
wire core_siphash_word_108_; 
wire core_siphash_word_109_; 
wire core_siphash_word_10_; 
wire core_siphash_word_110_; 
wire core_siphash_word_111_; 
wire core_siphash_word_112_; 
wire core_siphash_word_113_; 
wire core_siphash_word_114_; 
wire core_siphash_word_115_; 
wire core_siphash_word_116_; 
wire core_siphash_word_117_; 
wire core_siphash_word_118_; 
wire core_siphash_word_119_; 
wire core_siphash_word_11_; 
wire core_siphash_word_120_; 
wire core_siphash_word_121_; 
wire core_siphash_word_122_; 
wire core_siphash_word_123_; 
wire core_siphash_word_124_; 
wire core_siphash_word_125_; 
wire core_siphash_word_126_; 
wire core_siphash_word_127_; 
wire core_siphash_word_12_; 
wire core_siphash_word_13_; 
wire core_siphash_word_14_; 
wire core_siphash_word_15_; 
wire core_siphash_word_16_; 
wire core_siphash_word_17_; 
wire core_siphash_word_18_; 
wire core_siphash_word_19_; 
wire core_siphash_word_1_; 
wire core_siphash_word_20_; 
wire core_siphash_word_21_; 
wire core_siphash_word_22_; 
wire core_siphash_word_23_; 
wire core_siphash_word_24_; 
wire core_siphash_word_25_; 
wire core_siphash_word_26_; 
wire core_siphash_word_27_; 
wire core_siphash_word_28_; 
wire core_siphash_word_29_; 
wire core_siphash_word_2_; 
wire core_siphash_word_30_; 
wire core_siphash_word_31_; 
wire core_siphash_word_32_; 
wire core_siphash_word_33_; 
wire core_siphash_word_34_; 
wire core_siphash_word_35_; 
wire core_siphash_word_36_; 
wire core_siphash_word_37_; 
wire core_siphash_word_38_; 
wire core_siphash_word_39_; 
wire core_siphash_word_3_; 
wire core_siphash_word_40_; 
wire core_siphash_word_41_; 
wire core_siphash_word_42_; 
wire core_siphash_word_43_; 
wire core_siphash_word_44_; 
wire core_siphash_word_45_; 
wire core_siphash_word_46_; 
wire core_siphash_word_47_; 
wire core_siphash_word_48_; 
wire core_siphash_word_49_; 
wire core_siphash_word_4_; 
wire core_siphash_word_50_; 
wire core_siphash_word_51_; 
wire core_siphash_word_52_; 
wire core_siphash_word_53_; 
wire core_siphash_word_54_; 
wire core_siphash_word_55_; 
wire core_siphash_word_56_; 
wire core_siphash_word_57_; 
wire core_siphash_word_58_; 
wire core_siphash_word_59_; 
wire core_siphash_word_5_; 
wire core_siphash_word_60_; 
wire core_siphash_word_61_; 
wire core_siphash_word_62_; 
wire core_siphash_word_63_; 
wire core_siphash_word_64_; 
wire core_siphash_word_65_; 
wire core_siphash_word_66_; 
wire core_siphash_word_67_; 
wire core_siphash_word_68_; 
wire core_siphash_word_69_; 
wire core_siphash_word_6_; 
wire core_siphash_word_70_; 
wire core_siphash_word_71_; 
wire core_siphash_word_72_; 
wire core_siphash_word_73_; 
wire core_siphash_word_74_; 
wire core_siphash_word_75_; 
wire core_siphash_word_76_; 
wire core_siphash_word_77_; 
wire core_siphash_word_78_; 
wire core_siphash_word_79_; 
wire core_siphash_word_7_; 
wire core_siphash_word_80_; 
wire core_siphash_word_81_; 
wire core_siphash_word_82_; 
wire core_siphash_word_83_; 
wire core_siphash_word_84_; 
wire core_siphash_word_85_; 
wire core_siphash_word_86_; 
wire core_siphash_word_87_; 
wire core_siphash_word_88_; 
wire core_siphash_word_89_; 
wire core_siphash_word_8_; 
wire core_siphash_word_90_; 
wire core_siphash_word_91_; 
wire core_siphash_word_92_; 
wire core_siphash_word_93_; 
wire core_siphash_word_94_; 
wire core_siphash_word_95_; 
wire core_siphash_word_96_; 
wire core_siphash_word_97_; 
wire core_siphash_word_98_; 
wire core_siphash_word_99_; 
wire core_siphash_word_9_; 
wire core_v0_reg_0_; 
wire core_v0_reg_10_; 
wire core_v0_reg_11_; 
wire core_v0_reg_12_; 
wire core_v0_reg_13_; 
wire core_v0_reg_14_; 
wire core_v0_reg_15_; 
wire core_v0_reg_16_; 
wire core_v0_reg_17_; 
wire core_v0_reg_18_; 
wire core_v0_reg_19_; 
wire core_v0_reg_1_; 
wire core_v0_reg_20_; 
wire core_v0_reg_21_; 
wire core_v0_reg_22_; 
wire core_v0_reg_23_; 
wire core_v0_reg_24_; 
wire core_v0_reg_25_; 
wire core_v0_reg_26_; 
wire core_v0_reg_27_; 
wire core_v0_reg_28_; 
wire core_v0_reg_29_; 
wire core_v0_reg_2_; 
wire core_v0_reg_30_; 
wire core_v0_reg_31_; 
wire core_v0_reg_32_; 
wire core_v0_reg_33_; 
wire core_v0_reg_34_; 
wire core_v0_reg_35_; 
wire core_v0_reg_36_; 
wire core_v0_reg_37_; 
wire core_v0_reg_38_; 
wire core_v0_reg_39_; 
wire core_v0_reg_3_; 
wire core_v0_reg_40_; 
wire core_v0_reg_41_; 
wire core_v0_reg_42_; 
wire core_v0_reg_43_; 
wire core_v0_reg_44_; 
wire core_v0_reg_45_; 
wire core_v0_reg_46_; 
wire core_v0_reg_47_; 
wire core_v0_reg_48_; 
wire core_v0_reg_49_; 
wire core_v0_reg_4_; 
wire core_v0_reg_50_; 
wire core_v0_reg_51_; 
wire core_v0_reg_52_; 
wire core_v0_reg_53_; 
wire core_v0_reg_54_; 
wire core_v0_reg_55_; 
wire core_v0_reg_56_; 
wire core_v0_reg_57_; 
wire core_v0_reg_58_; 
wire core_v0_reg_59_; 
wire core_v0_reg_5_; 
wire core_v0_reg_60_; 
wire core_v0_reg_61_; 
wire core_v0_reg_62_; 
wire core_v0_reg_63_; 
wire core_v0_reg_6_; 
wire core_v0_reg_7_; 
wire core_v0_reg_8_; 
wire core_v0_reg_9_; 
wire core_v1_reg_0_; 
wire core_v1_reg_10_; 
wire core_v1_reg_11_; 
wire core_v1_reg_12_; 
wire core_v1_reg_13_; 
wire core_v1_reg_14_; 
wire core_v1_reg_15_; 
wire core_v1_reg_16_; 
wire core_v1_reg_17_; 
wire core_v1_reg_18_; 
wire core_v1_reg_19_; 
wire core_v1_reg_1_; 
wire core_v1_reg_20_; 
wire core_v1_reg_21_; 
wire core_v1_reg_22_; 
wire core_v1_reg_23_; 
wire core_v1_reg_24_; 
wire core_v1_reg_25_; 
wire core_v1_reg_26_; 
wire core_v1_reg_27_; 
wire core_v1_reg_28_; 
wire core_v1_reg_29_; 
wire core_v1_reg_2_; 
wire core_v1_reg_30_; 
wire core_v1_reg_31_; 
wire core_v1_reg_32_; 
wire core_v1_reg_33_; 
wire core_v1_reg_34_; 
wire core_v1_reg_35_; 
wire core_v1_reg_36_; 
wire core_v1_reg_37_; 
wire core_v1_reg_38_; 
wire core_v1_reg_39_; 
wire core_v1_reg_3_; 
wire core_v1_reg_40_; 
wire core_v1_reg_41_; 
wire core_v1_reg_42_; 
wire core_v1_reg_43_; 
wire core_v1_reg_44_; 
wire core_v1_reg_45_; 
wire core_v1_reg_46_; 
wire core_v1_reg_47_; 
wire core_v1_reg_48_; 
wire core_v1_reg_49_; 
wire core_v1_reg_4_; 
wire core_v1_reg_50_; 
wire core_v1_reg_51_; 
wire core_v1_reg_52_; 
wire core_v1_reg_53_; 
wire core_v1_reg_54_; 
wire core_v1_reg_55_; 
wire core_v1_reg_56_; 
wire core_v1_reg_57_; 
wire core_v1_reg_58_; 
wire core_v1_reg_59_; 
wire core_v1_reg_5_; 
wire core_v1_reg_60_; 
wire core_v1_reg_61_; 
wire core_v1_reg_62_; 
wire core_v1_reg_63_; 
wire core_v1_reg_6_; 
wire core_v1_reg_7_; 
wire core_v1_reg_8_; 
wire core_v1_reg_9_; 
wire core_v2_reg_0_; 
wire core_v2_reg_10_; 
wire core_v2_reg_11_; 
wire core_v2_reg_12_; 
wire core_v2_reg_13_; 
wire core_v2_reg_14_; 
wire core_v2_reg_15_; 
wire core_v2_reg_16_; 
wire core_v2_reg_17_; 
wire core_v2_reg_18_; 
wire core_v2_reg_19_; 
wire core_v2_reg_1_; 
wire core_v2_reg_20_; 
wire core_v2_reg_21_; 
wire core_v2_reg_22_; 
wire core_v2_reg_23_; 
wire core_v2_reg_24_; 
wire core_v2_reg_25_; 
wire core_v2_reg_26_; 
wire core_v2_reg_27_; 
wire core_v2_reg_28_; 
wire core_v2_reg_29_; 
wire core_v2_reg_2_; 
wire core_v2_reg_30_; 
wire core_v2_reg_31_; 
wire core_v2_reg_32_; 
wire core_v2_reg_33_; 
wire core_v2_reg_34_; 
wire core_v2_reg_35_; 
wire core_v2_reg_36_; 
wire core_v2_reg_37_; 
wire core_v2_reg_38_; 
wire core_v2_reg_39_; 
wire core_v2_reg_3_; 
wire core_v2_reg_40_; 
wire core_v2_reg_41_; 
wire core_v2_reg_42_; 
wire core_v2_reg_43_; 
wire core_v2_reg_44_; 
wire core_v2_reg_45_; 
wire core_v2_reg_46_; 
wire core_v2_reg_47_; 
wire core_v2_reg_48_; 
wire core_v2_reg_49_; 
wire core_v2_reg_4_; 
wire core_v2_reg_50_; 
wire core_v2_reg_51_; 
wire core_v2_reg_52_; 
wire core_v2_reg_53_; 
wire core_v2_reg_54_; 
wire core_v2_reg_55_; 
wire core_v2_reg_56_; 
wire core_v2_reg_57_; 
wire core_v2_reg_58_; 
wire core_v2_reg_59_; 
wire core_v2_reg_5_; 
wire core_v2_reg_60_; 
wire core_v2_reg_61_; 
wire core_v2_reg_62_; 
wire core_v2_reg_63_; 
wire core_v2_reg_6_; 
wire core_v2_reg_7_; 
wire core_v2_reg_8_; 
wire core_v2_reg_9_; 
wire core_v3_reg_0_; 
wire core_v3_reg_10_; 
wire core_v3_reg_11_; 
wire core_v3_reg_12_; 
wire core_v3_reg_13_; 
wire core_v3_reg_14_; 
wire core_v3_reg_15_; 
wire core_v3_reg_16_; 
wire core_v3_reg_17_; 
wire core_v3_reg_18_; 
wire core_v3_reg_19_; 
wire core_v3_reg_1_; 
wire core_v3_reg_20_; 
wire core_v3_reg_21_; 
wire core_v3_reg_22_; 
wire core_v3_reg_23_; 
wire core_v3_reg_24_; 
wire core_v3_reg_25_; 
wire core_v3_reg_26_; 
wire core_v3_reg_27_; 
wire core_v3_reg_28_; 
wire core_v3_reg_29_; 
wire core_v3_reg_2_; 
wire core_v3_reg_30_; 
wire core_v3_reg_31_; 
wire core_v3_reg_32_; 
wire core_v3_reg_33_; 
wire core_v3_reg_34_; 
wire core_v3_reg_35_; 
wire core_v3_reg_36_; 
wire core_v3_reg_37_; 
wire core_v3_reg_38_; 
wire core_v3_reg_39_; 
wire core_v3_reg_3_; 
wire core_v3_reg_40_; 
wire core_v3_reg_41_; 
wire core_v3_reg_42_; 
wire core_v3_reg_43_; 
wire core_v3_reg_44_; 
wire core_v3_reg_45_; 
wire core_v3_reg_46_; 
wire core_v3_reg_47_; 
wire core_v3_reg_48_; 
wire core_v3_reg_49_; 
wire core_v3_reg_4_; 
wire core_v3_reg_50_; 
wire core_v3_reg_51_; 
wire core_v3_reg_52_; 
wire core_v3_reg_53_; 
wire core_v3_reg_54_; 
wire core_v3_reg_55_; 
wire core_v3_reg_56_; 
wire core_v3_reg_57_; 
wire core_v3_reg_58_; 
wire core_v3_reg_59_; 
wire core_v3_reg_5_; 
wire core_v3_reg_60_; 
wire core_v3_reg_61_; 
wire core_v3_reg_62_; 
wire core_v3_reg_63_; 
wire core_v3_reg_6_; 
wire core_v3_reg_7_; 
wire core_v3_reg_8_; 
wire core_v3_reg_9_; 
input cs;
output \read_data[0] ;
output \read_data[10] ;
output \read_data[11] ;
output \read_data[12] ;
output \read_data[13] ;
output \read_data[14] ;
output \read_data[15] ;
output \read_data[16] ;
output \read_data[17] ;
output \read_data[18] ;
output \read_data[19] ;
output \read_data[1] ;
output \read_data[20] ;
output \read_data[21] ;
output \read_data[22] ;
output \read_data[23] ;
output \read_data[24] ;
output \read_data[25] ;
output \read_data[26] ;
output \read_data[27] ;
output \read_data[28] ;
output \read_data[29] ;
output \read_data[2] ;
output \read_data[30] ;
output \read_data[31] ;
output \read_data[3] ;
output \read_data[4] ;
output \read_data[5] ;
output \read_data[6] ;
output \read_data[7] ;
output \read_data[8] ;
output \read_data[9] ;
input reset_n;
wire reset_n_bF_buf0; 
wire reset_n_bF_buf1; 
wire reset_n_bF_buf10; 
wire reset_n_bF_buf11; 
wire reset_n_bF_buf12; 
wire reset_n_bF_buf13; 
wire reset_n_bF_buf14; 
wire reset_n_bF_buf15; 
wire reset_n_bF_buf16; 
wire reset_n_bF_buf17; 
wire reset_n_bF_buf18; 
wire reset_n_bF_buf19; 
wire reset_n_bF_buf2; 
wire reset_n_bF_buf20; 
wire reset_n_bF_buf21; 
wire reset_n_bF_buf22; 
wire reset_n_bF_buf23; 
wire reset_n_bF_buf24; 
wire reset_n_bF_buf25; 
wire reset_n_bF_buf26; 
wire reset_n_bF_buf27; 
wire reset_n_bF_buf28; 
wire reset_n_bF_buf29; 
wire reset_n_bF_buf3; 
wire reset_n_bF_buf30; 
wire reset_n_bF_buf31; 
wire reset_n_bF_buf32; 
wire reset_n_bF_buf33; 
wire reset_n_bF_buf34; 
wire reset_n_bF_buf35; 
wire reset_n_bF_buf36; 
wire reset_n_bF_buf37; 
wire reset_n_bF_buf38; 
wire reset_n_bF_buf39; 
wire reset_n_bF_buf4; 
wire reset_n_bF_buf40; 
wire reset_n_bF_buf41; 
wire reset_n_bF_buf42; 
wire reset_n_bF_buf43; 
wire reset_n_bF_buf44; 
wire reset_n_bF_buf45; 
wire reset_n_bF_buf46; 
wire reset_n_bF_buf47; 
wire reset_n_bF_buf48; 
wire reset_n_bF_buf49; 
wire reset_n_bF_buf5; 
wire reset_n_bF_buf50; 
wire reset_n_bF_buf51; 
wire reset_n_bF_buf52; 
wire reset_n_bF_buf53; 
wire reset_n_bF_buf54; 
wire reset_n_bF_buf55; 
wire reset_n_bF_buf56; 
wire reset_n_bF_buf57; 
wire reset_n_bF_buf58; 
wire reset_n_bF_buf59; 
wire reset_n_bF_buf6; 
wire reset_n_bF_buf60; 
wire reset_n_bF_buf61; 
wire reset_n_bF_buf62; 
wire reset_n_bF_buf63; 
wire reset_n_bF_buf64; 
wire reset_n_bF_buf65; 
wire reset_n_bF_buf66; 
wire reset_n_bF_buf67; 
wire reset_n_bF_buf68; 
wire reset_n_bF_buf69; 
wire reset_n_bF_buf7; 
wire reset_n_bF_buf8; 
wire reset_n_bF_buf9; 
wire reset_n_hier0_bF_buf0; 
wire reset_n_hier0_bF_buf1; 
wire reset_n_hier0_bF_buf2; 
wire reset_n_hier0_bF_buf3; 
wire reset_n_hier0_bF_buf4; 
wire reset_n_hier0_bF_buf5; 
wire reset_n_hier0_bF_buf6; 
wire reset_n_hier0_bF_buf7; 
input we;
wire word0_reg_0_; 
wire word0_reg_10_; 
wire word0_reg_11_; 
wire word0_reg_12_; 
wire word0_reg_13_; 
wire word0_reg_14_; 
wire word0_reg_15_; 
wire word0_reg_16_; 
wire word0_reg_17_; 
wire word0_reg_18_; 
wire word0_reg_19_; 
wire word0_reg_1_; 
wire word0_reg_20_; 
wire word0_reg_21_; 
wire word0_reg_22_; 
wire word0_reg_23_; 
wire word0_reg_24_; 
wire word0_reg_25_; 
wire word0_reg_26_; 
wire word0_reg_27_; 
wire word0_reg_28_; 
wire word0_reg_29_; 
wire word0_reg_2_; 
wire word0_reg_30_; 
wire word0_reg_31_; 
wire word0_reg_3_; 
wire word0_reg_4_; 
wire word0_reg_5_; 
wire word0_reg_6_; 
wire word0_reg_7_; 
wire word0_reg_8_; 
wire word0_reg_9_; 
wire word1_reg_0_; 
wire word1_reg_10_; 
wire word1_reg_11_; 
wire word1_reg_12_; 
wire word1_reg_13_; 
wire word1_reg_14_; 
wire word1_reg_15_; 
wire word1_reg_16_; 
wire word1_reg_17_; 
wire word1_reg_18_; 
wire word1_reg_19_; 
wire word1_reg_1_; 
wire word1_reg_20_; 
wire word1_reg_21_; 
wire word1_reg_22_; 
wire word1_reg_23_; 
wire word1_reg_24_; 
wire word1_reg_25_; 
wire word1_reg_26_; 
wire word1_reg_27_; 
wire word1_reg_28_; 
wire word1_reg_29_; 
wire word1_reg_2_; 
wire word1_reg_30_; 
wire word1_reg_31_; 
wire word1_reg_3_; 
wire word1_reg_4_; 
wire word1_reg_5_; 
wire word1_reg_6_; 
wire word1_reg_7_; 
wire word1_reg_8_; 
wire word1_reg_9_; 
wire word2_reg_0_; 
wire word2_reg_10_; 
wire word2_reg_11_; 
wire word2_reg_12_; 
wire word2_reg_13_; 
wire word2_reg_14_; 
wire word2_reg_15_; 
wire word2_reg_16_; 
wire word2_reg_17_; 
wire word2_reg_18_; 
wire word2_reg_19_; 
wire word2_reg_1_; 
wire word2_reg_20_; 
wire word2_reg_21_; 
wire word2_reg_22_; 
wire word2_reg_23_; 
wire word2_reg_24_; 
wire word2_reg_25_; 
wire word2_reg_26_; 
wire word2_reg_27_; 
wire word2_reg_28_; 
wire word2_reg_29_; 
wire word2_reg_2_; 
wire word2_reg_30_; 
wire word2_reg_31_; 
wire word2_reg_3_; 
wire word2_reg_4_; 
wire word2_reg_5_; 
wire word2_reg_6_; 
wire word2_reg_7_; 
wire word2_reg_8_; 
wire word2_reg_9_; 
wire word3_reg_0_; 
wire word3_reg_10_; 
wire word3_reg_11_; 
wire word3_reg_12_; 
wire word3_reg_13_; 
wire word3_reg_14_; 
wire word3_reg_15_; 
wire word3_reg_16_; 
wire word3_reg_17_; 
wire word3_reg_18_; 
wire word3_reg_19_; 
wire word3_reg_1_; 
wire word3_reg_20_; 
wire word3_reg_21_; 
wire word3_reg_22_; 
wire word3_reg_23_; 
wire word3_reg_24_; 
wire word3_reg_25_; 
wire word3_reg_26_; 
wire word3_reg_27_; 
wire word3_reg_28_; 
wire word3_reg_29_; 
wire word3_reg_2_; 
wire word3_reg_30_; 
wire word3_reg_31_; 
wire word3_reg_3_; 
wire word3_reg_4_; 
wire word3_reg_5_; 
wire word3_reg_6_; 
wire word3_reg_7_; 
wire word3_reg_8_; 
wire word3_reg_9_; 
input \write_data[0] ;
input \write_data[10] ;
input \write_data[11] ;
input \write_data[12] ;
input \write_data[13] ;
input \write_data[14] ;
input \write_data[15] ;
input \write_data[16] ;
input \write_data[17] ;
input \write_data[18] ;
input \write_data[19] ;
input \write_data[1] ;
input \write_data[20] ;
input \write_data[21] ;
input \write_data[22] ;
input \write_data[23] ;
input \write_data[24] ;
input \write_data[25] ;
input \write_data[26] ;
input \write_data[27] ;
input \write_data[28] ;
input \write_data[29] ;
input \write_data[2] ;
input \write_data[30] ;
input \write_data[31] ;
input \write_data[3] ;
input \write_data[4] ;
input \write_data[5] ;
input \write_data[6] ;
input \write_data[7] ;
input \write_data[8] ;
input \write_data[9] ;
AND2X2 AND2X2_1 ( .A(_abc_19873_new_n875_), .B(_abc_19873_new_n876_), .Y(_abc_19873_new_n877_));
AND2X2 AND2X2_10 ( .A(core_v1_reg_9_), .B(core_v0_reg_9_), .Y(core__abc_21302_new_n1302_));
AND2X2 AND2X2_100 ( .A(core__abc_21302_new_n3296_), .B(core__abc_21302_new_n1751_), .Y(core__abc_21302_new_n3297_));
AND2X2 AND2X2_101 ( .A(core__abc_21302_new_n2639__bF_buf6), .B(core_key_81_), .Y(core__abc_21302_new_n3328_));
AND2X2 AND2X2_102 ( .A(core__abc_21302_new_n3353_), .B(core__abc_21302_new_n1905_), .Y(core__abc_21302_new_n3354_));
AND2X2 AND2X2_103 ( .A(core__abc_21302_new_n3382_), .B(core__abc_21302_new_n3377_), .Y(core__abc_21302_new_n3391_));
AND2X2 AND2X2_104 ( .A(core__abc_21302_new_n3389_), .B(core__abc_21302_new_n3393_), .Y(core__abc_21302_new_n3394_));
AND2X2 AND2X2_105 ( .A(core__abc_21302_new_n3420_), .B(core__abc_21302_new_n1424_), .Y(core__abc_21302_new_n3426_));
AND2X2 AND2X2_106 ( .A(core__abc_21302_new_n3427_), .B(core__abc_21302_new_n3423_), .Y(core__abc_21302_new_n3432_));
AND2X2 AND2X2_107 ( .A(core__abc_21302_new_n3353_), .B(core__abc_21302_new_n3441_), .Y(core__abc_21302_new_n3442_));
AND2X2 AND2X2_108 ( .A(core__abc_21302_new_n3541_), .B(core__abc_21302_new_n3538_), .Y(core__abc_21302_new_n3544_));
AND2X2 AND2X2_109 ( .A(core__abc_21302_new_n3549_), .B(core__abc_21302_new_n2575_), .Y(core__abc_21302_new_n3550_));
AND2X2 AND2X2_11 ( .A(core_v1_reg_10_), .B(core_v0_reg_10_), .Y(core__abc_21302_new_n1313_));
AND2X2 AND2X2_110 ( .A(core__abc_21302_new_n3552_), .B(core__abc_21302_new_n3555_), .Y(core__abc_21302_new_n3556_));
AND2X2 AND2X2_111 ( .A(core__abc_21302_new_n3557_), .B(core__abc_21302_new_n3561_), .Y(core__abc_21302_new_n3562_));
AND2X2 AND2X2_112 ( .A(core__abc_21302_new_n3536_), .B(core__abc_21302_new_n3562_), .Y(core__abc_21302_new_n3563_));
AND2X2 AND2X2_113 ( .A(core__abc_21302_new_n2639__bF_buf5), .B(core_key_87_), .Y(core__abc_21302_new_n3598_));
AND2X2 AND2X2_114 ( .A(core__abc_21302_new_n2548_), .B(core__abc_21302_new_n3633_), .Y(core__abc_21302_new_n3634_));
AND2X2 AND2X2_115 ( .A(core__abc_21302_new_n3646_), .B(core__abc_21302_new_n2745_), .Y(core__abc_21302_new_n3647_));
AND2X2 AND2X2_116 ( .A(core__abc_21302_new_n3658_), .B(core__abc_21302_new_n3659_), .Y(core__abc_21302_new_n3674_));
AND2X2 AND2X2_117 ( .A(core__abc_21302_new_n3704_), .B(core__abc_21302_new_n2551_), .Y(core__abc_21302_new_n3706_));
AND2X2 AND2X2_118 ( .A(core__abc_21302_new_n3709_), .B(core__abc_21302_new_n3707_), .Y(core__abc_21302_new_n3710_));
AND2X2 AND2X2_119 ( .A(core__abc_21302_new_n3717_), .B(core__abc_21302_new_n2807_), .Y(core__abc_21302_new_n3718_));
AND2X2 AND2X2_12 ( .A(core_v1_reg_11_), .B(core_v0_reg_11_), .Y(core__abc_21302_new_n1325_));
AND2X2 AND2X2_120 ( .A(core__abc_21302_new_n3725_), .B(core__abc_21302_new_n3710_), .Y(core__abc_21302_new_n3726_));
AND2X2 AND2X2_121 ( .A(core__abc_21302_new_n3738_), .B(core__abc_21302_new_n3741_), .Y(core__abc_21302_new_n3742_));
AND2X2 AND2X2_122 ( .A(core__abc_21302_new_n3747_), .B(core__abc_21302_new_n3743_), .Y(core__abc_21302_new_n3748_));
AND2X2 AND2X2_123 ( .A(core__abc_21302_new_n1874_), .B(core__abc_21302_new_n1887_), .Y(core__abc_21302_new_n3769_));
AND2X2 AND2X2_124 ( .A(core__abc_21302_new_n3767_), .B(core__abc_21302_new_n3779_), .Y(core__abc_21302_new_n3780_));
AND2X2 AND2X2_125 ( .A(core__abc_21302_new_n3821_), .B(core__abc_21302_new_n2940_), .Y(core__abc_21302_new_n3822_));
AND2X2 AND2X2_126 ( .A(core__abc_21302_new_n3833_), .B(core__abc_21302_new_n3831_), .Y(core__abc_21302_new_n3835_));
AND2X2 AND2X2_127 ( .A(core__abc_21302_new_n3837_), .B(core__abc_21302_new_n1551_), .Y(core__abc_21302_new_n3839_));
AND2X2 AND2X2_128 ( .A(core__abc_21302_new_n3840_), .B(core__abc_21302_new_n3847_), .Y(core__abc_21302_new_n3848_));
AND2X2 AND2X2_129 ( .A(core__abc_21302_new_n3815_), .B(core__abc_21302_new_n3812_), .Y(core__abc_21302_new_n3860_));
AND2X2 AND2X2_13 ( .A(core__abc_21302_new_n1340_), .B(core__abc_21302_new_n1337_), .Y(core__abc_21302_new_n1341_));
AND2X2 AND2X2_130 ( .A(core__abc_21302_new_n3849_), .B(core__abc_21302_new_n3853_), .Y(core__abc_21302_new_n3866_));
AND2X2 AND2X2_131 ( .A(core__abc_21302_new_n3869_), .B(core__abc_21302_new_n2971_), .Y(core__abc_21302_new_n3870_));
AND2X2 AND2X2_132 ( .A(core__abc_21302_new_n3886_), .B(core__abc_21302_new_n3889_), .Y(core__abc_21302_new_n3890_));
AND2X2 AND2X2_133 ( .A(core__abc_21302_new_n2639__bF_buf4), .B(core_key_95_), .Y(core__abc_21302_new_n3902_));
AND2X2 AND2X2_134 ( .A(core__abc_21302_new_n3926_), .B(core__abc_21302_new_n1211_), .Y(core__abc_21302_new_n3927_));
AND2X2 AND2X2_135 ( .A(core__abc_21302_new_n3924_), .B(core__abc_21302_new_n1568_), .Y(core__abc_21302_new_n3950_));
AND2X2 AND2X2_136 ( .A(core__abc_21302_new_n3951_), .B(core__abc_21302_new_n3953_), .Y(core__abc_21302_new_n3956_));
AND2X2 AND2X2_137 ( .A(core__abc_21302_new_n2639__bF_buf3), .B(core_key_98_), .Y(core__abc_21302_new_n3970_));
AND2X2 AND2X2_138 ( .A(core__abc_21302_new_n3990_), .B(core__abc_21302_new_n3993_), .Y(core__abc_21302_new_n3994_));
AND2X2 AND2X2_139 ( .A(core__abc_21302_new_n2639__bF_buf2), .B(core_key_100_), .Y(core__abc_21302_new_n4031_));
AND2X2 AND2X2_14 ( .A(core_v1_reg_13_), .B(core_v0_reg_13_), .Y(core__abc_21302_new_n1347_));
AND2X2 AND2X2_140 ( .A(core__abc_21302_new_n2639__bF_buf0), .B(core_key_104_), .Y(core__abc_21302_new_n4154_));
AND2X2 AND2X2_141 ( .A(core__abc_21302_new_n4177_), .B(core__abc_21302_new_n4178_), .Y(core__abc_21302_new_n4179_));
AND2X2 AND2X2_142 ( .A(core__abc_21302_new_n4222_), .B(core__abc_21302_new_n4221_), .Y(core__abc_21302_new_n4223_));
AND2X2 AND2X2_143 ( .A(core__abc_21302_new_n4227_), .B(core__abc_21302_new_n4230_), .Y(core__abc_21302_new_n4231_));
AND2X2 AND2X2_144 ( .A(core__abc_21302_new_n4284_), .B(core__abc_21302_new_n2482_), .Y(core__abc_21302_new_n4333_));
AND2X2 AND2X2_145 ( .A(core__abc_21302_new_n4386_), .B(core__abc_21302_new_n4323_), .Y(core__abc_21302_new_n4387_));
AND2X2 AND2X2_146 ( .A(core__abc_21302_new_n4421_), .B(core__abc_21302_new_n4395_), .Y(core__abc_21302_new_n4422_));
AND2X2 AND2X2_147 ( .A(core__abc_21302_new_n2420_), .B(core__abc_21302_new_n2431_), .Y(core__abc_21302_new_n4445_));
AND2X2 AND2X2_148 ( .A(core__abc_21302_new_n4451_), .B(core__abc_21302_new_n4452_), .Y(core__abc_21302_new_n4453_));
AND2X2 AND2X2_149 ( .A(core__abc_21302_new_n4476_), .B(core__abc_21302_new_n4477_), .Y(core__abc_21302_new_n4478_));
AND2X2 AND2X2_15 ( .A(core__abc_21302_new_n1352_), .B(core__abc_21302_new_n1349_), .Y(core__abc_21302_new_n1353_));
AND2X2 AND2X2_150 ( .A(core__abc_21302_new_n2639__bF_buf5), .B(core_key_116_), .Y(core__abc_21302_new_n4492_));
AND2X2 AND2X2_151 ( .A(core__abc_21302_new_n2639__bF_buf3), .B(core_key_120_), .Y(core__abc_21302_new_n4593_));
AND2X2 AND2X2_152 ( .A(core__abc_21302_new_n4653_), .B(core__abc_21302_new_n4656_), .Y(core__abc_21302_new_n4657_));
AND2X2 AND2X2_153 ( .A(core__abc_21302_new_n4650_), .B(core__abc_21302_new_n1497_), .Y(core__abc_21302_new_n4676_));
AND2X2 AND2X2_154 ( .A(core__abc_21302_new_n4598_), .B(core__abc_21302_new_n4601_), .Y(core__abc_21302_new_n4734_));
AND2X2 AND2X2_155 ( .A(core__abc_21302_new_n4713_), .B(core__abc_21302_new_n4717_), .Y(core__abc_21302_new_n4739_));
AND2X2 AND2X2_156 ( .A(core__abc_21302_new_n4858_), .B(core__abc_21302_new_n4860_), .Y(core__abc_21302_new_n4861_));
AND2X2 AND2X2_157 ( .A(core__abc_21302_new_n4865_), .B(core__abc_21302_new_n4863_), .Y(core__abc_21302_new_n4866_));
AND2X2 AND2X2_158 ( .A(core__abc_21302_new_n4885_), .B(core__abc_21302_new_n4829_), .Y(core__abc_21302_new_n4886_));
AND2X2 AND2X2_159 ( .A(core__abc_21302_new_n4910_), .B(core__abc_21302_new_n4914_), .Y(core__abc_21302_new_n4915_));
AND2X2 AND2X2_16 ( .A(core_v1_reg_14_), .B(core_v0_reg_14_), .Y(core__abc_21302_new_n1359_));
AND2X2 AND2X2_160 ( .A(core__abc_21302_new_n4972_), .B(core__abc_21302_new_n4973_), .Y(core__abc_21302_new_n4974_));
AND2X2 AND2X2_161 ( .A(core__abc_21302_new_n4998_), .B(core__abc_21302_new_n4997_), .Y(core__abc_21302_new_n4999_));
AND2X2 AND2X2_162 ( .A(core__abc_21302_new_n4963_), .B(core__abc_21302_new_n5071_), .Y(core__abc_21302_new_n5072_));
AND2X2 AND2X2_163 ( .A(core__abc_21302_new_n5075_), .B(core__abc_21302_new_n5076_), .Y(core__abc_21302_new_n5077_));
AND2X2 AND2X2_164 ( .A(core__abc_21302_new_n5094_), .B(core__abc_21302_new_n4888_), .Y(core__abc_21302_new_n5095_));
AND2X2 AND2X2_165 ( .A(core__abc_21302_new_n5117_), .B(core__abc_21302_new_n5119_), .Y(core__abc_21302_new_n5120_));
AND2X2 AND2X2_166 ( .A(core__abc_21302_new_n5129_), .B(reset_n_bF_buf68), .Y(core__0v2_reg_63_0__2_));
AND2X2 AND2X2_167 ( .A(core__abc_21302_new_n5197_), .B(core__abc_21302_new_n5198_), .Y(core__abc_21302_new_n5199_));
AND2X2 AND2X2_168 ( .A(core__abc_21302_new_n5272_), .B(core__abc_21302_new_n5273_), .Y(core__abc_21302_new_n5274_));
AND2X2 AND2X2_169 ( .A(core__abc_21302_new_n5289_), .B(core__abc_21302_new_n5292_), .Y(core__abc_21302_new_n5293_));
AND2X2 AND2X2_17 ( .A(core__abc_21302_new_n1364_), .B(core__abc_21302_new_n1361_), .Y(core__abc_21302_new_n1365_));
AND2X2 AND2X2_170 ( .A(core__abc_21302_new_n5310_), .B(core__abc_21302_new_n5347_), .Y(core__abc_21302_new_n5348_));
AND2X2 AND2X2_171 ( .A(core__abc_21302_new_n5355_), .B(core__abc_21302_new_n5352_), .Y(core__abc_21302_new_n5356_));
AND2X2 AND2X2_172 ( .A(core__abc_21302_new_n5390_), .B(core__abc_21302_new_n5394_), .Y(core__abc_21302_new_n5415_));
AND2X2 AND2X2_173 ( .A(core__abc_21302_new_n5482_), .B(core__abc_21302_new_n5483_), .Y(core__abc_21302_new_n5484_));
AND2X2 AND2X2_174 ( .A(core__abc_21302_new_n5546_), .B(core__abc_21302_new_n5470_), .Y(core__abc_21302_new_n5547_));
AND2X2 AND2X2_175 ( .A(core__abc_21302_new_n3210_), .B(core__abc_21302_new_n5572_), .Y(core__abc_21302_new_n5573_));
AND2X2 AND2X2_176 ( .A(core__abc_21302_new_n5648_), .B(core__abc_21302_new_n5649_), .Y(core__abc_21302_new_n5652_));
AND2X2 AND2X2_177 ( .A(core__abc_21302_new_n2639__bF_buf6), .B(core_key_33_), .Y(core__abc_21302_new_n5707_));
AND2X2 AND2X2_178 ( .A(core__abc_21302_new_n5710_), .B(core__abc_21302_new_n2634__bF_buf7), .Y(core__abc_21302_new_n5711_));
AND2X2 AND2X2_179 ( .A(core__abc_21302_new_n5104__bF_buf5), .B(core__abc_21302_new_n5793_), .Y(core__abc_21302_new_n5794_));
AND2X2 AND2X2_18 ( .A(core_v1_reg_15_), .B(core_v0_reg_15_), .Y(core__abc_21302_new_n1371_));
AND2X2 AND2X2_180 ( .A(core__abc_21302_new_n2639__bF_buf2), .B(core_key_47_), .Y(core__abc_21302_new_n5827_));
AND2X2 AND2X2_181 ( .A(core__abc_21302_new_n5879_), .B(core__abc_21302_new_n5890_), .Y(core__abc_21302_new_n5891_));
AND2X2 AND2X2_182 ( .A(core__abc_21302_new_n5104__bF_buf0), .B(core__abc_21302_new_n5933_), .Y(core__abc_21302_new_n5934_));
AND2X2 AND2X2_183 ( .A(core__abc_21302_new_n5423_), .B(core__abc_21302_new_n6015_), .Y(core__abc_21302_new_n6016_));
AND2X2 AND2X2_184 ( .A(core__abc_21302_new_n6054_), .B(core__abc_21302_new_n6055_), .Y(core__abc_21302_new_n6056_));
AND2X2 AND2X2_185 ( .A(core__abc_21302_new_n5783_), .B(core__abc_21302_new_n5572_), .Y(core__abc_21302_new_n6075_));
AND2X2 AND2X2_186 ( .A(core__abc_21302_new_n5804_), .B(core__abc_21302_new_n5603_), .Y(core__abc_21302_new_n6088_));
AND2X2 AND2X2_187 ( .A(core__abc_21302_new_n5842_), .B(core__abc_21302_new_n5687_), .Y(core__abc_21302_new_n6113_));
AND2X2 AND2X2_188 ( .A(core__abc_21302_new_n5903_), .B(core__abc_21302_new_n5030_), .Y(core__abc_21302_new_n6153_));
AND2X2 AND2X2_189 ( .A(core__abc_21302_new_n5938_), .B(core__abc_21302_new_n5010_), .Y(core__abc_21302_new_n6181_));
AND2X2 AND2X2_19 ( .A(core_v1_reg_16_), .B(core_v0_reg_16_), .Y(core__abc_21302_new_n1383_));
AND2X2 AND2X2_190 ( .A(core__abc_21302_new_n5242_), .B(core__abc_21302_new_n6274_), .Y(core__abc_21302_new_n6275_));
AND2X2 AND2X2_191 ( .A(core__abc_21302_new_n5485_), .B(core__abc_21302_new_n5155_), .Y(core__abc_21302_new_n6359_));
AND2X2 AND2X2_192 ( .A(core__abc_21302_new_n2658_), .B(core__abc_21302_new_n2634__bF_buf6), .Y(core__abc_21302_new_n6457_));
AND2X2 AND2X2_193 ( .A(core__abc_21302_new_n2947_), .B(core__abc_21302_new_n2634__bF_buf4), .Y(core__abc_21302_new_n6506_));
AND2X2 AND2X2_194 ( .A(core__abc_21302_new_n3025_), .B(core__abc_21302_new_n2634__bF_buf3), .Y(core__abc_21302_new_n6521_));
AND2X2 AND2X2_195 ( .A(core__abc_21302_new_n3062_), .B(core__abc_21302_new_n2634__bF_buf2), .Y(core__abc_21302_new_n6528_));
AND2X2 AND2X2_196 ( .A(core__abc_21302_new_n3110_), .B(core__abc_21302_new_n2634__bF_buf1), .Y(core__abc_21302_new_n6535_));
AND2X2 AND2X2_197 ( .A(core__abc_21302_new_n3154_), .B(core__abc_21302_new_n2634__bF_buf0), .Y(core__abc_21302_new_n6543_));
AND2X2 AND2X2_198 ( .A(core__abc_21302_new_n3310_), .B(core__abc_21302_new_n2634__bF_buf8), .Y(core__abc_21302_new_n6564_));
AND2X2 AND2X2_199 ( .A(core__abc_21302_new_n3565_), .B(core__abc_21302_new_n2634__bF_buf7), .Y(core__abc_21302_new_n6607_));
AND2X2 AND2X2_2 ( .A(_abc_19873_new_n903_), .B(_abc_19873_new_n904_), .Y(_abc_19873_new_n905_));
AND2X2 AND2X2_20 ( .A(core_v1_reg_17_), .B(core_v0_reg_17_), .Y(core__abc_21302_new_n1394_));
AND2X2 AND2X2_200 ( .A(core__abc_21302_new_n6449__bF_buf6), .B(core__abc_21302_new_n6621_), .Y(core__abc_21302_new_n6622_));
AND2X2 AND2X2_201 ( .A(core__abc_21302_new_n3717_), .B(core__abc_21302_new_n2634__bF_buf6), .Y(core__abc_21302_new_n6636_));
AND2X2 AND2X2_202 ( .A(core__abc_21302_new_n3782_), .B(core__abc_21302_new_n2634__bF_buf5), .Y(core__abc_21302_new_n6652_));
AND2X2 AND2X2_203 ( .A(core__abc_21302_new_n3869_), .B(core__abc_21302_new_n2634__bF_buf4), .Y(core__abc_21302_new_n6666_));
AND2X2 AND2X2_204 ( .A(core__abc_21302_new_n3995_), .B(core__abc_21302_new_n2634__bF_buf3), .Y(core__abc_21302_new_n6692_));
AND2X2 AND2X2_205 ( .A(core__abc_21302_new_n4056_), .B(core__abc_21302_new_n2634__bF_buf2), .Y(core__abc_21302_new_n6706_));
AND2X2 AND2X2_206 ( .A(core__abc_21302_new_n6449__bF_buf6), .B(core__abc_21302_new_n6733_), .Y(core__abc_21302_new_n6734_));
AND2X2 AND2X2_207 ( .A(core__abc_21302_new_n4241_), .B(core__abc_21302_new_n2634__bF_buf1), .Y(core__abc_21302_new_n6747_));
AND2X2 AND2X2_208 ( .A(core__abc_21302_new_n4291_), .B(core__abc_21302_new_n2634__bF_buf0), .Y(core__abc_21302_new_n6761_));
AND2X2 AND2X2_209 ( .A(core__abc_21302_new_n6449__bF_buf6), .B(core__abc_21302_new_n6789_), .Y(core__abc_21302_new_n6790_));
AND2X2 AND2X2_21 ( .A(core_v1_reg_18_), .B(core_v0_reg_18_), .Y(core__abc_21302_new_n1406_));
AND2X2 AND2X2_210 ( .A(core__abc_21302_new_n4508_), .B(core__abc_21302_new_n2634__bF_buf8), .Y(core__abc_21302_new_n6816_));
AND2X2 AND2X2_211 ( .A(core__abc_21302_new_n4556_), .B(core__abc_21302_new_n2634__bF_buf7), .Y(core__abc_21302_new_n6831_));
AND2X2 AND2X2_212 ( .A(core__abc_21302_new_n4610_), .B(core__abc_21302_new_n2634__bF_buf6), .Y(core__abc_21302_new_n6845_));
AND2X2 AND2X2_213 ( .A(core__abc_21302_new_n4723_), .B(core__abc_21302_new_n2634__bF_buf5), .Y(core__abc_21302_new_n6876_));
AND2X2 AND2X2_22 ( .A(core_v1_reg_19_), .B(core_v0_reg_19_), .Y(core__abc_21302_new_n1418_));
AND2X2 AND2X2_23 ( .A(core_v1_reg_20_), .B(core_v0_reg_20_), .Y(core__abc_21302_new_n1430_));
AND2X2 AND2X2_24 ( .A(core_v1_reg_21_), .B(core_v0_reg_21_), .Y(core__abc_21302_new_n1442_));
AND2X2 AND2X2_25 ( .A(core_v1_reg_22_), .B(core_v0_reg_22_), .Y(core__abc_21302_new_n1454_));
AND2X2 AND2X2_26 ( .A(core_v1_reg_23_), .B(core_v0_reg_23_), .Y(core__abc_21302_new_n1466_));
AND2X2 AND2X2_27 ( .A(core_v1_reg_24_), .B(core_v0_reg_24_), .Y(core__abc_21302_new_n1474_));
AND2X2 AND2X2_28 ( .A(core__abc_21302_new_n1489_), .B(core__abc_21302_new_n1486_), .Y(core__abc_21302_new_n1490_));
AND2X2 AND2X2_29 ( .A(core_v1_reg_26_), .B(core_v0_reg_26_), .Y(core__abc_21302_new_n1496_));
AND2X2 AND2X2_3 ( .A(core_v1_reg_2_), .B(core_v0_reg_2_), .Y(core__abc_21302_new_n1232_));
AND2X2 AND2X2_30 ( .A(core_v1_reg_27_), .B(core_v0_reg_27_), .Y(core__abc_21302_new_n1508_));
AND2X2 AND2X2_31 ( .A(core_v1_reg_28_), .B(core_v0_reg_28_), .Y(core__abc_21302_new_n1520_));
AND2X2 AND2X2_32 ( .A(core_v1_reg_30_), .B(core_v0_reg_30_), .Y(core__abc_21302_new_n1545_));
AND2X2 AND2X2_33 ( .A(core_v1_reg_31_), .B(core_v0_reg_31_), .Y(core__abc_21302_new_n1557_));
AND2X2 AND2X2_34 ( .A(core_v1_reg_35_), .B(core_v0_reg_35_), .Y(core__abc_21302_new_n1603_));
AND2X2 AND2X2_35 ( .A(core_v1_reg_36_), .B(core_v0_reg_36_), .Y(core__abc_21302_new_n1615_));
AND2X2 AND2X2_36 ( .A(core_v1_reg_39_), .B(core_v0_reg_39_), .Y(core__abc_21302_new_n1648_));
AND2X2 AND2X2_37 ( .A(core_v1_reg_40_), .B(core_v0_reg_40_), .Y(core__abc_21302_new_n1659_));
AND2X2 AND2X2_38 ( .A(core_v1_reg_41_), .B(core_v0_reg_41_), .Y(core__abc_21302_new_n1670_));
AND2X2 AND2X2_39 ( .A(core_v1_reg_42_), .B(core_v0_reg_42_), .Y(core__abc_21302_new_n1681_));
AND2X2 AND2X2_4 ( .A(core_v2_reg_2_), .B(core_v3_reg_2_), .Y(core__abc_21302_new_n1235_));
AND2X2 AND2X2_40 ( .A(core_v1_reg_43_), .B(core_v0_reg_43_), .Y(core__abc_21302_new_n1692_));
AND2X2 AND2X2_41 ( .A(core_v1_reg_47_), .B(core_v0_reg_47_), .Y(core__abc_21302_new_n1738_));
AND2X2 AND2X2_42 ( .A(core_v2_reg_51_), .B(core_v3_reg_51_), .Y(core__abc_21302_new_n1787_));
AND2X2 AND2X2_43 ( .A(core_v2_reg_53_), .B(core_v3_reg_53_), .Y(core__abc_21302_new_n1813_));
AND2X2 AND2X2_44 ( .A(core_v1_reg_3_), .B(core_v0_reg_3_), .Y(core__abc_21302_new_n2373_));
AND2X2 AND2X2_45 ( .A(core_v1_reg_6_), .B(core_v0_reg_6_), .Y(core__abc_21302_new_n2380_));
AND2X2 AND2X2_46 ( .A(core_v1_reg_7_), .B(core_v0_reg_7_), .Y(core__abc_21302_new_n2383_));
AND2X2 AND2X2_47 ( .A(core_v1_reg_5_), .B(core_v0_reg_5_), .Y(core__abc_21302_new_n2388_));
AND2X2 AND2X2_48 ( .A(core__abc_21302_new_n1407_), .B(core__abc_21302_new_n1419_), .Y(core__abc_21302_new_n2432_));
AND2X2 AND2X2_49 ( .A(core__abc_21302_new_n1360_), .B(core__abc_21302_new_n1372_), .Y(core__abc_21302_new_n2481_));
AND2X2 AND2X2_5 ( .A(core_v2_reg_3_), .B(core_v3_reg_3_), .Y(core__abc_21302_new_n1244_));
AND2X2 AND2X2_50 ( .A(core__abc_21302_new_n1336_), .B(core__abc_21302_new_n1348_), .Y(core__abc_21302_new_n2482_));
AND2X2 AND2X2_51 ( .A(core__abc_21302_new_n1314_), .B(core__abc_21302_new_n1326_), .Y(core__abc_21302_new_n2484_));
AND2X2 AND2X2_52 ( .A(core__abc_21302_new_n2423_), .B(core__abc_21302_new_n2426_), .Y(core__abc_21302_new_n2493_));
AND2X2 AND2X2_53 ( .A(core__abc_21302_new_n2530_), .B(core__abc_21302_new_n2531_), .Y(core__abc_21302_new_n2532_));
AND2X2 AND2X2_54 ( .A(core__abc_21302_new_n1318_), .B(core__abc_21302_new_n1315_), .Y(core__abc_21302_new_n2534_));
AND2X2 AND2X2_55 ( .A(core__abc_21302_new_n1330_), .B(core__abc_21302_new_n1327_), .Y(core__abc_21302_new_n2535_));
AND2X2 AND2X2_56 ( .A(core__abc_21302_new_n1501_), .B(core__abc_21302_new_n1498_), .Y(core__abc_21302_new_n2551_));
AND2X2 AND2X2_57 ( .A(core__abc_21302_new_n1513_), .B(core__abc_21302_new_n1510_), .Y(core__abc_21302_new_n2552_));
AND2X2 AND2X2_58 ( .A(core__abc_21302_new_n2558_), .B(core__abc_21302_new_n2557_), .Y(core__abc_21302_new_n2559_));
AND2X2 AND2X2_59 ( .A(core__abc_21302_new_n1411_), .B(core__abc_21302_new_n1408_), .Y(core__abc_21302_new_n2560_));
AND2X2 AND2X2_6 ( .A(core_v2_reg_4_), .B(core_v3_reg_4_), .Y(core__abc_21302_new_n1254_));
AND2X2 AND2X2_60 ( .A(core__abc_21302_new_n1423_), .B(core__abc_21302_new_n1420_), .Y(core__abc_21302_new_n2561_));
AND2X2 AND2X2_61 ( .A(core__abc_21302_new_n1399_), .B(core__abc_21302_new_n1396_), .Y(core__abc_21302_new_n2563_));
AND2X2 AND2X2_62 ( .A(core__abc_21302_new_n2548_), .B(core__abc_21302_new_n2567_), .Y(core__abc_21302_new_n2568_));
AND2X2 AND2X2_63 ( .A(core__abc_21302_new_n2666_), .B(core__abc_21302_new_n2667_), .Y(core__abc_21302_new_n2670_));
AND2X2 AND2X2_64 ( .A(core__abc_21302_new_n2762_), .B(core__abc_21302_new_n2763_), .Y(core__abc_21302_new_n2764_));
AND2X2 AND2X2_65 ( .A(core__abc_21302_new_n2767_), .B(core__abc_21302_new_n1616_), .Y(core__abc_21302_new_n2768_));
AND2X2 AND2X2_66 ( .A(core__abc_21302_new_n2789_), .B(core__abc_21302_new_n2781_), .Y(core__abc_21302_new_n2790_));
AND2X2 AND2X2_67 ( .A(core__abc_21302_new_n2816_), .B(core__abc_21302_new_n2609_), .Y(core__abc_21302_new_n2817_));
AND2X2 AND2X2_68 ( .A(core__abc_21302_new_n2819_), .B(core__abc_21302_new_n2821_), .Y(core__abc_21302_new_n2822_));
AND2X2 AND2X2_69 ( .A(core__abc_21302_new_n2823_), .B(core__abc_21302_new_n2822_), .Y(core__abc_21302_new_n2824_));
AND2X2 AND2X2_7 ( .A(core_v2_reg_5_), .B(core_v3_reg_5_), .Y(core__abc_21302_new_n1266_));
AND2X2 AND2X2_70 ( .A(core__abc_21302_new_n2813_), .B(core__abc_21302_new_n2830_), .Y(core__abc_21302_new_n2831_));
AND2X2 AND2X2_71 ( .A(core__abc_21302_new_n2800_), .B(core__abc_21302_new_n1616_), .Y(core__abc_21302_new_n2841_));
AND2X2 AND2X2_72 ( .A(core__abc_21302_new_n2842_), .B(core__abc_21302_new_n1638_), .Y(core__abc_21302_new_n2844_));
AND2X2 AND2X2_73 ( .A(core__abc_21302_new_n2868_), .B(core_v3_reg_33_), .Y(core__abc_21302_new_n2870_));
AND2X2 AND2X2_74 ( .A(core_v1_reg_38_), .B(core_v0_reg_38_), .Y(core__abc_21302_new_n2879_));
AND2X2 AND2X2_75 ( .A(core__abc_21302_new_n2900_), .B(core__abc_21302_new_n2895_), .Y(core__abc_21302_new_n2901_));
AND2X2 AND2X2_76 ( .A(core__abc_21302_new_n2894_), .B(core__abc_21302_new_n2906_), .Y(core__abc_21302_new_n2907_));
AND2X2 AND2X2_77 ( .A(core__abc_21302_new_n2924_), .B(core__abc_21302_new_n2923_), .Y(core__abc_21302_new_n2925_));
AND2X2 AND2X2_78 ( .A(core__abc_21302_new_n2942_), .B(core__abc_21302_new_n2943_), .Y(core__abc_21302_new_n2944_));
AND2X2 AND2X2_79 ( .A(core__abc_21302_new_n2919_), .B(core__abc_21302_new_n2944_), .Y(core__abc_21302_new_n2946_));
AND2X2 AND2X2_8 ( .A(core_v2_reg_6_), .B(core_v3_reg_6_), .Y(core__abc_21302_new_n1276_));
AND2X2 AND2X2_80 ( .A(core__abc_21302_new_n2965_), .B(core__abc_21302_new_n2967_), .Y(core__abc_21302_new_n2973_));
AND2X2 AND2X2_81 ( .A(core__abc_21302_new_n2979_), .B(core__abc_21302_new_n2991_), .Y(core__abc_21302_new_n2992_));
AND2X2 AND2X2_82 ( .A(core__abc_21302_new_n3012_), .B(core__abc_21302_new_n3006_), .Y(core__abc_21302_new_n3014_));
AND2X2 AND2X2_83 ( .A(core__abc_21302_new_n2522_), .B(core__abc_21302_new_n2519_), .Y(core__abc_21302_new_n3015_));
AND2X2 AND2X2_84 ( .A(core__abc_21302_new_n3023_), .B(core__abc_21302_new_n3020_), .Y(core__abc_21302_new_n3024_));
AND2X2 AND2X2_85 ( .A(core__abc_21302_new_n3051_), .B(core__abc_21302_new_n3052_), .Y(core__abc_21302_new_n3053_));
AND2X2 AND2X2_86 ( .A(core__abc_21302_new_n3055_), .B(core__abc_21302_new_n3054_), .Y(core__abc_21302_new_n3056_));
AND2X2 AND2X2_87 ( .A(core__abc_21302_new_n2639__bF_buf2), .B(core_key_76_), .Y(core__abc_21302_new_n3082_));
AND2X2 AND2X2_88 ( .A(core__abc_21302_new_n3139_), .B(core__abc_21302_new_n3140_), .Y(core__abc_21302_new_n3141_));
AND2X2 AND2X2_89 ( .A(core__abc_21302_new_n3151_), .B(core__abc_21302_new_n3149_), .Y(core__abc_21302_new_n3153_));
AND2X2 AND2X2_9 ( .A(core_v2_reg_7_), .B(core_v3_reg_7_), .Y(core__abc_21302_new_n1286_));
AND2X2 AND2X2_90 ( .A(core__abc_21302_new_n3190_), .B(core__abc_21302_new_n3186_), .Y(core__abc_21302_new_n3191_));
AND2X2 AND2X2_91 ( .A(core__abc_21302_new_n3196_), .B(core__abc_21302_new_n3194_), .Y(core__abc_21302_new_n3201_));
AND2X2 AND2X2_92 ( .A(core__abc_21302_new_n3202_), .B(core__abc_21302_new_n3198_), .Y(core__abc_21302_new_n3203_));
AND2X2 AND2X2_93 ( .A(core__abc_21302_new_n1853_), .B(core__abc_21302_new_n1865_), .Y(core__abc_21302_new_n3207_));
AND2X2 AND2X2_94 ( .A(core__abc_21302_new_n3229_), .B(core__abc_21302_new_n3227_), .Y(core__abc_21302_new_n3230_));
AND2X2 AND2X2_95 ( .A(core__abc_21302_new_n3231_), .B(core__abc_21302_new_n3234_), .Y(core__abc_21302_new_n3235_));
AND2X2 AND2X2_96 ( .A(core__abc_21302_new_n3248_), .B(core__abc_21302_new_n1879_), .Y(core__abc_21302_new_n3250_));
AND2X2 AND2X2_97 ( .A(core__abc_21302_new_n2639__bF_buf1), .B(core_key_79_), .Y(core__abc_21302_new_n3259_));
AND2X2 AND2X2_98 ( .A(core__abc_21302_new_n2639__bF_buf0), .B(core_key_80_), .Y(core__abc_21302_new_n3266_));
AND2X2 AND2X2_99 ( .A(core__abc_21302_new_n3142_), .B(core__abc_21302_new_n3144_), .Y(core__abc_21302_new_n3270_));
AOI21X1 AOI21X1_1 ( .A(_abc_19873_new_n908_), .B(_abc_19873_new_n926_), .C(_abc_19873_new_n928__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_27087_0_));
AOI21X1 AOI21X1_10 ( .A(_abc_19873_new_n1106_), .B(_abc_19873_new_n1115_), .C(_abc_19873_new_n928__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_27087_9_));
AOI21X1 AOI21X1_100 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1694_), .C(_abc_19873_new_n1695_), .Y(_0word1_reg_31_0__2_));
AOI21X1 AOI21X1_1000 ( .A(core__abc_21302_new_n6443_), .B(core__abc_21302_new_n6445_), .C(core__abc_21302_new_n6446_), .Y(core__0v1_reg_63_0__63_));
AOI21X1 AOI21X1_1001 ( .A(core__abc_21302_new_n6455_), .B(core__abc_21302_new_n6451_), .C(core__abc_21302_new_n1185__bF_buf2), .Y(core__0v0_reg_63_0__0_));
AOI21X1 AOI21X1_1002 ( .A(core__abc_21302_new_n6461_), .B(core__abc_21302_new_n6462_), .C(core__abc_21302_new_n1185__bF_buf1), .Y(core__0v0_reg_63_0__1_));
AOI21X1 AOI21X1_1003 ( .A(core__abc_21302_new_n6469_), .B(core__abc_21302_new_n6470_), .C(core__abc_21302_new_n1185__bF_buf0), .Y(core__0v0_reg_63_0__2_));
AOI21X1 AOI21X1_1004 ( .A(core__abc_21302_new_n6476_), .B(core__abc_21302_new_n6472_), .C(core__abc_21302_new_n1185__bF_buf13), .Y(core__0v0_reg_63_0__3_));
AOI21X1 AOI21X1_1005 ( .A(core__abc_21302_new_n6482_), .B(core__abc_21302_new_n6483_), .C(core__abc_21302_new_n1185__bF_buf12), .Y(core__0v0_reg_63_0__4_));
AOI21X1 AOI21X1_1006 ( .A(core__abc_21302_new_n6489_), .B(core__abc_21302_new_n6490_), .C(core__abc_21302_new_n1185__bF_buf11), .Y(core__0v0_reg_63_0__5_));
AOI21X1 AOI21X1_1007 ( .A(core__abc_21302_new_n6496_), .B(core__abc_21302_new_n6497_), .C(core__abc_21302_new_n1185__bF_buf10), .Y(core__0v0_reg_63_0__6_));
AOI21X1 AOI21X1_1008 ( .A(core__abc_21302_new_n6503_), .B(core__abc_21302_new_n6504_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v0_reg_63_0__7_));
AOI21X1 AOI21X1_1009 ( .A(core__abc_21302_new_n6510_), .B(core__abc_21302_new_n6511_), .C(core__abc_21302_new_n1185__bF_buf8), .Y(core__0v0_reg_63_0__8_));
AOI21X1 AOI21X1_101 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1697_), .C(_abc_19873_new_n1698_), .Y(_0word1_reg_31_0__3_));
AOI21X1 AOI21X1_1010 ( .A(core__abc_21302_new_n6518_), .B(core__abc_21302_new_n6519_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0v0_reg_63_0__9_));
AOI21X1 AOI21X1_1011 ( .A(core__abc_21302_new_n6525_), .B(core__abc_21302_new_n6526_), .C(core__abc_21302_new_n1185__bF_buf6), .Y(core__0v0_reg_63_0__10_));
AOI21X1 AOI21X1_1012 ( .A(core__abc_21302_new_n6532_), .B(core__abc_21302_new_n6533_), .C(core__abc_21302_new_n1185__bF_buf5), .Y(core__0v0_reg_63_0__11_));
AOI21X1 AOI21X1_1013 ( .A(core__abc_21302_new_n6540_), .B(core__abc_21302_new_n6541_), .C(core__abc_21302_new_n1185__bF_buf4), .Y(core__0v0_reg_63_0__12_));
AOI21X1 AOI21X1_1014 ( .A(core__abc_21302_new_n6547_), .B(core__abc_21302_new_n6548_), .C(core__abc_21302_new_n1185__bF_buf3), .Y(core__0v0_reg_63_0__13_));
AOI21X1 AOI21X1_1015 ( .A(core__abc_21302_new_n6554_), .B(core__abc_21302_new_n6555_), .C(core__abc_21302_new_n1185__bF_buf2), .Y(core__0v0_reg_63_0__14_));
AOI21X1 AOI21X1_1016 ( .A(core__abc_21302_new_n3243_), .B(core__abc_21302_new_n3244_), .C(core__abc_21302_new_n2673__bF_buf4), .Y(core__abc_21302_new_n6557_));
AOI21X1 AOI21X1_1017 ( .A(core__abc_21302_new_n6561_), .B(core__abc_21302_new_n6562_), .C(core__abc_21302_new_n1185__bF_buf1), .Y(core__0v0_reg_63_0__15_));
AOI21X1 AOI21X1_1018 ( .A(core__abc_21302_new_n6568_), .B(core__abc_21302_new_n6569_), .C(core__abc_21302_new_n1185__bF_buf0), .Y(core__0v0_reg_63_0__16_));
AOI21X1 AOI21X1_1019 ( .A(core__abc_21302_new_n6575_), .B(core__abc_21302_new_n6576_), .C(core__abc_21302_new_n1185__bF_buf13), .Y(core__0v0_reg_63_0__17_));
AOI21X1 AOI21X1_102 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1700_), .C(_abc_19873_new_n1701_), .Y(_0word1_reg_31_0__4_));
AOI21X1 AOI21X1_1020 ( .A(core__abc_21302_new_n6583_), .B(core__abc_21302_new_n6584_), .C(core__abc_21302_new_n1185__bF_buf12), .Y(core__0v0_reg_63_0__18_));
AOI21X1 AOI21X1_1021 ( .A(core__abc_21302_new_n3436_), .B(core__abc_21302_new_n3437_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n6586_));
AOI21X1 AOI21X1_1022 ( .A(core__abc_21302_new_n6590_), .B(core__abc_21302_new_n6591_), .C(core__abc_21302_new_n1185__bF_buf11), .Y(core__0v0_reg_63_0__19_));
AOI21X1 AOI21X1_1023 ( .A(core__abc_21302_new_n6597_), .B(core__abc_21302_new_n6598_), .C(core__abc_21302_new_n1185__bF_buf10), .Y(core__0v0_reg_63_0__20_));
AOI21X1 AOI21X1_1024 ( .A(core__abc_21302_new_n6604_), .B(core__abc_21302_new_n6605_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v0_reg_63_0__21_));
AOI21X1 AOI21X1_1025 ( .A(core__abc_21302_new_n6611_), .B(core__abc_21302_new_n6612_), .C(core__abc_21302_new_n1185__bF_buf8), .Y(core__0v0_reg_63_0__22_));
AOI21X1 AOI21X1_1026 ( .A(core__abc_21302_new_n3594_), .B(core__abc_21302_new_n3593_), .C(core__abc_21302_new_n2673__bF_buf10), .Y(core__abc_21302_new_n6614_));
AOI21X1 AOI21X1_1027 ( .A(core__abc_21302_new_n6618_), .B(core__abc_21302_new_n6619_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0v0_reg_63_0__23_));
AOI21X1 AOI21X1_1028 ( .A(core__abc_21302_new_n6625_), .B(core__abc_21302_new_n6626_), .C(core__abc_21302_new_n1185__bF_buf6), .Y(core__0v0_reg_63_0__24_));
AOI21X1 AOI21X1_1029 ( .A(core__abc_21302_new_n6633_), .B(core__abc_21302_new_n6634_), .C(core__abc_21302_new_n1185__bF_buf5), .Y(core__0v0_reg_63_0__25_));
AOI21X1 AOI21X1_103 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1035_), .C(_abc_19873_new_n1703_), .Y(_0word1_reg_31_0__5_));
AOI21X1 AOI21X1_1030 ( .A(core__abc_21302_new_n6641_), .B(core__abc_21302_new_n6642_), .C(core__abc_21302_new_n1185__bF_buf4), .Y(core__0v0_reg_63_0__26_));
AOI21X1 AOI21X1_1031 ( .A(core__abc_21302_new_n3750_), .B(core__abc_21302_new_n3749_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n6644_));
AOI21X1 AOI21X1_1032 ( .A(core__abc_21302_new_n6649_), .B(core__abc_21302_new_n6650_), .C(core__abc_21302_new_n1185__bF_buf3), .Y(core__0v0_reg_63_0__27_));
AOI21X1 AOI21X1_1033 ( .A(core__abc_21302_new_n6656_), .B(core__abc_21302_new_n6657_), .C(core__abc_21302_new_n1185__bF_buf2), .Y(core__0v0_reg_63_0__28_));
AOI21X1 AOI21X1_1034 ( .A(core__abc_21302_new_n6663_), .B(core__abc_21302_new_n6664_), .C(core__abc_21302_new_n1185__bF_buf1), .Y(core__0v0_reg_63_0__29_));
AOI21X1 AOI21X1_1035 ( .A(core__abc_21302_new_n6670_), .B(core__abc_21302_new_n6671_), .C(core__abc_21302_new_n1185__bF_buf0), .Y(core__0v0_reg_63_0__30_));
AOI21X1 AOI21X1_1036 ( .A(core__abc_21302_new_n3896_), .B(core__abc_21302_new_n3898_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n6673_));
AOI21X1 AOI21X1_1037 ( .A(core__abc_21302_new_n6677_), .B(core__abc_21302_new_n6678_), .C(core__abc_21302_new_n1185__bF_buf13), .Y(core__0v0_reg_63_0__31_));
AOI21X1 AOI21X1_1038 ( .A(core__abc_21302_new_n6683_), .B(core__abc_21302_new_n6684_), .C(core__abc_21302_new_n1185__bF_buf12), .Y(core__0v0_reg_63_0__32_));
AOI21X1 AOI21X1_1039 ( .A(core__abc_21302_new_n6689_), .B(core__abc_21302_new_n6690_), .C(core__abc_21302_new_n1185__bF_buf11), .Y(core__0v0_reg_63_0__33_));
AOI21X1 AOI21X1_104 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1705_), .C(_abc_19873_new_n1706_), .Y(_0word1_reg_31_0__6_));
AOI21X1 AOI21X1_1040 ( .A(core__abc_21302_new_n6696_), .B(core__abc_21302_new_n6697_), .C(core__abc_21302_new_n1185__bF_buf10), .Y(core__0v0_reg_63_0__34_));
AOI21X1 AOI21X1_1041 ( .A(core__abc_21302_new_n4019_), .B(core__abc_21302_new_n4020_), .C(core__abc_21302_new_n2673__bF_buf2), .Y(core__abc_21302_new_n6699_));
AOI21X1 AOI21X1_1042 ( .A(core__abc_21302_new_n6703_), .B(core__abc_21302_new_n6704_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v0_reg_63_0__35_));
AOI21X1 AOI21X1_1043 ( .A(core__abc_21302_new_n6710_), .B(core__abc_21302_new_n6711_), .C(core__abc_21302_new_n1185__bF_buf8), .Y(core__0v0_reg_63_0__36_));
AOI21X1 AOI21X1_1044 ( .A(core__abc_21302_new_n6716_), .B(core__abc_21302_new_n6717_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0v0_reg_63_0__37_));
AOI21X1 AOI21X1_1045 ( .A(core__abc_21302_new_n6723_), .B(core__abc_21302_new_n6724_), .C(core__abc_21302_new_n1185__bF_buf6), .Y(core__0v0_reg_63_0__38_));
AOI21X1 AOI21X1_1046 ( .A(core__abc_21302_new_n4142_), .B(core__abc_21302_new_n4140_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n6726_));
AOI21X1 AOI21X1_1047 ( .A(core__abc_21302_new_n6730_), .B(core__abc_21302_new_n6731_), .C(core__abc_21302_new_n1185__bF_buf5), .Y(core__0v0_reg_63_0__39_));
AOI21X1 AOI21X1_1048 ( .A(core__abc_21302_new_n6736_), .B(core__abc_21302_new_n6737_), .C(core__abc_21302_new_n1185__bF_buf4), .Y(core__0v0_reg_63_0__40_));
AOI21X1 AOI21X1_1049 ( .A(core__abc_21302_new_n6744_), .B(core__abc_21302_new_n6745_), .C(core__abc_21302_new_n1185__bF_buf3), .Y(core__0v0_reg_63_0__41_));
AOI21X1 AOI21X1_105 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1708_), .C(_abc_19873_new_n1709_), .Y(_0word1_reg_31_0__7_));
AOI21X1 AOI21X1_1050 ( .A(core__abc_21302_new_n6751_), .B(core__abc_21302_new_n6752_), .C(core__abc_21302_new_n1185__bF_buf2), .Y(core__0v0_reg_63_0__42_));
AOI21X1 AOI21X1_1051 ( .A(core__abc_21302_new_n4263_), .B(core__abc_21302_new_n4261_), .C(core__abc_21302_new_n2673__bF_buf8), .Y(core__abc_21302_new_n6754_));
AOI21X1 AOI21X1_1052 ( .A(core__abc_21302_new_n6758_), .B(core__abc_21302_new_n6759_), .C(core__abc_21302_new_n1185__bF_buf1), .Y(core__0v0_reg_63_0__43_));
AOI21X1 AOI21X1_1053 ( .A(core__abc_21302_new_n6765_), .B(core__abc_21302_new_n6766_), .C(core__abc_21302_new_n1185__bF_buf0), .Y(core__0v0_reg_63_0__44_));
AOI21X1 AOI21X1_1054 ( .A(core__abc_21302_new_n6772_), .B(core__abc_21302_new_n6773_), .C(core__abc_21302_new_n1185__bF_buf13), .Y(core__0v0_reg_63_0__45_));
AOI21X1 AOI21X1_1055 ( .A(core__abc_21302_new_n6779_), .B(core__abc_21302_new_n6780_), .C(core__abc_21302_new_n1185__bF_buf12), .Y(core__0v0_reg_63_0__46_));
AOI21X1 AOI21X1_1056 ( .A(core__abc_21302_new_n6786_), .B(core__abc_21302_new_n6787_), .C(core__abc_21302_new_n1185__bF_buf11), .Y(core__0v0_reg_63_0__47_));
AOI21X1 AOI21X1_1057 ( .A(core__abc_21302_new_n6792_), .B(core__abc_21302_new_n6793_), .C(core__abc_21302_new_n1185__bF_buf10), .Y(core__0v0_reg_63_0__48_));
AOI21X1 AOI21X1_1058 ( .A(core__abc_21302_new_n6799_), .B(core__abc_21302_new_n6800_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v0_reg_63_0__49_));
AOI21X1 AOI21X1_1059 ( .A(core__abc_21302_new_n6806_), .B(core__abc_21302_new_n6807_), .C(core__abc_21302_new_n1185__bF_buf8), .Y(core__0v0_reg_63_0__50_));
AOI21X1 AOI21X1_106 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1084_), .C(_abc_19873_new_n1711_), .Y(_0word1_reg_31_0__8_));
AOI21X1 AOI21X1_1060 ( .A(core__abc_21302_new_n4479_), .B(core__abc_21302_new_n4481_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n6809_));
AOI21X1 AOI21X1_1061 ( .A(core__abc_21302_new_n6813_), .B(core__abc_21302_new_n6814_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0v0_reg_63_0__51_));
AOI21X1 AOI21X1_1062 ( .A(core__abc_21302_new_n6821_), .B(core__abc_21302_new_n6822_), .C(core__abc_21302_new_n1185__bF_buf6), .Y(core__0v0_reg_63_0__52_));
AOI21X1 AOI21X1_1063 ( .A(core__abc_21302_new_n4528_), .B(core__abc_21302_new_n4526_), .C(core__abc_21302_new_n2673__bF_buf0), .Y(core__abc_21302_new_n6824_));
AOI21X1 AOI21X1_1064 ( .A(core__abc_21302_new_n6828_), .B(core__abc_21302_new_n6829_), .C(core__abc_21302_new_n1185__bF_buf5), .Y(core__0v0_reg_63_0__53_));
AOI21X1 AOI21X1_1065 ( .A(core__abc_21302_new_n6835_), .B(core__abc_21302_new_n6836_), .C(core__abc_21302_new_n1185__bF_buf4), .Y(core__0v0_reg_63_0__54_));
AOI21X1 AOI21X1_1066 ( .A(core__abc_21302_new_n4578_), .B(core__abc_21302_new_n4581_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n6838_));
AOI21X1 AOI21X1_1067 ( .A(core__abc_21302_new_n6842_), .B(core__abc_21302_new_n6843_), .C(core__abc_21302_new_n1185__bF_buf3), .Y(core__0v0_reg_63_0__55_));
AOI21X1 AOI21X1_1068 ( .A(core__abc_21302_new_n6849_), .B(core__abc_21302_new_n6850_), .C(core__abc_21302_new_n1185__bF_buf2), .Y(core__0v0_reg_63_0__56_));
AOI21X1 AOI21X1_1069 ( .A(core__abc_21302_new_n6857_), .B(core__abc_21302_new_n6858_), .C(core__abc_21302_new_n1185__bF_buf1), .Y(core__0v0_reg_63_0__57_));
AOI21X1 AOI21X1_107 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1103_), .C(_abc_19873_new_n1713_), .Y(_0word1_reg_31_0__9_));
AOI21X1 AOI21X1_1070 ( .A(core__abc_21302_new_n6865_), .B(core__abc_21302_new_n6866_), .C(core__abc_21302_new_n1185__bF_buf0), .Y(core__0v0_reg_63_0__58_));
AOI21X1 AOI21X1_1071 ( .A(core__abc_21302_new_n4683_), .B(core__abc_21302_new_n4686_), .C(core__abc_21302_new_n2673__bF_buf8), .Y(core__abc_21302_new_n6868_));
AOI21X1 AOI21X1_1072 ( .A(core__abc_21302_new_n6873_), .B(core__abc_21302_new_n6874_), .C(core__abc_21302_new_n1185__bF_buf13), .Y(core__0v0_reg_63_0__59_));
AOI21X1 AOI21X1_1073 ( .A(core__abc_21302_new_n6880_), .B(core__abc_21302_new_n6881_), .C(core__abc_21302_new_n1185__bF_buf12), .Y(core__0v0_reg_63_0__60_));
AOI21X1 AOI21X1_1074 ( .A(core__abc_21302_new_n4749_), .B(core__abc_21302_new_n4752_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n6883_));
AOI21X1 AOI21X1_1075 ( .A(core__abc_21302_new_n6887_), .B(core__abc_21302_new_n6888_), .C(core__abc_21302_new_n1185__bF_buf11), .Y(core__0v0_reg_63_0__61_));
AOI21X1 AOI21X1_1076 ( .A(core__abc_21302_new_n6895_), .B(core__abc_21302_new_n6896_), .C(core__abc_21302_new_n1185__bF_buf10), .Y(core__0v0_reg_63_0__62_));
AOI21X1 AOI21X1_1077 ( .A(core__abc_21302_new_n4809_), .B(core__abc_21302_new_n4807_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n6898_));
AOI21X1 AOI21X1_1078 ( .A(core__abc_21302_new_n6902_), .B(core__abc_21302_new_n6903_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v0_reg_63_0__63_));
AOI21X1 AOI21X1_1079 ( .A(core__abc_21302_new_n6912_), .B(core__abc_21302_new_n1150_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0siphash_valid_reg_0_0_));
AOI21X1 AOI21X1_108 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1122_), .C(_abc_19873_new_n1715_), .Y(_0word1_reg_31_0__10_));
AOI21X1 AOI21X1_109 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1717_), .C(_abc_19873_new_n1718_), .Y(_0word1_reg_31_0__11_));
AOI21X1 AOI21X1_11 ( .A(_abc_19873_new_n1125_), .B(_abc_19873_new_n1134_), .C(_abc_19873_new_n928__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_27087_10_));
AOI21X1 AOI21X1_110 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1720_), .C(_abc_19873_new_n1721_), .Y(_0word1_reg_31_0__12_));
AOI21X1 AOI21X1_111 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1723_), .C(_abc_19873_new_n1724_), .Y(_0word1_reg_31_0__13_));
AOI21X1 AOI21X1_112 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1726_), .C(_abc_19873_new_n1727_), .Y(_0word1_reg_31_0__14_));
AOI21X1 AOI21X1_113 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1215_), .C(_abc_19873_new_n1729_), .Y(_0word1_reg_31_0__15_));
AOI21X1 AOI21X1_114 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1731_), .C(_abc_19873_new_n1732_), .Y(_0word1_reg_31_0__16_));
AOI21X1 AOI21X1_115 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1734_), .C(_abc_19873_new_n1735_), .Y(_0word1_reg_31_0__17_));
AOI21X1 AOI21X1_116 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1737_), .C(_abc_19873_new_n1738_), .Y(_0word1_reg_31_0__18_));
AOI21X1 AOI21X1_117 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1740_), .C(_abc_19873_new_n1741_), .Y(_0word1_reg_31_0__19_));
AOI21X1 AOI21X1_118 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1743_), .C(_abc_19873_new_n1744_), .Y(_0word1_reg_31_0__20_));
AOI21X1 AOI21X1_119 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1746_), .C(_abc_19873_new_n1747_), .Y(_0word1_reg_31_0__21_));
AOI21X1 AOI21X1_12 ( .A(_abc_19873_new_n1153_), .B(_abc_19873_new_n1142_), .C(_abc_19873_new_n928__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_27087_11_));
AOI21X1 AOI21X1_120 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1749_), .C(_abc_19873_new_n1750_), .Y(_0word1_reg_31_0__22_));
AOI21X1 AOI21X1_121 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1361_), .C(_abc_19873_new_n1752_), .Y(_0word1_reg_31_0__23_));
AOI21X1 AOI21X1_122 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1754_), .C(_abc_19873_new_n1755_), .Y(_0word1_reg_31_0__24_));
AOI21X1 AOI21X1_123 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1757_), .C(_abc_19873_new_n1758_), .Y(_0word1_reg_31_0__25_));
AOI21X1 AOI21X1_124 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1416_), .C(_abc_19873_new_n1760_), .Y(_0word1_reg_31_0__26_));
AOI21X1 AOI21X1_125 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1435_), .C(_abc_19873_new_n1762_), .Y(_0word1_reg_31_0__27_));
AOI21X1 AOI21X1_126 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1764_), .C(_abc_19873_new_n1765_), .Y(_0word1_reg_31_0__28_));
AOI21X1 AOI21X1_127 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1467_), .C(_abc_19873_new_n1767_), .Y(_0word1_reg_31_0__29_));
AOI21X1 AOI21X1_128 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1769_), .C(_abc_19873_new_n1770_), .Y(_0word1_reg_31_0__30_));
AOI21X1 AOI21X1_129 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1510_), .C(_abc_19873_new_n1772_), .Y(_0word1_reg_31_0__31_));
AOI21X1 AOI21X1_13 ( .A(_abc_19873_new_n1172_), .B(_abc_19873_new_n1161_), .C(_abc_19873_new_n928__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_27087_12_));
AOI21X1 AOI21X1_130 ( .A(_abc_19873_new_n1774_), .B(_abc_19873_new_n1524__bF_buf14), .C(_abc_19873_new_n1775_), .Y(_0word0_reg_31_0__0_));
AOI21X1 AOI21X1_131 ( .A(_abc_19873_new_n1777_), .B(_abc_19873_new_n1524__bF_buf12), .C(_abc_19873_new_n1778_), .Y(_0word0_reg_31_0__1_));
AOI21X1 AOI21X1_132 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1780_), .C(_abc_19873_new_n1781_), .Y(_0word0_reg_31_0__2_));
AOI21X1 AOI21X1_133 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1783_), .C(_abc_19873_new_n1784_), .Y(_0word0_reg_31_0__3_));
AOI21X1 AOI21X1_134 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1786_), .C(_abc_19873_new_n1787_), .Y(_0word0_reg_31_0__4_));
AOI21X1 AOI21X1_135 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1789_), .C(_abc_19873_new_n1790_), .Y(_0word0_reg_31_0__5_));
AOI21X1 AOI21X1_136 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1792_), .C(_abc_19873_new_n1793_), .Y(_0word0_reg_31_0__6_));
AOI21X1 AOI21X1_137 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1062_), .C(_abc_19873_new_n1795_), .Y(_0word0_reg_31_0__7_));
AOI21X1 AOI21X1_138 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1085_), .C(_abc_19873_new_n1797_), .Y(_0word0_reg_31_0__8_));
AOI21X1 AOI21X1_139 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1104_), .C(_abc_19873_new_n1799_), .Y(_0word0_reg_31_0__9_));
AOI21X1 AOI21X1_14 ( .A(_abc_19873_new_n1190_), .B(_abc_19873_new_n1182_), .C(_abc_19873_new_n928__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_27087_13_));
AOI21X1 AOI21X1_140 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1123_), .C(_abc_19873_new_n1801_), .Y(_0word0_reg_31_0__10_));
AOI21X1 AOI21X1_141 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1150_), .C(_abc_19873_new_n1803_), .Y(_0word0_reg_31_0__11_));
AOI21X1 AOI21X1_142 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1169_), .C(_abc_19873_new_n1805_), .Y(_0word0_reg_31_0__12_));
AOI21X1 AOI21X1_143 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1807_), .C(_abc_19873_new_n1808_), .Y(_0word0_reg_31_0__13_));
AOI21X1 AOI21X1_144 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1198_), .C(_abc_19873_new_n1810_), .Y(_0word0_reg_31_0__14_));
AOI21X1 AOI21X1_145 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1216_), .C(_abc_19873_new_n1812_), .Y(_0word0_reg_31_0__15_));
AOI21X1 AOI21X1_146 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1235_), .C(_abc_19873_new_n1814_), .Y(_0word0_reg_31_0__16_));
AOI21X1 AOI21X1_147 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1250_), .C(_abc_19873_new_n1816_), .Y(_0word0_reg_31_0__17_));
AOI21X1 AOI21X1_148 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1279_), .C(_abc_19873_new_n1818_), .Y(_0word0_reg_31_0__18_));
AOI21X1 AOI21X1_149 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1290_), .C(_abc_19873_new_n1820_), .Y(_0word0_reg_31_0__19_));
AOI21X1 AOI21X1_15 ( .A(_abc_19873_new_n1208_), .B(_abc_19873_new_n1197_), .C(_abc_19873_new_n928__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_27087_14_));
AOI21X1 AOI21X1_150 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1315_), .C(_abc_19873_new_n1822_), .Y(_0word0_reg_31_0__20_));
AOI21X1 AOI21X1_151 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1824_), .C(_abc_19873_new_n1825_), .Y(_0word0_reg_31_0__21_));
AOI21X1 AOI21X1_152 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1344_), .C(_abc_19873_new_n1827_), .Y(_0word0_reg_31_0__22_));
AOI21X1 AOI21X1_153 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1362_), .C(_abc_19873_new_n1829_), .Y(_0word0_reg_31_0__23_));
AOI21X1 AOI21X1_154 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1381_), .C(_abc_19873_new_n1831_), .Y(_0word0_reg_31_0__24_));
AOI21X1 AOI21X1_155 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1399_), .C(_abc_19873_new_n1833_), .Y(_0word0_reg_31_0__25_));
AOI21X1 AOI21X1_156 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1417_), .C(_abc_19873_new_n1835_), .Y(_0word0_reg_31_0__26_));
AOI21X1 AOI21X1_157 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1436_), .C(_abc_19873_new_n1837_), .Y(_0word0_reg_31_0__27_));
AOI21X1 AOI21X1_158 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1455_), .C(_abc_19873_new_n1839_), .Y(_0word0_reg_31_0__28_));
AOI21X1 AOI21X1_159 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1468_), .C(_abc_19873_new_n1841_), .Y(_0word0_reg_31_0__29_));
AOI21X1 AOI21X1_16 ( .A(_abc_19873_new_n1218_), .B(_abc_19873_new_n1227_), .C(_abc_19873_new_n928__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_27087_15_));
AOI21X1 AOI21X1_160 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1493_), .C(_abc_19873_new_n1843_), .Y(_0word0_reg_31_0__30_));
AOI21X1 AOI21X1_161 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1511_), .C(_abc_19873_new_n1845_), .Y(_0word0_reg_31_0__31_));
AOI21X1 AOI21X1_162 ( .A(_abc_19873_new_n1847_), .B(_abc_19873_new_n1849__bF_buf6), .C(_abc_19873_new_n1850_), .Y(_0mi1_reg_31_0__0_));
AOI21X1 AOI21X1_163 ( .A(_abc_19873_new_n1852_), .B(_abc_19873_new_n1849__bF_buf4), .C(_abc_19873_new_n1853_), .Y(_0mi1_reg_31_0__1_));
AOI21X1 AOI21X1_164 ( .A(_abc_19873_new_n967_), .B(_abc_19873_new_n1849__bF_buf2), .C(_abc_19873_new_n1855_), .Y(_0mi1_reg_31_0__2_));
AOI21X1 AOI21X1_165 ( .A(_abc_19873_new_n978_), .B(_abc_19873_new_n1849__bF_buf0), .C(_abc_19873_new_n1857_), .Y(_0mi1_reg_31_0__3_));
AOI21X1 AOI21X1_166 ( .A(_abc_19873_new_n999_), .B(_abc_19873_new_n1849__bF_buf6), .C(_abc_19873_new_n1859_), .Y(_0mi1_reg_31_0__4_));
AOI21X1 AOI21X1_167 ( .A(_abc_19873_new_n1861_), .B(_abc_19873_new_n1849__bF_buf4), .C(_abc_19873_new_n1862_), .Y(_0mi1_reg_31_0__5_));
AOI21X1 AOI21X1_168 ( .A(_abc_19873_new_n1041_), .B(_abc_19873_new_n1849__bF_buf2), .C(_abc_19873_new_n1864_), .Y(_0mi1_reg_31_0__6_));
AOI21X1 AOI21X1_169 ( .A(_abc_19873_new_n1063_), .B(_abc_19873_new_n1849__bF_buf0), .C(_abc_19873_new_n1866_), .Y(_0mi1_reg_31_0__7_));
AOI21X1 AOI21X1_17 ( .A(_abc_19873_new_n1245_), .B(_abc_19873_new_n1234_), .C(_abc_19873_new_n928__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_27087_16_));
AOI21X1 AOI21X1_170 ( .A(_abc_19873_new_n1093_), .B(_abc_19873_new_n1849__bF_buf6), .C(_abc_19873_new_n1868_), .Y(_0mi1_reg_31_0__8_));
AOI21X1 AOI21X1_171 ( .A(_abc_19873_new_n1112_), .B(_abc_19873_new_n1849__bF_buf4), .C(_abc_19873_new_n1870_), .Y(_0mi1_reg_31_0__9_));
AOI21X1 AOI21X1_172 ( .A(_abc_19873_new_n1131_), .B(_abc_19873_new_n1849__bF_buf2), .C(_abc_19873_new_n1872_), .Y(_0mi1_reg_31_0__10_));
AOI21X1 AOI21X1_173 ( .A(_abc_19873_new_n1151_), .B(_abc_19873_new_n1849__bF_buf0), .C(_abc_19873_new_n1874_), .Y(_0mi1_reg_31_0__11_));
AOI21X1 AOI21X1_174 ( .A(_abc_19873_new_n1170_), .B(_abc_19873_new_n1849__bF_buf6), .C(_abc_19873_new_n1876_), .Y(_0mi1_reg_31_0__12_));
AOI21X1 AOI21X1_175 ( .A(_abc_19873_new_n1183_), .B(_abc_19873_new_n1849__bF_buf4), .C(_abc_19873_new_n1878_), .Y(_0mi1_reg_31_0__13_));
AOI21X1 AOI21X1_176 ( .A(_abc_19873_new_n1880_), .B(_abc_19873_new_n1849__bF_buf2), .C(_abc_19873_new_n1881_), .Y(_0mi1_reg_31_0__14_));
AOI21X1 AOI21X1_177 ( .A(_abc_19873_new_n1224_), .B(_abc_19873_new_n1849__bF_buf0), .C(_abc_19873_new_n1883_), .Y(_0mi1_reg_31_0__15_));
AOI21X1 AOI21X1_178 ( .A(_abc_19873_new_n1885_), .B(_abc_19873_new_n1849__bF_buf6), .C(_abc_19873_new_n1886_), .Y(_0mi1_reg_31_0__16_));
AOI21X1 AOI21X1_179 ( .A(_abc_19873_new_n1251_), .B(_abc_19873_new_n1849__bF_buf4), .C(_abc_19873_new_n1888_), .Y(_0mi1_reg_31_0__17_));
AOI21X1 AOI21X1_18 ( .A(_abc_19873_new_n1264_), .B(_abc_19873_new_n1253_), .C(_abc_19873_new_n928__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_27087_17_));
AOI21X1 AOI21X1_180 ( .A(_abc_19873_new_n1280_), .B(_abc_19873_new_n1849__bF_buf2), .C(_abc_19873_new_n1890_), .Y(_0mi1_reg_31_0__18_));
AOI21X1 AOI21X1_181 ( .A(_abc_19873_new_n1892_), .B(_abc_19873_new_n1849__bF_buf0), .C(_abc_19873_new_n1893_), .Y(_0mi1_reg_31_0__19_));
AOI21X1 AOI21X1_182 ( .A(_abc_19873_new_n1316_), .B(_abc_19873_new_n1849__bF_buf6), .C(_abc_19873_new_n1895_), .Y(_0mi1_reg_31_0__20_));
AOI21X1 AOI21X1_183 ( .A(_abc_19873_new_n1329_), .B(_abc_19873_new_n1849__bF_buf4), .C(_abc_19873_new_n1897_), .Y(_0mi1_reg_31_0__21_));
AOI21X1 AOI21X1_184 ( .A(_abc_19873_new_n1899_), .B(_abc_19873_new_n1849__bF_buf2), .C(_abc_19873_new_n1900_), .Y(_0mi1_reg_31_0__22_));
AOI21X1 AOI21X1_185 ( .A(_abc_19873_new_n1370_), .B(_abc_19873_new_n1849__bF_buf0), .C(_abc_19873_new_n1902_), .Y(_0mi1_reg_31_0__23_));
AOI21X1 AOI21X1_186 ( .A(_abc_19873_new_n1904_), .B(_abc_19873_new_n1849__bF_buf6), .C(_abc_19873_new_n1905_), .Y(_0mi1_reg_31_0__24_));
AOI21X1 AOI21X1_187 ( .A(_abc_19873_new_n1907_), .B(_abc_19873_new_n1849__bF_buf4), .C(_abc_19873_new_n1908_), .Y(_0mi1_reg_31_0__25_));
AOI21X1 AOI21X1_188 ( .A(_abc_19873_new_n1425_), .B(_abc_19873_new_n1849__bF_buf2), .C(_abc_19873_new_n1910_), .Y(_0mi1_reg_31_0__26_));
AOI21X1 AOI21X1_189 ( .A(_abc_19873_new_n1444_), .B(_abc_19873_new_n1849__bF_buf0), .C(_abc_19873_new_n1912_), .Y(_0mi1_reg_31_0__27_));
AOI21X1 AOI21X1_19 ( .A(_abc_19873_new_n1282_), .B(_abc_19873_new_n1271_), .C(_abc_19873_new_n928__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_27087_18_));
AOI21X1 AOI21X1_190 ( .A(_abc_19873_new_n1914_), .B(_abc_19873_new_n1849__bF_buf6), .C(_abc_19873_new_n1915_), .Y(_0mi1_reg_31_0__28_));
AOI21X1 AOI21X1_191 ( .A(_abc_19873_new_n1917_), .B(_abc_19873_new_n1849__bF_buf4), .C(_abc_19873_new_n1918_), .Y(_0mi1_reg_31_0__29_));
AOI21X1 AOI21X1_192 ( .A(_abc_19873_new_n1920_), .B(_abc_19873_new_n1849__bF_buf2), .C(_abc_19873_new_n1921_), .Y(_0mi1_reg_31_0__30_));
AOI21X1 AOI21X1_193 ( .A(_abc_19873_new_n1519_), .B(_abc_19873_new_n1849__bF_buf0), .C(_abc_19873_new_n1923_), .Y(_0mi1_reg_31_0__31_));
AOI21X1 AOI21X1_194 ( .A(_abc_19873_new_n909_), .B(_abc_19873_new_n1925__bF_buf6), .C(_abc_19873_new_n1926_), .Y(_0mi0_reg_31_0__0_));
AOI21X1 AOI21X1_195 ( .A(_abc_19873_new_n941_), .B(_abc_19873_new_n1925__bF_buf4), .C(_abc_19873_new_n1928_), .Y(_0mi0_reg_31_0__1_));
AOI21X1 AOI21X1_196 ( .A(_abc_19873_new_n968_), .B(_abc_19873_new_n1925__bF_buf2), .C(_abc_19873_new_n1930_), .Y(_0mi0_reg_31_0__2_));
AOI21X1 AOI21X1_197 ( .A(_abc_19873_new_n979_), .B(_abc_19873_new_n1925__bF_buf0), .C(_abc_19873_new_n1932_), .Y(_0mi0_reg_31_0__3_));
AOI21X1 AOI21X1_198 ( .A(_abc_19873_new_n1000_), .B(_abc_19873_new_n1925__bF_buf6), .C(_abc_19873_new_n1934_), .Y(_0mi0_reg_31_0__4_));
AOI21X1 AOI21X1_199 ( .A(_abc_19873_new_n1031_), .B(_abc_19873_new_n1925__bF_buf4), .C(_abc_19873_new_n1936_), .Y(_0mi0_reg_31_0__5_));
AOI21X1 AOI21X1_2 ( .A(_abc_19873_new_n940_), .B(_abc_19873_new_n950_), .C(_abc_19873_new_n928__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_27087_1_));
AOI21X1 AOI21X1_20 ( .A(_abc_19873_new_n1300_), .B(_abc_19873_new_n1289_), .C(_abc_19873_new_n928__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_27087_19_));
AOI21X1 AOI21X1_200 ( .A(_abc_19873_new_n1042_), .B(_abc_19873_new_n1925__bF_buf2), .C(_abc_19873_new_n1938_), .Y(_0mi0_reg_31_0__6_));
AOI21X1 AOI21X1_201 ( .A(_abc_19873_new_n1074_), .B(_abc_19873_new_n1925__bF_buf0), .C(_abc_19873_new_n1940_), .Y(_0mi0_reg_31_0__7_));
AOI21X1 AOI21X1_202 ( .A(_abc_19873_new_n1094_), .B(_abc_19873_new_n1925__bF_buf6), .C(_abc_19873_new_n1942_), .Y(_0mi0_reg_31_0__8_));
AOI21X1 AOI21X1_203 ( .A(_abc_19873_new_n1113_), .B(_abc_19873_new_n1925__bF_buf4), .C(_abc_19873_new_n1944_), .Y(_0mi0_reg_31_0__9_));
AOI21X1 AOI21X1_204 ( .A(_abc_19873_new_n1132_), .B(_abc_19873_new_n1925__bF_buf2), .C(_abc_19873_new_n1946_), .Y(_0mi0_reg_31_0__10_));
AOI21X1 AOI21X1_205 ( .A(_abc_19873_new_n1136_), .B(_abc_19873_new_n1925__bF_buf0), .C(_abc_19873_new_n1948_), .Y(_0mi0_reg_31_0__11_));
AOI21X1 AOI21X1_206 ( .A(_abc_19873_new_n1155_), .B(_abc_19873_new_n1925__bF_buf6), .C(_abc_19873_new_n1950_), .Y(_0mi0_reg_31_0__12_));
AOI21X1 AOI21X1_207 ( .A(_abc_19873_new_n1184_), .B(_abc_19873_new_n1925__bF_buf4), .C(_abc_19873_new_n1952_), .Y(_0mi0_reg_31_0__13_));
AOI21X1 AOI21X1_208 ( .A(_abc_19873_new_n1192_), .B(_abc_19873_new_n1925__bF_buf2), .C(_abc_19873_new_n1954_), .Y(_0mi0_reg_31_0__14_));
AOI21X1 AOI21X1_209 ( .A(_abc_19873_new_n1225_), .B(_abc_19873_new_n1925__bF_buf0), .C(_abc_19873_new_n1956_), .Y(_0mi0_reg_31_0__15_));
AOI21X1 AOI21X1_21 ( .A(_abc_19873_new_n1318_), .B(_abc_19873_new_n1307_), .C(_abc_19873_new_n928__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_27087_20_));
AOI21X1 AOI21X1_210 ( .A(_abc_19873_new_n1229_), .B(_abc_19873_new_n1925__bF_buf6), .C(_abc_19873_new_n1958_), .Y(_0mi0_reg_31_0__16_));
AOI21X1 AOI21X1_211 ( .A(_abc_19873_new_n1960_), .B(_abc_19873_new_n1925__bF_buf4), .C(_abc_19873_new_n1961_), .Y(_0mi0_reg_31_0__17_));
AOI21X1 AOI21X1_212 ( .A(_abc_19873_new_n1266_), .B(_abc_19873_new_n1925__bF_buf2), .C(_abc_19873_new_n1963_), .Y(_0mi0_reg_31_0__18_));
AOI21X1 AOI21X1_213 ( .A(_abc_19873_new_n1284_), .B(_abc_19873_new_n1925__bF_buf0), .C(_abc_19873_new_n1965_), .Y(_0mi0_reg_31_0__19_));
AOI21X1 AOI21X1_214 ( .A(_abc_19873_new_n1302_), .B(_abc_19873_new_n1925__bF_buf6), .C(_abc_19873_new_n1967_), .Y(_0mi0_reg_31_0__20_));
AOI21X1 AOI21X1_215 ( .A(_abc_19873_new_n1330_), .B(_abc_19873_new_n1925__bF_buf4), .C(_abc_19873_new_n1969_), .Y(_0mi0_reg_31_0__21_));
AOI21X1 AOI21X1_216 ( .A(_abc_19873_new_n1338_), .B(_abc_19873_new_n1925__bF_buf2), .C(_abc_19873_new_n1971_), .Y(_0mi0_reg_31_0__22_));
AOI21X1 AOI21X1_217 ( .A(_abc_19873_new_n1371_), .B(_abc_19873_new_n1925__bF_buf0), .C(_abc_19873_new_n1973_), .Y(_0mi0_reg_31_0__23_));
AOI21X1 AOI21X1_218 ( .A(_abc_19873_new_n1375_), .B(_abc_19873_new_n1925__bF_buf6), .C(_abc_19873_new_n1975_), .Y(_0mi0_reg_31_0__24_));
AOI21X1 AOI21X1_219 ( .A(_abc_19873_new_n1393_), .B(_abc_19873_new_n1925__bF_buf4), .C(_abc_19873_new_n1977_), .Y(_0mi0_reg_31_0__25_));
AOI21X1 AOI21X1_22 ( .A(_abc_19873_new_n1336_), .B(_abc_19873_new_n1328_), .C(_abc_19873_new_n928__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_27087_21_));
AOI21X1 AOI21X1_220 ( .A(_abc_19873_new_n1426_), .B(_abc_19873_new_n1925__bF_buf2), .C(_abc_19873_new_n1979_), .Y(_0mi0_reg_31_0__26_));
AOI21X1 AOI21X1_221 ( .A(_abc_19873_new_n1445_), .B(_abc_19873_new_n1925__bF_buf0), .C(_abc_19873_new_n1981_), .Y(_0mi0_reg_31_0__27_));
AOI21X1 AOI21X1_222 ( .A(_abc_19873_new_n1449_), .B(_abc_19873_new_n1925__bF_buf6), .C(_abc_19873_new_n1983_), .Y(_0mi0_reg_31_0__28_));
AOI21X1 AOI21X1_223 ( .A(_abc_19873_new_n1985_), .B(_abc_19873_new_n1925__bF_buf4), .C(_abc_19873_new_n1986_), .Y(_0mi0_reg_31_0__29_));
AOI21X1 AOI21X1_224 ( .A(_abc_19873_new_n1487_), .B(_abc_19873_new_n1925__bF_buf2), .C(_abc_19873_new_n1988_), .Y(_0mi0_reg_31_0__30_));
AOI21X1 AOI21X1_225 ( .A(_abc_19873_new_n1520_), .B(_abc_19873_new_n1925__bF_buf0), .C(_abc_19873_new_n1990_), .Y(_0mi0_reg_31_0__31_));
AOI21X1 AOI21X1_226 ( .A(_abc_19873_new_n910_), .B(_abc_19873_new_n1992__bF_buf6), .C(_abc_19873_new_n1993_), .Y(_0key3_reg_31_0__0_));
AOI21X1 AOI21X1_227 ( .A(_abc_19873_new_n942_), .B(_abc_19873_new_n1992__bF_buf4), .C(_abc_19873_new_n1995_), .Y(_0key3_reg_31_0__1_));
AOI21X1 AOI21X1_228 ( .A(_abc_19873_new_n955_), .B(_abc_19873_new_n1992__bF_buf2), .C(_abc_19873_new_n1997_), .Y(_0key3_reg_31_0__2_));
AOI21X1 AOI21X1_229 ( .A(_abc_19873_new_n992_), .B(_abc_19873_new_n1992__bF_buf0), .C(_abc_19873_new_n1999_), .Y(_0key3_reg_31_0__3_));
AOI21X1 AOI21X1_23 ( .A(_abc_19873_new_n1354_), .B(_abc_19873_new_n1343_), .C(_abc_19873_new_n928__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_27087_22_));
AOI21X1 AOI21X1_230 ( .A(_abc_19873_new_n1013_), .B(_abc_19873_new_n1992__bF_buf6), .C(_abc_19873_new_n2001_), .Y(_0key3_reg_31_0__4_));
AOI21X1 AOI21X1_231 ( .A(_abc_19873_new_n1032_), .B(_abc_19873_new_n1992__bF_buf4), .C(_abc_19873_new_n2003_), .Y(_0key3_reg_31_0__5_));
AOI21X1 AOI21X1_232 ( .A(_abc_19873_new_n1052_), .B(_abc_19873_new_n1992__bF_buf2), .C(_abc_19873_new_n2005_), .Y(_0key3_reg_31_0__6_));
AOI21X1 AOI21X1_233 ( .A(_abc_19873_new_n1075_), .B(_abc_19873_new_n1992__bF_buf0), .C(_abc_19873_new_n2007_), .Y(_0key3_reg_31_0__7_));
AOI21X1 AOI21X1_234 ( .A(_abc_19873_new_n1081_), .B(_abc_19873_new_n1992__bF_buf6), .C(_abc_19873_new_n2009_), .Y(_0key3_reg_31_0__8_));
AOI21X1 AOI21X1_235 ( .A(_abc_19873_new_n1100_), .B(_abc_19873_new_n1992__bF_buf4), .C(_abc_19873_new_n2011_), .Y(_0key3_reg_31_0__9_));
AOI21X1 AOI21X1_236 ( .A(_abc_19873_new_n1119_), .B(_abc_19873_new_n1992__bF_buf2), .C(_abc_19873_new_n2013_), .Y(_0key3_reg_31_0__10_));
AOI21X1 AOI21X1_237 ( .A(_abc_19873_new_n1137_), .B(_abc_19873_new_n1992__bF_buf0), .C(_abc_19873_new_n2015_), .Y(_0key3_reg_31_0__11_));
AOI21X1 AOI21X1_238 ( .A(_abc_19873_new_n1156_), .B(_abc_19873_new_n1992__bF_buf6), .C(_abc_19873_new_n2017_), .Y(_0key3_reg_31_0__12_));
AOI21X1 AOI21X1_239 ( .A(_abc_19873_new_n1179_), .B(_abc_19873_new_n1992__bF_buf4), .C(_abc_19873_new_n2019_), .Y(_0key3_reg_31_0__13_));
AOI21X1 AOI21X1_24 ( .A(_abc_19873_new_n1364_), .B(_abc_19873_new_n1373_), .C(_abc_19873_new_n928__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_27087_23_));
AOI21X1 AOI21X1_240 ( .A(_abc_19873_new_n1193_), .B(_abc_19873_new_n1992__bF_buf2), .C(_abc_19873_new_n2021_), .Y(_0key3_reg_31_0__14_));
AOI21X1 AOI21X1_241 ( .A(_abc_19873_new_n1212_), .B(_abc_19873_new_n1992__bF_buf0), .C(_abc_19873_new_n2023_), .Y(_0key3_reg_31_0__15_));
AOI21X1 AOI21X1_242 ( .A(_abc_19873_new_n1230_), .B(_abc_19873_new_n1992__bF_buf6), .C(_abc_19873_new_n2025_), .Y(_0key3_reg_31_0__16_));
AOI21X1 AOI21X1_243 ( .A(_abc_19873_new_n1261_), .B(_abc_19873_new_n1992__bF_buf4), .C(_abc_19873_new_n2027_), .Y(_0key3_reg_31_0__17_));
AOI21X1 AOI21X1_244 ( .A(_abc_19873_new_n1267_), .B(_abc_19873_new_n1992__bF_buf2), .C(_abc_19873_new_n2029_), .Y(_0key3_reg_31_0__18_));
AOI21X1 AOI21X1_245 ( .A(_abc_19873_new_n1285_), .B(_abc_19873_new_n1992__bF_buf0), .C(_abc_19873_new_n2031_), .Y(_0key3_reg_31_0__19_));
AOI21X1 AOI21X1_246 ( .A(_abc_19873_new_n1303_), .B(_abc_19873_new_n1992__bF_buf6), .C(_abc_19873_new_n2033_), .Y(_0key3_reg_31_0__20_));
AOI21X1 AOI21X1_247 ( .A(_abc_19873_new_n1325_), .B(_abc_19873_new_n1992__bF_buf4), .C(_abc_19873_new_n2035_), .Y(_0key3_reg_31_0__21_));
AOI21X1 AOI21X1_248 ( .A(_abc_19873_new_n1339_), .B(_abc_19873_new_n1992__bF_buf2), .C(_abc_19873_new_n2037_), .Y(_0key3_reg_31_0__22_));
AOI21X1 AOI21X1_249 ( .A(_abc_19873_new_n1358_), .B(_abc_19873_new_n1992__bF_buf0), .C(_abc_19873_new_n2039_), .Y(_0key3_reg_31_0__23_));
AOI21X1 AOI21X1_25 ( .A(_abc_19873_new_n1391_), .B(_abc_19873_new_n1380_), .C(_abc_19873_new_n928__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_27087_24_));
AOI21X1 AOI21X1_250 ( .A(_abc_19873_new_n1376_), .B(_abc_19873_new_n1992__bF_buf6), .C(_abc_19873_new_n2041_), .Y(_0key3_reg_31_0__24_));
AOI21X1 AOI21X1_251 ( .A(_abc_19873_new_n1394_), .B(_abc_19873_new_n1992__bF_buf4), .C(_abc_19873_new_n2043_), .Y(_0key3_reg_31_0__25_));
AOI21X1 AOI21X1_252 ( .A(_abc_19873_new_n1413_), .B(_abc_19873_new_n1992__bF_buf2), .C(_abc_19873_new_n2045_), .Y(_0key3_reg_31_0__26_));
AOI21X1 AOI21X1_253 ( .A(_abc_19873_new_n1432_), .B(_abc_19873_new_n1992__bF_buf0), .C(_abc_19873_new_n2047_), .Y(_0key3_reg_31_0__27_));
AOI21X1 AOI21X1_254 ( .A(_abc_19873_new_n1450_), .B(_abc_19873_new_n1992__bF_buf6), .C(_abc_19873_new_n2049_), .Y(_0key3_reg_31_0__28_));
AOI21X1 AOI21X1_255 ( .A(_abc_19873_new_n2051_), .B(_abc_19873_new_n1992__bF_buf4), .C(_abc_19873_new_n2052_), .Y(_0key3_reg_31_0__29_));
AOI21X1 AOI21X1_256 ( .A(_abc_19873_new_n1488_), .B(_abc_19873_new_n1992__bF_buf2), .C(_abc_19873_new_n2054_), .Y(_0key3_reg_31_0__30_));
AOI21X1 AOI21X1_257 ( .A(_abc_19873_new_n1507_), .B(_abc_19873_new_n1992__bF_buf0), .C(_abc_19873_new_n2056_), .Y(_0key3_reg_31_0__31_));
AOI21X1 AOI21X1_258 ( .A(_abc_19873_new_n884_), .B(_abc_19873_new_n2058__bF_buf6), .C(_abc_19873_new_n2059_), .Y(_0key2_reg_31_0__0_));
AOI21X1 AOI21X1_259 ( .A(_abc_19873_new_n933_), .B(_abc_19873_new_n2058__bF_buf4), .C(_abc_19873_new_n2061_), .Y(_0key2_reg_31_0__1_));
AOI21X1 AOI21X1_26 ( .A(_abc_19873_new_n1409_), .B(_abc_19873_new_n1398_), .C(_abc_19873_new_n928__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_27087_25_));
AOI21X1 AOI21X1_260 ( .A(_abc_19873_new_n956_), .B(_abc_19873_new_n2058__bF_buf2), .C(_abc_19873_new_n2063_), .Y(_0key2_reg_31_0__2_));
AOI21X1 AOI21X1_261 ( .A(_abc_19873_new_n993_), .B(_abc_19873_new_n2058__bF_buf0), .C(_abc_19873_new_n2065_), .Y(_0key2_reg_31_0__3_));
AOI21X1 AOI21X1_262 ( .A(_abc_19873_new_n1014_), .B(_abc_19873_new_n2058__bF_buf6), .C(_abc_19873_new_n2067_), .Y(_0key2_reg_31_0__4_));
AOI21X1 AOI21X1_263 ( .A(_abc_19873_new_n1020_), .B(_abc_19873_new_n2058__bF_buf4), .C(_abc_19873_new_n2069_), .Y(_0key2_reg_31_0__5_));
AOI21X1 AOI21X1_264 ( .A(_abc_19873_new_n2071_), .B(_abc_19873_new_n2058__bF_buf2), .C(_abc_19873_new_n2072_), .Y(_0key2_reg_31_0__6_));
AOI21X1 AOI21X1_265 ( .A(_abc_19873_new_n2074_), .B(_abc_19873_new_n2058__bF_buf0), .C(_abc_19873_new_n2075_), .Y(_0key2_reg_31_0__7_));
AOI21X1 AOI21X1_266 ( .A(_abc_19873_new_n1082_), .B(_abc_19873_new_n2058__bF_buf6), .C(_abc_19873_new_n2077_), .Y(_0key2_reg_31_0__8_));
AOI21X1 AOI21X1_267 ( .A(_abc_19873_new_n1101_), .B(_abc_19873_new_n2058__bF_buf4), .C(_abc_19873_new_n2079_), .Y(_0key2_reg_31_0__9_));
AOI21X1 AOI21X1_268 ( .A(_abc_19873_new_n1120_), .B(_abc_19873_new_n2058__bF_buf2), .C(_abc_19873_new_n2081_), .Y(_0key2_reg_31_0__10_));
AOI21X1 AOI21X1_269 ( .A(_abc_19873_new_n1139_), .B(_abc_19873_new_n2058__bF_buf0), .C(_abc_19873_new_n2083_), .Y(_0key2_reg_31_0__11_));
AOI21X1 AOI21X1_27 ( .A(_abc_19873_new_n1419_), .B(_abc_19873_new_n1428_), .C(_abc_19873_new_n928__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_27087_26_));
AOI21X1 AOI21X1_270 ( .A(_abc_19873_new_n1158_), .B(_abc_19873_new_n2058__bF_buf6), .C(_abc_19873_new_n2085_), .Y(_0key2_reg_31_0__12_));
AOI21X1 AOI21X1_271 ( .A(_abc_19873_new_n1180_), .B(_abc_19873_new_n2058__bF_buf4), .C(_abc_19873_new_n2087_), .Y(_0key2_reg_31_0__13_));
AOI21X1 AOI21X1_272 ( .A(_abc_19873_new_n1195_), .B(_abc_19873_new_n2058__bF_buf2), .C(_abc_19873_new_n2089_), .Y(_0key2_reg_31_0__14_));
AOI21X1 AOI21X1_273 ( .A(_abc_19873_new_n1213_), .B(_abc_19873_new_n2058__bF_buf0), .C(_abc_19873_new_n2091_), .Y(_0key2_reg_31_0__15_));
AOI21X1 AOI21X1_274 ( .A(_abc_19873_new_n1232_), .B(_abc_19873_new_n2058__bF_buf6), .C(_abc_19873_new_n2093_), .Y(_0key2_reg_31_0__16_));
AOI21X1 AOI21X1_275 ( .A(_abc_19873_new_n1254_), .B(_abc_19873_new_n2058__bF_buf4), .C(_abc_19873_new_n2095_), .Y(_0key2_reg_31_0__17_));
AOI21X1 AOI21X1_276 ( .A(_abc_19873_new_n1269_), .B(_abc_19873_new_n2058__bF_buf2), .C(_abc_19873_new_n2097_), .Y(_0key2_reg_31_0__18_));
AOI21X1 AOI21X1_277 ( .A(_abc_19873_new_n1287_), .B(_abc_19873_new_n2058__bF_buf0), .C(_abc_19873_new_n2099_), .Y(_0key2_reg_31_0__19_));
AOI21X1 AOI21X1_278 ( .A(_abc_19873_new_n1305_), .B(_abc_19873_new_n2058__bF_buf6), .C(_abc_19873_new_n2101_), .Y(_0key2_reg_31_0__20_));
AOI21X1 AOI21X1_279 ( .A(_abc_19873_new_n1326_), .B(_abc_19873_new_n2058__bF_buf4), .C(_abc_19873_new_n2103_), .Y(_0key2_reg_31_0__21_));
AOI21X1 AOI21X1_28 ( .A(_abc_19873_new_n1438_), .B(_abc_19873_new_n1447_), .C(_abc_19873_new_n928__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_27087_27_));
AOI21X1 AOI21X1_280 ( .A(_abc_19873_new_n1341_), .B(_abc_19873_new_n2058__bF_buf2), .C(_abc_19873_new_n2105_), .Y(_0key2_reg_31_0__22_));
AOI21X1 AOI21X1_281 ( .A(_abc_19873_new_n1359_), .B(_abc_19873_new_n2058__bF_buf0), .C(_abc_19873_new_n2107_), .Y(_0key2_reg_31_0__23_));
AOI21X1 AOI21X1_282 ( .A(_abc_19873_new_n1378_), .B(_abc_19873_new_n2058__bF_buf6), .C(_abc_19873_new_n2109_), .Y(_0key2_reg_31_0__24_));
AOI21X1 AOI21X1_283 ( .A(_abc_19873_new_n1396_), .B(_abc_19873_new_n2058__bF_buf4), .C(_abc_19873_new_n2111_), .Y(_0key2_reg_31_0__25_));
AOI21X1 AOI21X1_284 ( .A(_abc_19873_new_n1414_), .B(_abc_19873_new_n2058__bF_buf2), .C(_abc_19873_new_n2113_), .Y(_0key2_reg_31_0__26_));
AOI21X1 AOI21X1_285 ( .A(_abc_19873_new_n1433_), .B(_abc_19873_new_n2058__bF_buf0), .C(_abc_19873_new_n2115_), .Y(_0key2_reg_31_0__27_));
AOI21X1 AOI21X1_286 ( .A(_abc_19873_new_n1452_), .B(_abc_19873_new_n2058__bF_buf6), .C(_abc_19873_new_n2117_), .Y(_0key2_reg_31_0__28_));
AOI21X1 AOI21X1_287 ( .A(_abc_19873_new_n1477_), .B(_abc_19873_new_n2058__bF_buf4), .C(_abc_19873_new_n2119_), .Y(_0key2_reg_31_0__29_));
AOI21X1 AOI21X1_288 ( .A(_abc_19873_new_n1490_), .B(_abc_19873_new_n2058__bF_buf2), .C(_abc_19873_new_n2121_), .Y(_0key2_reg_31_0__30_));
AOI21X1 AOI21X1_289 ( .A(_abc_19873_new_n1508_), .B(_abc_19873_new_n2058__bF_buf0), .C(_abc_19873_new_n2123_), .Y(_0key2_reg_31_0__31_));
AOI21X1 AOI21X1_29 ( .A(_abc_19873_new_n1465_), .B(_abc_19873_new_n1454_), .C(_abc_19873_new_n928__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_27087_28_));
AOI21X1 AOI21X1_290 ( .A(_abc_19873_new_n885_), .B(_abc_19873_new_n2125__bF_buf6), .C(_abc_19873_new_n2126_), .Y(_0key1_reg_31_0__0_));
AOI21X1 AOI21X1_291 ( .A(_abc_19873_new_n934_), .B(_abc_19873_new_n2125__bF_buf4), .C(_abc_19873_new_n2128_), .Y(_0key1_reg_31_0__1_));
AOI21X1 AOI21X1_292 ( .A(_abc_19873_new_n958_), .B(_abc_19873_new_n2125__bF_buf2), .C(_abc_19873_new_n2130_), .Y(_0key1_reg_31_0__2_));
AOI21X1 AOI21X1_293 ( .A(_abc_19873_new_n2132_), .B(_abc_19873_new_n2125__bF_buf0), .C(_abc_19873_new_n2133_), .Y(_0key1_reg_31_0__3_));
AOI21X1 AOI21X1_294 ( .A(_abc_19873_new_n2135_), .B(_abc_19873_new_n2125__bF_buf6), .C(_abc_19873_new_n2136_), .Y(_0key1_reg_31_0__4_));
AOI21X1 AOI21X1_295 ( .A(_abc_19873_new_n2138_), .B(_abc_19873_new_n2125__bF_buf4), .C(_abc_19873_new_n2139_), .Y(_0key1_reg_31_0__5_));
AOI21X1 AOI21X1_296 ( .A(_abc_19873_new_n1055_), .B(_abc_19873_new_n2125__bF_buf2), .C(_abc_19873_new_n2141_), .Y(_0key1_reg_31_0__6_));
AOI21X1 AOI21X1_297 ( .A(_abc_19873_new_n1060_), .B(_abc_19873_new_n2125__bF_buf0), .C(_abc_19873_new_n2143_), .Y(_0key1_reg_31_0__7_));
AOI21X1 AOI21X1_298 ( .A(_abc_19873_new_n1090_), .B(_abc_19873_new_n2125__bF_buf6), .C(_abc_19873_new_n2145_), .Y(_0key1_reg_31_0__8_));
AOI21X1 AOI21X1_299 ( .A(_abc_19873_new_n1109_), .B(_abc_19873_new_n2125__bF_buf4), .C(_abc_19873_new_n2147_), .Y(_0key1_reg_31_0__9_));
AOI21X1 AOI21X1_3 ( .A(_abc_19873_new_n974_), .B(_abc_19873_new_n962_), .C(_abc_19873_new_n928__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_27087_2_));
AOI21X1 AOI21X1_30 ( .A(_abc_19873_new_n880_), .B(_abc_19873_new_n871_), .C(_abc_19873_new_n890_), .Y(_abc_19873_new_n1480_));
AOI21X1 AOI21X1_300 ( .A(_abc_19873_new_n1128_), .B(_abc_19873_new_n2125__bF_buf2), .C(_abc_19873_new_n2149_), .Y(_0key1_reg_31_0__10_));
AOI21X1 AOI21X1_301 ( .A(_abc_19873_new_n2151_), .B(_abc_19873_new_n2125__bF_buf0), .C(_abc_19873_new_n2152_), .Y(_0key1_reg_31_0__11_));
AOI21X1 AOI21X1_302 ( .A(_abc_19873_new_n2154_), .B(_abc_19873_new_n2125__bF_buf6), .C(_abc_19873_new_n2155_), .Y(_0key1_reg_31_0__12_));
AOI21X1 AOI21X1_303 ( .A(_abc_19873_new_n1174_), .B(_abc_19873_new_n2125__bF_buf4), .C(_abc_19873_new_n2157_), .Y(_0key1_reg_31_0__13_));
AOI21X1 AOI21X1_304 ( .A(_abc_19873_new_n1205_), .B(_abc_19873_new_n2125__bF_buf2), .C(_abc_19873_new_n2159_), .Y(_0key1_reg_31_0__14_));
AOI21X1 AOI21X1_305 ( .A(_abc_19873_new_n1221_), .B(_abc_19873_new_n2125__bF_buf0), .C(_abc_19873_new_n2161_), .Y(_0key1_reg_31_0__15_));
AOI21X1 AOI21X1_306 ( .A(_abc_19873_new_n1242_), .B(_abc_19873_new_n2125__bF_buf6), .C(_abc_19873_new_n2163_), .Y(_0key1_reg_31_0__16_));
AOI21X1 AOI21X1_307 ( .A(_abc_19873_new_n1255_), .B(_abc_19873_new_n2125__bF_buf4), .C(_abc_19873_new_n2165_), .Y(_0key1_reg_31_0__17_));
AOI21X1 AOI21X1_308 ( .A(_abc_19873_new_n2167_), .B(_abc_19873_new_n2125__bF_buf2), .C(_abc_19873_new_n2168_), .Y(_0key1_reg_31_0__18_));
AOI21X1 AOI21X1_309 ( .A(_abc_19873_new_n1297_), .B(_abc_19873_new_n2125__bF_buf0), .C(_abc_19873_new_n2170_), .Y(_0key1_reg_31_0__19_));
AOI21X1 AOI21X1_31 ( .A(_abc_19873_new_n1485_), .B(_abc_19873_new_n1473_), .C(_abc_19873_new_n928__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_27087_29_));
AOI21X1 AOI21X1_310 ( .A(_abc_19873_new_n2172_), .B(_abc_19873_new_n2125__bF_buf6), .C(_abc_19873_new_n2173_), .Y(_0key1_reg_31_0__20_));
AOI21X1 AOI21X1_311 ( .A(_abc_19873_new_n1322_), .B(_abc_19873_new_n2125__bF_buf4), .C(_abc_19873_new_n2175_), .Y(_0key1_reg_31_0__21_));
AOI21X1 AOI21X1_312 ( .A(_abc_19873_new_n1351_), .B(_abc_19873_new_n2125__bF_buf2), .C(_abc_19873_new_n2177_), .Y(_0key1_reg_31_0__22_));
AOI21X1 AOI21X1_313 ( .A(_abc_19873_new_n1367_), .B(_abc_19873_new_n2125__bF_buf0), .C(_abc_19873_new_n2179_), .Y(_0key1_reg_31_0__23_));
AOI21X1 AOI21X1_314 ( .A(_abc_19873_new_n1388_), .B(_abc_19873_new_n2125__bF_buf6), .C(_abc_19873_new_n2181_), .Y(_0key1_reg_31_0__24_));
AOI21X1 AOI21X1_315 ( .A(_abc_19873_new_n1406_), .B(_abc_19873_new_n2125__bF_buf4), .C(_abc_19873_new_n2183_), .Y(_0key1_reg_31_0__25_));
AOI21X1 AOI21X1_316 ( .A(_abc_19873_new_n1422_), .B(_abc_19873_new_n2125__bF_buf2), .C(_abc_19873_new_n2185_), .Y(_0key1_reg_31_0__26_));
AOI21X1 AOI21X1_317 ( .A(_abc_19873_new_n1441_), .B(_abc_19873_new_n2125__bF_buf0), .C(_abc_19873_new_n2187_), .Y(_0key1_reg_31_0__27_));
AOI21X1 AOI21X1_318 ( .A(_abc_19873_new_n1462_), .B(_abc_19873_new_n2125__bF_buf6), .C(_abc_19873_new_n2189_), .Y(_0key1_reg_31_0__28_));
AOI21X1 AOI21X1_319 ( .A(_abc_19873_new_n1478_), .B(_abc_19873_new_n2125__bF_buf4), .C(_abc_19873_new_n2191_), .Y(_0key1_reg_31_0__29_));
AOI21X1 AOI21X1_32 ( .A(_abc_19873_new_n1503_), .B(_abc_19873_new_n1492_), .C(_abc_19873_new_n928__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_27087_30_));
AOI21X1 AOI21X1_320 ( .A(_abc_19873_new_n1500_), .B(_abc_19873_new_n2125__bF_buf2), .C(_abc_19873_new_n2193_), .Y(_0key1_reg_31_0__30_));
AOI21X1 AOI21X1_321 ( .A(_abc_19873_new_n1516_), .B(_abc_19873_new_n2125__bF_buf0), .C(_abc_19873_new_n2195_), .Y(_0key1_reg_31_0__31_));
AOI21X1 AOI21X1_322 ( .A(_abc_19873_new_n2197_), .B(_abc_19873_new_n2198__bF_buf6), .C(_abc_19873_new_n2199_), .Y(_0key0_reg_31_0__0_));
AOI21X1 AOI21X1_323 ( .A(_abc_19873_new_n2201_), .B(_abc_19873_new_n2198__bF_buf4), .C(_abc_19873_new_n2202_), .Y(_0key0_reg_31_0__1_));
AOI21X1 AOI21X1_324 ( .A(_abc_19873_new_n959_), .B(_abc_19873_new_n2198__bF_buf2), .C(_abc_19873_new_n2204_), .Y(_0key0_reg_31_0__2_));
AOI21X1 AOI21X1_325 ( .A(_abc_19873_new_n989_), .B(_abc_19873_new_n2198__bF_buf0), .C(_abc_19873_new_n2206_), .Y(_0key0_reg_31_0__3_));
AOI21X1 AOI21X1_326 ( .A(_abc_19873_new_n1010_), .B(_abc_19873_new_n2198__bF_buf6), .C(_abc_19873_new_n2208_), .Y(_0key0_reg_31_0__4_));
AOI21X1 AOI21X1_327 ( .A(_abc_19873_new_n1028_), .B(_abc_19873_new_n2198__bF_buf4), .C(_abc_19873_new_n2210_), .Y(_0key0_reg_31_0__5_));
AOI21X1 AOI21X1_328 ( .A(_abc_19873_new_n1044_), .B(_abc_19873_new_n2198__bF_buf2), .C(_abc_19873_new_n2212_), .Y(_0key0_reg_31_0__6_));
AOI21X1 AOI21X1_329 ( .A(_abc_19873_new_n1059_), .B(_abc_19873_new_n2198__bF_buf0), .C(_abc_19873_new_n2214_), .Y(_0key0_reg_31_0__7_));
AOI21X1 AOI21X1_33 ( .A(_abc_19873_new_n1513_), .B(_abc_19873_new_n1522_), .C(_abc_19873_new_n928__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_27087_31_));
AOI21X1 AOI21X1_330 ( .A(_abc_19873_new_n1091_), .B(_abc_19873_new_n2198__bF_buf6), .C(_abc_19873_new_n2216_), .Y(_0key0_reg_31_0__8_));
AOI21X1 AOI21X1_331 ( .A(_abc_19873_new_n1110_), .B(_abc_19873_new_n2198__bF_buf4), .C(_abc_19873_new_n2218_), .Y(_0key0_reg_31_0__9_));
AOI21X1 AOI21X1_332 ( .A(_abc_19873_new_n1129_), .B(_abc_19873_new_n2198__bF_buf2), .C(_abc_19873_new_n2220_), .Y(_0key0_reg_31_0__10_));
AOI21X1 AOI21X1_333 ( .A(_abc_19873_new_n1147_), .B(_abc_19873_new_n2198__bF_buf0), .C(_abc_19873_new_n2222_), .Y(_0key0_reg_31_0__11_));
AOI21X1 AOI21X1_334 ( .A(_abc_19873_new_n1166_), .B(_abc_19873_new_n2198__bF_buf6), .C(_abc_19873_new_n2224_), .Y(_0key0_reg_31_0__12_));
AOI21X1 AOI21X1_335 ( .A(_abc_19873_new_n1175_), .B(_abc_19873_new_n2198__bF_buf4), .C(_abc_19873_new_n2226_), .Y(_0key0_reg_31_0__13_));
AOI21X1 AOI21X1_336 ( .A(_abc_19873_new_n1206_), .B(_abc_19873_new_n2198__bF_buf2), .C(_abc_19873_new_n2228_), .Y(_0key0_reg_31_0__14_));
AOI21X1 AOI21X1_337 ( .A(_abc_19873_new_n1222_), .B(_abc_19873_new_n2198__bF_buf0), .C(_abc_19873_new_n2230_), .Y(_0key0_reg_31_0__15_));
AOI21X1 AOI21X1_338 ( .A(_abc_19873_new_n1243_), .B(_abc_19873_new_n2198__bF_buf6), .C(_abc_19873_new_n2232_), .Y(_0key0_reg_31_0__16_));
AOI21X1 AOI21X1_339 ( .A(_abc_19873_new_n1247_), .B(_abc_19873_new_n2198__bF_buf4), .C(_abc_19873_new_n2234_), .Y(_0key0_reg_31_0__17_));
AOI21X1 AOI21X1_34 ( .A(_abc_19873_new_n921_), .B(_abc_19873_new_n1524__bF_buf14), .C(_abc_19873_new_n1525_), .Y(_0word3_reg_31_0__0_));
AOI21X1 AOI21X1_340 ( .A(_abc_19873_new_n1276_), .B(_abc_19873_new_n2198__bF_buf2), .C(_abc_19873_new_n2236_), .Y(_0key0_reg_31_0__18_));
AOI21X1 AOI21X1_341 ( .A(_abc_19873_new_n1298_), .B(_abc_19873_new_n2198__bF_buf0), .C(_abc_19873_new_n2238_), .Y(_0key0_reg_31_0__19_));
AOI21X1 AOI21X1_342 ( .A(_abc_19873_new_n1312_), .B(_abc_19873_new_n2198__bF_buf6), .C(_abc_19873_new_n2240_), .Y(_0key0_reg_31_0__20_));
AOI21X1 AOI21X1_343 ( .A(_abc_19873_new_n1323_), .B(_abc_19873_new_n2198__bF_buf4), .C(_abc_19873_new_n2242_), .Y(_0key0_reg_31_0__21_));
AOI21X1 AOI21X1_344 ( .A(_abc_19873_new_n1352_), .B(_abc_19873_new_n2198__bF_buf2), .C(_abc_19873_new_n2244_), .Y(_0key0_reg_31_0__22_));
AOI21X1 AOI21X1_345 ( .A(_abc_19873_new_n1368_), .B(_abc_19873_new_n2198__bF_buf0), .C(_abc_19873_new_n2246_), .Y(_0key0_reg_31_0__23_));
AOI21X1 AOI21X1_346 ( .A(_abc_19873_new_n1389_), .B(_abc_19873_new_n2198__bF_buf6), .C(_abc_19873_new_n2248_), .Y(_0key0_reg_31_0__24_));
AOI21X1 AOI21X1_347 ( .A(_abc_19873_new_n1407_), .B(_abc_19873_new_n2198__bF_buf4), .C(_abc_19873_new_n2250_), .Y(_0key0_reg_31_0__25_));
AOI21X1 AOI21X1_348 ( .A(_abc_19873_new_n1423_), .B(_abc_19873_new_n2198__bF_buf2), .C(_abc_19873_new_n2252_), .Y(_0key0_reg_31_0__26_));
AOI21X1 AOI21X1_349 ( .A(_abc_19873_new_n1442_), .B(_abc_19873_new_n2198__bF_buf0), .C(_abc_19873_new_n2254_), .Y(_0key0_reg_31_0__27_));
AOI21X1 AOI21X1_35 ( .A(_abc_19873_new_n947_), .B(_abc_19873_new_n1524__bF_buf12), .C(_abc_19873_new_n1527_), .Y(_0word3_reg_31_0__1_));
AOI21X1 AOI21X1_350 ( .A(_abc_19873_new_n1463_), .B(_abc_19873_new_n2198__bF_buf6), .C(_abc_19873_new_n2256_), .Y(_0key0_reg_31_0__28_));
AOI21X1 AOI21X1_351 ( .A(_abc_19873_new_n2258_), .B(_abc_19873_new_n2198__bF_buf4), .C(_abc_19873_new_n2259_), .Y(_0key0_reg_31_0__29_));
AOI21X1 AOI21X1_352 ( .A(_abc_19873_new_n1501_), .B(_abc_19873_new_n2198__bF_buf2), .C(_abc_19873_new_n2261_), .Y(_0key0_reg_31_0__30_));
AOI21X1 AOI21X1_353 ( .A(_abc_19873_new_n1517_), .B(_abc_19873_new_n2198__bF_buf0), .C(_abc_19873_new_n2263_), .Y(_0key0_reg_31_0__31_));
AOI21X1 AOI21X1_354 ( .A(_abc_19873_new_n916_), .B(_abc_19873_new_n2266_), .C(_abc_19873_new_n2267_), .Y(_0param_reg_7_0__0_));
AOI21X1 AOI21X1_355 ( .A(_abc_19873_new_n2265_), .B(\write_data[1] ), .C(_abc_19873_new_n2269_), .Y(_abc_19873_new_n2270_));
AOI21X1 AOI21X1_356 ( .A(_abc_19873_new_n971_), .B(_abc_19873_new_n2266_), .C(_abc_19873_new_n2272_), .Y(_0param_reg_7_0__2_));
AOI21X1 AOI21X1_357 ( .A(_abc_19873_new_n981_), .B(_abc_19873_new_n2266_), .C(_abc_19873_new_n2274_), .Y(_0param_reg_7_0__3_));
AOI21X1 AOI21X1_358 ( .A(_abc_19873_new_n1002_), .B(_abc_19873_new_n2266_), .C(_abc_19873_new_n2276_), .Y(_0param_reg_7_0__4_));
AOI21X1 AOI21X1_359 ( .A(_abc_19873_new_n1021_), .B(_abc_19873_new_n2266_), .C(_abc_19873_new_n2278_), .Y(_0param_reg_7_0__5_));
AOI21X1 AOI21X1_36 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1529_), .C(_abc_19873_new_n1530_), .Y(_0word3_reg_31_0__2_));
AOI21X1 AOI21X1_360 ( .A(_abc_19873_new_n2265_), .B(\write_data[6] ), .C(_abc_19873_new_n2269_), .Y(_abc_19873_new_n2280_));
AOI21X1 AOI21X1_361 ( .A(_abc_19873_new_n1071_), .B(_abc_19873_new_n2266_), .C(_abc_19873_new_n2282_), .Y(_0param_reg_7_0__7_));
AOI21X1 AOI21X1_362 ( .A(_abc_19873_new_n2293_), .B(_abc_19873_new_n2295_), .C(_abc_19873_new_n2296_), .Y(_0long_reg_0_0_));
AOI21X1 AOI21X1_363 ( .A(core_final_rounds_0_), .B(core_loop_ctr_reg_0_), .C(core__abc_21302_new_n1169_), .Y(core__abc_21302_new_n1170_));
AOI21X1 AOI21X1_364 ( .A(core__abc_21302_new_n1175_), .B(core__abc_21302_new_n1153_), .C(core__abc_21302_new_n1177_), .Y(core__abc_21302_new_n1178_));
AOI21X1 AOI21X1_365 ( .A(core__abc_21302_new_n1217_), .B(core_siphash_word1_we_bF_buf8), .C(core__abc_21302_new_n1218_), .Y(core__0siphash_word1_reg_63_0__0_));
AOI21X1 AOI21X1_366 ( .A(core__abc_21302_new_n1229_), .B(core_siphash_word1_we_bF_buf6), .C(core__abc_21302_new_n1230_), .Y(core__0siphash_word1_reg_63_0__1_));
AOI21X1 AOI21X1_367 ( .A(core__abc_21302_new_n1238_), .B(core_siphash_word1_we_bF_buf4), .C(core__abc_21302_new_n1239_), .Y(core__0siphash_word1_reg_63_0__2_));
AOI21X1 AOI21X1_368 ( .A(core__abc_21302_new_n1248_), .B(core_siphash_word1_we_bF_buf2), .C(core__abc_21302_new_n1249_), .Y(core__0siphash_word1_reg_63_0__3_));
AOI21X1 AOI21X1_369 ( .A(core__abc_21302_new_n1258_), .B(core_siphash_word1_we_bF_buf0), .C(core__abc_21302_new_n1259_), .Y(core__0siphash_word1_reg_63_0__4_));
AOI21X1 AOI21X1_37 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n976_), .C(_abc_19873_new_n1532_), .Y(_0word3_reg_31_0__3_));
AOI21X1 AOI21X1_370 ( .A(core__abc_21302_new_n1270_), .B(core_siphash_word1_we_bF_buf9), .C(core__abc_21302_new_n1271_), .Y(core__0siphash_word1_reg_63_0__5_));
AOI21X1 AOI21X1_371 ( .A(core__abc_21302_new_n1280_), .B(core_siphash_word1_we_bF_buf7), .C(core__abc_21302_new_n1281_), .Y(core__0siphash_word1_reg_63_0__6_));
AOI21X1 AOI21X1_372 ( .A(core__abc_21302_new_n1290_), .B(core_siphash_word1_we_bF_buf5), .C(core__abc_21302_new_n1291_), .Y(core__0siphash_word1_reg_63_0__7_));
AOI21X1 AOI21X1_373 ( .A(core__abc_21302_new_n1298_), .B(core_siphash_word1_we_bF_buf3), .C(core__abc_21302_new_n1299_), .Y(core__0siphash_word1_reg_63_0__8_));
AOI21X1 AOI21X1_374 ( .A(core__abc_21302_new_n1309_), .B(core_siphash_word1_we_bF_buf1), .C(core__abc_21302_new_n1310_), .Y(core__0siphash_word1_reg_63_0__9_));
AOI21X1 AOI21X1_375 ( .A(core__abc_21302_new_n1321_), .B(core_siphash_word1_we_bF_buf10), .C(core__abc_21302_new_n1322_), .Y(core__0siphash_word1_reg_63_0__10_));
AOI21X1 AOI21X1_376 ( .A(core__abc_21302_new_n1333_), .B(core_siphash_word1_we_bF_buf8), .C(core__abc_21302_new_n1334_), .Y(core__0siphash_word1_reg_63_0__11_));
AOI21X1 AOI21X1_377 ( .A(core__abc_21302_new_n1343_), .B(core_siphash_word1_we_bF_buf6), .C(core__abc_21302_new_n1344_), .Y(core__0siphash_word1_reg_63_0__12_));
AOI21X1 AOI21X1_378 ( .A(core__abc_21302_new_n1355_), .B(core_siphash_word1_we_bF_buf4), .C(core__abc_21302_new_n1356_), .Y(core__0siphash_word1_reg_63_0__13_));
AOI21X1 AOI21X1_379 ( .A(core__abc_21302_new_n1367_), .B(core_siphash_word1_we_bF_buf2), .C(core__abc_21302_new_n1368_), .Y(core__0siphash_word1_reg_63_0__14_));
AOI21X1 AOI21X1_38 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n997_), .C(_abc_19873_new_n1534_), .Y(_0word3_reg_31_0__4_));
AOI21X1 AOI21X1_380 ( .A(core__abc_21302_new_n1379_), .B(core_siphash_word1_we_bF_buf0), .C(core__abc_21302_new_n1380_), .Y(core__0siphash_word1_reg_63_0__15_));
AOI21X1 AOI21X1_381 ( .A(core__abc_21302_new_n1390_), .B(core_siphash_word1_we_bF_buf9), .C(core__abc_21302_new_n1391_), .Y(core__0siphash_word1_reg_63_0__16_));
AOI21X1 AOI21X1_382 ( .A(core__abc_21302_new_n1402_), .B(core_siphash_word1_we_bF_buf7), .C(core__abc_21302_new_n1403_), .Y(core__0siphash_word1_reg_63_0__17_));
AOI21X1 AOI21X1_383 ( .A(core__abc_21302_new_n1414_), .B(core_siphash_word1_we_bF_buf5), .C(core__abc_21302_new_n1415_), .Y(core__0siphash_word1_reg_63_0__18_));
AOI21X1 AOI21X1_384 ( .A(core__abc_21302_new_n1426_), .B(core_siphash_word1_we_bF_buf3), .C(core__abc_21302_new_n1427_), .Y(core__0siphash_word1_reg_63_0__19_));
AOI21X1 AOI21X1_385 ( .A(core__abc_21302_new_n1438_), .B(core_siphash_word1_we_bF_buf1), .C(core__abc_21302_new_n1439_), .Y(core__0siphash_word1_reg_63_0__20_));
AOI21X1 AOI21X1_386 ( .A(core__abc_21302_new_n1450_), .B(core_siphash_word1_we_bF_buf10), .C(core__abc_21302_new_n1451_), .Y(core__0siphash_word1_reg_63_0__21_));
AOI21X1 AOI21X1_387 ( .A(core__abc_21302_new_n1462_), .B(core_siphash_word1_we_bF_buf8), .C(core__abc_21302_new_n1463_), .Y(core__0siphash_word1_reg_63_0__22_));
AOI21X1 AOI21X1_388 ( .A(core__abc_21302_new_n1470_), .B(core_siphash_word1_we_bF_buf6), .C(core__abc_21302_new_n1471_), .Y(core__0siphash_word1_reg_63_0__23_));
AOI21X1 AOI21X1_389 ( .A(core__abc_21302_new_n1482_), .B(core_siphash_word1_we_bF_buf4), .C(core__abc_21302_new_n1483_), .Y(core__0siphash_word1_reg_63_0__24_));
AOI21X1 AOI21X1_39 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1034_), .C(_abc_19873_new_n1536_), .Y(_0word3_reg_31_0__5_));
AOI21X1 AOI21X1_390 ( .A(core__abc_21302_new_n1492_), .B(core_siphash_word1_we_bF_buf2), .C(core__abc_21302_new_n1493_), .Y(core__0siphash_word1_reg_63_0__25_));
AOI21X1 AOI21X1_391 ( .A(core__abc_21302_new_n1504_), .B(core_siphash_word1_we_bF_buf0), .C(core__abc_21302_new_n1505_), .Y(core__0siphash_word1_reg_63_0__26_));
AOI21X1 AOI21X1_392 ( .A(core__abc_21302_new_n1516_), .B(core_siphash_word1_we_bF_buf9), .C(core__abc_21302_new_n1517_), .Y(core__0siphash_word1_reg_63_0__27_));
AOI21X1 AOI21X1_393 ( .A(core__abc_21302_new_n1528_), .B(core_siphash_word1_we_bF_buf7), .C(core__abc_21302_new_n1529_), .Y(core__0siphash_word1_reg_63_0__28_));
AOI21X1 AOI21X1_394 ( .A(core__abc_21302_new_n1541_), .B(core_siphash_word1_we_bF_buf5), .C(core__abc_21302_new_n1542_), .Y(core__0siphash_word1_reg_63_0__29_));
AOI21X1 AOI21X1_395 ( .A(core__abc_21302_new_n1553_), .B(core_siphash_word1_we_bF_buf3), .C(core__abc_21302_new_n1554_), .Y(core__0siphash_word1_reg_63_0__30_));
AOI21X1 AOI21X1_396 ( .A(core__abc_21302_new_n1561_), .B(core_siphash_word1_we_bF_buf1), .C(core__abc_21302_new_n1562_), .Y(core__0siphash_word1_reg_63_0__31_));
AOI21X1 AOI21X1_397 ( .A(core__abc_21302_new_n1573_), .B(core_siphash_word1_we_bF_buf10), .C(core__abc_21302_new_n1574_), .Y(core__0siphash_word1_reg_63_0__32_));
AOI21X1 AOI21X1_398 ( .A(core__abc_21302_new_n1585_), .B(core_siphash_word1_we_bF_buf8), .C(core__abc_21302_new_n1586_), .Y(core__0siphash_word1_reg_63_0__33_));
AOI21X1 AOI21X1_399 ( .A(core__abc_21302_new_n1599_), .B(core_siphash_word1_we_bF_buf6), .C(core__abc_21302_new_n1600_), .Y(core__0siphash_word1_reg_63_0__34_));
AOI21X1 AOI21X1_4 ( .A(_abc_19873_new_n995_), .B(_abc_19873_new_n984_), .C(_abc_19873_new_n928__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_27087_3_));
AOI21X1 AOI21X1_40 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1039_), .C(_abc_19873_new_n1538_), .Y(_0word3_reg_31_0__6_));
AOI21X1 AOI21X1_400 ( .A(core__abc_21302_new_n1611_), .B(core_siphash_word1_we_bF_buf4), .C(core__abc_21302_new_n1612_), .Y(core__0siphash_word1_reg_63_0__35_));
AOI21X1 AOI21X1_401 ( .A(core__abc_21302_new_n1622_), .B(core_siphash_word1_we_bF_buf2), .C(core__abc_21302_new_n1623_), .Y(core__0siphash_word1_reg_63_0__36_));
AOI21X1 AOI21X1_402 ( .A(core__abc_21302_new_n1635_), .B(core_siphash_word1_we_bF_buf0), .C(core__abc_21302_new_n1636_), .Y(core__0siphash_word1_reg_63_0__37_));
AOI21X1 AOI21X1_403 ( .A(core__abc_21302_new_n1644_), .B(core_siphash_word1_we_bF_buf9), .C(core__abc_21302_new_n1645_), .Y(core__0siphash_word1_reg_63_0__38_));
AOI21X1 AOI21X1_404 ( .A(core__abc_21302_new_n1655_), .B(core_siphash_word1_we_bF_buf7), .C(core__abc_21302_new_n1656_), .Y(core__0siphash_word1_reg_63_0__39_));
AOI21X1 AOI21X1_405 ( .A(core__abc_21302_new_n1666_), .B(core_siphash_word1_we_bF_buf5), .C(core__abc_21302_new_n1667_), .Y(core__0siphash_word1_reg_63_0__40_));
AOI21X1 AOI21X1_406 ( .A(core__abc_21302_new_n1677_), .B(core_siphash_word1_we_bF_buf3), .C(core__abc_21302_new_n1678_), .Y(core__0siphash_word1_reg_63_0__41_));
AOI21X1 AOI21X1_407 ( .A(core__abc_21302_new_n1688_), .B(core_siphash_word1_we_bF_buf1), .C(core__abc_21302_new_n1689_), .Y(core__0siphash_word1_reg_63_0__42_));
AOI21X1 AOI21X1_408 ( .A(core__abc_21302_new_n1699_), .B(core_siphash_word1_we_bF_buf10), .C(core__abc_21302_new_n1700_), .Y(core__0siphash_word1_reg_63_0__43_));
AOI21X1 AOI21X1_409 ( .A(core__abc_21302_new_n1711_), .B(core_siphash_word1_we_bF_buf8), .C(core__abc_21302_new_n1712_), .Y(core__0siphash_word1_reg_63_0__44_));
AOI21X1 AOI21X1_41 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1540_), .C(_abc_19873_new_n1541_), .Y(_0word3_reg_31_0__7_));
AOI21X1 AOI21X1_410 ( .A(core__abc_21302_new_n1722_), .B(core_siphash_word1_we_bF_buf6), .C(core__abc_21302_new_n1723_), .Y(core__0siphash_word1_reg_63_0__45_));
AOI21X1 AOI21X1_411 ( .A(core__abc_21302_new_n1734_), .B(core_siphash_word1_we_bF_buf4), .C(core__abc_21302_new_n1735_), .Y(core__0siphash_word1_reg_63_0__46_));
AOI21X1 AOI21X1_412 ( .A(core__abc_21302_new_n1745_), .B(core_siphash_word1_we_bF_buf2), .C(core__abc_21302_new_n1746_), .Y(core__0siphash_word1_reg_63_0__47_));
AOI21X1 AOI21X1_413 ( .A(core__abc_21302_new_n1758_), .B(core_siphash_word1_we_bF_buf0), .C(core__abc_21302_new_n1759_), .Y(core__0siphash_word1_reg_63_0__48_));
AOI21X1 AOI21X1_414 ( .A(core__abc_21302_new_n1767_), .B(core_siphash_word1_we_bF_buf9), .C(core__abc_21302_new_n1768_), .Y(core__0siphash_word1_reg_63_0__49_));
AOI21X1 AOI21X1_415 ( .A(core__abc_21302_new_n1779_), .B(core_siphash_word1_we_bF_buf7), .C(core__abc_21302_new_n1780_), .Y(core__0siphash_word1_reg_63_0__50_));
AOI21X1 AOI21X1_416 ( .A(core__abc_21302_new_n1790_), .B(core_siphash_word1_we_bF_buf5), .C(core__abc_21302_new_n1791_), .Y(core__0siphash_word1_reg_63_0__51_));
AOI21X1 AOI21X1_417 ( .A(core__abc_21302_new_n1804_), .B(core_siphash_word1_we_bF_buf3), .C(core__abc_21302_new_n1805_), .Y(core__0siphash_word1_reg_63_0__52_));
AOI21X1 AOI21X1_418 ( .A(core__abc_21302_new_n1815_), .B(core_siphash_word1_we_bF_buf1), .C(core__abc_21302_new_n1816_), .Y(core__0siphash_word1_reg_63_0__53_));
AOI21X1 AOI21X1_419 ( .A(core__abc_21302_new_n1828_), .B(core_siphash_word1_we_bF_buf10), .C(core__abc_21302_new_n1829_), .Y(core__0siphash_word1_reg_63_0__54_));
AOI21X1 AOI21X1_42 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1088_), .C(_abc_19873_new_n1543_), .Y(_0word3_reg_31_0__8_));
AOI21X1 AOI21X1_420 ( .A(core__abc_21302_new_n1841_), .B(core_siphash_word1_we_bF_buf8), .C(core__abc_21302_new_n1842_), .Y(core__0siphash_word1_reg_63_0__55_));
AOI21X1 AOI21X1_421 ( .A(core__abc_21302_new_n1855_), .B(core_siphash_word1_we_bF_buf6), .C(core__abc_21302_new_n1856_), .Y(core__0siphash_word1_reg_63_0__56_));
AOI21X1 AOI21X1_422 ( .A(core__abc_21302_new_n1867_), .B(core_siphash_word1_we_bF_buf4), .C(core__abc_21302_new_n1868_), .Y(core__0siphash_word1_reg_63_0__57_));
AOI21X1 AOI21X1_423 ( .A(core__abc_21302_new_n1881_), .B(core_siphash_word1_we_bF_buf2), .C(core__abc_21302_new_n1882_), .Y(core__0siphash_word1_reg_63_0__58_));
AOI21X1 AOI21X1_424 ( .A(core__abc_21302_new_n1893_), .B(core_siphash_word1_we_bF_buf0), .C(core__abc_21302_new_n1894_), .Y(core__0siphash_word1_reg_63_0__59_));
AOI21X1 AOI21X1_425 ( .A(core__abc_21302_new_n1907_), .B(core_siphash_word1_we_bF_buf9), .C(core__abc_21302_new_n1908_), .Y(core__0siphash_word1_reg_63_0__60_));
AOI21X1 AOI21X1_426 ( .A(core__abc_21302_new_n1921_), .B(core_siphash_word1_we_bF_buf7), .C(core__abc_21302_new_n1922_), .Y(core__0siphash_word1_reg_63_0__61_));
AOI21X1 AOI21X1_427 ( .A(core__abc_21302_new_n1934_), .B(core_siphash_word1_we_bF_buf5), .C(core__abc_21302_new_n1935_), .Y(core__0siphash_word1_reg_63_0__62_));
AOI21X1 AOI21X1_428 ( .A(core__abc_21302_new_n1940_), .B(core_siphash_word1_we_bF_buf3), .C(core__abc_21302_new_n1941_), .Y(core__0siphash_word1_reg_63_0__63_));
AOI21X1 AOI21X1_429 ( .A(core__abc_21302_new_n2149_), .B(core__abc_21302_new_n2151_), .C(core__abc_21302_new_n2152_), .Y(core__0loop_ctr_reg_3_0__1_));
AOI21X1 AOI21X1_43 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1098_), .C(_abc_19873_new_n1545_), .Y(_0word3_reg_31_0__9_));
AOI21X1 AOI21X1_430 ( .A(core__abc_21302_new_n2149_), .B(core__abc_21302_new_n2154_), .C(core_loop_ctr_reg_2_), .Y(core__abc_21302_new_n2155_));
AOI21X1 AOI21X1_431 ( .A(core__abc_21302_new_n2144_), .B(core__abc_21302_new_n2142_), .C(core__abc_21302_new_n2157_), .Y(core__abc_21302_new_n2158_));
AOI21X1 AOI21X1_432 ( .A(core__abc_21302_new_n2161_), .B(core_loop_ctr_reg_3_), .C(core__abc_21302_new_n2162_), .Y(core__0loop_ctr_reg_3_0__3_));
AOI21X1 AOI21X1_433 ( .A(core__abc_21302_new_n2164_), .B(core__abc_21302_new_n2168__bF_buf11), .C(core__abc_21302_new_n2169_), .Y(core__0mi_reg_63_0__0_));
AOI21X1 AOI21X1_434 ( .A(core__abc_21302_new_n2171_), .B(core__abc_21302_new_n2168__bF_buf9), .C(core__abc_21302_new_n2172_), .Y(core__0mi_reg_63_0__1_));
AOI21X1 AOI21X1_435 ( .A(core__abc_21302_new_n2174_), .B(core__abc_21302_new_n2168__bF_buf7), .C(core__abc_21302_new_n2175_), .Y(core__0mi_reg_63_0__2_));
AOI21X1 AOI21X1_436 ( .A(core__abc_21302_new_n2177_), .B(core__abc_21302_new_n2168__bF_buf5), .C(core__abc_21302_new_n2178_), .Y(core__0mi_reg_63_0__3_));
AOI21X1 AOI21X1_437 ( .A(core__abc_21302_new_n2180_), .B(core__abc_21302_new_n2168__bF_buf3), .C(core__abc_21302_new_n2181_), .Y(core__0mi_reg_63_0__4_));
AOI21X1 AOI21X1_438 ( .A(core__abc_21302_new_n2183_), .B(core__abc_21302_new_n2168__bF_buf1), .C(core__abc_21302_new_n2184_), .Y(core__0mi_reg_63_0__5_));
AOI21X1 AOI21X1_439 ( .A(core__abc_21302_new_n2186_), .B(core__abc_21302_new_n2168__bF_buf12), .C(core__abc_21302_new_n2187_), .Y(core__0mi_reg_63_0__6_));
AOI21X1 AOI21X1_44 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1126_), .C(_abc_19873_new_n1547_), .Y(_0word3_reg_31_0__10_));
AOI21X1 AOI21X1_440 ( .A(core__abc_21302_new_n2189_), .B(core__abc_21302_new_n2168__bF_buf10), .C(core__abc_21302_new_n2190_), .Y(core__0mi_reg_63_0__7_));
AOI21X1 AOI21X1_441 ( .A(core__abc_21302_new_n2192_), .B(core__abc_21302_new_n2168__bF_buf8), .C(core__abc_21302_new_n2193_), .Y(core__0mi_reg_63_0__8_));
AOI21X1 AOI21X1_442 ( .A(core__abc_21302_new_n2195_), .B(core__abc_21302_new_n2168__bF_buf6), .C(core__abc_21302_new_n2196_), .Y(core__0mi_reg_63_0__9_));
AOI21X1 AOI21X1_443 ( .A(core__abc_21302_new_n2198_), .B(core__abc_21302_new_n2168__bF_buf4), .C(core__abc_21302_new_n2199_), .Y(core__0mi_reg_63_0__10_));
AOI21X1 AOI21X1_444 ( .A(core__abc_21302_new_n2201_), .B(core__abc_21302_new_n2168__bF_buf2), .C(core__abc_21302_new_n2202_), .Y(core__0mi_reg_63_0__11_));
AOI21X1 AOI21X1_445 ( .A(core__abc_21302_new_n2204_), .B(core__abc_21302_new_n2168__bF_buf0), .C(core__abc_21302_new_n2205_), .Y(core__0mi_reg_63_0__12_));
AOI21X1 AOI21X1_446 ( .A(core__abc_21302_new_n2207_), .B(core__abc_21302_new_n2168__bF_buf11), .C(core__abc_21302_new_n2208_), .Y(core__0mi_reg_63_0__13_));
AOI21X1 AOI21X1_447 ( .A(core__abc_21302_new_n2210_), .B(core__abc_21302_new_n2168__bF_buf9), .C(core__abc_21302_new_n2211_), .Y(core__0mi_reg_63_0__14_));
AOI21X1 AOI21X1_448 ( .A(core__abc_21302_new_n2213_), .B(core__abc_21302_new_n2168__bF_buf7), .C(core__abc_21302_new_n2214_), .Y(core__0mi_reg_63_0__15_));
AOI21X1 AOI21X1_449 ( .A(core__abc_21302_new_n2216_), .B(core__abc_21302_new_n2168__bF_buf5), .C(core__abc_21302_new_n2217_), .Y(core__0mi_reg_63_0__16_));
AOI21X1 AOI21X1_45 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1549_), .C(_abc_19873_new_n1550_), .Y(_0word3_reg_31_0__11_));
AOI21X1 AOI21X1_450 ( .A(core__abc_21302_new_n2219_), .B(core__abc_21302_new_n2168__bF_buf3), .C(core__abc_21302_new_n2220_), .Y(core__0mi_reg_63_0__17_));
AOI21X1 AOI21X1_451 ( .A(core__abc_21302_new_n2222_), .B(core__abc_21302_new_n2168__bF_buf1), .C(core__abc_21302_new_n2223_), .Y(core__0mi_reg_63_0__18_));
AOI21X1 AOI21X1_452 ( .A(core__abc_21302_new_n2225_), .B(core__abc_21302_new_n2168__bF_buf12), .C(core__abc_21302_new_n2226_), .Y(core__0mi_reg_63_0__19_));
AOI21X1 AOI21X1_453 ( .A(core__abc_21302_new_n2228_), .B(core__abc_21302_new_n2168__bF_buf10), .C(core__abc_21302_new_n2229_), .Y(core__0mi_reg_63_0__20_));
AOI21X1 AOI21X1_454 ( .A(core__abc_21302_new_n2231_), .B(core__abc_21302_new_n2168__bF_buf8), .C(core__abc_21302_new_n2232_), .Y(core__0mi_reg_63_0__21_));
AOI21X1 AOI21X1_455 ( .A(core__abc_21302_new_n2234_), .B(core__abc_21302_new_n2168__bF_buf6), .C(core__abc_21302_new_n2235_), .Y(core__0mi_reg_63_0__22_));
AOI21X1 AOI21X1_456 ( .A(core__abc_21302_new_n2237_), .B(core__abc_21302_new_n2168__bF_buf4), .C(core__abc_21302_new_n2238_), .Y(core__0mi_reg_63_0__23_));
AOI21X1 AOI21X1_457 ( .A(core__abc_21302_new_n2240_), .B(core__abc_21302_new_n2168__bF_buf2), .C(core__abc_21302_new_n2241_), .Y(core__0mi_reg_63_0__24_));
AOI21X1 AOI21X1_458 ( .A(core__abc_21302_new_n2243_), .B(core__abc_21302_new_n2168__bF_buf0), .C(core__abc_21302_new_n2244_), .Y(core__0mi_reg_63_0__25_));
AOI21X1 AOI21X1_459 ( .A(core__abc_21302_new_n2246_), .B(core__abc_21302_new_n2168__bF_buf11), .C(core__abc_21302_new_n2247_), .Y(core__0mi_reg_63_0__26_));
AOI21X1 AOI21X1_46 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1552_), .C(_abc_19873_new_n1553_), .Y(_0word3_reg_31_0__12_));
AOI21X1 AOI21X1_460 ( .A(core__abc_21302_new_n2249_), .B(core__abc_21302_new_n2168__bF_buf9), .C(core__abc_21302_new_n2250_), .Y(core__0mi_reg_63_0__27_));
AOI21X1 AOI21X1_461 ( .A(core__abc_21302_new_n2252_), .B(core__abc_21302_new_n2168__bF_buf7), .C(core__abc_21302_new_n2253_), .Y(core__0mi_reg_63_0__28_));
AOI21X1 AOI21X1_462 ( .A(core__abc_21302_new_n2255_), .B(core__abc_21302_new_n2168__bF_buf5), .C(core__abc_21302_new_n2256_), .Y(core__0mi_reg_63_0__29_));
AOI21X1 AOI21X1_463 ( .A(core__abc_21302_new_n2258_), .B(core__abc_21302_new_n2168__bF_buf3), .C(core__abc_21302_new_n2259_), .Y(core__0mi_reg_63_0__30_));
AOI21X1 AOI21X1_464 ( .A(core__abc_21302_new_n2261_), .B(core__abc_21302_new_n2168__bF_buf1), .C(core__abc_21302_new_n2262_), .Y(core__0mi_reg_63_0__31_));
AOI21X1 AOI21X1_465 ( .A(core__abc_21302_new_n2264_), .B(core__abc_21302_new_n2168__bF_buf12), .C(core__abc_21302_new_n2265_), .Y(core__0mi_reg_63_0__32_));
AOI21X1 AOI21X1_466 ( .A(core__abc_21302_new_n2267_), .B(core__abc_21302_new_n2168__bF_buf10), .C(core__abc_21302_new_n2268_), .Y(core__0mi_reg_63_0__33_));
AOI21X1 AOI21X1_467 ( .A(core__abc_21302_new_n2270_), .B(core__abc_21302_new_n2168__bF_buf8), .C(core__abc_21302_new_n2271_), .Y(core__0mi_reg_63_0__34_));
AOI21X1 AOI21X1_468 ( .A(core__abc_21302_new_n2273_), .B(core__abc_21302_new_n2168__bF_buf6), .C(core__abc_21302_new_n2274_), .Y(core__0mi_reg_63_0__35_));
AOI21X1 AOI21X1_469 ( .A(core__abc_21302_new_n2276_), .B(core__abc_21302_new_n2168__bF_buf4), .C(core__abc_21302_new_n2277_), .Y(core__0mi_reg_63_0__36_));
AOI21X1 AOI21X1_47 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1555_), .C(_abc_19873_new_n1556_), .Y(_0word3_reg_31_0__13_));
AOI21X1 AOI21X1_470 ( .A(core__abc_21302_new_n2279_), .B(core__abc_21302_new_n2168__bF_buf2), .C(core__abc_21302_new_n2280_), .Y(core__0mi_reg_63_0__37_));
AOI21X1 AOI21X1_471 ( .A(core__abc_21302_new_n2282_), .B(core__abc_21302_new_n2168__bF_buf0), .C(core__abc_21302_new_n2283_), .Y(core__0mi_reg_63_0__38_));
AOI21X1 AOI21X1_472 ( .A(core__abc_21302_new_n2285_), .B(core__abc_21302_new_n2168__bF_buf11), .C(core__abc_21302_new_n2286_), .Y(core__0mi_reg_63_0__39_));
AOI21X1 AOI21X1_473 ( .A(core__abc_21302_new_n2288_), .B(core__abc_21302_new_n2168__bF_buf9), .C(core__abc_21302_new_n2289_), .Y(core__0mi_reg_63_0__40_));
AOI21X1 AOI21X1_474 ( .A(core__abc_21302_new_n2291_), .B(core__abc_21302_new_n2168__bF_buf7), .C(core__abc_21302_new_n2292_), .Y(core__0mi_reg_63_0__41_));
AOI21X1 AOI21X1_475 ( .A(core__abc_21302_new_n2294_), .B(core__abc_21302_new_n2168__bF_buf5), .C(core__abc_21302_new_n2295_), .Y(core__0mi_reg_63_0__42_));
AOI21X1 AOI21X1_476 ( .A(core__abc_21302_new_n2297_), .B(core__abc_21302_new_n2168__bF_buf3), .C(core__abc_21302_new_n2298_), .Y(core__0mi_reg_63_0__43_));
AOI21X1 AOI21X1_477 ( .A(core__abc_21302_new_n2300_), .B(core__abc_21302_new_n2168__bF_buf1), .C(core__abc_21302_new_n2301_), .Y(core__0mi_reg_63_0__44_));
AOI21X1 AOI21X1_478 ( .A(core__abc_21302_new_n2303_), .B(core__abc_21302_new_n2168__bF_buf12), .C(core__abc_21302_new_n2304_), .Y(core__0mi_reg_63_0__45_));
AOI21X1 AOI21X1_479 ( .A(core__abc_21302_new_n2306_), .B(core__abc_21302_new_n2168__bF_buf10), .C(core__abc_21302_new_n2307_), .Y(core__0mi_reg_63_0__46_));
AOI21X1 AOI21X1_48 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1558_), .C(_abc_19873_new_n1559_), .Y(_0word3_reg_31_0__14_));
AOI21X1 AOI21X1_480 ( .A(core__abc_21302_new_n2309_), .B(core__abc_21302_new_n2168__bF_buf8), .C(core__abc_21302_new_n2310_), .Y(core__0mi_reg_63_0__47_));
AOI21X1 AOI21X1_481 ( .A(core__abc_21302_new_n2312_), .B(core__abc_21302_new_n2168__bF_buf6), .C(core__abc_21302_new_n2313_), .Y(core__0mi_reg_63_0__48_));
AOI21X1 AOI21X1_482 ( .A(core__abc_21302_new_n2315_), .B(core__abc_21302_new_n2168__bF_buf4), .C(core__abc_21302_new_n2316_), .Y(core__0mi_reg_63_0__49_));
AOI21X1 AOI21X1_483 ( .A(core__abc_21302_new_n2318_), .B(core__abc_21302_new_n2168__bF_buf2), .C(core__abc_21302_new_n2319_), .Y(core__0mi_reg_63_0__50_));
AOI21X1 AOI21X1_484 ( .A(core__abc_21302_new_n2321_), .B(core__abc_21302_new_n2168__bF_buf0), .C(core__abc_21302_new_n2322_), .Y(core__0mi_reg_63_0__51_));
AOI21X1 AOI21X1_485 ( .A(core__abc_21302_new_n2324_), .B(core__abc_21302_new_n2168__bF_buf11), .C(core__abc_21302_new_n2325_), .Y(core__0mi_reg_63_0__52_));
AOI21X1 AOI21X1_486 ( .A(core__abc_21302_new_n2327_), .B(core__abc_21302_new_n2168__bF_buf9), .C(core__abc_21302_new_n2328_), .Y(core__0mi_reg_63_0__53_));
AOI21X1 AOI21X1_487 ( .A(core__abc_21302_new_n2330_), .B(core__abc_21302_new_n2168__bF_buf7), .C(core__abc_21302_new_n2331_), .Y(core__0mi_reg_63_0__54_));
AOI21X1 AOI21X1_488 ( .A(core__abc_21302_new_n2333_), .B(core__abc_21302_new_n2168__bF_buf5), .C(core__abc_21302_new_n2334_), .Y(core__0mi_reg_63_0__55_));
AOI21X1 AOI21X1_489 ( .A(core__abc_21302_new_n2336_), .B(core__abc_21302_new_n2168__bF_buf3), .C(core__abc_21302_new_n2337_), .Y(core__0mi_reg_63_0__56_));
AOI21X1 AOI21X1_49 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1210_), .C(_abc_19873_new_n1561_), .Y(_0word3_reg_31_0__15_));
AOI21X1 AOI21X1_490 ( .A(core__abc_21302_new_n2339_), .B(core__abc_21302_new_n2168__bF_buf1), .C(core__abc_21302_new_n2340_), .Y(core__0mi_reg_63_0__57_));
AOI21X1 AOI21X1_491 ( .A(core__abc_21302_new_n2342_), .B(core__abc_21302_new_n2168__bF_buf12), .C(core__abc_21302_new_n2343_), .Y(core__0mi_reg_63_0__58_));
AOI21X1 AOI21X1_492 ( .A(core__abc_21302_new_n2345_), .B(core__abc_21302_new_n2168__bF_buf10), .C(core__abc_21302_new_n2346_), .Y(core__0mi_reg_63_0__59_));
AOI21X1 AOI21X1_493 ( .A(core__abc_21302_new_n2348_), .B(core__abc_21302_new_n2168__bF_buf8), .C(core__abc_21302_new_n2349_), .Y(core__0mi_reg_63_0__60_));
AOI21X1 AOI21X1_494 ( .A(core__abc_21302_new_n2351_), .B(core__abc_21302_new_n2168__bF_buf6), .C(core__abc_21302_new_n2352_), .Y(core__0mi_reg_63_0__61_));
AOI21X1 AOI21X1_495 ( .A(core__abc_21302_new_n2354_), .B(core__abc_21302_new_n2168__bF_buf4), .C(core__abc_21302_new_n2355_), .Y(core__0mi_reg_63_0__62_));
AOI21X1 AOI21X1_496 ( .A(core__abc_21302_new_n2357_), .B(core__abc_21302_new_n2168__bF_buf2), .C(core__abc_21302_new_n2358_), .Y(core__0mi_reg_63_0__63_));
AOI21X1 AOI21X1_497 ( .A(core__abc_21302_new_n1241_), .B(core__abc_21302_new_n1232_), .C(core__abc_21302_new_n2373_), .Y(core__abc_21302_new_n2377_));
AOI21X1 AOI21X1_498 ( .A(core__abc_21302_new_n2391_), .B(core__abc_21302_new_n2378_), .C(core__abc_21302_new_n2396_), .Y(core__abc_21302_new_n2397_));
AOI21X1 AOI21X1_499 ( .A(core__abc_21302_new_n1372_), .B(core__abc_21302_new_n1359_), .C(core__abc_21302_new_n1371_), .Y(core__abc_21302_new_n2417_));
AOI21X1 AOI21X1_5 ( .A(_abc_19873_new_n1016_), .B(_abc_19873_new_n1005_), .C(_abc_19873_new_n928__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_27087_4_));
AOI21X1 AOI21X1_50 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1563_), .C(_abc_19873_new_n1564_), .Y(_0word3_reg_31_0__16_));
AOI21X1 AOI21X1_500 ( .A(core__abc_21302_new_n2412_), .B(core__abc_21302_new_n2400_), .C(core__abc_21302_new_n2418_), .Y(core__abc_21302_new_n2419_));
AOI21X1 AOI21X1_501 ( .A(core__abc_21302_new_n1467_), .B(core__abc_21302_new_n1454_), .C(core__abc_21302_new_n1466_), .Y(core__abc_21302_new_n2450_));
AOI21X1 AOI21X1_502 ( .A(core__abc_21302_new_n2445_), .B(core__abc_21302_new_n2430_), .C(core__abc_21302_new_n2451_), .Y(core__abc_21302_new_n2452_));
AOI21X1 AOI21X1_503 ( .A(core__abc_21302_new_n1509_), .B(core__abc_21302_new_n1496_), .C(core__abc_21302_new_n1508_), .Y(core__abc_21302_new_n2458_));
AOI21X1 AOI21X1_504 ( .A(core__abc_21302_new_n1558_), .B(core__abc_21302_new_n1545_), .C(core__abc_21302_new_n1557_), .Y(core__abc_21302_new_n2460_));
AOI21X1 AOI21X1_505 ( .A(core__abc_21302_new_n2423_), .B(core__abc_21302_new_n2459_), .C(core__abc_21302_new_n2464_), .Y(core__abc_21302_new_n2465_));
AOI21X1 AOI21X1_506 ( .A(core__abc_21302_new_n2420_), .B(core__abc_21302_new_n2434_), .C(core__abc_21302_new_n2466_), .Y(core__abc_21302_new_n2467_));
AOI21X1 AOI21X1_507 ( .A(core__abc_21302_new_n2470_), .B(core__abc_21302_new_n2472_), .C(core__abc_21302_new_n1243_), .Y(core__abc_21302_new_n2473_));
AOI21X1 AOI21X1_508 ( .A(core__abc_21302_new_n2473_), .B(core__abc_21302_new_n2375_), .C(core__abc_21302_new_n2474_), .Y(core__abc_21302_new_n2475_));
AOI21X1 AOI21X1_509 ( .A(core__abc_21302_new_n2476_), .B(core__abc_21302_new_n2392_), .C(core__abc_21302_new_n2394_), .Y(core__abc_21302_new_n2479_));
AOI21X1 AOI21X1_51 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1566_), .C(_abc_19873_new_n1567_), .Y(_0word3_reg_31_0__17_));
AOI21X1 AOI21X1_510 ( .A(core__abc_21302_new_n2480_), .B(core__abc_21302_new_n2486_), .C(core__abc_21302_new_n2491_), .Y(core__abc_21302_new_n2492_));
AOI21X1 AOI21X1_511 ( .A(core__abc_21302_new_n2500_), .B(core__abc_21302_new_n2493_), .C(core__abc_21302_new_n2503_), .Y(core__abc_21302_new_n2504_));
AOI21X1 AOI21X1_512 ( .A(core__abc_21302_new_n2515_), .B(core__abc_21302_new_n1235_), .C(core__abc_21302_new_n1244_), .Y(core__abc_21302_new_n2516_));
AOI21X1 AOI21X1_513 ( .A(core__abc_21302_new_n1268_), .B(core__abc_21302_new_n1254_), .C(core__abc_21302_new_n1266_), .Y(core__abc_21302_new_n2523_));
AOI21X1 AOI21X1_514 ( .A(core__abc_21302_new_n1288_), .B(core__abc_21302_new_n1276_), .C(core__abc_21302_new_n1286_), .Y(core__abc_21302_new_n2524_));
AOI21X1 AOI21X1_515 ( .A(core__abc_21302_new_n2519_), .B(core__abc_21302_new_n2522_), .C(core__abc_21302_new_n2525_), .Y(core__abc_21302_new_n2526_));
AOI21X1 AOI21X1_516 ( .A(core__abc_21302_new_n1328_), .B(core__abc_21302_new_n1329_), .C(core__abc_21302_new_n1315_), .Y(core__abc_21302_new_n2539_));
AOI21X1 AOI21X1_517 ( .A(core_v2_reg_11_), .B(core_v3_reg_11_), .C(core__abc_21302_new_n2539_), .Y(core__abc_21302_new_n2540_));
AOI21X1 AOI21X1_518 ( .A(core__abc_21302_new_n2541_), .B(core__abc_21302_new_n2529_), .C(core__abc_21302_new_n2546_), .Y(core__abc_21302_new_n2547_));
AOI21X1 AOI21X1_519 ( .A(core__abc_21302_new_n2571_), .B(core__abc_21302_new_n2570_), .C(core__abc_21302_new_n2572_), .Y(core__abc_21302_new_n2573_));
AOI21X1 AOI21X1_52 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1569_), .C(_abc_19873_new_n1570_), .Y(_0word3_reg_31_0__18_));
AOI21X1 AOI21X1_520 ( .A(core__abc_21302_new_n2576_), .B(core__abc_21302_new_n2580_), .C(core__abc_21302_new_n2583_), .Y(core__abc_21302_new_n2584_));
AOI21X1 AOI21X1_521 ( .A(core__abc_21302_new_n2595_), .B(core__abc_21302_new_n2593_), .C(core__abc_21302_new_n2596_), .Y(core__abc_21302_new_n2597_));
AOI21X1 AOI21X1_522 ( .A(core__abc_21302_new_n2607_), .B(core__abc_21302_new_n2611_), .C(core__abc_21302_new_n2612_), .Y(core__abc_21302_new_n2613_));
AOI21X1 AOI21X1_523 ( .A(core__abc_21302_new_n2615_), .B(core__abc_21302_new_n1641_), .C(core__abc_21302_new_n1651_), .Y(core__abc_21302_new_n2616_));
AOI21X1 AOI21X1_524 ( .A(core__abc_21302_new_n2610_), .B(core__abc_21302_new_n2620_), .C(core__abc_21302_new_n2622_), .Y(core__abc_21302_new_n2623_));
AOI21X1 AOI21X1_525 ( .A(core__abc_21302_new_n2627_), .B(core__abc_21302_new_n2625_), .C(core__abc_21302_new_n1512_), .Y(core__abc_21302_new_n2628_));
AOI21X1 AOI21X1_526 ( .A(core__abc_21302_new_n2630_), .B(core__abc_21302_new_n2629_), .C(core_v3_reg_27_), .Y(core__abc_21302_new_n2631_));
AOI21X1 AOI21X1_527 ( .A(core__abc_21302_new_n2512_), .B(core__abc_21302_new_n2632_), .C(core__abc_21302_new_n2635_), .Y(core__abc_21302_new_n2636_));
AOI21X1 AOI21X1_528 ( .A(core__abc_21302_new_n2360_), .B(core__abc_21302_new_n2370_), .C(core__abc_21302_new_n2645_), .Y(core__0v3_reg_63_0__0_));
AOI21X1 AOI21X1_529 ( .A(core__abc_21302_new_n2650_), .B(core__abc_21302_new_n2649_), .C(core__abc_21302_new_n2653_), .Y(core__abc_21302_new_n2654_));
AOI21X1 AOI21X1_53 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1572_), .C(_abc_19873_new_n1573_), .Y(_0word3_reg_31_0__19_));
AOI21X1 AOI21X1_530 ( .A(core__abc_21302_new_n1697_), .B(core__abc_21302_new_n1684_), .C(core__abc_21302_new_n1696_), .Y(core__abc_21302_new_n2661_));
AOI21X1 AOI21X1_531 ( .A(core__abc_21302_new_n2610_), .B(core__abc_21302_new_n2620_), .C(core__abc_21302_new_n2663_), .Y(core__abc_21302_new_n2664_));
AOI21X1 AOI21X1_532 ( .A(core__abc_21302_new_n2672_), .B(core__abc_21302_new_n2658_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n2674_));
AOI21X1 AOI21X1_533 ( .A(core__abc_21302_new_n2675_), .B(core__abc_21302_new_n2678_), .C(core__abc_21302_new_n2679_), .Y(core__0v3_reg_63_0__1_));
AOI21X1 AOI21X1_534 ( .A(core__abc_21302_new_n2710_), .B(core__abc_21302_new_n2700_), .C(core__abc_21302_new_n2673__bF_buf10), .Y(core__abc_21302_new_n2711_));
AOI21X1 AOI21X1_535 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n2713_), .C(core__abc_21302_new_n2715_), .Y(core__abc_21302_new_n2716_));
AOI21X1 AOI21X1_536 ( .A(core__abc_21302_new_n2712_), .B(core__abc_21302_new_n2716_), .C(core__abc_21302_new_n2717_), .Y(core__0v3_reg_63_0__2_));
AOI21X1 AOI21X1_537 ( .A(core__abc_21302_new_n2721_), .B(core__abc_21302_new_n2723_), .C(core__abc_21302_new_n1732_), .Y(core__abc_21302_new_n2724_));
AOI21X1 AOI21X1_538 ( .A(core__abc_21302_new_n2681_), .B(core__abc_21302_new_n2694_), .C(core__abc_21302_new_n2697_), .Y(core__abc_21302_new_n2734_));
AOI21X1 AOI21X1_539 ( .A(core__abc_21302_new_n2738_), .B(core__abc_21302_new_n2735_), .C(core__abc_21302_new_n2745_), .Y(core__abc_21302_new_n2748_));
AOI21X1 AOI21X1_54 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1575_), .C(_abc_19873_new_n1576_), .Y(_0word3_reg_31_0__20_));
AOI21X1 AOI21X1_540 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n2756_), .C(core__abc_21302_new_n2758_), .Y(core__abc_21302_new_n2759_));
AOI21X1 AOI21X1_541 ( .A(core__abc_21302_new_n2755_), .B(core__abc_21302_new_n2759_), .C(core__abc_21302_new_n2760_), .Y(core__0v3_reg_63_0__3_));
AOI21X1 AOI21X1_542 ( .A(core__abc_21302_new_n2737_), .B(core__abc_21302_new_n2736_), .C(core__abc_21302_new_n1603_), .Y(core__abc_21302_new_n2763_));
AOI21X1 AOI21X1_543 ( .A(core__abc_21302_new_n2782_), .B(core__abc_21302_new_n2784_), .C(core__abc_21302_new_n2588_), .Y(core__abc_21302_new_n2785_));
AOI21X1 AOI21X1_544 ( .A(core__abc_21302_new_n2786_), .B(core__abc_21302_new_n2787_), .C(core_v3_reg_31_), .Y(core__abc_21302_new_n2788_));
AOI21X1 AOI21X1_545 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n2792_), .C(core__abc_21302_new_n2793_), .Y(core__abc_21302_new_n2794_));
AOI21X1 AOI21X1_546 ( .A(core__abc_21302_new_n2519_), .B(core__abc_21302_new_n1256_), .C(core__abc_21302_new_n1254_), .Y(core__abc_21302_new_n2805_));
AOI21X1 AOI21X1_547 ( .A(core__abc_21302_new_n2814_), .B(core__abc_21302_new_n2722_), .C(core__abc_21302_new_n2820_), .Y(core__abc_21302_new_n2821_));
AOI21X1 AOI21X1_548 ( .A(core__abc_21302_new_n2818_), .B(core__abc_21302_new_n2824_), .C(core__abc_21302_new_n2827_), .Y(core__abc_21302_new_n2828_));
AOI21X1 AOI21X1_549 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n2833_), .C(core__abc_21302_new_n2834_), .Y(core__abc_21302_new_n2835_));
AOI21X1 AOI21X1_55 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1578_), .C(_abc_19873_new_n1579_), .Y(_0word3_reg_31_0__21_));
AOI21X1 AOI21X1_550 ( .A(core__abc_21302_new_n2767_), .B(core__abc_21302_new_n2841_), .C(core__abc_21302_new_n2840_), .Y(core__abc_21302_new_n2842_));
AOI21X1 AOI21X1_551 ( .A(core__abc_21302_new_n2811_), .B(core__abc_21302_new_n2808_), .C(core__abc_21302_new_n2779_), .Y(core__abc_21302_new_n2861_));
AOI21X1 AOI21X1_552 ( .A(core__abc_21302_new_n2861_), .B(core__abc_21302_new_n2780_), .C(core__abc_21302_new_n2860_), .Y(core__abc_21302_new_n2862_));
AOI21X1 AOI21X1_553 ( .A(core__abc_21302_new_n2863_), .B(core__abc_21302_new_n2871_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n2872_));
AOI21X1 AOI21X1_554 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n2874_), .C(core__abc_21302_new_n2875_), .Y(core__abc_21302_new_n2876_));
AOI21X1 AOI21X1_555 ( .A(core__abc_21302_new_n2873_), .B(core__abc_21302_new_n2876_), .C(core__abc_21302_new_n2877_), .Y(core__0v3_reg_63_0__6_));
AOI21X1 AOI21X1_556 ( .A(core__abc_21302_new_n2825_), .B(core__abc_21302_new_n2897_), .C(core__abc_21302_new_n2899_), .Y(core__abc_21302_new_n2900_));
AOI21X1 AOI21X1_557 ( .A(core_key_71_), .B(core__abc_21302_new_n2639__bF_buf5), .C(core__abc_21302_new_n2910_), .Y(core__abc_21302_new_n2911_));
AOI21X1 AOI21X1_558 ( .A(core__abc_21302_new_n2881_), .B(core__abc_21302_new_n2887_), .C(core__abc_21302_new_n2855_), .Y(core__abc_21302_new_n2917_));
AOI21X1 AOI21X1_559 ( .A(core__abc_21302_new_n2890_), .B(core__abc_21302_new_n2886_), .C(core__abc_21302_new_n2917_), .Y(core__abc_21302_new_n2918_));
AOI21X1 AOI21X1_56 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1581_), .C(_abc_19873_new_n1582_), .Y(_0word3_reg_31_0__22_));
AOI21X1 AOI21X1_560 ( .A(core__abc_21302_new_n2889_), .B(core__abc_21302_new_n2879_), .C(core__abc_21302_new_n1648_), .Y(core__abc_21302_new_n2924_));
AOI21X1 AOI21X1_561 ( .A(core__abc_21302_new_n2505_), .B(core__abc_21302_new_n2927_), .C(core__abc_21302_new_n2926_), .Y(core__abc_21302_new_n2928_));
AOI21X1 AOI21X1_562 ( .A(core__abc_21302_new_n2931_), .B(core__abc_21302_new_n2930_), .C(core__abc_21302_new_n2932_), .Y(core__abc_21302_new_n2933_));
AOI21X1 AOI21X1_563 ( .A(core__abc_21302_new_n2947_), .B(core__abc_21302_new_n2956_), .C(core__abc_21302_new_n2673__bF_buf6), .Y(core__abc_21302_new_n2957_));
AOI21X1 AOI21X1_564 ( .A(core__abc_21302_new_n2961_), .B(core__abc_21302_new_n2369__bF_buf7), .C(core__abc_21302_new_n2962_), .Y(core__0v3_reg_63_0__8_));
AOI21X1 AOI21X1_565 ( .A(core__abc_21302_new_n2818_), .B(core__abc_21302_new_n2824_), .C(core__abc_21302_new_n2982_), .Y(core__abc_21302_new_n2983_));
AOI21X1 AOI21X1_566 ( .A(core__abc_21302_new_n1788_), .B(core__abc_21302_new_n1776_), .C(core__abc_21302_new_n1787_), .Y(core__abc_21302_new_n2985_));
AOI21X1 AOI21X1_567 ( .A(core_key_73_), .B(core__abc_21302_new_n2639__bF_buf4), .C(core__abc_21302_new_n2995_), .Y(core__abc_21302_new_n2996_));
AOI21X1 AOI21X1_568 ( .A(core__abc_21302_new_n2977_), .B(core__abc_21302_new_n2975_), .C(core__abc_21302_new_n3003_), .Y(core__abc_21302_new_n3004_));
AOI21X1 AOI21X1_569 ( .A(core__abc_21302_new_n3009_), .B(core__abc_21302_new_n1659_), .C(core__abc_21302_new_n1670_), .Y(core__abc_21302_new_n3010_));
AOI21X1 AOI21X1_57 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1365_), .C(_abc_19873_new_n1584_), .Y(_0word3_reg_31_0__23_));
AOI21X1 AOI21X1_570 ( .A(core__abc_21302_new_n2935_), .B(core__abc_21302_new_n3008_), .C(core__abc_21302_new_n3011_), .Y(core__abc_21302_new_n3012_));
AOI21X1 AOI21X1_571 ( .A(core__abc_21302_new_n3025_), .B(core__abc_21302_new_n3034_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n3035_));
AOI21X1 AOI21X1_572 ( .A(core__abc_21302_new_n3039_), .B(core__abc_21302_new_n2369__bF_buf3), .C(core__abc_21302_new_n3040_), .Y(core__0v3_reg_63_0__10_));
AOI21X1 AOI21X1_573 ( .A(core__abc_21302_new_n1814_), .B(core__abc_21302_new_n1801_), .C(core__abc_21302_new_n1813_), .Y(core__abc_21302_new_n3065_));
AOI21X1 AOI21X1_574 ( .A(core__abc_21302_new_n3062_), .B(core__abc_21302_new_n3074_), .C(core__abc_21302_new_n2673__bF_buf4), .Y(core__abc_21302_new_n3075_));
AOI21X1 AOI21X1_575 ( .A(core_key_75_), .B(core__abc_21302_new_n2639__bF_buf3), .C(core__abc_21302_new_n3078_), .Y(core__abc_21302_new_n3079_));
AOI21X1 AOI21X1_576 ( .A(core__abc_21302_new_n3076_), .B(core__abc_21302_new_n3079_), .C(core__abc_21302_new_n3080_), .Y(core__0v3_reg_63_0__11_));
AOI21X1 AOI21X1_577 ( .A(core__abc_21302_new_n1693_), .B(core__abc_21302_new_n1681_), .C(core__abc_21302_new_n1692_), .Y(core__abc_21302_new_n3092_));
AOI21X1 AOI21X1_578 ( .A(core__abc_21302_new_n2935_), .B(core__abc_21302_new_n3095_), .C(core__abc_21302_new_n3093_), .Y(core__abc_21302_new_n3099_));
AOI21X1 AOI21X1_579 ( .A(core__abc_21302_new_n3110_), .B(core__abc_21302_new_n3121_), .C(core__abc_21302_new_n2673__bF_buf3), .Y(core__abc_21302_new_n3122_));
AOI21X1 AOI21X1_58 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1586_), .C(_abc_19873_new_n1587_), .Y(_0word3_reg_31_0__24_));
AOI21X1 AOI21X1_580 ( .A(core__abc_21302_new_n3126_), .B(core__abc_21302_new_n2369__bF_buf7), .C(core__abc_21302_new_n3127_), .Y(core__0v3_reg_63_0__12_));
AOI21X1 AOI21X1_581 ( .A(core__abc_21302_new_n1826_), .B(core__abc_21302_new_n1839_), .C(core__abc_21302_new_n3157_), .Y(core__abc_21302_new_n3158_));
AOI21X1 AOI21X1_582 ( .A(core__abc_21302_new_n3155_), .B(core__abc_21302_new_n3160_), .C(core__abc_21302_new_n3158_), .Y(core__abc_21302_new_n3161_));
AOI21X1 AOI21X1_583 ( .A(core__abc_21302_new_n3154_), .B(core__abc_21302_new_n3167_), .C(core__abc_21302_new_n2673__bF_buf2), .Y(core__abc_21302_new_n3168_));
AOI21X1 AOI21X1_584 ( .A(core__abc_21302_new_n3172_), .B(core__abc_21302_new_n2369__bF_buf5), .C(core__abc_21302_new_n3173_), .Y(core__0v3_reg_63_0__13_));
AOI21X1 AOI21X1_585 ( .A(core__abc_21302_new_n3097_), .B(core__abc_21302_new_n3180_), .C(core__abc_21302_new_n3178_), .Y(core__abc_21302_new_n3181_));
AOI21X1 AOI21X1_586 ( .A(core__abc_21302_new_n3188_), .B(core__abc_21302_new_n3102_), .C(core__abc_21302_new_n2528_), .Y(core__abc_21302_new_n3189_));
AOI21X1 AOI21X1_587 ( .A(core__abc_21302_new_n1852_), .B(core__abc_21302_new_n1865_), .C(core__abc_21302_new_n3209_), .Y(core__abc_21302_new_n3210_));
AOI21X1 AOI21X1_588 ( .A(core__abc_21302_new_n3205_), .B(core__abc_21302_new_n3215_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n3216_));
AOI21X1 AOI21X1_589 ( .A(core__abc_21302_new_n3220_), .B(core__abc_21302_new_n2369__bF_buf3), .C(core__abc_21302_new_n3221_), .Y(core__0v3_reg_63_0__14_));
AOI21X1 AOI21X1_59 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1589_), .C(_abc_19873_new_n1590_), .Y(_0word3_reg_31_0__25_));
AOI21X1 AOI21X1_590 ( .A(core__abc_21302_new_n3199_), .B(core__abc_21302_new_n1726_), .C(core__abc_21302_new_n1739_), .Y(core__abc_21302_new_n3239_));
AOI21X1 AOI21X1_591 ( .A(core__abc_21302_new_n1865_), .B(core__abc_21302_new_n1852_), .C(core__abc_21302_new_n1864_), .Y(core__abc_21302_new_n3247_));
AOI21X1 AOI21X1_592 ( .A(core__abc_21302_new_n3245_), .B(core__abc_21302_new_n3256_), .C(core__abc_21302_new_n2673__bF_buf0), .Y(core__abc_21302_new_n3257_));
AOI21X1 AOI21X1_593 ( .A(core__abc_21302_new_n3258_), .B(core__abc_21302_new_n3262_), .C(core__abc_21302_new_n3263_), .Y(core__0v3_reg_63_0__15_));
AOI21X1 AOI21X1_594 ( .A(core__abc_21302_new_n3146_), .B(core__abc_21302_new_n3278_), .C(core__abc_21302_new_n3148_), .Y(core__abc_21302_new_n3279_));
AOI21X1 AOI21X1_595 ( .A(core__abc_21302_new_n1739_), .B(core__abc_21302_new_n1727_), .C(core__abc_21302_new_n1738_), .Y(core__abc_21302_new_n3290_));
AOI21X1 AOI21X1_596 ( .A(core__abc_21302_new_n3093_), .B(core__abc_21302_new_n3287_), .C(core__abc_21302_new_n3291_), .Y(core__abc_21302_new_n3292_));
AOI21X1 AOI21X1_597 ( .A(core__abc_21302_new_n2926_), .B(core__abc_21302_new_n3289_), .C(core__abc_21302_new_n3293_), .Y(core__abc_21302_new_n3294_));
AOI21X1 AOI21X1_598 ( .A(core__abc_21302_new_n3315_), .B(core__abc_21302_new_n3314_), .C(core__abc_21302_new_n3311_), .Y(core__abc_21302_new_n3316_));
AOI21X1 AOI21X1_599 ( .A(core__abc_21302_new_n3253_), .B(core__abc_21302_new_n3312_), .C(core__abc_21302_new_n3313_), .Y(core__abc_21302_new_n3319_));
AOI21X1 AOI21X1_6 ( .A(_abc_19873_new_n1027_), .B(_abc_19873_new_n1037_), .C(_abc_19873_new_n928__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_27087_5_));
AOI21X1 AOI21X1_60 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1420_), .C(_abc_19873_new_n1592_), .Y(_0word3_reg_31_0__26_));
AOI21X1 AOI21X1_600 ( .A(core__abc_21302_new_n3326_), .B(core__abc_21302_new_n3265_), .C(core__abc_21302_new_n1185__bF_buf12), .Y(core__0v3_reg_63_0__16_));
AOI21X1 AOI21X1_601 ( .A(core__abc_21302_new_n2505_), .B(core__abc_21302_new_n3330_), .C(core__abc_21302_new_n3329_), .Y(core__abc_21302_new_n3331_));
AOI21X1 AOI21X1_602 ( .A(core__abc_21302_new_n3307_), .B(core__abc_21302_new_n3304_), .C(core__abc_21302_new_n3346_), .Y(core__abc_21302_new_n3349_));
AOI21X1 AOI21X1_603 ( .A(core__abc_21302_new_n1891_), .B(core__abc_21302_new_n1878_), .C(core__abc_21302_new_n1890_), .Y(core__abc_21302_new_n3352_));
AOI21X1 AOI21X1_604 ( .A(core__abc_21302_new_n3351_), .B(core__abc_21302_new_n3360_), .C(core__abc_21302_new_n2673__bF_buf10), .Y(core__abc_21302_new_n3361_));
AOI21X1 AOI21X1_605 ( .A(core__abc_21302_new_n3365_), .B(core__abc_21302_new_n2369__bF_buf7), .C(core__abc_21302_new_n3366_), .Y(core__0v3_reg_63_0__17_));
AOI21X1 AOI21X1_606 ( .A(core__abc_21302_new_n3370_), .B(core__abc_21302_new_n3373_), .C(core__abc_21302_new_n3372_), .Y(core__abc_21302_new_n3374_));
AOI21X1 AOI21X1_607 ( .A(core__abc_21302_new_n3296_), .B(core__abc_21302_new_n3378_), .C(core__abc_21302_new_n3381_), .Y(core__abc_21302_new_n3382_));
AOI21X1 AOI21X1_608 ( .A(core__abc_21302_new_n2548_), .B(core__abc_21302_new_n3385_), .C(core__abc_21302_new_n2571_), .Y(core__abc_21302_new_n3386_));
AOI21X1 AOI21X1_609 ( .A(core__abc_21302_new_n3396_), .B(core__abc_21302_new_n3407_), .C(core__abc_21302_new_n2673__bF_buf9), .Y(core__abc_21302_new_n3408_));
AOI21X1 AOI21X1_61 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1430_), .C(_abc_19873_new_n1594_), .Y(_0word3_reg_31_0__27_));
AOI21X1 AOI21X1_610 ( .A(core__abc_21302_new_n3412_), .B(core__abc_21302_new_n2369__bF_buf5), .C(core__abc_21302_new_n3413_), .Y(core__0v3_reg_63_0__18_));
AOI21X1 AOI21X1_611 ( .A(core__abc_21302_new_n3417_), .B(core__abc_21302_new_n3419_), .C(core__abc_21302_new_n3428_), .Y(core__abc_21302_new_n3429_));
AOI21X1 AOI21X1_612 ( .A(core__abc_21302_new_n3430_), .B(core__abc_21302_new_n3431_), .C(core__abc_21302_new_n3432_), .Y(core__abc_21302_new_n3433_));
AOI21X1 AOI21X1_613 ( .A(core__abc_21302_new_n3444_), .B(core__abc_21302_new_n3445_), .C(core_v3_reg_46_), .Y(core__abc_21302_new_n3446_));
AOI21X1 AOI21X1_614 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n3451_), .C(core__abc_21302_new_n3453_), .Y(core__abc_21302_new_n3454_));
AOI21X1 AOI21X1_615 ( .A(core__abc_21302_new_n3417_), .B(core__abc_21302_new_n3419_), .C(core__abc_21302_new_n3432_), .Y(core__abc_21302_new_n3462_));
AOI21X1 AOI21X1_616 ( .A(core__abc_21302_new_n3344_), .B(core__abc_21302_new_n3342_), .C(core__abc_21302_new_n3305_), .Y(core__abc_21302_new_n3465_));
AOI21X1 AOI21X1_617 ( .A(core__abc_21302_new_n3285_), .B(core__abc_21302_new_n3467_), .C(core__abc_21302_new_n3464_), .Y(core__abc_21302_new_n3468_));
AOI21X1 AOI21X1_618 ( .A(core__abc_21302_new_n1785_), .B(core__abc_21302_new_n1772_), .C(core__abc_21302_new_n1784_), .Y(core__abc_21302_new_n3471_));
AOI21X1 AOI21X1_619 ( .A(core__abc_21302_new_n3296_), .B(core__abc_21302_new_n3474_), .C(core__abc_21302_new_n3472_), .Y(core__abc_21302_new_n3475_));
AOI21X1 AOI21X1_62 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1596_), .C(_abc_19873_new_n1597_), .Y(_0word3_reg_31_0__28_));
AOI21X1 AOI21X1_620 ( .A(core__abc_21302_new_n2548_), .B(core__abc_21302_new_n2565_), .C(core__abc_21302_new_n3477_), .Y(core__abc_21302_new_n3478_));
AOI21X1 AOI21X1_621 ( .A(core__abc_21302_new_n3491_), .B(core__abc_21302_new_n3488_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n3492_));
AOI21X1 AOI21X1_622 ( .A(core__abc_21302_new_n3493_), .B(core__abc_21302_new_n3496_), .C(core__abc_21302_new_n3497_), .Y(core__0v3_reg_63_0__20_));
AOI21X1 AOI21X1_623 ( .A(core__abc_21302_new_n3501_), .B(core__abc_21302_new_n1797_), .C(core__abc_21302_new_n1796_), .Y(core__abc_21302_new_n3502_));
AOI21X1 AOI21X1_624 ( .A(core__abc_21302_new_n3506_), .B(core__abc_21302_new_n3503_), .C(core__abc_21302_new_n3516_), .Y(core__abc_21302_new_n3517_));
AOI21X1 AOI21X1_625 ( .A(core__abc_21302_new_n3512_), .B(core__abc_21302_new_n3515_), .C(core__abc_21302_new_n3518_), .Y(core__abc_21302_new_n3519_));
AOI21X1 AOI21X1_626 ( .A(core__abc_21302_new_n3523_), .B(core__abc_21302_new_n2510_), .C(core__abc_21302_new_n2673__bF_buf6), .Y(core__abc_21302_new_n3524_));
AOI21X1 AOI21X1_627 ( .A(core__abc_21302_new_n3528_), .B(core__abc_21302_new_n2369__bF_buf0), .C(core__abc_21302_new_n3529_), .Y(core__0v3_reg_63_0__21_));
AOI21X1 AOI21X1_628 ( .A(core__abc_21302_new_n3533_), .B(core__abc_21302_new_n3483_), .C(core__abc_21302_new_n3517_), .Y(core__abc_21302_new_n3534_));
AOI21X1 AOI21X1_629 ( .A(core__abc_21302_new_n3565_), .B(core__abc_21302_new_n2653_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n3566_));
AOI21X1 AOI21X1_63 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1470_), .C(_abc_19873_new_n1599_), .Y(_0word3_reg_31_0__29_));
AOI21X1 AOI21X1_630 ( .A(core__abc_21302_new_n3570_), .B(core__abc_21302_new_n2369__bF_buf6), .C(core__abc_21302_new_n3571_), .Y(core__0v3_reg_63_0__22_));
AOI21X1 AOI21X1_631 ( .A(core__abc_21302_new_n3579_), .B(core__abc_21302_new_n3577_), .C(core__abc_21302_new_n3587_), .Y(core__abc_21302_new_n3588_));
AOI21X1 AOI21X1_632 ( .A(core__abc_21302_new_n3595_), .B(core__abc_21302_new_n3573_), .C(core__abc_21302_new_n2673__bF_buf4), .Y(core__abc_21302_new_n3596_));
AOI21X1 AOI21X1_633 ( .A(core__abc_21302_new_n3597_), .B(core__abc_21302_new_n3601_), .C(core__abc_21302_new_n3602_), .Y(core__0v3_reg_63_0__23_));
AOI21X1 AOI21X1_634 ( .A(core__abc_21302_new_n3610_), .B(core__abc_21302_new_n3574_), .C(core__abc_21302_new_n3591_), .Y(core__abc_21302_new_n3611_));
AOI21X1 AOI21X1_635 ( .A(core__abc_21302_new_n3285_), .B(core__abc_21302_new_n3615_), .C(core__abc_21302_new_n3612_), .Y(core__abc_21302_new_n3616_));
AOI21X1 AOI21X1_636 ( .A(core__abc_21302_new_n1834_), .B(core__abc_21302_new_n1820_), .C(core__abc_21302_new_n1833_), .Y(core__abc_21302_new_n3623_));
AOI21X1 AOI21X1_637 ( .A(core__abc_21302_new_n3296_), .B(core__abc_21302_new_n3621_), .C(core__abc_21302_new_n3625_), .Y(core__abc_21302_new_n3626_));
AOI21X1 AOI21X1_638 ( .A(core__abc_21302_new_n2548_), .B(core__abc_21302_new_n3633_), .C(core__abc_21302_new_n3632_), .Y(core__abc_21302_new_n3636_));
AOI21X1 AOI21X1_639 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n3649_), .C(core__abc_21302_new_n3650_), .Y(core__abc_21302_new_n3651_));
AOI21X1 AOI21X1_64 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1601_), .C(_abc_19873_new_n1602_), .Y(_0word3_reg_31_0__30_));
AOI21X1 AOI21X1_640 ( .A(core__abc_21302_new_n3678_), .B(core__abc_21302_new_n2775_), .C(core__abc_21302_new_n2673__bF_buf3), .Y(core__abc_21302_new_n3679_));
AOI21X1 AOI21X1_641 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n3681_), .C(core__abc_21302_new_n3683_), .Y(core__abc_21302_new_n3684_));
AOI21X1 AOI21X1_642 ( .A(core__abc_21302_new_n3680_), .B(core__abc_21302_new_n3684_), .C(core__abc_21302_new_n3685_), .Y(core__0v3_reg_63_0__25_));
AOI21X1 AOI21X1_643 ( .A(core__abc_21302_new_n3630_), .B(core__abc_21302_new_n3695_), .C(core__abc_21302_new_n3697_), .Y(core__abc_21302_new_n3712_));
AOI21X1 AOI21X1_644 ( .A(core__abc_21302_new_n3722_), .B(core__abc_21302_new_n2369__bF_buf6), .C(core__abc_21302_new_n3723_), .Y(core__0v3_reg_63_0__26_));
AOI21X1 AOI21X1_645 ( .A(core__abc_21302_new_n3700_), .B(core__abc_21302_new_n3730_), .C(core__abc_21302_new_n1887_), .Y(core__abc_21302_new_n3745_));
AOI21X1 AOI21X1_646 ( .A(core__abc_21302_new_n3751_), .B(core__abc_21302_new_n2854_), .C(core__abc_21302_new_n2673__bF_buf2), .Y(core__abc_21302_new_n3752_));
AOI21X1 AOI21X1_647 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n3754_), .C(core__abc_21302_new_n3755_), .Y(core__abc_21302_new_n3756_));
AOI21X1 AOI21X1_648 ( .A(core__abc_21302_new_n3753_), .B(core__abc_21302_new_n3756_), .C(core__abc_21302_new_n3757_), .Y(core__0v3_reg_63_0__27_));
AOI21X1 AOI21X1_649 ( .A(core__abc_21302_new_n3733_), .B(core__abc_21302_new_n3731_), .C(core__abc_21302_new_n3742_), .Y(core__abc_21302_new_n3762_));
AOI21X1 AOI21X1_65 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1505_), .C(_abc_19873_new_n1604_), .Y(_0word3_reg_31_0__31_));
AOI21X1 AOI21X1_650 ( .A(core__abc_21302_new_n3726_), .B(core__abc_21302_new_n3743_), .C(core__abc_21302_new_n3762_), .Y(core__abc_21302_new_n3763_));
AOI21X1 AOI21X1_651 ( .A(core__abc_21302_new_n3697_), .B(core__abc_21302_new_n3769_), .C(core__abc_21302_new_n3771_), .Y(core__abc_21302_new_n3772_));
AOI21X1 AOI21X1_652 ( .A(core__abc_21302_new_n3783_), .B(core__abc_21302_new_n3784_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n3785_));
AOI21X1 AOI21X1_653 ( .A(core__abc_21302_new_n3788_), .B(core__abc_21302_new_n3759_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v3_reg_63_0__28_));
AOI21X1 AOI21X1_654 ( .A(core__abc_21302_new_n3774_), .B(core__abc_21302_new_n3778_), .C(core__abc_21302_new_n3780_), .Y(core__abc_21302_new_n3790_));
AOI21X1 AOI21X1_655 ( .A(core__abc_21302_new_n2376_), .B(core__abc_21302_new_n2377_), .C(core__abc_21302_new_n2478_), .Y(core__abc_21302_new_n3794_));
AOI21X1 AOI21X1_656 ( .A(core__abc_21302_new_n3795_), .B(core__abc_21302_new_n2419_), .C(core__abc_21302_new_n2497_), .Y(core__abc_21302_new_n3796_));
AOI21X1 AOI21X1_657 ( .A(core__abc_21302_new_n3797_), .B(core__abc_21302_new_n3294_), .C(core__abc_21302_new_n3628_), .Y(core__abc_21302_new_n3798_));
AOI21X1 AOI21X1_658 ( .A(core__abc_21302_new_n3800_), .B(core__abc_21302_new_n3772_), .C(core__abc_21302_new_n3803_), .Y(core__abc_21302_new_n3804_));
AOI21X1 AOI21X1_659 ( .A(core__abc_21302_new_n3792_), .B(core__abc_21302_new_n3793_), .C(core__abc_21302_new_n3804_), .Y(core__abc_21302_new_n3805_));
AOI21X1 AOI21X1_66 ( .A(_abc_19873_new_n1606_), .B(_abc_19873_new_n1524__bF_buf14), .C(_abc_19873_new_n1607_), .Y(_0word2_reg_31_0__0_));
AOI21X1 AOI21X1_660 ( .A(core__abc_21302_new_n3808_), .B(core__abc_21302_new_n1522_), .C(core__abc_21302_new_n3806_), .Y(core__abc_21302_new_n3814_));
AOI21X1 AOI21X1_661 ( .A(core__abc_21302_new_n3805_), .B(core__abc_21302_new_n3791_), .C(core__abc_21302_new_n3816_), .Y(core__abc_21302_new_n3817_));
AOI21X1 AOI21X1_662 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n3824_), .C(core__abc_21302_new_n3825_), .Y(core__abc_21302_new_n3826_));
AOI21X1 AOI21X1_663 ( .A(core__abc_21302_new_n3773_), .B(core__abc_21302_new_n3802_), .C(core__abc_21302_new_n3832_), .Y(core__abc_21302_new_n3833_));
AOI21X1 AOI21X1_664 ( .A(core__abc_21302_new_n3843_), .B(core__abc_21302_new_n2597_), .C(core__abc_21302_new_n3842_), .Y(core__abc_21302_new_n3844_));
AOI21X1 AOI21X1_665 ( .A(core__abc_21302_new_n3864_), .B(core__abc_21302_new_n3857_), .C(core__abc_21302_new_n3854_), .Y(core__abc_21302_new_n3865_));
AOI21X1 AOI21X1_666 ( .A(core__abc_21302_new_n3874_), .B(core__abc_21302_new_n2369__bF_buf0), .C(core__abc_21302_new_n3875_), .Y(core__0v3_reg_63_0__30_));
AOI21X1 AOI21X1_667 ( .A(core__abc_21302_new_n3899_), .B(core__abc_21302_new_n3022_), .C(core__abc_21302_new_n2673__bF_buf0), .Y(core__abc_21302_new_n3900_));
AOI21X1 AOI21X1_668 ( .A(core__abc_21302_new_n3901_), .B(core__abc_21302_new_n3905_), .C(core__abc_21302_new_n3906_), .Y(core__0v3_reg_63_0__31_));
AOI21X1 AOI21X1_669 ( .A(core__abc_21302_new_n3086_), .B(core__abc_21302_new_n3274_), .C(core__abc_21302_new_n3283_), .Y(core__abc_21302_new_n3909_));
AOI21X1 AOI21X1_67 ( .A(_abc_19873_new_n1609_), .B(_abc_19873_new_n1524__bF_buf12), .C(_abc_19873_new_n1610_), .Y(_0word2_reg_31_0__1_));
AOI21X1 AOI21X1_670 ( .A(core__abc_21302_new_n3275_), .B(core__abc_21302_new_n3909_), .C(core__abc_21302_new_n3912_), .Y(core__abc_21302_new_n3913_));
AOI21X1 AOI21X1_671 ( .A(core__abc_21302_new_n3764_), .B(core__abc_21302_new_n3911_), .C(core__abc_21302_new_n3918_), .Y(core__abc_21302_new_n3919_));
AOI21X1 AOI21X1_672 ( .A(core__abc_21302_new_n3935_), .B(core__abc_21302_new_n3934_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n3936_));
AOI21X1 AOI21X1_673 ( .A(core__abc_21302_new_n3940_), .B(core__abc_21302_new_n3908_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0v3_reg_63_0__32_));
AOI21X1 AOI21X1_674 ( .A(core__abc_21302_new_n3967_), .B(core__abc_21302_new_n3942_), .C(core__abc_21302_new_n1185__bF_buf6), .Y(core__0v3_reg_63_0__33_));
AOI21X1 AOI21X1_675 ( .A(core__abc_21302_new_n3999_), .B(core__abc_21302_new_n3969_), .C(core__abc_21302_new_n1185__bF_buf5), .Y(core__0v3_reg_63_0__34_));
AOI21X1 AOI21X1_676 ( .A(core__abc_21302_new_n4021_), .B(core__abc_21302_new_n3201_), .C(core__abc_21302_new_n2673__bF_buf8), .Y(core__abc_21302_new_n4022_));
AOI21X1 AOI21X1_677 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n4024_), .C(core__abc_21302_new_n4026_), .Y(core__abc_21302_new_n4027_));
AOI21X1 AOI21X1_678 ( .A(core__abc_21302_new_n4023_), .B(core__abc_21302_new_n4027_), .C(core__abc_21302_new_n4028_), .Y(core__0v3_reg_63_0__35_));
AOI21X1 AOI21X1_679 ( .A(core__abc_21302_new_n4010_), .B(core__abc_21302_new_n4013_), .C(core__abc_21302_new_n4016_), .Y(core__abc_21302_new_n4034_));
AOI21X1 AOI21X1_68 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n952_), .C(_abc_19873_new_n1612_), .Y(_0word2_reg_31_0__2_));
AOI21X1 AOI21X1_680 ( .A(core__abc_21302_new_n4017_), .B(core__abc_21302_new_n4033_), .C(core__abc_21302_new_n4034_), .Y(core__abc_21302_new_n4035_));
AOI21X1 AOI21X1_681 ( .A(core__abc_21302_new_n4060_), .B(core__abc_21302_new_n4030_), .C(core__abc_21302_new_n1185__bF_buf4), .Y(core__0v3_reg_63_0__36_));
AOI21X1 AOI21X1_682 ( .A(core__abc_21302_new_n4045_), .B(core__abc_21302_new_n4048_), .C(core__abc_21302_new_n1619_), .Y(core__abc_21302_new_n4067_));
AOI21X1 AOI21X1_683 ( .A(core__abc_21302_new_n4071_), .B(core__abc_21302_new_n4074_), .C(core__abc_21302_new_n4065_), .Y(core__abc_21302_new_n4077_));
AOI21X1 AOI21X1_684 ( .A(core__abc_21302_new_n4084_), .B(core__abc_21302_new_n4082_), .C(core__abc_21302_new_n2673__bF_buf6), .Y(core__abc_21302_new_n4085_));
AOI21X1 AOI21X1_685 ( .A(core__abc_21302_new_n4088_), .B(core__abc_21302_new_n4062_), .C(core__abc_21302_new_n1185__bF_buf3), .Y(core__0v3_reg_63_0__37_));
AOI21X1 AOI21X1_686 ( .A(core__abc_21302_new_n2378_), .B(core__abc_21302_new_n2477_), .C(core__abc_21302_new_n2392_), .Y(core__abc_21302_new_n4096_));
AOI21X1 AOI21X1_687 ( .A(core__abc_21302_new_n4045_), .B(core__abc_21302_new_n2604_), .C(core__abc_21302_new_n2617_), .Y(core__abc_21302_new_n4100_));
AOI21X1 AOI21X1_688 ( .A(core__abc_21302_new_n4119_), .B(core__abc_21302_new_n4118_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n4120_));
AOI21X1 AOI21X1_689 ( .A(core__abc_21302_new_n4123_), .B(core__abc_21302_new_n4090_), .C(core__abc_21302_new_n1185__bF_buf2), .Y(core__0v3_reg_63_0__38_));
AOI21X1 AOI21X1_69 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1614_), .C(_abc_19873_new_n1615_), .Y(_0word2_reg_31_0__3_));
AOI21X1 AOI21X1_690 ( .A(core__abc_21302_new_n4131_), .B(core__abc_21302_new_n4132_), .C(core__abc_21302_new_n2582_), .Y(core__abc_21302_new_n4136_));
AOI21X1 AOI21X1_691 ( .A(core__abc_21302_new_n4128_), .B(core__abc_21302_new_n4129_), .C(core_v3_reg_23_), .Y(core__abc_21302_new_n4137_));
AOI21X1 AOI21X1_692 ( .A(core__abc_21302_new_n4114_), .B(core__abc_21302_new_n4111_), .C(core__abc_21302_new_n4139_), .Y(core__abc_21302_new_n4141_));
AOI21X1 AOI21X1_693 ( .A(core__abc_21302_new_n4146_), .B(core__abc_21302_new_n4150_), .C(core__abc_21302_new_n4151_), .Y(core__0v3_reg_63_0__39_));
AOI21X1 AOI21X1_694 ( .A(core__abc_21302_new_n4138_), .B(core__abc_21302_new_n4134_), .C(core__abc_21302_new_n4112_), .Y(core__abc_21302_new_n4155_));
AOI21X1 AOI21X1_695 ( .A(core__abc_21302_new_n3893_), .B(core__abc_21302_new_n3892_), .C(core__abc_21302_new_n3894_), .Y(core__abc_21302_new_n4164_));
AOI21X1 AOI21X1_696 ( .A(core__abc_21302_new_n3612_), .B(core__abc_21302_new_n4162_), .C(core__abc_21302_new_n4169_), .Y(core__abc_21302_new_n4170_));
AOI21X1 AOI21X1_697 ( .A(core__abc_21302_new_n4170_), .B(core__abc_21302_new_n4163_), .C(core__abc_21302_new_n4171_), .Y(core__abc_21302_new_n4172_));
AOI21X1 AOI21X1_698 ( .A(core__abc_21302_new_n4188_), .B(core__abc_21302_new_n4153_), .C(core__abc_21302_new_n1185__bF_buf1), .Y(core__0v3_reg_63_0__40_));
AOI21X1 AOI21X1_699 ( .A(core__abc_21302_new_n4174_), .B(core__abc_21302_new_n4196_), .C(core__abc_21302_new_n1662_), .Y(core__abc_21302_new_n4197_));
AOI21X1 AOI21X1_7 ( .A(_abc_19873_new_n1057_), .B(_abc_19873_new_n1047_), .C(_abc_19873_new_n928__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_27087_6_));
AOI21X1 AOI21X1_70 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1617_), .C(_abc_19873_new_n1618_), .Y(_0word2_reg_31_0__4_));
AOI21X1 AOI21X1_700 ( .A(core__abc_21302_new_n4210_), .B(core__abc_21302_new_n4209_), .C(core__abc_21302_new_n2673__bF_buf3), .Y(core__abc_21302_new_n4211_));
AOI21X1 AOI21X1_701 ( .A(core__abc_21302_new_n4215_), .B(core__abc_21302_new_n4190_), .C(core__abc_21302_new_n1185__bF_buf0), .Y(core__0v3_reg_63_0__41_));
AOI21X1 AOI21X1_702 ( .A(core__abc_21302_new_n4242_), .B(core__abc_21302_new_n4240_), .C(core__abc_21302_new_n2673__bF_buf2), .Y(core__abc_21302_new_n4243_));
AOI21X1 AOI21X1_703 ( .A(core__abc_21302_new_n4246_), .B(core__abc_21302_new_n4217_), .C(core__abc_21302_new_n1185__bF_buf13), .Y(core__0v3_reg_63_0__42_));
AOI21X1 AOI21X1_704 ( .A(core__abc_21302_new_n4264_), .B(core__abc_21302_new_n3560_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n4265_));
AOI21X1 AOI21X1_705 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n4267_), .C(core__abc_21302_new_n4269_), .Y(core__abc_21302_new_n4270_));
AOI21X1 AOI21X1_706 ( .A(core__abc_21302_new_n4266_), .B(core__abc_21302_new_n4270_), .C(core__abc_21302_new_n4271_), .Y(core__0v3_reg_63_0__43_));
AOI21X1 AOI21X1_707 ( .A(core__abc_21302_new_n4256_), .B(core__abc_21302_new_n4254_), .C(core__abc_21302_new_n4257_), .Y(core__abc_21302_new_n4275_));
AOI21X1 AOI21X1_708 ( .A(core__abc_21302_new_n4262_), .B(core__abc_21302_new_n4258_), .C(core__abc_21302_new_n4275_), .Y(core__abc_21302_new_n4276_));
AOI21X1 AOI21X1_709 ( .A(core__abc_21302_new_n4280_), .B(core__abc_21302_new_n4278_), .C(core__abc_21302_new_n4281_), .Y(core__abc_21302_new_n4282_));
AOI21X1 AOI21X1_71 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1620_), .C(_abc_19873_new_n1621_), .Y(_0word2_reg_31_0__5_));
AOI21X1 AOI21X1_710 ( .A(core__abc_21302_new_n4297_), .B(core__abc_21302_new_n4273_), .C(core__abc_21302_new_n1185__bF_buf12), .Y(core__0v3_reg_63_0__44_));
AOI21X1 AOI21X1_711 ( .A(core__abc_21302_new_n4312_), .B(core__abc_21302_new_n4316_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n4317_));
AOI21X1 AOI21X1_712 ( .A(core__abc_21302_new_n4320_), .B(core__abc_21302_new_n4299_), .C(core__abc_21302_new_n1185__bF_buf11), .Y(core__0v3_reg_63_0__45_));
AOI21X1 AOI21X1_713 ( .A(core__abc_21302_new_n4308_), .B(core__abc_21302_new_n4306_), .C(core__abc_21302_new_n4289_), .Y(core__abc_21302_new_n4323_));
AOI21X1 AOI21X1_714 ( .A(core__abc_21302_new_n4287_), .B(core__abc_21302_new_n4325_), .C(core__abc_21302_new_n4327_), .Y(core__abc_21302_new_n4328_));
AOI21X1 AOI21X1_715 ( .A(core__abc_21302_new_n4284_), .B(core__abc_21302_new_n2482_), .C(core__abc_21302_new_n2415_), .Y(core__abc_21302_new_n4335_));
AOI21X1 AOI21X1_716 ( .A(core__abc_21302_new_n4347_), .B(core__abc_21302_new_n4345_), .C(core__abc_21302_new_n4324_), .Y(core__abc_21302_new_n4348_));
AOI21X1 AOI21X1_717 ( .A(core__abc_21302_new_n4344_), .B(core__abc_21302_new_n4351_), .C(core__abc_21302_new_n2673__bF_buf10), .Y(core__abc_21302_new_n4352_));
AOI21X1 AOI21X1_718 ( .A(core__abc_21302_new_n4355_), .B(core__abc_21302_new_n4322_), .C(core__abc_21302_new_n1185__bF_buf10), .Y(core__0v3_reg_63_0__46_));
AOI21X1 AOI21X1_719 ( .A(core__abc_21302_new_n4370_), .B(core__abc_21302_new_n4329_), .C(core__abc_21302_new_n4341_), .Y(core__abc_21302_new_n4371_));
AOI21X1 AOI21X1_72 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1623_), .C(_abc_19873_new_n1624_), .Y(_0word2_reg_31_0__6_));
AOI21X1 AOI21X1_720 ( .A(core__abc_21302_new_n4374_), .B(core__abc_21302_new_n4377_), .C(core__abc_21302_new_n2673__bF_buf9), .Y(core__abc_21302_new_n4378_));
AOI21X1 AOI21X1_721 ( .A(core__abc_21302_new_n4382_), .B(core__abc_21302_new_n4357_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v3_reg_63_0__47_));
AOI21X1 AOI21X1_722 ( .A(core__abc_21302_new_n4366_), .B(core__abc_21302_new_n4364_), .C(core__abc_21302_new_n4341_), .Y(core__abc_21302_new_n4386_));
AOI21X1 AOI21X1_723 ( .A(core__abc_21302_new_n4161_), .B(core__abc_21302_new_n4390_), .C(core__abc_21302_new_n4394_), .Y(core__abc_21302_new_n4395_));
AOI21X1 AOI21X1_724 ( .A(core__abc_21302_new_n4408_), .B(core__abc_21302_new_n4384_), .C(core__abc_21302_new_n1185__bF_buf8), .Y(core__0v3_reg_63_0__48_));
AOI21X1 AOI21X1_725 ( .A(core__abc_21302_new_n4170_), .B(core__abc_21302_new_n4163_), .C(core__abc_21302_new_n4388_), .Y(core__abc_21302_new_n4426_));
AOI21X1 AOI21X1_726 ( .A(core__abc_21302_new_n4435_), .B(core__abc_21302_new_n4433_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n4436_));
AOI21X1 AOI21X1_727 ( .A(core__abc_21302_new_n4440_), .B(core__abc_21302_new_n4410_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0v3_reg_63_0__49_));
AOI21X1 AOI21X1_728 ( .A(core__abc_21302_new_n4399_), .B(core__abc_21302_new_n4417_), .C(core__abc_21302_new_n4415_), .Y(core__abc_21302_new_n4443_));
AOI21X1 AOI21X1_729 ( .A(core__abc_21302_new_n2420_), .B(core__abc_21302_new_n2431_), .C(core__abc_21302_new_n4444_), .Y(core__abc_21302_new_n4447_));
AOI21X1 AOI21X1_73 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1626_), .C(_abc_19873_new_n1627_), .Y(_0word2_reg_31_0__7_));
AOI21X1 AOI21X1_730 ( .A(core__abc_21302_new_n4431_), .B(core__abc_21302_new_n4443_), .C(core__abc_21302_new_n4454_), .Y(core__abc_21302_new_n4455_));
AOI21X1 AOI21X1_731 ( .A(core__abc_21302_new_n4462_), .B(core__abc_21302_new_n4463_), .C(core__abc_21302_new_n2673__bF_buf6), .Y(core__abc_21302_new_n4464_));
AOI21X1 AOI21X1_732 ( .A(core__abc_21302_new_n4467_), .B(core__abc_21302_new_n4442_), .C(core__abc_21302_new_n1185__bF_buf6), .Y(core__0v3_reg_63_0__50_));
AOI21X1 AOI21X1_733 ( .A(core__abc_21302_new_n2954_), .B(core__abc_21302_new_n2955_), .C(core__abc_21302_new_n4474_), .Y(core__abc_21302_new_n4475_));
AOI21X1 AOI21X1_734 ( .A(core__abc_21302_new_n4483_), .B(core__abc_21302_new_n4484_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n4485_));
AOI21X1 AOI21X1_735 ( .A(core__abc_21302_new_n4489_), .B(core__abc_21302_new_n4469_), .C(core__abc_21302_new_n1185__bF_buf5), .Y(core__0v3_reg_63_0__51_));
AOI21X1 AOI21X1_736 ( .A(core__abc_21302_new_n4477_), .B(core__abc_21302_new_n4450_), .C(core__abc_21302_new_n4475_), .Y(core__abc_21302_new_n4494_));
AOI21X1 AOI21X1_737 ( .A(core__abc_21302_new_n4512_), .B(core__abc_21302_new_n4491_), .C(core__abc_21302_new_n1185__bF_buf4), .Y(core__0v3_reg_63_0__52_));
AOI21X1 AOI21X1_738 ( .A(core__abc_21302_new_n4421_), .B(core__abc_21302_new_n4395_), .C(core__abc_21302_new_n4498_), .Y(core__abc_21302_new_n4515_));
AOI21X1 AOI21X1_739 ( .A(core__abc_21302_new_n3031_), .B(core__abc_21302_new_n3032_), .C(core__abc_21302_new_n4521_), .Y(core__abc_21302_new_n4524_));
AOI21X1 AOI21X1_74 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1079_), .C(_abc_19873_new_n1629_), .Y(_0word2_reg_31_0__8_));
AOI21X1 AOI21X1_740 ( .A(core__abc_21302_new_n4532_), .B(core__abc_21302_new_n4529_), .C(core__abc_21302_new_n2673__bF_buf3), .Y(core__abc_21302_new_n4533_));
AOI21X1 AOI21X1_741 ( .A(core__abc_21302_new_n4536_), .B(core__abc_21302_new_n4514_), .C(core__abc_21302_new_n1185__bF_buf3), .Y(core__0v3_reg_63_0__53_));
AOI21X1 AOI21X1_742 ( .A(core__abc_21302_new_n4540_), .B(core__abc_21302_new_n4543_), .C(core__abc_21302_new_n4551_), .Y(core__abc_21302_new_n4552_));
AOI21X1 AOI21X1_743 ( .A(core__abc_21302_new_n4557_), .B(core__abc_21302_new_n4555_), .C(core__abc_21302_new_n2673__bF_buf2), .Y(core__abc_21302_new_n4558_));
AOI21X1 AOI21X1_744 ( .A(core__abc_21302_new_n4561_), .B(core__abc_21302_new_n4538_), .C(core__abc_21302_new_n1185__bF_buf2), .Y(core__0v3_reg_63_0__54_));
AOI21X1 AOI21X1_745 ( .A(core__abc_21302_new_n4582_), .B(core__abc_21302_new_n4585_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n4586_));
AOI21X1 AOI21X1_746 ( .A(core__abc_21302_new_n4590_), .B(core__abc_21302_new_n4563_), .C(core__abc_21302_new_n1185__bF_buf1), .Y(core__0v3_reg_63_0__55_));
AOI21X1 AOI21X1_747 ( .A(core__abc_21302_new_n4574_), .B(core__abc_21302_new_n4576_), .C(core__abc_21302_new_n4551_), .Y(core__abc_21302_new_n4595_));
AOI21X1 AOI21X1_748 ( .A(core__abc_21302_new_n4421_), .B(core__abc_21302_new_n4395_), .C(core__abc_21302_new_n4596_), .Y(core__abc_21302_new_n4597_));
AOI21X1 AOI21X1_749 ( .A(core__abc_21302_new_n2420_), .B(core__abc_21302_new_n2496_), .C(core__abc_21302_new_n2500_), .Y(core__abc_21302_new_n4606_));
AOI21X1 AOI21X1_75 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1107_), .C(_abc_19873_new_n1631_), .Y(_0word2_reg_31_0__9_));
AOI21X1 AOI21X1_750 ( .A(core__abc_21302_new_n4614_), .B(core__abc_21302_new_n4592_), .C(core__abc_21302_new_n1185__bF_buf0), .Y(core__0v3_reg_63_0__56_));
AOI21X1 AOI21X1_751 ( .A(core__abc_21302_new_n4621_), .B(core__abc_21302_new_n4622_), .C(core__abc_21302_new_n4624_), .Y(core__abc_21302_new_n4625_));
AOI21X1 AOI21X1_752 ( .A(core__abc_21302_new_n3211_), .B(core__abc_21302_new_n3214_), .C(core__abc_21302_new_n4626_), .Y(core__abc_21302_new_n4627_));
AOI21X1 AOI21X1_753 ( .A(core__abc_21302_new_n4634_), .B(core__abc_21302_new_n4632_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n4635_));
AOI21X1 AOI21X1_754 ( .A(core__abc_21302_new_n4639_), .B(core__abc_21302_new_n4616_), .C(core__abc_21302_new_n1185__bF_buf13), .Y(core__0v3_reg_63_0__57_));
AOI21X1 AOI21X1_755 ( .A(core__abc_21302_new_n4649_), .B(core__abc_21302_new_n4646_), .C(core__abc_21302_new_n4658_), .Y(core__abc_21302_new_n4659_));
AOI21X1 AOI21X1_756 ( .A(core__abc_21302_new_n4663_), .B(core__abc_21302_new_n4665_), .C(core__abc_21302_new_n2673__bF_buf10), .Y(core__abc_21302_new_n4666_));
AOI21X1 AOI21X1_757 ( .A(core__abc_21302_new_n4669_), .B(core__abc_21302_new_n4641_), .C(core__abc_21302_new_n1185__bF_buf12), .Y(core__0v3_reg_63_0__58_));
AOI21X1 AOI21X1_758 ( .A(core__abc_21302_new_n4650_), .B(core__abc_21302_new_n1497_), .C(core__abc_21302_new_n1496_), .Y(core__abc_21302_new_n4674_));
AOI21X1 AOI21X1_759 ( .A(core__abc_21302_new_n4683_), .B(core__abc_21302_new_n4686_), .C(core__abc_21302_new_n4671_), .Y(core__abc_21302_new_n4688_));
AOI21X1 AOI21X1_76 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1117_), .C(_abc_19873_new_n1633_), .Y(_0word2_reg_31_0__10_));
AOI21X1 AOI21X1_760 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n4691_), .C(core__abc_21302_new_n4693_), .Y(core__abc_21302_new_n4694_));
AOI21X1 AOI21X1_761 ( .A(core__abc_21302_new_n4690_), .B(core__abc_21302_new_n4694_), .C(core__abc_21302_new_n4695_), .Y(core__0v3_reg_63_0__59_));
AOI21X1 AOI21X1_762 ( .A(core__abc_21302_new_n4699_), .B(core__abc_21302_new_n4704_), .C(core__abc_21302_new_n4703_), .Y(core__abc_21302_new_n4705_));
AOI21X1 AOI21X1_763 ( .A(core__abc_21302_new_n4702_), .B(core__abc_21302_new_n4705_), .C(core__abc_21302_new_n4718_), .Y(core__abc_21302_new_n4719_));
AOI21X1 AOI21X1_764 ( .A(core__abc_21302_new_n4724_), .B(core__abc_21302_new_n4722_), .C(core__abc_21302_new_n2673__bF_buf8), .Y(core__abc_21302_new_n4725_));
AOI21X1 AOI21X1_765 ( .A(core__abc_21302_new_n4728_), .B(core__abc_21302_new_n4697_), .C(core__abc_21302_new_n1185__bF_buf11), .Y(core__0v3_reg_63_0__60_));
AOI21X1 AOI21X1_766 ( .A(core__abc_21302_new_n4733_), .B(core__abc_21302_new_n4734_), .C(core__abc_21302_new_n4735_), .Y(core__abc_21302_new_n4736_));
AOI21X1 AOI21X1_767 ( .A(core__abc_21302_new_n3406_), .B(core__abc_21302_new_n3402_), .C(core__abc_21302_new_n4744_), .Y(core__abc_21302_new_n4747_));
AOI21X1 AOI21X1_768 ( .A(core__abc_21302_new_n4753_), .B(core__abc_21302_new_n4756_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n4757_));
AOI21X1 AOI21X1_769 ( .A(core__abc_21302_new_n4760_), .B(core__abc_21302_new_n4730_), .C(core__abc_21302_new_n1185__bF_buf10), .Y(core__0v3_reg_63_0__61_));
AOI21X1 AOI21X1_77 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1635_), .C(_abc_19873_new_n1636_), .Y(_0word2_reg_31_0__11_));
AOI21X1 AOI21X1_770 ( .A(core__abc_21302_new_n4707_), .B(core__abc_21302_new_n4706_), .C(core__abc_21302_new_n2422_), .Y(core__abc_21302_new_n4768_));
AOI21X1 AOI21X1_771 ( .A(core__abc_21302_new_n4702_), .B(core__abc_21302_new_n4705_), .C(core__abc_21302_new_n4783_), .Y(core__abc_21302_new_n4784_));
AOI21X1 AOI21X1_772 ( .A(core__abc_21302_new_n4789_), .B(core__abc_21302_new_n4786_), .C(core__abc_21302_new_n2673__bF_buf6), .Y(core__abc_21302_new_n4790_));
AOI21X1 AOI21X1_773 ( .A(core__abc_21302_new_n4793_), .B(core__abc_21302_new_n4762_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v3_reg_63_0__62_));
AOI21X1 AOI21X1_774 ( .A(core__abc_21302_new_n2167_), .B(core__abc_21302_new_n4816_), .C(core__abc_21302_new_n4818_), .Y(core__abc_21302_new_n4819_));
AOI21X1 AOI21X1_775 ( .A(core__abc_21302_new_n4815_), .B(core__abc_21302_new_n4819_), .C(core__abc_21302_new_n4820_), .Y(core__0v3_reg_63_0__63_));
AOI21X1 AOI21X1_776 ( .A(core__abc_21302_new_n4801_), .B(core__abc_21302_new_n4799_), .C(core__abc_21302_new_n4824_), .Y(core__abc_21302_new_n4827_));
AOI21X1 AOI21X1_777 ( .A(core__abc_21302_new_n4853_), .B(core__abc_21302_new_n4878_), .C(core__abc_21302_new_n4887_), .Y(core__abc_21302_new_n4888_));
AOI21X1 AOI21X1_778 ( .A(core__abc_21302_new_n4898_), .B(core__abc_21302_new_n4897_), .C(core_v1_reg_10_), .Y(core__abc_21302_new_n4902_));
AOI21X1 AOI21X1_779 ( .A(core__abc_21302_new_n4572_), .B(core__abc_21302_new_n4570_), .C(core__abc_21302_new_n4248_), .Y(core__abc_21302_new_n4903_));
AOI21X1 AOI21X1_78 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1638_), .C(_abc_19873_new_n1639_), .Y(_0word2_reg_31_0__12_));
AOI21X1 AOI21X1_780 ( .A(core__abc_21302_new_n4960_), .B(core__abc_21302_new_n4904_), .C(core__abc_21302_new_n4959_), .Y(core__abc_21302_new_n4961_));
AOI21X1 AOI21X1_781 ( .A(core__abc_21302_new_n4955_), .B(core__abc_21302_new_n4928_), .C(core__abc_21302_new_n4962_), .Y(core__abc_21302_new_n4963_));
AOI21X1 AOI21X1_782 ( .A(core__abc_21302_new_n4967_), .B(core__abc_21302_new_n3230_), .C(core__abc_21302_new_n4972_), .Y(core__abc_21302_new_n4985_));
AOI21X1 AOI21X1_783 ( .A(core__abc_21302_new_n3233_), .B(core__abc_21302_new_n4984_), .C(core__abc_21302_new_n4985_), .Y(core__abc_21302_new_n4986_));
AOI21X1 AOI21X1_784 ( .A(core__abc_21302_new_n5009_), .B(core__abc_21302_new_n5015_), .C(core__abc_21302_new_n5006_), .Y(core__abc_21302_new_n5016_));
AOI21X1 AOI21X1_785 ( .A(core__abc_21302_new_n5023_), .B(core__abc_21302_new_n5026_), .C(core__abc_21302_new_n5021_), .Y(core__abc_21302_new_n5027_));
AOI21X1 AOI21X1_786 ( .A(core__abc_21302_new_n5044_), .B(core__abc_21302_new_n5043_), .C(core__abc_21302_new_n2651_), .Y(core__abc_21302_new_n5045_));
AOI21X1 AOI21X1_787 ( .A(core__abc_21302_new_n5048_), .B(core__abc_21302_new_n5049_), .C(core__abc_21302_new_n5045_), .Y(core__abc_21302_new_n5050_));
AOI21X1 AOI21X1_788 ( .A(core__abc_21302_new_n5053_), .B(core__abc_21302_new_n5040_), .C(core__abc_21302_new_n5039_), .Y(core__abc_21302_new_n5054_));
AOI21X1 AOI21X1_789 ( .A(core__abc_21302_new_n5016_), .B(core__abc_21302_new_n5063_), .C(core__abc_21302_new_n4994_), .Y(core__abc_21302_new_n5064_));
AOI21X1 AOI21X1_79 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1177_), .C(_abc_19873_new_n1641_), .Y(_0word2_reg_31_0__13_));
AOI21X1 AOI21X1_790 ( .A(core__abc_21302_new_n5083_), .B(core__abc_21302_new_n5086_), .C(core__abc_21302_new_n1185__bF_buf8), .Y(core__0v2_reg_63_0__0_));
AOI21X1 AOI21X1_791 ( .A(core__abc_21302_new_n5101_), .B(core__abc_21302_new_n5102_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0v2_reg_63_0__1_));
AOI21X1 AOI21X1_792 ( .A(core__abc_21302_new_n5148_), .B(core__abc_21302_new_n5149_), .C(core__abc_21302_new_n1185__bF_buf6), .Y(core__0v2_reg_63_0__3_));
AOI21X1 AOI21X1_793 ( .A(core__abc_21302_new_n5162_), .B(core__abc_21302_new_n5160_), .C(core__abc_21302_new_n5154_), .Y(core__abc_21302_new_n5163_));
AOI21X1 AOI21X1_794 ( .A(core__abc_21302_new_n5184_), .B(core__abc_21302_new_n5185_), .C(core__abc_21302_new_n1185__bF_buf4), .Y(core__0v2_reg_63_0__5_));
AOI21X1 AOI21X1_795 ( .A(core__abc_21302_new_n5166_), .B(core__abc_21302_new_n5194_), .C(core__abc_21302_new_n5193_), .Y(core__abc_21302_new_n5195_));
AOI21X1 AOI21X1_796 ( .A(core__abc_21302_new_n5202_), .B(core__abc_21302_new_n5203_), .C(core__abc_21302_new_n1185__bF_buf3), .Y(core__0v2_reg_63_0__6_));
AOI21X1 AOI21X1_797 ( .A(core__abc_21302_new_n5217_), .B(core__abc_21302_new_n5219_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n5220_));
AOI21X1 AOI21X1_798 ( .A(core__abc_21302_new_n5223_), .B(core__abc_21302_new_n5224_), .C(core__abc_21302_new_n1185__bF_buf2), .Y(core__0v2_reg_63_0__7_));
AOI21X1 AOI21X1_799 ( .A(core__abc_21302_new_n5212_), .B(core__abc_21302_new_n5215_), .C(core__abc_21302_new_n5192_), .Y(core__abc_21302_new_n5226_));
AOI21X1 AOI21X1_8 ( .A(_abc_19873_new_n1077_), .B(_abc_19873_new_n1066_), .C(_abc_19873_new_n928__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_27087_7_));
AOI21X1 AOI21X1_80 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1643_), .C(_abc_19873_new_n1644_), .Y(_0word2_reg_31_0__14_));
AOI21X1 AOI21X1_800 ( .A(core__abc_21302_new_n5073_), .B(core__abc_21302_new_n5228_), .C(core__abc_21302_new_n5234_), .Y(core__abc_21302_new_n5235_));
AOI21X1 AOI21X1_801 ( .A(core__abc_21302_new_n5242_), .B(core__abc_21302_new_n2634__bF_buf2), .C(core__abc_21302_new_n5244_), .Y(core__abc_21302_new_n5245_));
AOI21X1 AOI21X1_802 ( .A(core__abc_21302_new_n5259_), .B(core__abc_21302_new_n5104__bF_buf3), .C(core__abc_21302_new_n5260_), .Y(core__0v2_reg_63_0__9_));
AOI21X1 AOI21X1_803 ( .A(core__abc_21302_new_n5253_), .B(core__abc_21302_new_n5239_), .C(core__abc_21302_new_n5264_), .Y(core__abc_21302_new_n5265_));
AOI21X1 AOI21X1_804 ( .A(core__abc_21302_new_n5279_), .B(core__abc_21302_new_n2634__bF_buf0), .C(core__abc_21302_new_n5281_), .Y(core__abc_21302_new_n5282_));
AOI21X1 AOI21X1_805 ( .A(core__abc_21302_new_n5292_), .B(core__abc_21302_new_n5304_), .C(core__abc_21302_new_n5305_), .Y(core__abc_21302_new_n5306_));
AOI21X1 AOI21X1_806 ( .A(core__abc_21302_new_n5319_), .B(core__abc_21302_new_n5104__bF_buf6), .C(core__abc_21302_new_n5320_), .Y(core__0v2_reg_63_0__12_));
AOI21X1 AOI21X1_807 ( .A(core__abc_21302_new_n5337_), .B(core__abc_21302_new_n5339_), .C(core__abc_21302_new_n5340_), .Y(core__0v2_reg_63_0__13_));
AOI21X1 AOI21X1_808 ( .A(core__abc_21302_new_n5342_), .B(core__abc_21302_new_n5313_), .C(core__abc_21302_new_n5344_), .Y(core__abc_21302_new_n5345_));
AOI21X1 AOI21X1_809 ( .A(core__abc_21302_new_n3226_), .B(core__abc_21302_new_n3224_), .C(core__abc_21302_new_n1588_), .Y(core__abc_21302_new_n5370_));
AOI21X1 AOI21X1_81 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1219_), .C(_abc_19873_new_n1646_), .Y(_0word2_reg_31_0__15_));
AOI21X1 AOI21X1_810 ( .A(core__abc_21302_new_n5359_), .B(core__abc_21302_new_n5358_), .C(core__abc_21302_new_n5360_), .Y(core__abc_21302_new_n5379_));
AOI21X1 AOI21X1_811 ( .A(core__abc_21302_new_n5374_), .B(core__abc_21302_new_n5371_), .C(core__abc_21302_new_n5360_), .Y(core__abc_21302_new_n5388_));
AOI21X1 AOI21X1_812 ( .A(core__abc_21302_new_n5378_), .B(core__abc_21302_new_n5393_), .C(core__abc_21302_new_n5392_), .Y(core__abc_21302_new_n5394_));
AOI21X1 AOI21X1_813 ( .A(core__abc_21302_new_n5397_), .B(core__abc_21302_new_n5234_), .C(core__abc_21302_new_n5395_), .Y(core__abc_21302_new_n5398_));
AOI21X1 AOI21X1_814 ( .A(core__abc_21302_new_n5412_), .B(core__abc_21302_new_n5104__bF_buf1), .C(core__abc_21302_new_n5413_), .Y(core__0v2_reg_63_0__16_));
AOI21X1 AOI21X1_815 ( .A(core__abc_21302_new_n5094_), .B(core__abc_21302_new_n4888_), .C(core__abc_21302_new_n5402_), .Y(core__abc_21302_new_n5418_));
AOI21X1 AOI21X1_816 ( .A(core__abc_21302_new_n5428_), .B(core__abc_21302_new_n5431_), .C(core__abc_21302_new_n5432_), .Y(core__0v2_reg_63_0__17_));
AOI21X1 AOI21X1_817 ( .A(core__abc_21302_new_n5449_), .B(core__abc_21302_new_n5451_), .C(core__abc_21302_new_n5452_), .Y(core__0v2_reg_63_0__18_));
AOI21X1 AOI21X1_818 ( .A(core__abc_21302_new_n5472_), .B(core__abc_21302_new_n5398_), .C(core__abc_21302_new_n5475_), .Y(core__abc_21302_new_n5476_));
AOI21X1 AOI21X1_819 ( .A(core__abc_21302_new_n5486_), .B(core__abc_21302_new_n5489_), .C(core__abc_21302_new_n5490_), .Y(core__0v2_reg_63_0__20_));
AOI21X1 AOI21X1_82 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1648_), .C(_abc_19873_new_n1649_), .Y(_0word2_reg_31_0__16_));
AOI21X1 AOI21X1_820 ( .A(core__abc_21302_new_n5516_), .B(core__abc_21302_new_n5518_), .C(core__abc_21302_new_n5513_), .Y(core__abc_21302_new_n5519_));
AOI21X1 AOI21X1_821 ( .A(core__abc_21302_new_n5539_), .B(core__abc_21302_new_n5542_), .C(core__abc_21302_new_n5543_), .Y(core__0v2_reg_63_0__23_));
AOI21X1 AOI21X1_822 ( .A(core__abc_21302_new_n5533_), .B(core__abc_21302_new_n5536_), .C(core__abc_21302_new_n5548_), .Y(core__abc_21302_new_n5549_));
AOI21X1 AOI21X1_823 ( .A(core__abc_21302_new_n5472_), .B(core__abc_21302_new_n5398_), .C(core__abc_21302_new_n5552_), .Y(core__abc_21302_new_n5553_));
AOI21X1 AOI21X1_824 ( .A(core__abc_21302_new_n5578_), .B(core__abc_21302_new_n5580_), .C(core__abc_21302_new_n5581_), .Y(core__0v2_reg_63_0__25_));
AOI21X1 AOI21X1_825 ( .A(core__abc_21302_new_n5576_), .B(core__abc_21302_new_n5555_), .C(core__abc_21302_new_n5573_), .Y(core__abc_21302_new_n5591_));
AOI21X1 AOI21X1_826 ( .A(core__abc_21302_new_n5590_), .B(core__abc_21302_new_n5591_), .C(core__abc_21302_new_n5587_), .Y(core__abc_21302_new_n5592_));
AOI21X1 AOI21X1_827 ( .A(core__abc_21302_new_n5612_), .B(core__abc_21302_new_n5614_), .C(core__abc_21302_new_n5615_), .Y(core__0v2_reg_63_0__27_));
AOI21X1 AOI21X1_828 ( .A(core__abc_21302_new_n5633_), .B(core__abc_21302_new_n5631_), .C(core__abc_21302_new_n5618_), .Y(core__abc_21302_new_n5634_));
AOI21X1 AOI21X1_829 ( .A(core__abc_21302_new_n5620_), .B(core__abc_21302_new_n5624_), .C(core__abc_21302_new_n5654_), .Y(core__abc_21302_new_n5655_));
AOI21X1 AOI21X1_83 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1651_), .C(_abc_19873_new_n1652_), .Y(_0word2_reg_31_0__17_));
AOI21X1 AOI21X1_830 ( .A(core__abc_21302_new_n5637_), .B(core__abc_21302_new_n5653_), .C(core__abc_21302_new_n5655_), .Y(core__abc_21302_new_n5656_));
AOI21X1 AOI21X1_831 ( .A(core__abc_21302_new_n5664_), .B(core__abc_21302_new_n5666_), .C(core__abc_21302_new_n5674_), .Y(core__abc_21302_new_n5691_));
AOI21X1 AOI21X1_832 ( .A(core__abc_21302_new_n5693_), .B(core__abc_21302_new_n5696_), .C(core__abc_21302_new_n5697_), .Y(core__0v2_reg_63_0__31_));
AOI21X1 AOI21X1_833 ( .A(core__abc_21302_new_n5703_), .B(core__abc_21302_new_n5704_), .C(core__abc_21302_new_n1185__bF_buf4), .Y(core__0v2_reg_63_0__32_));
AOI21X1 AOI21X1_834 ( .A(core__abc_21302_new_n5712_), .B(core__abc_21302_new_n5706_), .C(core__abc_21302_new_n1185__bF_buf3), .Y(core__0v2_reg_63_0__33_));
AOI21X1 AOI21X1_835 ( .A(core__abc_21302_new_n5715_), .B(core__abc_21302_new_n5717_), .C(core__abc_21302_new_n5718_), .Y(core__0v2_reg_63_0__34_));
AOI21X1 AOI21X1_836 ( .A(core__abc_21302_new_n5722_), .B(core__abc_21302_new_n5725_), .C(core__abc_21302_new_n5726_), .Y(core__0v2_reg_63_0__35_));
AOI21X1 AOI21X1_837 ( .A(core__abc_21302_new_n5728_), .B(core__abc_21302_new_n5085__bF_buf3), .C(core__abc_21302_new_n5735_), .Y(core__0v2_reg_63_0__36_));
AOI21X1 AOI21X1_838 ( .A(core__abc_21302_new_n5742_), .B(core__abc_21302_new_n5104__bF_buf4), .C(core__abc_21302_new_n5743_), .Y(core__0v2_reg_63_0__37_));
AOI21X1 AOI21X1_839 ( .A(core__abc_21302_new_n5746_), .B(core__abc_21302_new_n5749_), .C(core__abc_21302_new_n5750_), .Y(core__0v2_reg_63_0__38_));
AOI21X1 AOI21X1_84 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1654_), .C(_abc_19873_new_n1655_), .Y(_0word2_reg_31_0__18_));
AOI21X1 AOI21X1_840 ( .A(core__abc_21302_new_n5757_), .B(core__abc_21302_new_n5761_), .C(core__abc_21302_new_n5762_), .Y(core__0v2_reg_63_0__39_));
AOI21X1 AOI21X1_841 ( .A(core__abc_21302_new_n5765_), .B(core__abc_21302_new_n5769_), .C(core__abc_21302_new_n5770_), .Y(core__0v2_reg_63_0__40_));
AOI21X1 AOI21X1_842 ( .A(core__abc_21302_new_n5779_), .B(core__abc_21302_new_n5104__bF_buf7), .C(core__abc_21302_new_n5780_), .Y(core__0v2_reg_63_0__41_));
AOI21X1 AOI21X1_843 ( .A(core__abc_21302_new_n5059_), .B(core__abc_21302_new_n5062_), .C(core__abc_21302_new_n5015_), .Y(core__abc_21302_new_n5782_));
AOI21X1 AOI21X1_844 ( .A(core__abc_21302_new_n5784_), .B(core__abc_21302_new_n5787_), .C(core__abc_21302_new_n5788_), .Y(core__0v2_reg_63_0__42_));
AOI21X1 AOI21X1_845 ( .A(core__abc_21302_new_n5792_), .B(core__abc_21302_new_n5794_), .C(core__abc_21302_new_n5795_), .Y(core__0v2_reg_63_0__43_));
AOI21X1 AOI21X1_846 ( .A(core__abc_21302_new_n5805_), .B(core__abc_21302_new_n5808_), .C(core__abc_21302_new_n5809_), .Y(core__0v2_reg_63_0__44_));
AOI21X1 AOI21X1_847 ( .A(core__abc_21302_new_n5816_), .B(core__abc_21302_new_n5104__bF_buf1), .C(core__abc_21302_new_n5817_), .Y(core__0v2_reg_63_0__45_));
AOI21X1 AOI21X1_848 ( .A(core__abc_21302_new_n5821_), .B(core__abc_21302_new_n5824_), .C(core__abc_21302_new_n5825_), .Y(core__0v2_reg_63_0__46_));
AOI21X1 AOI21X1_849 ( .A(core__abc_21302_new_n5835_), .B(core__abc_21302_new_n5104__bF_buf6), .C(core__abc_21302_new_n5836_), .Y(core__0v2_reg_63_0__47_));
AOI21X1 AOI21X1_85 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1657_), .C(_abc_19873_new_n1658_), .Y(_0word2_reg_31_0__19_));
AOI21X1 AOI21X1_850 ( .A(core__abc_21302_new_n5843_), .B(core__abc_21302_new_n5846_), .C(core__abc_21302_new_n5847_), .Y(core__0v2_reg_63_0__48_));
AOI21X1 AOI21X1_851 ( .A(core__abc_21302_new_n5864_), .B(core__abc_21302_new_n5868_), .C(core__abc_21302_new_n5869_), .Y(core__0v2_reg_63_0__50_));
AOI21X1 AOI21X1_852 ( .A(core__abc_21302_new_n5875_), .B(core__abc_21302_new_n5104__bF_buf1), .C(core__abc_21302_new_n5876_), .Y(core__0v2_reg_63_0__51_));
AOI21X1 AOI21X1_853 ( .A(core__abc_21302_new_n5886_), .B(core__abc_21302_new_n5104__bF_buf7), .C(core__abc_21302_new_n5887_), .Y(core__0v2_reg_63_0__52_));
AOI21X1 AOI21X1_854 ( .A(core__abc_21302_new_n5896_), .B(core__abc_21302_new_n5104__bF_buf5), .C(core__abc_21302_new_n5897_), .Y(core__0v2_reg_63_0__53_));
AOI21X1 AOI21X1_855 ( .A(core__abc_21302_new_n5924_), .B(core__abc_21302_new_n2634__bF_buf0), .C(core__abc_21302_new_n5926_), .Y(core__abc_21302_new_n5927_));
AOI21X1 AOI21X1_856 ( .A(core__abc_21302_new_n5932_), .B(core__abc_21302_new_n5934_), .C(core__abc_21302_new_n5935_), .Y(core__0v2_reg_63_0__57_));
AOI21X1 AOI21X1_857 ( .A(core__abc_21302_new_n5941_), .B(core__abc_21302_new_n5104__bF_buf5), .C(core__abc_21302_new_n5942_), .Y(core__0v2_reg_63_0__58_));
AOI21X1 AOI21X1_858 ( .A(core__abc_21302_new_n5950_), .B(core__abc_21302_new_n5104__bF_buf3), .C(core__abc_21302_new_n5951_), .Y(core__0v2_reg_63_0__59_));
AOI21X1 AOI21X1_859 ( .A(core__abc_21302_new_n5959_), .B(core__abc_21302_new_n5962_), .C(core__abc_21302_new_n5963_), .Y(core__0v2_reg_63_0__60_));
AOI21X1 AOI21X1_86 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1660_), .C(_abc_19873_new_n1661_), .Y(_0word2_reg_31_0__20_));
AOI21X1 AOI21X1_860 ( .A(core__abc_21302_new_n5992_), .B(core__abc_21302_new_n5104__bF_buf6), .C(core__abc_21302_new_n5993_), .Y(core__0v2_reg_63_0__63_));
AOI21X1 AOI21X1_861 ( .A(core__abc_21302_new_n6004_), .B(core__abc_21302_new_n5996_), .C(core__abc_21302_new_n1185__bF_buf11), .Y(core__0v1_reg_63_0__0_));
AOI21X1 AOI21X1_862 ( .A(core__abc_21302_new_n5405_), .B(core__abc_21302_new_n5710_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n6006_));
AOI21X1 AOI21X1_863 ( .A(core__abc_21302_new_n2639__bF_buf4), .B(core__abc_21302_new_n6008_), .C(core__abc_21302_new_n6010_), .Y(core__abc_21302_new_n6011_));
AOI21X1 AOI21X1_864 ( .A(core__abc_21302_new_n6007_), .B(core__abc_21302_new_n6011_), .C(core__abc_21302_new_n6012_), .Y(core__0v1_reg_63_0__1_));
AOI21X1 AOI21X1_865 ( .A(core__abc_21302_new_n6020_), .B(core__abc_21302_new_n6014_), .C(core__abc_21302_new_n1185__bF_buf10), .Y(core__0v1_reg_63_0__2_));
AOI21X1 AOI21X1_866 ( .A(core__abc_21302_new_n2634__bF_buf4), .B(core__abc_21302_new_n6023_), .C(core__abc_21302_new_n5435_), .Y(core__abc_21302_new_n6024_));
AOI21X1 AOI21X1_867 ( .A(core__abc_21302_new_n5435_), .B(core__abc_21302_new_n5722_), .C(core__abc_21302_new_n6024_), .Y(core__abc_21302_new_n6025_));
AOI21X1 AOI21X1_868 ( .A(core__abc_21302_new_n6028_), .B(core__abc_21302_new_n6022_), .C(core__abc_21302_new_n1185__bF_buf9), .Y(core__0v1_reg_63_0__3_));
AOI21X1 AOI21X1_869 ( .A(core__abc_21302_new_n5466_), .B(core__abc_21302_new_n5731_), .C(core__abc_21302_new_n6033_), .Y(core__abc_21302_new_n6034_));
AOI21X1 AOI21X1_87 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1320_), .C(_abc_19873_new_n1663_), .Y(_0word2_reg_31_0__21_));
AOI21X1 AOI21X1_870 ( .A(core__abc_21302_new_n6036_), .B(core__abc_21302_new_n6030_), .C(core__abc_21302_new_n1185__bF_buf8), .Y(core__0v1_reg_63_0__4_));
AOI21X1 AOI21X1_871 ( .A(core__abc_21302_new_n6038_), .B(core__abc_21302_new_n5479_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n6039_));
AOI21X1 AOI21X1_872 ( .A(core__abc_21302_new_n2639__bF_buf1), .B(core__abc_21302_new_n6041_), .C(core__abc_21302_new_n6042_), .Y(core__abc_21302_new_n6043_));
AOI21X1 AOI21X1_873 ( .A(core__abc_21302_new_n6040_), .B(core__abc_21302_new_n6043_), .C(core__abc_21302_new_n6044_), .Y(core__0v1_reg_63_0__5_));
AOI21X1 AOI21X1_874 ( .A(core__abc_21302_new_n6051_), .B(core__abc_21302_new_n6046_), .C(core__abc_21302_new_n1185__bF_buf7), .Y(core__0v1_reg_63_0__6_));
AOI21X1 AOI21X1_875 ( .A(core__abc_21302_new_n6059_), .B(core__abc_21302_new_n6053_), .C(core__abc_21302_new_n1185__bF_buf6), .Y(core__0v1_reg_63_0__7_));
AOI21X1 AOI21X1_876 ( .A(core__abc_21302_new_n6065_), .B(core__abc_21302_new_n6009__bF_buf4), .C(core__abc_21302_new_n6066_), .Y(core__0v1_reg_63_0__8_));
AOI21X1 AOI21X1_877 ( .A(core__abc_21302_new_n5554_), .B(core__abc_21302_new_n5776_), .C(core__abc_21302_new_n6069_), .Y(core__abc_21302_new_n6070_));
AOI21X1 AOI21X1_878 ( .A(core__abc_21302_new_n5998__bF_buf1), .B(core_v1_reg_9_), .C(core__abc_21302_new_n6068_), .Y(core__abc_21302_new_n6071_));
AOI21X1 AOI21X1_879 ( .A(core__abc_21302_new_n4906_), .B(core__abc_21302_new_n6068_), .C(core__abc_21302_new_n6073_), .Y(core__0v1_reg_63_0__9_));
AOI21X1 AOI21X1_88 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1665_), .C(_abc_19873_new_n1666_), .Y(_0word2_reg_31_0__22_));
AOI21X1 AOI21X1_880 ( .A(core__abc_21302_new_n6078_), .B(core__abc_21302_new_n6009__bF_buf1), .C(core__abc_21302_new_n6079_), .Y(core__0v1_reg_63_0__10_));
AOI21X1 AOI21X1_881 ( .A(core__abc_21302_new_n6081_), .B(core__abc_21302_new_n5791_), .C(core__abc_21302_new_n6082_), .Y(core__abc_21302_new_n6083_));
AOI21X1 AOI21X1_882 ( .A(core__abc_21302_new_n5998__bF_buf0), .B(core_v1_reg_11_), .C(core__abc_21302_new_n6068_), .Y(core__abc_21302_new_n6084_));
AOI21X1 AOI21X1_883 ( .A(core__abc_21302_new_n4871_), .B(core__abc_21302_new_n6068_), .C(core__abc_21302_new_n6086_), .Y(core__0v1_reg_63_0__11_));
AOI21X1 AOI21X1_884 ( .A(core__abc_21302_new_n6091_), .B(core__abc_21302_new_n6009__bF_buf9), .C(core__abc_21302_new_n6092_), .Y(core__0v1_reg_63_0__12_));
AOI21X1 AOI21X1_885 ( .A(core__abc_21302_new_n5625_), .B(core__abc_21302_new_n5813_), .C(core__abc_21302_new_n6094_), .Y(core__abc_21302_new_n6095_));
AOI21X1 AOI21X1_886 ( .A(core__abc_21302_new_n5998__bF_buf3), .B(core_v1_reg_13_), .C(core__abc_21302_new_n6068_), .Y(core__abc_21302_new_n6096_));
AOI21X1 AOI21X1_887 ( .A(core__abc_21302_new_n5820_), .B(core__abc_21302_new_n6100_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n6101_));
AOI21X1 AOI21X1_888 ( .A(core__abc_21302_new_n6104_), .B(core__abc_21302_new_n6009__bF_buf6), .C(core__abc_21302_new_n6105_), .Y(core__0v1_reg_63_0__14_));
AOI21X1 AOI21X1_889 ( .A(core__abc_21302_new_n5832_), .B(core__abc_21302_new_n5670_), .C(core__abc_21302_new_n2673__bF_buf6), .Y(core__abc_21302_new_n6107_));
AOI21X1 AOI21X1_89 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1356_), .C(_abc_19873_new_n1668_), .Y(_0word2_reg_31_0__23_));
AOI21X1 AOI21X1_890 ( .A(core__abc_21302_new_n6110_), .B(core__abc_21302_new_n6009__bF_buf4), .C(core__abc_21302_new_n6111_), .Y(core__0v1_reg_63_0__15_));
AOI21X1 AOI21X1_891 ( .A(core__abc_21302_new_n6116_), .B(core__abc_21302_new_n6009__bF_buf2), .C(core__abc_21302_new_n6117_), .Y(core__0v1_reg_63_0__16_));
AOI21X1 AOI21X1_892 ( .A(core__abc_21302_new_n5851_), .B(core__abc_21302_new_n5047_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n6119_));
AOI21X1 AOI21X1_893 ( .A(core__abc_21302_new_n6122_), .B(core__abc_21302_new_n6009__bF_buf0), .C(core__abc_21302_new_n6123_), .Y(core__0v1_reg_63_0__17_));
AOI21X1 AOI21X1_894 ( .A(core__abc_21302_new_n5863_), .B(core__abc_21302_new_n6125_), .C(core__abc_21302_new_n2673__bF_buf4), .Y(core__abc_21302_new_n6126_));
AOI21X1 AOI21X1_895 ( .A(core__abc_21302_new_n6129_), .B(core__abc_21302_new_n6009__bF_buf8), .C(core__abc_21302_new_n6130_), .Y(core__0v1_reg_63_0__18_));
AOI21X1 AOI21X1_896 ( .A(core__abc_21302_new_n5872_), .B(core__abc_21302_new_n6132_), .C(core__abc_21302_new_n2673__bF_buf3), .Y(core__abc_21302_new_n6133_));
AOI21X1 AOI21X1_897 ( .A(core_v1_reg_19_), .B(core__abc_21302_new_n5998__bF_buf2), .C(core__abc_21302_new_n6135_), .Y(core__abc_21302_new_n6136_));
AOI21X1 AOI21X1_898 ( .A(core__abc_21302_new_n6134_), .B(core__abc_21302_new_n6136_), .C(core__abc_21302_new_n6137_), .Y(core__0v1_reg_63_0__19_));
AOI21X1 AOI21X1_899 ( .A(core_key_84_), .B(core__abc_21302_new_n2639__bF_buf0), .C(core__abc_21302_new_n6143_), .Y(core__abc_21302_new_n6144_));
AOI21X1 AOI21X1_9 ( .A(_abc_19873_new_n1087_), .B(_abc_19873_new_n1096_), .C(_abc_19873_new_n928__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_27087_8_));
AOI21X1 AOI21X1_90 ( .A(_abc_19873_new_n1524__bF_buf14), .B(_abc_19873_new_n1670_), .C(_abc_19873_new_n1671_), .Y(_0word2_reg_31_0__24_));
AOI21X1 AOI21X1_900 ( .A(core__abc_21302_new_n6141_), .B(core__abc_21302_new_n6144_), .C(core__abc_21302_new_n6145_), .Y(core__0v1_reg_63_0__20_));
AOI21X1 AOI21X1_901 ( .A(core__abc_21302_new_n5892_), .B(core__abc_21302_new_n5035_), .C(core__abc_21302_new_n2673__bF_buf2), .Y(core__abc_21302_new_n6147_));
AOI21X1 AOI21X1_902 ( .A(core__abc_21302_new_n6150_), .B(core__abc_21302_new_n6009__bF_buf2), .C(core__abc_21302_new_n6151_), .Y(core__0v1_reg_63_0__21_));
AOI21X1 AOI21X1_903 ( .A(core__abc_21302_new_n6157_), .B(core__abc_21302_new_n6009__bF_buf0), .C(core__abc_21302_new_n6158_), .Y(core__0v1_reg_63_0__22_));
AOI21X1 AOI21X1_904 ( .A(core__abc_21302_new_n5914_), .B(core__abc_21302_new_n5025_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n6160_));
AOI21X1 AOI21X1_905 ( .A(core__abc_21302_new_n6161_), .B(core__abc_21302_new_n6164_), .C(core__abc_21302_new_n6165_), .Y(core__0v1_reg_63_0__23_));
AOI21X1 AOI21X1_906 ( .A(core_key_88_), .B(core__abc_21302_new_n2639__bF_buf6), .C(core__abc_21302_new_n6170_), .Y(core__abc_21302_new_n6171_));
AOI21X1 AOI21X1_907 ( .A(core__abc_21302_new_n6169_), .B(core__abc_21302_new_n6171_), .C(core__abc_21302_new_n6172_), .Y(core__0v1_reg_63_0__24_));
AOI21X1 AOI21X1_908 ( .A(core__abc_21302_new_n5931_), .B(core__abc_21302_new_n5012_), .C(core__abc_21302_new_n2673__bF_buf0), .Y(core__abc_21302_new_n6174_));
AOI21X1 AOI21X1_909 ( .A(core__abc_21302_new_n3682_), .B(core__abc_21302_new_n2639__bF_buf5), .C(core__abc_21302_new_n6177_), .Y(core__abc_21302_new_n6178_));
AOI21X1 AOI21X1_91 ( .A(_abc_19873_new_n1524__bF_buf12), .B(_abc_19873_new_n1673_), .C(_abc_19873_new_n1674_), .Y(_0word2_reg_31_0__25_));
AOI21X1 AOI21X1_910 ( .A(core__abc_21302_new_n6175_), .B(core__abc_21302_new_n6178_), .C(core__abc_21302_new_n6179_), .Y(core__0v1_reg_63_0__25_));
AOI21X1 AOI21X1_911 ( .A(core__abc_21302_new_n3687_), .B(core__abc_21302_new_n2639__bF_buf4), .C(core__abc_21302_new_n6183_), .Y(core__abc_21302_new_n6184_));
AOI21X1 AOI21X1_912 ( .A(core__abc_21302_new_n5947_), .B(core__abc_21302_new_n5001_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n6188_));
AOI21X1 AOI21X1_913 ( .A(core_v1_reg_27_), .B(core__abc_21302_new_n5998__bF_buf1), .C(core__abc_21302_new_n6190_), .Y(core__abc_21302_new_n6191_));
AOI21X1 AOI21X1_914 ( .A(core__abc_21302_new_n6189_), .B(core__abc_21302_new_n6191_), .C(core__abc_21302_new_n6192_), .Y(core__0v1_reg_63_0__27_));
AOI21X1 AOI21X1_915 ( .A(core_key_92_), .B(core__abc_21302_new_n2639__bF_buf3), .C(core__abc_21302_new_n6197_), .Y(core__abc_21302_new_n6198_));
AOI21X1 AOI21X1_916 ( .A(core__abc_21302_new_n6196_), .B(core__abc_21302_new_n6198_), .C(core__abc_21302_new_n6199_), .Y(core__0v1_reg_63_0__28_));
AOI21X1 AOI21X1_917 ( .A(core__abc_21302_new_n5970_), .B(core__abc_21302_new_n4979_), .C(core__abc_21302_new_n2673__bF_buf10), .Y(core__abc_21302_new_n6201_));
AOI21X1 AOI21X1_918 ( .A(core_v1_reg_29_), .B(core__abc_21302_new_n5998__bF_buf0), .C(core__abc_21302_new_n6203_), .Y(core__abc_21302_new_n6204_));
AOI21X1 AOI21X1_919 ( .A(core__abc_21302_new_n6202_), .B(core__abc_21302_new_n6204_), .C(core__abc_21302_new_n6205_), .Y(core__0v1_reg_63_0__29_));
AOI21X1 AOI21X1_92 ( .A(_abc_19873_new_n1524__bF_buf10), .B(_abc_19873_new_n1411_), .C(_abc_19873_new_n1676_), .Y(_0word2_reg_31_0__26_));
AOI21X1 AOI21X1_920 ( .A(core__abc_21302_new_n5979_), .B(core__abc_21302_new_n4977_), .C(core__abc_21302_new_n2673__bF_buf9), .Y(core__abc_21302_new_n6208_));
AOI21X1 AOI21X1_921 ( .A(core__abc_21302_new_n6211_), .B(core__abc_21302_new_n6009__bF_buf4), .C(core__abc_21302_new_n6212_), .Y(core__0v1_reg_63_0__30_));
AOI21X1 AOI21X1_922 ( .A(core__abc_21302_new_n5989_), .B(core__abc_21302_new_n4971_), .C(core__abc_21302_new_n2673__bF_buf8), .Y(core__abc_21302_new_n6214_));
AOI21X1 AOI21X1_923 ( .A(core__abc_21302_new_n6215_), .B(core__abc_21302_new_n6217_), .C(core__abc_21302_new_n6218_), .Y(core__0v1_reg_63_0__31_));
AOI21X1 AOI21X1_924 ( .A(core__abc_21302_new_n3937_), .B(core__abc_21302_new_n2639__bF_buf2), .C(core__abc_21302_new_n6223_), .Y(core__abc_21302_new_n6224_));
AOI21X1 AOI21X1_925 ( .A(core__abc_21302_new_n6222_), .B(core__abc_21302_new_n6224_), .C(core__abc_21302_new_n6225_), .Y(core__0v1_reg_63_0__32_));
AOI21X1 AOI21X1_926 ( .A(core__abc_21302_new_n5097_), .B(core__abc_21302_new_n4946_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n6227_));
AOI21X1 AOI21X1_927 ( .A(core_key_97_), .B(core__abc_21302_new_n2639__bF_buf1), .C(core__abc_21302_new_n6229_), .Y(core__abc_21302_new_n6230_));
AOI21X1 AOI21X1_928 ( .A(core__abc_21302_new_n6228_), .B(core__abc_21302_new_n6230_), .C(core__abc_21302_new_n6231_), .Y(core__0v1_reg_63_0__33_));
AOI21X1 AOI21X1_929 ( .A(core__abc_21302_new_n5124_), .B(core__abc_21302_new_n4945_), .C(core__abc_21302_new_n2673__bF_buf6), .Y(core__abc_21302_new_n6233_));
AOI21X1 AOI21X1_93 ( .A(_abc_19873_new_n1524__bF_buf8), .B(_abc_19873_new_n1439_), .C(_abc_19873_new_n1678_), .Y(_0word2_reg_31_0__27_));
AOI21X1 AOI21X1_930 ( .A(core__abc_21302_new_n6236_), .B(core__abc_21302_new_n6009__bF_buf6), .C(core__abc_21302_new_n6237_), .Y(core__0v1_reg_63_0__34_));
AOI21X1 AOI21X1_931 ( .A(core__abc_21302_new_n5145_), .B(core__abc_21302_new_n4930_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n6239_));
AOI21X1 AOI21X1_932 ( .A(core_v1_reg_35_), .B(core__abc_21302_new_n5998__bF_buf3), .C(core__abc_21302_new_n6241_), .Y(core__abc_21302_new_n6242_));
AOI21X1 AOI21X1_933 ( .A(core__abc_21302_new_n6240_), .B(core__abc_21302_new_n6242_), .C(core__abc_21302_new_n6243_), .Y(core__0v1_reg_63_0__35_));
AOI21X1 AOI21X1_934 ( .A(core__abc_21302_new_n5168_), .B(core__abc_21302_new_n6245_), .C(core__abc_21302_new_n2673__bF_buf4), .Y(core__abc_21302_new_n6246_));
AOI21X1 AOI21X1_935 ( .A(core__abc_21302_new_n6249_), .B(core__abc_21302_new_n6009__bF_buf2), .C(core__abc_21302_new_n6250_), .Y(core__0v1_reg_63_0__36_));
AOI21X1 AOI21X1_936 ( .A(core__abc_21302_new_n5181_), .B(core__abc_21302_new_n4925_), .C(core__abc_21302_new_n2673__bF_buf3), .Y(core__abc_21302_new_n6252_));
AOI21X1 AOI21X1_937 ( .A(core_v1_reg_37_), .B(core__abc_21302_new_n5998__bF_buf2), .C(core__abc_21302_new_n6254_), .Y(core__abc_21302_new_n6255_));
AOI21X1 AOI21X1_938 ( .A(core__abc_21302_new_n6253_), .B(core__abc_21302_new_n6255_), .C(core__abc_21302_new_n6256_), .Y(core__0v1_reg_63_0__37_));
AOI21X1 AOI21X1_939 ( .A(core_v1_reg_38_), .B(core__abc_21302_new_n5998__bF_buf1), .C(core__abc_21302_new_n6261_), .Y(core__abc_21302_new_n6262_));
AOI21X1 AOI21X1_94 ( .A(_abc_19873_new_n1524__bF_buf6), .B(_abc_19873_new_n1680_), .C(_abc_19873_new_n1681_), .Y(_0word2_reg_31_0__28_));
AOI21X1 AOI21X1_940 ( .A(core__abc_21302_new_n6260_), .B(core__abc_21302_new_n6262_), .C(core__abc_21302_new_n6263_), .Y(core__0v1_reg_63_0__38_));
AOI21X1 AOI21X1_941 ( .A(core_key_103_), .B(core__abc_21302_new_n2639__bF_buf0), .C(core__abc_21302_new_n6270_), .Y(core__abc_21302_new_n6271_));
AOI21X1 AOI21X1_942 ( .A(core__abc_21302_new_n6269_), .B(core__abc_21302_new_n6271_), .C(core__abc_21302_new_n6272_), .Y(core__0v1_reg_63_0__39_));
AOI21X1 AOI21X1_943 ( .A(core__abc_21302_new_n6279_), .B(core__abc_21302_new_n6009__bF_buf4), .C(core__abc_21302_new_n6280_), .Y(core__0v1_reg_63_0__40_));
AOI21X1 AOI21X1_944 ( .A(core__abc_21302_new_n5256_), .B(core__abc_21302_new_n6282_), .C(core__abc_21302_new_n2673__bF_buf2), .Y(core__abc_21302_new_n6283_));
AOI21X1 AOI21X1_945 ( .A(core__abc_21302_new_n4212_), .B(core__abc_21302_new_n2639__bF_buf6), .C(core__abc_21302_new_n6285_), .Y(core__abc_21302_new_n6286_));
AOI21X1 AOI21X1_946 ( .A(core__abc_21302_new_n6284_), .B(core__abc_21302_new_n6286_), .C(core__abc_21302_new_n6287_), .Y(core__0v1_reg_63_0__41_));
AOI21X1 AOI21X1_947 ( .A(core__abc_21302_new_n5278_), .B(core__abc_21302_new_n4869_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n6289_));
AOI21X1 AOI21X1_948 ( .A(core_key_106_), .B(core__abc_21302_new_n2639__bF_buf5), .C(core__abc_21302_new_n6291_), .Y(core__abc_21302_new_n6292_));
AOI21X1 AOI21X1_949 ( .A(core__abc_21302_new_n6290_), .B(core__abc_21302_new_n6292_), .C(core__abc_21302_new_n6293_), .Y(core__0v1_reg_63_0__42_));
AOI21X1 AOI21X1_95 ( .A(_abc_19873_new_n1524__bF_buf4), .B(_abc_19873_new_n1471_), .C(_abc_19873_new_n1683_), .Y(_0word2_reg_31_0__29_));
AOI21X1 AOI21X1_950 ( .A(core__abc_21302_new_n5296_), .B(core__abc_21302_new_n4864_), .C(core__abc_21302_new_n2673__bF_buf0), .Y(core__abc_21302_new_n6295_));
AOI21X1 AOI21X1_951 ( .A(core_v1_reg_43_), .B(core__abc_21302_new_n5998__bF_buf3), .C(core__abc_21302_new_n6297_), .Y(core__abc_21302_new_n6298_));
AOI21X1 AOI21X1_952 ( .A(core__abc_21302_new_n6296_), .B(core__abc_21302_new_n6298_), .C(core__abc_21302_new_n6299_), .Y(core__0v1_reg_63_0__43_));
AOI21X1 AOI21X1_953 ( .A(core__abc_21302_new_n4294_), .B(core__abc_21302_new_n2639__bF_buf4), .C(core__abc_21302_new_n6305_), .Y(core__abc_21302_new_n6306_));
AOI21X1 AOI21X1_954 ( .A(core__abc_21302_new_n6303_), .B(core__abc_21302_new_n6306_), .C(core__abc_21302_new_n6307_), .Y(core__0v1_reg_63_0__44_));
AOI21X1 AOI21X1_955 ( .A(core_v1_reg_45_), .B(core__abc_21302_new_n5998__bF_buf2), .C(core__abc_21302_new_n6312_), .Y(core__abc_21302_new_n6313_));
AOI21X1 AOI21X1_956 ( .A(core__abc_21302_new_n6311_), .B(core__abc_21302_new_n6313_), .C(core__abc_21302_new_n6314_), .Y(core__0v1_reg_63_0__45_));
AOI21X1 AOI21X1_957 ( .A(core__abc_21302_new_n5362_), .B(core__abc_21302_new_n6317_), .C(core__abc_21302_new_n2673__bF_buf11), .Y(core__abc_21302_new_n6318_));
AOI21X1 AOI21X1_958 ( .A(core_v1_reg_46_), .B(core__abc_21302_new_n5998__bF_buf1), .C(core__abc_21302_new_n6320_), .Y(core__abc_21302_new_n6321_));
AOI21X1 AOI21X1_959 ( .A(core__abc_21302_new_n6319_), .B(core__abc_21302_new_n6321_), .C(core__abc_21302_new_n6322_), .Y(core__0v1_reg_63_0__46_));
AOI21X1 AOI21X1_96 ( .A(_abc_19873_new_n1524__bF_buf2), .B(_abc_19873_new_n1685_), .C(_abc_19873_new_n1686_), .Y(_0word2_reg_31_0__30_));
AOI21X1 AOI21X1_960 ( .A(core__abc_21302_new_n5381_), .B(core__abc_21302_new_n4836_), .C(core__abc_21302_new_n2673__bF_buf10), .Y(core__abc_21302_new_n6324_));
AOI21X1 AOI21X1_961 ( .A(core_v1_reg_47_), .B(core__abc_21302_new_n5998__bF_buf0), .C(core__abc_21302_new_n6326_), .Y(core__abc_21302_new_n6327_));
AOI21X1 AOI21X1_962 ( .A(core__abc_21302_new_n6325_), .B(core__abc_21302_new_n6327_), .C(core__abc_21302_new_n6328_), .Y(core__0v1_reg_63_0__47_));
AOI21X1 AOI21X1_963 ( .A(core__abc_21302_new_n6334_), .B(core__abc_21302_new_n6009__bF_buf8), .C(core__abc_21302_new_n6335_), .Y(core__0v1_reg_63_0__48_));
AOI21X1 AOI21X1_964 ( .A(core__abc_21302_new_n5427_), .B(core__abc_21302_new_n6337_), .C(core__abc_21302_new_n2673__bF_buf9), .Y(core__abc_21302_new_n6338_));
AOI21X1 AOI21X1_965 ( .A(core__abc_21302_new_n4437_), .B(core__abc_21302_new_n2639__bF_buf3), .C(core__abc_21302_new_n6340_), .Y(core__abc_21302_new_n6341_));
AOI21X1 AOI21X1_966 ( .A(core__abc_21302_new_n6339_), .B(core__abc_21302_new_n6341_), .C(core__abc_21302_new_n6342_), .Y(core__0v1_reg_63_0__49_));
AOI21X1 AOI21X1_967 ( .A(core_v1_reg_50_), .B(core__abc_21302_new_n5998__bF_buf3), .C(core__abc_21302_new_n6348_), .Y(core__abc_21302_new_n6349_));
AOI21X1 AOI21X1_968 ( .A(core__abc_21302_new_n6347_), .B(core__abc_21302_new_n6349_), .C(core__abc_21302_new_n6350_), .Y(core__0v1_reg_63_0__50_));
AOI21X1 AOI21X1_969 ( .A(core__abc_21302_new_n5459_), .B(core__abc_21302_new_n5133_), .C(core__abc_21302_new_n2673__bF_buf8), .Y(core__abc_21302_new_n6352_));
AOI21X1 AOI21X1_97 ( .A(_abc_19873_new_n1524__bF_buf0), .B(_abc_19873_new_n1514_), .C(_abc_19873_new_n1688_), .Y(_0word2_reg_31_0__31_));
AOI21X1 AOI21X1_970 ( .A(core__abc_21302_new_n4486_), .B(core__abc_21302_new_n2639__bF_buf2), .C(core__abc_21302_new_n6355_), .Y(core__abc_21302_new_n6356_));
AOI21X1 AOI21X1_971 ( .A(core__abc_21302_new_n6353_), .B(core__abc_21302_new_n6356_), .C(core__abc_21302_new_n6357_), .Y(core__0v1_reg_63_0__51_));
AOI21X1 AOI21X1_972 ( .A(core__abc_21302_new_n5501_), .B(core__abc_21302_new_n5151_), .C(core__abc_21302_new_n2673__bF_buf7), .Y(core__abc_21302_new_n6366_));
AOI21X1 AOI21X1_973 ( .A(core_v1_reg_53_), .B(core__abc_21302_new_n5998__bF_buf2), .C(core__abc_21302_new_n6368_), .Y(core__abc_21302_new_n6369_));
AOI21X1 AOI21X1_974 ( .A(core__abc_21302_new_n6367_), .B(core__abc_21302_new_n6369_), .C(core__abc_21302_new_n6370_), .Y(core__0v1_reg_63_0__53_));
AOI21X1 AOI21X1_975 ( .A(core__abc_21302_new_n5522_), .B(core__abc_21302_new_n5176_), .C(core__abc_21302_new_n2673__bF_buf6), .Y(core__abc_21302_new_n6372_));
AOI21X1 AOI21X1_976 ( .A(core_v1_reg_54_), .B(core__abc_21302_new_n5998__bF_buf1), .C(core__abc_21302_new_n6374_), .Y(core__abc_21302_new_n6375_));
AOI21X1 AOI21X1_977 ( .A(core__abc_21302_new_n6373_), .B(core__abc_21302_new_n6375_), .C(core__abc_21302_new_n6376_), .Y(core__0v1_reg_63_0__54_));
AOI21X1 AOI21X1_978 ( .A(core_key_119_), .B(core__abc_21302_new_n2639__bF_buf1), .C(core__abc_21302_new_n6383_), .Y(core__abc_21302_new_n6384_));
AOI21X1 AOI21X1_979 ( .A(core__abc_21302_new_n6382_), .B(core__abc_21302_new_n6384_), .C(core__abc_21302_new_n6385_), .Y(core__0v1_reg_63_0__55_));
AOI21X1 AOI21X1_98 ( .A(_abc_19873_new_n922_), .B(_abc_19873_new_n1524__bF_buf14), .C(_abc_19873_new_n1690_), .Y(_0word1_reg_31_0__0_));
AOI21X1 AOI21X1_980 ( .A(core__abc_21302_new_n5563_), .B(core__abc_21302_new_n5231_), .C(core__abc_21302_new_n2673__bF_buf5), .Y(core__abc_21302_new_n6387_));
AOI21X1 AOI21X1_981 ( .A(core__abc_21302_new_n6388_), .B(core__abc_21302_new_n6390_), .C(core__abc_21302_new_n6391_), .Y(core__0v1_reg_63_0__56_));
AOI21X1 AOI21X1_982 ( .A(core__abc_21302_new_n6395_), .B(core__abc_21302_new_n5237_), .C(core__abc_21302_new_n2673__bF_buf4), .Y(core__abc_21302_new_n6396_));
AOI21X1 AOI21X1_983 ( .A(core_key_121_), .B(core__abc_21302_new_n2639__bF_buf0), .C(core__abc_21302_new_n6398_), .Y(core__abc_21302_new_n6399_));
AOI21X1 AOI21X1_984 ( .A(core__abc_21302_new_n6397_), .B(core__abc_21302_new_n6399_), .C(core__abc_21302_new_n6400_), .Y(core__0v1_reg_63_0__57_));
AOI21X1 AOI21X1_985 ( .A(core__abc_21302_new_n5595_), .B(core__abc_21302_new_n5252_), .C(core__abc_21302_new_n2673__bF_buf3), .Y(core__abc_21302_new_n6402_));
AOI21X1 AOI21X1_986 ( .A(core_v1_reg_58_), .B(core__abc_21302_new_n5998__bF_buf0), .C(core__abc_21302_new_n6404_), .Y(core__abc_21302_new_n6405_));
AOI21X1 AOI21X1_987 ( .A(core__abc_21302_new_n6403_), .B(core__abc_21302_new_n6405_), .C(core__abc_21302_new_n6406_), .Y(core__0v1_reg_63_0__58_));
AOI21X1 AOI21X1_988 ( .A(core_v1_reg_59_), .B(core__abc_21302_new_n5998__bF_buf3), .C(core__abc_21302_new_n6414_), .Y(core__abc_21302_new_n6415_));
AOI21X1 AOI21X1_989 ( .A(core__abc_21302_new_n6413_), .B(core__abc_21302_new_n6415_), .C(core__abc_21302_new_n6416_), .Y(core__0v1_reg_63_0__59_));
AOI21X1 AOI21X1_99 ( .A(_abc_19873_new_n948_), .B(_abc_19873_new_n1524__bF_buf12), .C(_abc_19873_new_n1692_), .Y(_0word1_reg_31_0__1_));
AOI21X1 AOI21X1_990 ( .A(core__abc_21302_new_n5638_), .B(core__abc_21302_new_n6419_), .C(core__abc_21302_new_n2673__bF_buf2), .Y(core__abc_21302_new_n6420_));
AOI21X1 AOI21X1_991 ( .A(core_v1_reg_60_), .B(core__abc_21302_new_n5998__bF_buf2), .C(core__abc_21302_new_n6423_), .Y(core__abc_21302_new_n6424_));
AOI21X1 AOI21X1_992 ( .A(core__abc_21302_new_n6421_), .B(core__abc_21302_new_n6424_), .C(core__abc_21302_new_n6425_), .Y(core__0v1_reg_63_0__60_));
AOI21X1 AOI21X1_993 ( .A(core__abc_21302_new_n5657_), .B(core__abc_21302_new_n5312_), .C(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n6427_));
AOI21X1 AOI21X1_994 ( .A(core_v1_reg_61_), .B(core__abc_21302_new_n5998__bF_buf1), .C(core__abc_21302_new_n6429_), .Y(core__abc_21302_new_n6430_));
AOI21X1 AOI21X1_995 ( .A(core__abc_21302_new_n6428_), .B(core__abc_21302_new_n6430_), .C(core__abc_21302_new_n6431_), .Y(core__0v1_reg_63_0__61_));
AOI21X1 AOI21X1_996 ( .A(core__abc_21302_new_n5677_), .B(core__abc_21302_new_n5328_), .C(core__abc_21302_new_n2673__bF_buf0), .Y(core__abc_21302_new_n6433_));
AOI21X1 AOI21X1_997 ( .A(core_v1_reg_62_), .B(core__abc_21302_new_n5998__bF_buf0), .C(core__abc_21302_new_n6435_), .Y(core__abc_21302_new_n6436_));
AOI21X1 AOI21X1_998 ( .A(core__abc_21302_new_n6434_), .B(core__abc_21302_new_n6436_), .C(core__abc_21302_new_n6437_), .Y(core__0v1_reg_63_0__62_));
AOI21X1 AOI21X1_999 ( .A(core_key_127_), .B(core__abc_21302_new_n2639__bF_buf6), .C(core__abc_21302_new_n6444_), .Y(core__abc_21302_new_n6445_));
AOI22X1 AOI22X1_1 ( .A(core_loop_ctr_reg_0_), .B(core_compression_rounds_0_), .C(core__abc_21302_new_n1135_), .D(core__abc_21302_new_n1132_), .Y(core__abc_21302_new_n1136_));
AOI22X1 AOI22X1_10 ( .A(core__abc_21302_new_n3891_), .B(core__abc_21302_new_n3916_), .C(core__abc_21302_new_n3856_), .D(core__abc_21302_new_n4166_), .Y(core__abc_21302_new_n4168_));
AOI22X1 AOI22X1_11 ( .A(core__abc_21302_new_n4392_), .B(core__abc_21302_new_n4391_), .C(core__abc_21302_new_n4328_), .D(core__abc_21302_new_n4386_), .Y(core__abc_21302_new_n4393_));
AOI22X1 AOI22X1_12 ( .A(core__abc_21302_new_n4599_), .B(core__abc_21302_new_n4600_), .C(core__abc_21302_new_n4542_), .D(core__abc_21302_new_n4595_), .Y(core__abc_21302_new_n4601_));
AOI22X1 AOI22X1_13 ( .A(core__abc_21302_new_n4776_), .B(core__abc_21302_new_n4778_), .C(core__abc_21302_new_n4767_), .D(core__abc_21302_new_n4765_), .Y(core__abc_21302_new_n4788_));
AOI22X1 AOI22X1_14 ( .A(core__abc_21302_new_n2365__bF_buf2), .B(core__abc_21302_new_n5169_), .C(core_key_4_), .D(core__abc_21302_new_n2639__bF_buf6), .Y(core__abc_21302_new_n5170_));
AOI22X1 AOI22X1_15 ( .A(core_v2_reg_4_), .B(core__abc_21302_new_n5085__bF_buf1), .C(core__abc_21302_new_n2362__bF_buf1), .D(core__abc_21302_new_n5171_), .Y(core__abc_21302_new_n5172_));
AOI22X1 AOI22X1_16 ( .A(core__abc_21302_new_n5230_), .B(core__abc_21302_new_n5232_), .C(core__abc_21302_new_n5226_), .D(core__abc_21302_new_n5193_), .Y(core__abc_21302_new_n5233_));
AOI22X1 AOI22X1_17 ( .A(core_v2_reg_8_), .B(core__abc_21302_new_n2365__bF_buf1), .C(core_key_8_), .D(core__abc_21302_new_n2639__bF_buf5), .Y(core__abc_21302_new_n5243_));
AOI22X1 AOI22X1_18 ( .A(core_v2_reg_9_), .B(core__abc_21302_new_n2365__bF_buf0), .C(core__abc_21302_new_n2634__bF_buf1), .D(core__abc_21302_new_n5256_), .Y(core__abc_21302_new_n5257_));
AOI22X1 AOI22X1_19 ( .A(core_v2_reg_10_), .B(core__abc_21302_new_n2365__bF_buf4), .C(core_key_10_), .D(core__abc_21302_new_n2639__bF_buf4), .Y(core__abc_21302_new_n5280_));
AOI22X1 AOI22X1_2 ( .A(core__abc_21302_new_n2138_), .B(core__abc_21302_new_n2361_), .C(core__abc_21302_new_n1183_), .D(core__abc_21302_new_n2165_), .Y(core__abc_21302_new_n2362_));
AOI22X1 AOI22X1_20 ( .A(core_v2_reg_12_), .B(core__abc_21302_new_n2365__bF_buf3), .C(core__abc_21302_new_n2634__bF_buf8), .D(core__abc_21302_new_n5316_), .Y(core__abc_21302_new_n5317_));
AOI22X1 AOI22X1_21 ( .A(core_v2_reg_16_), .B(core__abc_21302_new_n2365__bF_buf2), .C(core__abc_21302_new_n2634__bF_buf6), .D(core__abc_21302_new_n5409_), .Y(core__abc_21302_new_n5410_));
AOI22X1 AOI22X1_22 ( .A(core_v2_reg_43_), .B(core__abc_21302_new_n2365__bF_buf4), .C(core_key_43_), .D(core__abc_21302_new_n2639__bF_buf4), .Y(core__abc_21302_new_n5793_));
AOI22X1 AOI22X1_23 ( .A(core_v2_reg_51_), .B(core__abc_21302_new_n2365__bF_buf0), .C(core__abc_21302_new_n2634__bF_buf3), .D(core__abc_21302_new_n5872_), .Y(core__abc_21302_new_n5873_));
AOI22X1 AOI22X1_24 ( .A(core_v2_reg_52_), .B(core__abc_21302_new_n2365__bF_buf4), .C(core__abc_21302_new_n2634__bF_buf2), .D(core__abc_21302_new_n5883_), .Y(core__abc_21302_new_n5884_));
AOI22X1 AOI22X1_25 ( .A(core_v2_reg_53_), .B(core__abc_21302_new_n2365__bF_buf3), .C(core__abc_21302_new_n2634__bF_buf1), .D(core__abc_21302_new_n5893_), .Y(core__abc_21302_new_n5894_));
AOI22X1 AOI22X1_26 ( .A(core_v2_reg_56_), .B(core__abc_21302_new_n2365__bF_buf2), .C(core_key_56_), .D(core__abc_21302_new_n2639__bF_buf0), .Y(core__abc_21302_new_n5925_));
AOI22X1 AOI22X1_27 ( .A(core_v2_reg_57_), .B(core__abc_21302_new_n2365__bF_buf1), .C(core_key_57_), .D(core__abc_21302_new_n2639__bF_buf6), .Y(core__abc_21302_new_n5933_));
AOI22X1 AOI22X1_28 ( .A(core_v2_reg_58_), .B(core__abc_21302_new_n2365__bF_buf0), .C(core__abc_21302_new_n2634__bF_buf7), .D(core__abc_21302_new_n5938_), .Y(core__abc_21302_new_n5939_));
AOI22X1 AOI22X1_29 ( .A(core__abc_21302_new_n5998__bF_buf2), .B(core__abc_21302_new_n2471_), .C(core__abc_21302_new_n2639__bF_buf3), .D(core__abc_21302_new_n6017_), .Y(core__abc_21302_new_n6018_));
AOI22X1 AOI22X1_3 ( .A(core__abc_21302_new_n2410_), .B(core__abc_21302_new_n2488_), .C(core__abc_21302_new_n2484_), .D(core__abc_21302_new_n2487_), .Y(core__abc_21302_new_n2489_));
AOI22X1 AOI22X1_4 ( .A(core__abc_21302_new_n3538_), .B(core__abc_21302_new_n3541_), .C(core__abc_21302_new_n3540_), .D(core__abc_21302_new_n3501_), .Y(core__abc_21302_new_n3542_));
AOI22X1 AOI22X1_5 ( .A(core__abc_21302_new_n3582_), .B(core__abc_21302_new_n3586_), .C(core__abc_21302_new_n3589_), .D(core__abc_21302_new_n3590_), .Y(core__abc_21302_new_n3591_));
AOI22X1 AOI22X1_6 ( .A(core__abc_21302_new_n3673_), .B(core__abc_21302_new_n3692_), .C(core__abc_21302_new_n3691_), .D(core__abc_21302_new_n3689_), .Y(core__abc_21302_new_n3693_));
AOI22X1 AOI22X1_7 ( .A(core__abc_21302_new_n1538_), .B(core__abc_21302_new_n3836_), .C(core__abc_21302_new_n2550_), .D(core__abc_21302_new_n3776_), .Y(core__abc_21302_new_n3837_));
AOI22X1 AOI22X1_8 ( .A(core__abc_21302_new_n4158_), .B(core__abc_21302_new_n4159_), .C(core__abc_21302_new_n4095_), .D(core__abc_21302_new_n4155_), .Y(core__abc_21302_new_n4160_));
AOI22X1 AOI22X1_9 ( .A(core__abc_21302_new_n3886_), .B(core__abc_21302_new_n3889_), .C(core__abc_21302_new_n3880_), .D(core__abc_21302_new_n3882_), .Y(core__abc_21302_new_n4165_));
BUFX2 BUFX2_1 ( .A(_abc_19873_new_n905_), .Y(_abc_19873_new_n905__bF_buf2));
BUFX2 BUFX2_10 ( .A(_auto_iopadmap_cc_368_execute_27087_6_), .Y(\read_data[6] ));
BUFX2 BUFX2_11 ( .A(_auto_iopadmap_cc_368_execute_27087_7_), .Y(\read_data[7] ));
BUFX2 BUFX2_12 ( .A(_auto_iopadmap_cc_368_execute_27087_8_), .Y(\read_data[8] ));
BUFX2 BUFX2_13 ( .A(_auto_iopadmap_cc_368_execute_27087_9_), .Y(\read_data[9] ));
BUFX2 BUFX2_14 ( .A(_auto_iopadmap_cc_368_execute_27087_10_), .Y(\read_data[10] ));
BUFX2 BUFX2_15 ( .A(_auto_iopadmap_cc_368_execute_27087_11_), .Y(\read_data[11] ));
BUFX2 BUFX2_16 ( .A(_auto_iopadmap_cc_368_execute_27087_12_), .Y(\read_data[12] ));
BUFX2 BUFX2_17 ( .A(_auto_iopadmap_cc_368_execute_27087_13_), .Y(\read_data[13] ));
BUFX2 BUFX2_18 ( .A(_auto_iopadmap_cc_368_execute_27087_14_), .Y(\read_data[14] ));
BUFX2 BUFX2_19 ( .A(_auto_iopadmap_cc_368_execute_27087_15_), .Y(\read_data[15] ));
BUFX2 BUFX2_2 ( .A(_abc_19873_new_n905_), .Y(_abc_19873_new_n905__bF_buf1));
BUFX2 BUFX2_20 ( .A(_auto_iopadmap_cc_368_execute_27087_16_), .Y(\read_data[16] ));
BUFX2 BUFX2_21 ( .A(_auto_iopadmap_cc_368_execute_27087_17_), .Y(\read_data[17] ));
BUFX2 BUFX2_22 ( .A(_auto_iopadmap_cc_368_execute_27087_18_), .Y(\read_data[18] ));
BUFX2 BUFX2_23 ( .A(_auto_iopadmap_cc_368_execute_27087_19_), .Y(\read_data[19] ));
BUFX2 BUFX2_24 ( .A(_auto_iopadmap_cc_368_execute_27087_20_), .Y(\read_data[20] ));
BUFX2 BUFX2_25 ( .A(_auto_iopadmap_cc_368_execute_27087_21_), .Y(\read_data[21] ));
BUFX2 BUFX2_26 ( .A(_auto_iopadmap_cc_368_execute_27087_22_), .Y(\read_data[22] ));
BUFX2 BUFX2_27 ( .A(_auto_iopadmap_cc_368_execute_27087_23_), .Y(\read_data[23] ));
BUFX2 BUFX2_28 ( .A(_auto_iopadmap_cc_368_execute_27087_24_), .Y(\read_data[24] ));
BUFX2 BUFX2_29 ( .A(_auto_iopadmap_cc_368_execute_27087_25_), .Y(\read_data[25] ));
BUFX2 BUFX2_3 ( .A(_abc_19873_new_n905_), .Y(_abc_19873_new_n905__bF_buf0));
BUFX2 BUFX2_30 ( .A(_auto_iopadmap_cc_368_execute_27087_26_), .Y(\read_data[26] ));
BUFX2 BUFX2_31 ( .A(_auto_iopadmap_cc_368_execute_27087_27_), .Y(\read_data[27] ));
BUFX2 BUFX2_32 ( .A(_auto_iopadmap_cc_368_execute_27087_28_), .Y(\read_data[28] ));
BUFX2 BUFX2_33 ( .A(_auto_iopadmap_cc_368_execute_27087_29_), .Y(\read_data[29] ));
BUFX2 BUFX2_34 ( .A(_auto_iopadmap_cc_368_execute_27087_30_), .Y(\read_data[30] ));
BUFX2 BUFX2_35 ( .A(_auto_iopadmap_cc_368_execute_27087_31_), .Y(\read_data[31] ));
BUFX2 BUFX2_4 ( .A(_auto_iopadmap_cc_368_execute_27087_0_), .Y(\read_data[0] ));
BUFX2 BUFX2_5 ( .A(_auto_iopadmap_cc_368_execute_27087_1_), .Y(\read_data[1] ));
BUFX2 BUFX2_6 ( .A(_auto_iopadmap_cc_368_execute_27087_2_), .Y(\read_data[2] ));
BUFX2 BUFX2_7 ( .A(_auto_iopadmap_cc_368_execute_27087_3_), .Y(\read_data[3] ));
BUFX2 BUFX2_8 ( .A(_auto_iopadmap_cc_368_execute_27087_4_), .Y(\read_data[4] ));
BUFX2 BUFX2_9 ( .A(_auto_iopadmap_cc_368_execute_27087_5_), .Y(\read_data[5] ));
BUFX4 BUFX4_1 ( .A(clk), .Y(clk_hier0_bF_buf8));
BUFX4 BUFX4_10 ( .A(reset_n), .Y(reset_n_hier0_bF_buf7));
BUFX4 BUFX4_100 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf38));
BUFX4 BUFX4_101 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf37));
BUFX4 BUFX4_102 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf36));
BUFX4 BUFX4_103 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf35));
BUFX4 BUFX4_104 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf34));
BUFX4 BUFX4_105 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf33));
BUFX4 BUFX4_106 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf32));
BUFX4 BUFX4_107 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf31));
BUFX4 BUFX4_108 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf30));
BUFX4 BUFX4_109 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf29));
BUFX4 BUFX4_11 ( .A(reset_n), .Y(reset_n_hier0_bF_buf6));
BUFX4 BUFX4_110 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf28));
BUFX4 BUFX4_111 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf27));
BUFX4 BUFX4_112 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf26));
BUFX4 BUFX4_113 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf25));
BUFX4 BUFX4_114 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf24));
BUFX4 BUFX4_115 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf23));
BUFX4 BUFX4_116 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf22));
BUFX4 BUFX4_117 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf21));
BUFX4 BUFX4_118 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf20));
BUFX4 BUFX4_119 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf19));
BUFX4 BUFX4_12 ( .A(reset_n), .Y(reset_n_hier0_bF_buf5));
BUFX4 BUFX4_120 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf18));
BUFX4 BUFX4_121 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf17));
BUFX4 BUFX4_122 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf16));
BUFX4 BUFX4_123 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf15));
BUFX4 BUFX4_124 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf14));
BUFX4 BUFX4_125 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf13));
BUFX4 BUFX4_126 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf12));
BUFX4 BUFX4_127 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf11));
BUFX4 BUFX4_128 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf10));
BUFX4 BUFX4_129 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf9));
BUFX4 BUFX4_13 ( .A(reset_n), .Y(reset_n_hier0_bF_buf4));
BUFX4 BUFX4_130 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf8));
BUFX4 BUFX4_131 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf7));
BUFX4 BUFX4_132 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf6));
BUFX4 BUFX4_133 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf5));
BUFX4 BUFX4_134 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf4));
BUFX4 BUFX4_135 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf3));
BUFX4 BUFX4_136 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf2));
BUFX4 BUFX4_137 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf1));
BUFX4 BUFX4_138 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf0));
BUFX4 BUFX4_139 ( .A(_abc_19873_new_n895_), .Y(_abc_19873_new_n895__bF_buf4));
BUFX4 BUFX4_14 ( .A(reset_n), .Y(reset_n_hier0_bF_buf3));
BUFX4 BUFX4_140 ( .A(_abc_19873_new_n895_), .Y(_abc_19873_new_n895__bF_buf3));
BUFX4 BUFX4_141 ( .A(_abc_19873_new_n895_), .Y(_abc_19873_new_n895__bF_buf2));
BUFX4 BUFX4_142 ( .A(_abc_19873_new_n895_), .Y(_abc_19873_new_n895__bF_buf1));
BUFX4 BUFX4_143 ( .A(_abc_19873_new_n895_), .Y(_abc_19873_new_n895__bF_buf0));
BUFX4 BUFX4_144 ( .A(_abc_19873_new_n913_), .Y(_abc_19873_new_n913__bF_buf4));
BUFX4 BUFX4_145 ( .A(_abc_19873_new_n913_), .Y(_abc_19873_new_n913__bF_buf3));
BUFX4 BUFX4_146 ( .A(_abc_19873_new_n913_), .Y(_abc_19873_new_n913__bF_buf2));
BUFX4 BUFX4_147 ( .A(_abc_19873_new_n913_), .Y(_abc_19873_new_n913__bF_buf1));
BUFX4 BUFX4_148 ( .A(_abc_19873_new_n913_), .Y(_abc_19873_new_n913__bF_buf0));
BUFX4 BUFX4_149 ( .A(_abc_19873_new_n889_), .Y(_abc_19873_new_n889__bF_buf4));
BUFX4 BUFX4_15 ( .A(reset_n), .Y(reset_n_hier0_bF_buf2));
BUFX4 BUFX4_150 ( .A(_abc_19873_new_n889_), .Y(_abc_19873_new_n889__bF_buf3));
BUFX4 BUFX4_151 ( .A(_abc_19873_new_n889_), .Y(_abc_19873_new_n889__bF_buf2));
BUFX4 BUFX4_152 ( .A(_abc_19873_new_n889_), .Y(_abc_19873_new_n889__bF_buf1));
BUFX4 BUFX4_153 ( .A(_abc_19873_new_n889_), .Y(_abc_19873_new_n889__bF_buf0));
BUFX4 BUFX4_154 ( .A(_abc_19873_new_n1849_), .Y(_abc_19873_new_n1849__bF_buf7));
BUFX4 BUFX4_155 ( .A(_abc_19873_new_n1849_), .Y(_abc_19873_new_n1849__bF_buf6));
BUFX4 BUFX4_156 ( .A(_abc_19873_new_n1849_), .Y(_abc_19873_new_n1849__bF_buf5));
BUFX4 BUFX4_157 ( .A(_abc_19873_new_n1849_), .Y(_abc_19873_new_n1849__bF_buf4));
BUFX4 BUFX4_158 ( .A(_abc_19873_new_n1849_), .Y(_abc_19873_new_n1849__bF_buf3));
BUFX4 BUFX4_159 ( .A(_abc_19873_new_n1849_), .Y(_abc_19873_new_n1849__bF_buf2));
BUFX4 BUFX4_16 ( .A(reset_n), .Y(reset_n_hier0_bF_buf1));
BUFX4 BUFX4_160 ( .A(_abc_19873_new_n1849_), .Y(_abc_19873_new_n1849__bF_buf1));
BUFX4 BUFX4_161 ( .A(_abc_19873_new_n1849_), .Y(_abc_19873_new_n1849__bF_buf0));
BUFX4 BUFX4_162 ( .A(core__abc_21302_new_n2368_), .Y(core__abc_21302_new_n2368__bF_buf4));
BUFX4 BUFX4_163 ( .A(core__abc_21302_new_n2368_), .Y(core__abc_21302_new_n2368__bF_buf3));
BUFX4 BUFX4_164 ( .A(core__abc_21302_new_n2368_), .Y(core__abc_21302_new_n2368__bF_buf2));
BUFX4 BUFX4_165 ( .A(core__abc_21302_new_n2368_), .Y(core__abc_21302_new_n2368__bF_buf1));
BUFX4 BUFX4_166 ( .A(core__abc_21302_new_n2368_), .Y(core__abc_21302_new_n2368__bF_buf0));
BUFX4 BUFX4_167 ( .A(_abc_19873_new_n2058_), .Y(_abc_19873_new_n2058__bF_buf7));
BUFX4 BUFX4_168 ( .A(_abc_19873_new_n2058_), .Y(_abc_19873_new_n2058__bF_buf6));
BUFX4 BUFX4_169 ( .A(_abc_19873_new_n2058_), .Y(_abc_19873_new_n2058__bF_buf5));
BUFX4 BUFX4_17 ( .A(reset_n), .Y(reset_n_hier0_bF_buf0));
BUFX4 BUFX4_170 ( .A(_abc_19873_new_n2058_), .Y(_abc_19873_new_n2058__bF_buf4));
BUFX4 BUFX4_171 ( .A(_abc_19873_new_n2058_), .Y(_abc_19873_new_n2058__bF_buf3));
BUFX4 BUFX4_172 ( .A(_abc_19873_new_n2058_), .Y(_abc_19873_new_n2058__bF_buf2));
BUFX4 BUFX4_173 ( .A(_abc_19873_new_n2058_), .Y(_abc_19873_new_n2058__bF_buf1));
BUFX4 BUFX4_174 ( .A(_abc_19873_new_n2058_), .Y(_abc_19873_new_n2058__bF_buf0));
BUFX4 BUFX4_175 ( .A(core__abc_21302_new_n2365_), .Y(core__abc_21302_new_n2365__bF_buf4));
BUFX4 BUFX4_176 ( .A(core__abc_21302_new_n2365_), .Y(core__abc_21302_new_n2365__bF_buf3));
BUFX4 BUFX4_177 ( .A(core__abc_21302_new_n2365_), .Y(core__abc_21302_new_n2365__bF_buf2));
BUFX4 BUFX4_178 ( .A(core__abc_21302_new_n2365_), .Y(core__abc_21302_new_n2365__bF_buf1));
BUFX4 BUFX4_179 ( .A(core__abc_21302_new_n2365_), .Y(core__abc_21302_new_n2365__bF_buf0));
BUFX4 BUFX4_18 ( .A(_abc_19873_new_n969_), .Y(_abc_19873_new_n969__bF_buf3));
BUFX4 BUFX4_180 ( .A(_abc_19873_new_n901_), .Y(_abc_19873_new_n901__bF_buf7));
BUFX4 BUFX4_181 ( .A(_abc_19873_new_n901_), .Y(_abc_19873_new_n901__bF_buf6));
BUFX4 BUFX4_182 ( .A(_abc_19873_new_n901_), .Y(_abc_19873_new_n901__bF_buf5));
BUFX4 BUFX4_183 ( .A(_abc_19873_new_n901_), .Y(_abc_19873_new_n901__bF_buf4));
BUFX4 BUFX4_184 ( .A(_abc_19873_new_n901_), .Y(_abc_19873_new_n901__bF_buf3));
BUFX4 BUFX4_185 ( .A(_abc_19873_new_n901_), .Y(_abc_19873_new_n901__bF_buf2));
BUFX4 BUFX4_186 ( .A(_abc_19873_new_n901_), .Y(_abc_19873_new_n901__bF_buf1));
BUFX4 BUFX4_187 ( .A(_abc_19873_new_n901_), .Y(_abc_19873_new_n901__bF_buf0));
BUFX4 BUFX4_188 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf11));
BUFX4 BUFX4_189 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf10));
BUFX4 BUFX4_19 ( .A(_abc_19873_new_n969_), .Y(_abc_19873_new_n969__bF_buf2));
BUFX4 BUFX4_190 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf9));
BUFX4 BUFX4_191 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf8));
BUFX4 BUFX4_192 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf7));
BUFX4 BUFX4_193 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf6));
BUFX4 BUFX4_194 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf5));
BUFX4 BUFX4_195 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf4));
BUFX4 BUFX4_196 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf3));
BUFX4 BUFX4_197 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf2));
BUFX4 BUFX4_198 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf1));
BUFX4 BUFX4_199 ( .A(core__abc_21302_new_n2362_), .Y(core__abc_21302_new_n2362__bF_buf0));
BUFX4 BUFX4_2 ( .A(clk), .Y(clk_hier0_bF_buf7));
BUFX4 BUFX4_20 ( .A(_abc_19873_new_n969_), .Y(_abc_19873_new_n969__bF_buf1));
BUFX4 BUFX4_200 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf12));
BUFX4 BUFX4_201 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf11));
BUFX4 BUFX4_202 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf10));
BUFX4 BUFX4_203 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf9));
BUFX4 BUFX4_204 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf8));
BUFX4 BUFX4_205 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf7));
BUFX4 BUFX4_206 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf6));
BUFX4 BUFX4_207 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf5));
BUFX4 BUFX4_208 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf4));
BUFX4 BUFX4_209 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf3));
BUFX4 BUFX4_21 ( .A(_abc_19873_new_n969_), .Y(_abc_19873_new_n969__bF_buf0));
BUFX4 BUFX4_210 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf2));
BUFX4 BUFX4_211 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf1));
BUFX4 BUFX4_212 ( .A(core__abc_21302_new_n2168_), .Y(core__abc_21302_new_n2168__bF_buf0));
BUFX4 BUFX4_213 ( .A(_abc_19873_new_n1925_), .Y(_abc_19873_new_n1925__bF_buf7));
BUFX4 BUFX4_214 ( .A(_abc_19873_new_n1925_), .Y(_abc_19873_new_n1925__bF_buf6));
BUFX4 BUFX4_215 ( .A(_abc_19873_new_n1925_), .Y(_abc_19873_new_n1925__bF_buf5));
BUFX4 BUFX4_216 ( .A(_abc_19873_new_n1925_), .Y(_abc_19873_new_n1925__bF_buf4));
BUFX4 BUFX4_217 ( .A(_abc_19873_new_n1925_), .Y(_abc_19873_new_n1925__bF_buf3));
BUFX4 BUFX4_218 ( .A(_abc_19873_new_n1925_), .Y(_abc_19873_new_n1925__bF_buf2));
BUFX4 BUFX4_219 ( .A(_abc_19873_new_n1925_), .Y(_abc_19873_new_n1925__bF_buf1));
BUFX4 BUFX4_22 ( .A(core__abc_21302_new_n2639_), .Y(core__abc_21302_new_n2639__bF_buf6));
BUFX4 BUFX4_220 ( .A(_abc_19873_new_n1925_), .Y(_abc_19873_new_n1925__bF_buf0));
BUFX4 BUFX4_221 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf11));
BUFX4 BUFX4_222 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf10));
BUFX4 BUFX4_223 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf9));
BUFX4 BUFX4_224 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf8));
BUFX4 BUFX4_225 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf7));
BUFX4 BUFX4_226 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf6));
BUFX4 BUFX4_227 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf5));
BUFX4 BUFX4_228 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf4));
BUFX4 BUFX4_229 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf3));
BUFX4 BUFX4_23 ( .A(core__abc_21302_new_n2639_), .Y(core__abc_21302_new_n2639__bF_buf5));
BUFX4 BUFX4_230 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf2));
BUFX4 BUFX4_231 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf1));
BUFX4 BUFX4_232 ( .A(core__abc_21302_new_n2673_), .Y(core__abc_21302_new_n2673__bF_buf0));
BUFX4 BUFX4_233 ( .A(_abc_19873_new_n1064_), .Y(_abc_19873_new_n1064__bF_buf3));
BUFX4 BUFX4_234 ( .A(_abc_19873_new_n1064_), .Y(_abc_19873_new_n1064__bF_buf2));
BUFX4 BUFX4_235 ( .A(_abc_19873_new_n1064_), .Y(_abc_19873_new_n1064__bF_buf1));
BUFX4 BUFX4_236 ( .A(_abc_19873_new_n1064_), .Y(_abc_19873_new_n1064__bF_buf0));
BUFX4 BUFX4_237 ( .A(_abc_19873_new_n1992_), .Y(_abc_19873_new_n1992__bF_buf7));
BUFX4 BUFX4_238 ( .A(_abc_19873_new_n1992_), .Y(_abc_19873_new_n1992__bF_buf6));
BUFX4 BUFX4_239 ( .A(_abc_19873_new_n1992_), .Y(_abc_19873_new_n1992__bF_buf5));
BUFX4 BUFX4_24 ( .A(core__abc_21302_new_n2639_), .Y(core__abc_21302_new_n2639__bF_buf4));
BUFX4 BUFX4_240 ( .A(_abc_19873_new_n1992_), .Y(_abc_19873_new_n1992__bF_buf4));
BUFX4 BUFX4_241 ( .A(_abc_19873_new_n1992_), .Y(_abc_19873_new_n1992__bF_buf3));
BUFX4 BUFX4_242 ( .A(_abc_19873_new_n1992_), .Y(_abc_19873_new_n1992__bF_buf2));
BUFX4 BUFX4_243 ( .A(_abc_19873_new_n1992_), .Y(_abc_19873_new_n1992__bF_buf1));
BUFX4 BUFX4_244 ( .A(_abc_19873_new_n1992_), .Y(_abc_19873_new_n1992__bF_buf0));
BUFX4 BUFX4_245 ( .A(_abc_19873_new_n894_), .Y(_abc_19873_new_n894__bF_buf4));
BUFX4 BUFX4_246 ( .A(_abc_19873_new_n894_), .Y(_abc_19873_new_n894__bF_buf3));
BUFX4 BUFX4_247 ( .A(_abc_19873_new_n894_), .Y(_abc_19873_new_n894__bF_buf2));
BUFX4 BUFX4_248 ( .A(_abc_19873_new_n894_), .Y(_abc_19873_new_n894__bF_buf1));
BUFX4 BUFX4_249 ( .A(_abc_19873_new_n894_), .Y(_abc_19873_new_n894__bF_buf0));
BUFX4 BUFX4_25 ( .A(core__abc_21302_new_n2639_), .Y(core__abc_21302_new_n2639__bF_buf3));
BUFX4 BUFX4_250 ( .A(_abc_19873_new_n2125_), .Y(_abc_19873_new_n2125__bF_buf7));
BUFX4 BUFX4_251 ( .A(_abc_19873_new_n2125_), .Y(_abc_19873_new_n2125__bF_buf6));
BUFX4 BUFX4_252 ( .A(_abc_19873_new_n2125_), .Y(_abc_19873_new_n2125__bF_buf5));
BUFX4 BUFX4_253 ( .A(_abc_19873_new_n2125_), .Y(_abc_19873_new_n2125__bF_buf4));
BUFX4 BUFX4_254 ( .A(_abc_19873_new_n2125_), .Y(_abc_19873_new_n2125__bF_buf3));
BUFX4 BUFX4_255 ( .A(_abc_19873_new_n2125_), .Y(_abc_19873_new_n2125__bF_buf2));
BUFX4 BUFX4_256 ( .A(_abc_19873_new_n2125_), .Y(_abc_19873_new_n2125__bF_buf1));
BUFX4 BUFX4_257 ( .A(_abc_19873_new_n2125_), .Y(_abc_19873_new_n2125__bF_buf0));
BUFX4 BUFX4_258 ( .A(_abc_19873_new_n912_), .Y(_abc_19873_new_n912__bF_buf3));
BUFX4 BUFX4_259 ( .A(_abc_19873_new_n912_), .Y(_abc_19873_new_n912__bF_buf2));
BUFX4 BUFX4_26 ( .A(core__abc_21302_new_n2639_), .Y(core__abc_21302_new_n2639__bF_buf2));
BUFX4 BUFX4_260 ( .A(_abc_19873_new_n912_), .Y(_abc_19873_new_n912__bF_buf1));
BUFX4 BUFX4_261 ( .A(_abc_19873_new_n912_), .Y(_abc_19873_new_n912__bF_buf0));
BUFX4 BUFX4_262 ( .A(_abc_19873_new_n2198_), .Y(_abc_19873_new_n2198__bF_buf7));
BUFX4 BUFX4_263 ( .A(_abc_19873_new_n2198_), .Y(_abc_19873_new_n2198__bF_buf6));
BUFX4 BUFX4_264 ( .A(_abc_19873_new_n2198_), .Y(_abc_19873_new_n2198__bF_buf5));
BUFX4 BUFX4_265 ( .A(_abc_19873_new_n2198_), .Y(_abc_19873_new_n2198__bF_buf4));
BUFX4 BUFX4_266 ( .A(_abc_19873_new_n2198_), .Y(_abc_19873_new_n2198__bF_buf3));
BUFX4 BUFX4_267 ( .A(_abc_19873_new_n2198_), .Y(_abc_19873_new_n2198__bF_buf2));
BUFX4 BUFX4_268 ( .A(_abc_19873_new_n2198_), .Y(_abc_19873_new_n2198__bF_buf1));
BUFX4 BUFX4_269 ( .A(_abc_19873_new_n2198_), .Y(_abc_19873_new_n2198__bF_buf0));
BUFX4 BUFX4_27 ( .A(core__abc_21302_new_n2639_), .Y(core__abc_21302_new_n2639__bF_buf1));
BUFX4 BUFX4_270 ( .A(core__abc_21302_new_n6450_), .Y(core__abc_21302_new_n6450__bF_buf7));
BUFX4 BUFX4_271 ( .A(core__abc_21302_new_n6450_), .Y(core__abc_21302_new_n6450__bF_buf6));
BUFX4 BUFX4_272 ( .A(core__abc_21302_new_n6450_), .Y(core__abc_21302_new_n6450__bF_buf5));
BUFX4 BUFX4_273 ( .A(core__abc_21302_new_n6450_), .Y(core__abc_21302_new_n6450__bF_buf4));
BUFX4 BUFX4_274 ( .A(core__abc_21302_new_n6450_), .Y(core__abc_21302_new_n6450__bF_buf3));
BUFX4 BUFX4_275 ( .A(core__abc_21302_new_n6450_), .Y(core__abc_21302_new_n6450__bF_buf2));
BUFX4 BUFX4_276 ( .A(core__abc_21302_new_n6450_), .Y(core__abc_21302_new_n6450__bF_buf1));
BUFX4 BUFX4_277 ( .A(core__abc_21302_new_n6450_), .Y(core__abc_21302_new_n6450__bF_buf0));
BUFX4 BUFX4_278 ( .A(core__abc_21302_new_n2364_), .Y(core__abc_21302_new_n2364__bF_buf5));
BUFX4 BUFX4_279 ( .A(core__abc_21302_new_n2364_), .Y(core__abc_21302_new_n2364__bF_buf4));
BUFX4 BUFX4_28 ( .A(core__abc_21302_new_n2639_), .Y(core__abc_21302_new_n2639__bF_buf0));
BUFX4 BUFX4_280 ( .A(core__abc_21302_new_n2364_), .Y(core__abc_21302_new_n2364__bF_buf3));
BUFX4 BUFX4_281 ( .A(core__abc_21302_new_n2364_), .Y(core__abc_21302_new_n2364__bF_buf2));
BUFX4 BUFX4_282 ( .A(core__abc_21302_new_n2364_), .Y(core__abc_21302_new_n2364__bF_buf1));
BUFX4 BUFX4_283 ( .A(core__abc_21302_new_n2364_), .Y(core__abc_21302_new_n2364__bF_buf0));
BUFX4 BUFX4_284 ( .A(core__abc_21302_new_n5104_), .Y(core__abc_21302_new_n5104__bF_buf7));
BUFX4 BUFX4_285 ( .A(core__abc_21302_new_n5104_), .Y(core__abc_21302_new_n5104__bF_buf6));
BUFX4 BUFX4_286 ( .A(core__abc_21302_new_n5104_), .Y(core__abc_21302_new_n5104__bF_buf5));
BUFX4 BUFX4_287 ( .A(core__abc_21302_new_n5104_), .Y(core__abc_21302_new_n5104__bF_buf4));
BUFX4 BUFX4_288 ( .A(core__abc_21302_new_n5104_), .Y(core__abc_21302_new_n5104__bF_buf3));
BUFX4 BUFX4_289 ( .A(core__abc_21302_new_n5104_), .Y(core__abc_21302_new_n5104__bF_buf2));
BUFX4 BUFX4_29 ( .A(_abc_19873_new_n928_), .Y(_abc_19873_new_n928__bF_buf4));
BUFX4 BUFX4_290 ( .A(core__abc_21302_new_n5104_), .Y(core__abc_21302_new_n5104__bF_buf1));
BUFX4 BUFX4_291 ( .A(core__abc_21302_new_n5104_), .Y(core__abc_21302_new_n5104__bF_buf0));
BUFX4 BUFX4_292 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf10));
BUFX4 BUFX4_293 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf9));
BUFX4 BUFX4_294 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf8));
BUFX4 BUFX4_295 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf7));
BUFX4 BUFX4_296 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf6));
BUFX4 BUFX4_297 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf5));
BUFX4 BUFX4_298 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf4));
BUFX4 BUFX4_299 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf3));
BUFX4 BUFX4_3 ( .A(clk), .Y(clk_hier0_bF_buf6));
BUFX4 BUFX4_30 ( .A(_abc_19873_new_n928_), .Y(_abc_19873_new_n928__bF_buf3));
BUFX4 BUFX4_300 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf2));
BUFX4 BUFX4_301 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf1));
BUFX4 BUFX4_302 ( .A(core_siphash_word1_we), .Y(core_siphash_word1_we_bF_buf0));
BUFX4 BUFX4_303 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf69));
BUFX4 BUFX4_304 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf68));
BUFX4 BUFX4_305 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf67));
BUFX4 BUFX4_306 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf66));
BUFX4 BUFX4_307 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf65));
BUFX4 BUFX4_308 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf64));
BUFX4 BUFX4_309 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf63));
BUFX4 BUFX4_31 ( .A(_abc_19873_new_n928_), .Y(_abc_19873_new_n928__bF_buf2));
BUFX4 BUFX4_310 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf62));
BUFX4 BUFX4_311 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf61));
BUFX4 BUFX4_312 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf60));
BUFX4 BUFX4_313 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf59));
BUFX4 BUFX4_314 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf58));
BUFX4 BUFX4_315 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf57));
BUFX4 BUFX4_316 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf56));
BUFX4 BUFX4_317 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf55));
BUFX4 BUFX4_318 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf54));
BUFX4 BUFX4_319 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf53));
BUFX4 BUFX4_32 ( .A(_abc_19873_new_n928_), .Y(_abc_19873_new_n928__bF_buf1));
BUFX4 BUFX4_320 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf52));
BUFX4 BUFX4_321 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf51));
BUFX4 BUFX4_322 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf50));
BUFX4 BUFX4_323 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf49));
BUFX4 BUFX4_324 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf48));
BUFX4 BUFX4_325 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf47));
BUFX4 BUFX4_326 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf46));
BUFX4 BUFX4_327 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf45));
BUFX4 BUFX4_328 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf44));
BUFX4 BUFX4_329 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf43));
BUFX4 BUFX4_33 ( .A(_abc_19873_new_n928_), .Y(_abc_19873_new_n928__bF_buf0));
BUFX4 BUFX4_330 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf42));
BUFX4 BUFX4_331 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf41));
BUFX4 BUFX4_332 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf40));
BUFX4 BUFX4_333 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf39));
BUFX4 BUFX4_334 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf38));
BUFX4 BUFX4_335 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf37));
BUFX4 BUFX4_336 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf36));
BUFX4 BUFX4_337 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf35));
BUFX4 BUFX4_338 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf34));
BUFX4 BUFX4_339 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf33));
BUFX4 BUFX4_34 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf10));
BUFX4 BUFX4_340 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf32));
BUFX4 BUFX4_341 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf31));
BUFX4 BUFX4_342 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf30));
BUFX4 BUFX4_343 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf29));
BUFX4 BUFX4_344 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf28));
BUFX4 BUFX4_345 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf27));
BUFX4 BUFX4_346 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf26));
BUFX4 BUFX4_347 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf25));
BUFX4 BUFX4_348 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf24));
BUFX4 BUFX4_349 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf23));
BUFX4 BUFX4_35 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf9));
BUFX4 BUFX4_350 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf22));
BUFX4 BUFX4_351 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf21));
BUFX4 BUFX4_352 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf20));
BUFX4 BUFX4_353 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf19));
BUFX4 BUFX4_354 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf18));
BUFX4 BUFX4_355 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf17));
BUFX4 BUFX4_356 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf16));
BUFX4 BUFX4_357 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf15));
BUFX4 BUFX4_358 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf14));
BUFX4 BUFX4_359 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf13));
BUFX4 BUFX4_36 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf8));
BUFX4 BUFX4_360 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf12));
BUFX4 BUFX4_361 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf11));
BUFX4 BUFX4_362 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf10));
BUFX4 BUFX4_363 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf9));
BUFX4 BUFX4_364 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf8));
BUFX4 BUFX4_365 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf7));
BUFX4 BUFX4_366 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf6));
BUFX4 BUFX4_367 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf5));
BUFX4 BUFX4_368 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf4));
BUFX4 BUFX4_369 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf3));
BUFX4 BUFX4_37 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf7));
BUFX4 BUFX4_370 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf2));
BUFX4 BUFX4_371 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf1));
BUFX4 BUFX4_372 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf0));
BUFX4 BUFX4_373 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf13));
BUFX4 BUFX4_374 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf12));
BUFX4 BUFX4_375 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf11));
BUFX4 BUFX4_376 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf10));
BUFX4 BUFX4_377 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf9));
BUFX4 BUFX4_378 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf8));
BUFX4 BUFX4_379 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf7));
BUFX4 BUFX4_38 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf6));
BUFX4 BUFX4_380 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf6));
BUFX4 BUFX4_381 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf5));
BUFX4 BUFX4_382 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf4));
BUFX4 BUFX4_383 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf3));
BUFX4 BUFX4_384 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf2));
BUFX4 BUFX4_385 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf1));
BUFX4 BUFX4_386 ( .A(core__abc_21302_new_n1185_), .Y(core__abc_21302_new_n1185__bF_buf0));
BUFX4 BUFX4_387 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf11));
BUFX4 BUFX4_388 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf10));
BUFX4 BUFX4_389 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf9));
BUFX4 BUFX4_39 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf5));
BUFX4 BUFX4_390 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf8));
BUFX4 BUFX4_391 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf7));
BUFX4 BUFX4_392 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf6));
BUFX4 BUFX4_393 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf5));
BUFX4 BUFX4_394 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf4));
BUFX4 BUFX4_395 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf3));
BUFX4 BUFX4_396 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf2));
BUFX4 BUFX4_397 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf1));
BUFX4 BUFX4_398 ( .A(core__abc_21302_new_n2640_), .Y(core__abc_21302_new_n2640__bF_buf0));
BUFX4 BUFX4_399 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf9));
BUFX4 BUFX4_4 ( .A(clk), .Y(clk_hier0_bF_buf5));
BUFX4 BUFX4_40 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf4));
BUFX4 BUFX4_400 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf8));
BUFX4 BUFX4_401 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf7));
BUFX4 BUFX4_402 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf6));
BUFX4 BUFX4_403 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf5));
BUFX4 BUFX4_404 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf4));
BUFX4 BUFX4_405 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf3));
BUFX4 BUFX4_406 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf2));
BUFX4 BUFX4_407 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf1));
BUFX4 BUFX4_408 ( .A(core__abc_21302_new_n6009_), .Y(core__abc_21302_new_n6009__bF_buf0));
BUFX4 BUFX4_409 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf8));
BUFX4 BUFX4_41 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf3));
BUFX4 BUFX4_410 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf7));
BUFX4 BUFX4_411 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf6));
BUFX4 BUFX4_412 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf5));
BUFX4 BUFX4_413 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf4));
BUFX4 BUFX4_414 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf3));
BUFX4 BUFX4_415 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf2));
BUFX4 BUFX4_416 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf1));
BUFX4 BUFX4_417 ( .A(core__abc_21302_new_n2634_), .Y(core__abc_21302_new_n2634__bF_buf0));
BUFX4 BUFX4_418 ( .A(core__abc_21302_new_n5999_), .Y(core__abc_21302_new_n5999__bF_buf5));
BUFX4 BUFX4_419 ( .A(core__abc_21302_new_n5999_), .Y(core__abc_21302_new_n5999__bF_buf4));
BUFX4 BUFX4_42 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf2));
BUFX4 BUFX4_420 ( .A(core__abc_21302_new_n5999_), .Y(core__abc_21302_new_n5999__bF_buf3));
BUFX4 BUFX4_421 ( .A(core__abc_21302_new_n5999_), .Y(core__abc_21302_new_n5999__bF_buf2));
BUFX4 BUFX4_422 ( .A(core__abc_21302_new_n5999_), .Y(core__abc_21302_new_n5999__bF_buf1));
BUFX4 BUFX4_423 ( .A(core__abc_21302_new_n5999_), .Y(core__abc_21302_new_n5999__bF_buf0));
BUFX4 BUFX4_424 ( .A(_abc_19873_new_n896_), .Y(_abc_19873_new_n896__bF_buf4));
BUFX4 BUFX4_425 ( .A(_abc_19873_new_n896_), .Y(_abc_19873_new_n896__bF_buf3));
BUFX4 BUFX4_426 ( .A(_abc_19873_new_n896_), .Y(_abc_19873_new_n896__bF_buf2));
BUFX4 BUFX4_427 ( .A(_abc_19873_new_n896_), .Y(_abc_19873_new_n896__bF_buf1));
BUFX4 BUFX4_428 ( .A(_abc_19873_new_n896_), .Y(_abc_19873_new_n896__bF_buf0));
BUFX4 BUFX4_429 ( .A(_abc_19873_new_n914_), .Y(_abc_19873_new_n914__bF_buf4));
BUFX4 BUFX4_43 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf1));
BUFX4 BUFX4_430 ( .A(_abc_19873_new_n914_), .Y(_abc_19873_new_n914__bF_buf3));
BUFX4 BUFX4_431 ( .A(_abc_19873_new_n914_), .Y(_abc_19873_new_n914__bF_buf2));
BUFX4 BUFX4_432 ( .A(_abc_19873_new_n914_), .Y(_abc_19873_new_n914__bF_buf1));
BUFX4 BUFX4_433 ( .A(_abc_19873_new_n914_), .Y(_abc_19873_new_n914__bF_buf0));
BUFX4 BUFX4_434 ( .A(_abc_19873_new_n893_), .Y(_abc_19873_new_n893__bF_buf4));
BUFX4 BUFX4_435 ( .A(_abc_19873_new_n893_), .Y(_abc_19873_new_n893__bF_buf3));
BUFX4 BUFX4_436 ( .A(_abc_19873_new_n893_), .Y(_abc_19873_new_n893__bF_buf2));
BUFX4 BUFX4_437 ( .A(_abc_19873_new_n893_), .Y(_abc_19873_new_n893__bF_buf1));
BUFX4 BUFX4_438 ( .A(_abc_19873_new_n893_), .Y(_abc_19873_new_n893__bF_buf0));
BUFX4 BUFX4_439 ( .A(core__abc_21302_new_n6449_), .Y(core__abc_21302_new_n6449__bF_buf7));
BUFX4 BUFX4_44 ( .A(core__abc_21302_new_n1945_), .Y(core__abc_21302_new_n1945__bF_buf0));
BUFX4 BUFX4_440 ( .A(core__abc_21302_new_n6449_), .Y(core__abc_21302_new_n6449__bF_buf6));
BUFX4 BUFX4_441 ( .A(core__abc_21302_new_n6449_), .Y(core__abc_21302_new_n6449__bF_buf5));
BUFX4 BUFX4_442 ( .A(core__abc_21302_new_n6449_), .Y(core__abc_21302_new_n6449__bF_buf4));
BUFX4 BUFX4_443 ( .A(core__abc_21302_new_n6449_), .Y(core__abc_21302_new_n6449__bF_buf3));
BUFX4 BUFX4_444 ( .A(core__abc_21302_new_n6449_), .Y(core__abc_21302_new_n6449__bF_buf2));
BUFX4 BUFX4_445 ( .A(core__abc_21302_new_n6449_), .Y(core__abc_21302_new_n6449__bF_buf1));
BUFX4 BUFX4_446 ( .A(core__abc_21302_new_n6449_), .Y(core__abc_21302_new_n6449__bF_buf0));
BUFX4 BUFX4_447 ( .A(core__abc_21302_new_n2369_), .Y(core__abc_21302_new_n2369__bF_buf7));
BUFX4 BUFX4_448 ( .A(core__abc_21302_new_n2369_), .Y(core__abc_21302_new_n2369__bF_buf6));
BUFX4 BUFX4_449 ( .A(core__abc_21302_new_n2369_), .Y(core__abc_21302_new_n2369__bF_buf5));
BUFX4 BUFX4_45 ( .A(_abc_19873_new_n960_), .Y(_abc_19873_new_n960__bF_buf4));
BUFX4 BUFX4_450 ( .A(core__abc_21302_new_n2369_), .Y(core__abc_21302_new_n2369__bF_buf4));
BUFX4 BUFX4_451 ( .A(core__abc_21302_new_n2369_), .Y(core__abc_21302_new_n2369__bF_buf3));
BUFX4 BUFX4_452 ( .A(core__abc_21302_new_n2369_), .Y(core__abc_21302_new_n2369__bF_buf2));
BUFX4 BUFX4_453 ( .A(core__abc_21302_new_n2369_), .Y(core__abc_21302_new_n2369__bF_buf1));
BUFX4 BUFX4_454 ( .A(core__abc_21302_new_n2369_), .Y(core__abc_21302_new_n2369__bF_buf0));
BUFX4 BUFX4_455 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf15));
BUFX4 BUFX4_456 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf14));
BUFX4 BUFX4_457 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf13));
BUFX4 BUFX4_458 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf12));
BUFX4 BUFX4_459 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf11));
BUFX4 BUFX4_46 ( .A(_abc_19873_new_n960_), .Y(_abc_19873_new_n960__bF_buf3));
BUFX4 BUFX4_460 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf10));
BUFX4 BUFX4_461 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf9));
BUFX4 BUFX4_462 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf8));
BUFX4 BUFX4_463 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf7));
BUFX4 BUFX4_464 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf6));
BUFX4 BUFX4_465 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf5));
BUFX4 BUFX4_466 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf4));
BUFX4 BUFX4_467 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf3));
BUFX4 BUFX4_468 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf2));
BUFX4 BUFX4_469 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf1));
BUFX4 BUFX4_47 ( .A(_abc_19873_new_n960_), .Y(_abc_19873_new_n960__bF_buf2));
BUFX4 BUFX4_470 ( .A(_abc_19873_new_n1524_), .Y(_abc_19873_new_n1524__bF_buf0));
BUFX4 BUFX4_471 ( .A(_abc_19873_new_n905_), .Y(_abc_19873_new_n905__bF_buf3));
BUFX4 BUFX4_472 ( .A(core__abc_21302_new_n5085_), .Y(core__abc_21302_new_n5085__bF_buf5));
BUFX4 BUFX4_473 ( .A(core__abc_21302_new_n5085_), .Y(core__abc_21302_new_n5085__bF_buf4));
BUFX4 BUFX4_474 ( .A(core__abc_21302_new_n5085_), .Y(core__abc_21302_new_n5085__bF_buf3));
BUFX4 BUFX4_475 ( .A(core__abc_21302_new_n5085_), .Y(core__abc_21302_new_n5085__bF_buf2));
BUFX4 BUFX4_476 ( .A(core__abc_21302_new_n5085_), .Y(core__abc_21302_new_n5085__bF_buf1));
BUFX4 BUFX4_477 ( .A(core__abc_21302_new_n5085_), .Y(core__abc_21302_new_n5085__bF_buf0));
BUFX4 BUFX4_478 ( .A(core__abc_21302_new_n2363_), .Y(core__abc_21302_new_n2363__bF_buf5));
BUFX4 BUFX4_479 ( .A(core__abc_21302_new_n2363_), .Y(core__abc_21302_new_n2363__bF_buf4));
BUFX4 BUFX4_48 ( .A(_abc_19873_new_n960_), .Y(_abc_19873_new_n960__bF_buf1));
BUFX4 BUFX4_480 ( .A(core__abc_21302_new_n2363_), .Y(core__abc_21302_new_n2363__bF_buf3));
BUFX4 BUFX4_481 ( .A(core__abc_21302_new_n2363_), .Y(core__abc_21302_new_n2363__bF_buf2));
BUFX4 BUFX4_482 ( .A(core__abc_21302_new_n2363_), .Y(core__abc_21302_new_n2363__bF_buf1));
BUFX4 BUFX4_483 ( .A(core__abc_21302_new_n2363_), .Y(core__abc_21302_new_n2363__bF_buf0));
BUFX4 BUFX4_49 ( .A(_abc_19873_new_n960_), .Y(_abc_19873_new_n960__bF_buf0));
BUFX4 BUFX4_5 ( .A(clk), .Y(clk_hier0_bF_buf4));
BUFX4 BUFX4_50 ( .A(core__abc_21302_new_n5998_), .Y(core__abc_21302_new_n5998__bF_buf3));
BUFX4 BUFX4_51 ( .A(core__abc_21302_new_n5998_), .Y(core__abc_21302_new_n5998__bF_buf2));
BUFX4 BUFX4_52 ( .A(core__abc_21302_new_n5998_), .Y(core__abc_21302_new_n5998__bF_buf1));
BUFX4 BUFX4_53 ( .A(core__abc_21302_new_n5998_), .Y(core__abc_21302_new_n5998__bF_buf0));
BUFX4 BUFX4_54 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf84));
BUFX4 BUFX4_55 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf83));
BUFX4 BUFX4_56 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf82));
BUFX4 BUFX4_57 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf81));
BUFX4 BUFX4_58 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf80));
BUFX4 BUFX4_59 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf79));
BUFX4 BUFX4_6 ( .A(clk), .Y(clk_hier0_bF_buf3));
BUFX4 BUFX4_60 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf78));
BUFX4 BUFX4_61 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf77));
BUFX4 BUFX4_62 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf76));
BUFX4 BUFX4_63 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf75));
BUFX4 BUFX4_64 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf74));
BUFX4 BUFX4_65 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf73));
BUFX4 BUFX4_66 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf72));
BUFX4 BUFX4_67 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf71));
BUFX4 BUFX4_68 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf70));
BUFX4 BUFX4_69 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf69));
BUFX4 BUFX4_7 ( .A(clk), .Y(clk_hier0_bF_buf2));
BUFX4 BUFX4_70 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf68));
BUFX4 BUFX4_71 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf67));
BUFX4 BUFX4_72 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf66));
BUFX4 BUFX4_73 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf65));
BUFX4 BUFX4_74 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf64));
BUFX4 BUFX4_75 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf63));
BUFX4 BUFX4_76 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf62));
BUFX4 BUFX4_77 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf61));
BUFX4 BUFX4_78 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf60));
BUFX4 BUFX4_79 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf59));
BUFX4 BUFX4_8 ( .A(clk), .Y(clk_hier0_bF_buf1));
BUFX4 BUFX4_80 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf58));
BUFX4 BUFX4_81 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf57));
BUFX4 BUFX4_82 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf56));
BUFX4 BUFX4_83 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf55));
BUFX4 BUFX4_84 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf54));
BUFX4 BUFX4_85 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf53));
BUFX4 BUFX4_86 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf52));
BUFX4 BUFX4_87 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf51));
BUFX4 BUFX4_88 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf50));
BUFX4 BUFX4_89 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf49));
BUFX4 BUFX4_9 ( .A(clk), .Y(clk_hier0_bF_buf0));
BUFX4 BUFX4_90 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf48));
BUFX4 BUFX4_91 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf47));
BUFX4 BUFX4_92 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf46));
BUFX4 BUFX4_93 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf45));
BUFX4 BUFX4_94 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf44));
BUFX4 BUFX4_95 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf43));
BUFX4 BUFX4_96 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf42));
BUFX4 BUFX4_97 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf41));
BUFX4 BUFX4_98 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf40));
BUFX4 BUFX4_99 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf39));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf84), .D(_0ctrl_reg_2_0__0_), .Q(core_initalize));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf75), .D(_0param_reg_7_0__5_), .Q(core_final_rounds_1_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf70), .D(_0key2_reg_31_0__23_), .Q(core_key_87_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf69), .D(_0key2_reg_31_0__24_), .Q(core_key_88_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf68), .D(_0key2_reg_31_0__25_), .Q(core_key_89_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf67), .D(_0key2_reg_31_0__26_), .Q(core_key_90_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf66), .D(_0key2_reg_31_0__27_), .Q(core_key_91_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf65), .D(_0key2_reg_31_0__28_), .Q(core_key_92_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf64), .D(_0key2_reg_31_0__29_), .Q(core_key_93_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf63), .D(_0key2_reg_31_0__30_), .Q(core_key_94_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf62), .D(_0key2_reg_31_0__31_), .Q(core_key_95_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf61), .D(_0key3_reg_31_0__0_), .Q(core_key_96_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf74), .D(_0param_reg_7_0__6_), .Q(core_final_rounds_2_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf60), .D(_0key3_reg_31_0__1_), .Q(core_key_97_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf59), .D(_0key3_reg_31_0__2_), .Q(core_key_98_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf58), .D(_0key3_reg_31_0__3_), .Q(core_key_99_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf57), .D(_0key3_reg_31_0__4_), .Q(core_key_100_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf56), .D(_0key3_reg_31_0__5_), .Q(core_key_101_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf55), .D(_0key3_reg_31_0__6_), .Q(core_key_102_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf54), .D(_0key3_reg_31_0__7_), .Q(core_key_103_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf53), .D(_0key3_reg_31_0__8_), .Q(core_key_104_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf52), .D(_0key3_reg_31_0__9_), .Q(core_key_105_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf51), .D(_0key3_reg_31_0__10_), .Q(core_key_106_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf73), .D(_0param_reg_7_0__7_), .Q(core_final_rounds_3_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf50), .D(_0key3_reg_31_0__11_), .Q(core_key_107_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf49), .D(_0key3_reg_31_0__12_), .Q(core_key_108_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf48), .D(_0key3_reg_31_0__13_), .Q(core_key_109_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf47), .D(_0key3_reg_31_0__14_), .Q(core_key_110_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf46), .D(_0key3_reg_31_0__15_), .Q(core_key_111_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf45), .D(_0key3_reg_31_0__16_), .Q(core_key_112_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf44), .D(_0key3_reg_31_0__17_), .Q(core_key_113_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf43), .D(_0key3_reg_31_0__18_), .Q(core_key_114_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf42), .D(_0key3_reg_31_0__19_), .Q(core_key_115_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf41), .D(_0key3_reg_31_0__20_), .Q(core_key_116_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf72), .D(_0key0_reg_31_0__0_), .Q(core_key_0_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf40), .D(_0key3_reg_31_0__21_), .Q(core_key_117_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf39), .D(_0key3_reg_31_0__22_), .Q(core_key_118_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf38), .D(_0key3_reg_31_0__23_), .Q(core_key_119_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf37), .D(_0key3_reg_31_0__24_), .Q(core_key_120_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf36), .D(_0key3_reg_31_0__25_), .Q(core_key_121_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf35), .D(_0key3_reg_31_0__26_), .Q(core_key_122_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf34), .D(_0key3_reg_31_0__27_), .Q(core_key_123_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf33), .D(_0key3_reg_31_0__28_), .Q(core_key_124_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf32), .D(_0key3_reg_31_0__29_), .Q(core_key_125_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf31), .D(_0key3_reg_31_0__30_), .Q(core_key_126_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf71), .D(_0key0_reg_31_0__1_), .Q(core_key_1_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf30), .D(_0key3_reg_31_0__31_), .Q(core_key_127_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf29), .D(_0mi0_reg_31_0__0_), .Q(core_mi_0_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf28), .D(_0mi0_reg_31_0__1_), .Q(core_mi_1_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf27), .D(_0mi0_reg_31_0__2_), .Q(core_mi_2_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf26), .D(_0mi0_reg_31_0__3_), .Q(core_mi_3_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf25), .D(_0mi0_reg_31_0__4_), .Q(core_mi_4_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf24), .D(_0mi0_reg_31_0__5_), .Q(core_mi_5_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf23), .D(_0mi0_reg_31_0__6_), .Q(core_mi_6_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf22), .D(_0mi0_reg_31_0__7_), .Q(core_mi_7_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf21), .D(_0mi0_reg_31_0__8_), .Q(core_mi_8_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf70), .D(_0key0_reg_31_0__2_), .Q(core_key_2_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf20), .D(_0mi0_reg_31_0__9_), .Q(core_mi_9_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf19), .D(_0mi0_reg_31_0__10_), .Q(core_mi_10_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf18), .D(_0mi0_reg_31_0__11_), .Q(core_mi_11_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf17), .D(_0mi0_reg_31_0__12_), .Q(core_mi_12_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf16), .D(_0mi0_reg_31_0__13_), .Q(core_mi_13_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf15), .D(_0mi0_reg_31_0__14_), .Q(core_mi_14_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf14), .D(_0mi0_reg_31_0__15_), .Q(core_mi_15_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf13), .D(_0mi0_reg_31_0__16_), .Q(core_mi_16_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf12), .D(_0mi0_reg_31_0__17_), .Q(core_mi_17_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf11), .D(_0mi0_reg_31_0__18_), .Q(core_mi_18_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf69), .D(_0key0_reg_31_0__3_), .Q(core_key_3_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf10), .D(_0mi0_reg_31_0__19_), .Q(core_mi_19_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf9), .D(_0mi0_reg_31_0__20_), .Q(core_mi_20_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf8), .D(_0mi0_reg_31_0__21_), .Q(core_mi_21_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf7), .D(_0mi0_reg_31_0__22_), .Q(core_mi_22_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf6), .D(_0mi0_reg_31_0__23_), .Q(core_mi_23_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf5), .D(_0mi0_reg_31_0__24_), .Q(core_mi_24_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf4), .D(_0mi0_reg_31_0__25_), .Q(core_mi_25_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf3), .D(_0mi0_reg_31_0__26_), .Q(core_mi_26_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf2), .D(_0mi0_reg_31_0__27_), .Q(core_mi_27_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf1), .D(_0mi0_reg_31_0__28_), .Q(core_mi_28_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf68), .D(_0key0_reg_31_0__4_), .Q(core_key_4_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf0), .D(_0mi0_reg_31_0__29_), .Q(core_mi_29_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf84), .D(_0mi0_reg_31_0__30_), .Q(core_mi_30_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf83), .D(_0mi0_reg_31_0__31_), .Q(core_mi_31_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf82), .D(_0mi1_reg_31_0__0_), .Q(core_mi_32_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf81), .D(_0mi1_reg_31_0__1_), .Q(core_mi_33_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf80), .D(_0mi1_reg_31_0__2_), .Q(core_mi_34_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf79), .D(_0mi1_reg_31_0__3_), .Q(core_mi_35_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf78), .D(_0mi1_reg_31_0__4_), .Q(core_mi_36_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf77), .D(_0mi1_reg_31_0__5_), .Q(core_mi_37_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf76), .D(_0mi1_reg_31_0__6_), .Q(core_mi_38_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf67), .D(_0key0_reg_31_0__5_), .Q(core_key_5_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf75), .D(_0mi1_reg_31_0__7_), .Q(core_mi_39_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf74), .D(_0mi1_reg_31_0__8_), .Q(core_mi_40_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf73), .D(_0mi1_reg_31_0__9_), .Q(core_mi_41_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf72), .D(_0mi1_reg_31_0__10_), .Q(core_mi_42_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf71), .D(_0mi1_reg_31_0__11_), .Q(core_mi_43_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf70), .D(_0mi1_reg_31_0__12_), .Q(core_mi_44_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf69), .D(_0mi1_reg_31_0__13_), .Q(core_mi_45_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf68), .D(_0mi1_reg_31_0__14_), .Q(core_mi_46_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf67), .D(_0mi1_reg_31_0__15_), .Q(core_mi_47_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf66), .D(_0mi1_reg_31_0__16_), .Q(core_mi_48_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf66), .D(_0key0_reg_31_0__6_), .Q(core_key_6_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf65), .D(_0mi1_reg_31_0__17_), .Q(core_mi_49_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf64), .D(_0mi1_reg_31_0__18_), .Q(core_mi_50_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf63), .D(_0mi1_reg_31_0__19_), .Q(core_mi_51_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf62), .D(_0mi1_reg_31_0__20_), .Q(core_mi_52_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf61), .D(_0mi1_reg_31_0__21_), .Q(core_mi_53_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf60), .D(_0mi1_reg_31_0__22_), .Q(core_mi_54_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf59), .D(_0mi1_reg_31_0__23_), .Q(core_mi_55_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf58), .D(_0mi1_reg_31_0__24_), .Q(core_mi_56_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf57), .D(_0mi1_reg_31_0__25_), .Q(core_mi_57_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf56), .D(_0mi1_reg_31_0__26_), .Q(core_mi_58_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf83), .D(_0ctrl_reg_2_0__1_), .Q(core_compress));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf65), .D(_0key0_reg_31_0__7_), .Q(core_key_7_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf55), .D(_0mi1_reg_31_0__27_), .Q(core_mi_59_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf54), .D(_0mi1_reg_31_0__28_), .Q(core_mi_60_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf53), .D(_0mi1_reg_31_0__29_), .Q(core_mi_61_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf52), .D(_0mi1_reg_31_0__30_), .Q(core_mi_62_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf51), .D(_0mi1_reg_31_0__31_), .Q(core_mi_63_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf50), .D(_0word0_reg_31_0__0_), .Q(word0_reg_0_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf49), .D(_0word0_reg_31_0__1_), .Q(word0_reg_1_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf48), .D(_0word0_reg_31_0__2_), .Q(word0_reg_2_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf47), .D(_0word0_reg_31_0__3_), .Q(word0_reg_3_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf46), .D(_0word0_reg_31_0__4_), .Q(word0_reg_4_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf64), .D(_0key0_reg_31_0__8_), .Q(core_key_8_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf45), .D(_0word0_reg_31_0__5_), .Q(word0_reg_5_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf44), .D(_0word0_reg_31_0__6_), .Q(word0_reg_6_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf43), .D(_0word0_reg_31_0__7_), .Q(word0_reg_7_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf42), .D(_0word0_reg_31_0__8_), .Q(word0_reg_8_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf41), .D(_0word0_reg_31_0__9_), .Q(word0_reg_9_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf40), .D(_0word0_reg_31_0__10_), .Q(word0_reg_10_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf39), .D(_0word0_reg_31_0__11_), .Q(word0_reg_11_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf38), .D(_0word0_reg_31_0__12_), .Q(word0_reg_12_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf37), .D(_0word0_reg_31_0__13_), .Q(word0_reg_13_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf36), .D(_0word0_reg_31_0__14_), .Q(word0_reg_14_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf63), .D(_0key0_reg_31_0__9_), .Q(core_key_9_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf35), .D(_0word0_reg_31_0__15_), .Q(word0_reg_15_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf34), .D(_0word0_reg_31_0__16_), .Q(word0_reg_16_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf33), .D(_0word0_reg_31_0__17_), .Q(word0_reg_17_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf32), .D(_0word0_reg_31_0__18_), .Q(word0_reg_18_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf31), .D(_0word0_reg_31_0__19_), .Q(word0_reg_19_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf30), .D(_0word0_reg_31_0__20_), .Q(word0_reg_20_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf29), .D(_0word0_reg_31_0__21_), .Q(word0_reg_21_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf28), .D(_0word0_reg_31_0__22_), .Q(word0_reg_22_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf27), .D(_0word0_reg_31_0__23_), .Q(word0_reg_23_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf26), .D(_0word0_reg_31_0__24_), .Q(word0_reg_24_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf62), .D(_0key0_reg_31_0__10_), .Q(core_key_10_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf25), .D(_0word0_reg_31_0__25_), .Q(word0_reg_25_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf24), .D(_0word0_reg_31_0__26_), .Q(word0_reg_26_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf23), .D(_0word0_reg_31_0__27_), .Q(word0_reg_27_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf22), .D(_0word0_reg_31_0__28_), .Q(word0_reg_28_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf21), .D(_0word0_reg_31_0__29_), .Q(word0_reg_29_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf20), .D(_0word0_reg_31_0__30_), .Q(word0_reg_30_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf19), .D(_0word0_reg_31_0__31_), .Q(word0_reg_31_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf18), .D(_0word1_reg_31_0__0_), .Q(word1_reg_0_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf17), .D(_0word1_reg_31_0__1_), .Q(word1_reg_1_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf16), .D(_0word1_reg_31_0__2_), .Q(word1_reg_2_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf61), .D(_0key0_reg_31_0__11_), .Q(core_key_11_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf15), .D(_0word1_reg_31_0__3_), .Q(word1_reg_3_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf14), .D(_0word1_reg_31_0__4_), .Q(word1_reg_4_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf13), .D(_0word1_reg_31_0__5_), .Q(word1_reg_5_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf12), .D(_0word1_reg_31_0__6_), .Q(word1_reg_6_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf11), .D(_0word1_reg_31_0__7_), .Q(word1_reg_7_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf10), .D(_0word1_reg_31_0__8_), .Q(word1_reg_8_));
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf9), .D(_0word1_reg_31_0__9_), .Q(word1_reg_9_));
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf8), .D(_0word1_reg_31_0__10_), .Q(word1_reg_10_));
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf7), .D(_0word1_reg_31_0__11_), .Q(word1_reg_11_));
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf6), .D(_0word1_reg_31_0__12_), .Q(word1_reg_12_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf60), .D(_0key0_reg_31_0__12_), .Q(core_key_12_));
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf5), .D(_0word1_reg_31_0__13_), .Q(word1_reg_13_));
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf4), .D(_0word1_reg_31_0__14_), .Q(word1_reg_14_));
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf3), .D(_0word1_reg_31_0__15_), .Q(word1_reg_15_));
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf2), .D(_0word1_reg_31_0__16_), .Q(word1_reg_16_));
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf1), .D(_0word1_reg_31_0__17_), .Q(word1_reg_17_));
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf0), .D(_0word1_reg_31_0__18_), .Q(word1_reg_18_));
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf84), .D(_0word1_reg_31_0__19_), .Q(word1_reg_19_));
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf83), .D(_0word1_reg_31_0__20_), .Q(word1_reg_20_));
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf82), .D(_0word1_reg_31_0__21_), .Q(word1_reg_21_));
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf81), .D(_0word1_reg_31_0__22_), .Q(word1_reg_22_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf59), .D(_0key0_reg_31_0__13_), .Q(core_key_13_));
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf80), .D(_0word1_reg_31_0__23_), .Q(word1_reg_23_));
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf79), .D(_0word1_reg_31_0__24_), .Q(word1_reg_24_));
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf78), .D(_0word1_reg_31_0__25_), .Q(word1_reg_25_));
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf77), .D(_0word1_reg_31_0__26_), .Q(word1_reg_26_));
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf76), .D(_0word1_reg_31_0__27_), .Q(word1_reg_27_));
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf75), .D(_0word1_reg_31_0__28_), .Q(word1_reg_28_));
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf74), .D(_0word1_reg_31_0__29_), .Q(word1_reg_29_));
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf73), .D(_0word1_reg_31_0__30_), .Q(word1_reg_30_));
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf72), .D(_0word1_reg_31_0__31_), .Q(word1_reg_31_));
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf71), .D(_0word2_reg_31_0__0_), .Q(word2_reg_0_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf58), .D(_0key0_reg_31_0__14_), .Q(core_key_14_));
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf70), .D(_0word2_reg_31_0__1_), .Q(word2_reg_1_));
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf69), .D(_0word2_reg_31_0__2_), .Q(word2_reg_2_));
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf68), .D(_0word2_reg_31_0__3_), .Q(word2_reg_3_));
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf67), .D(_0word2_reg_31_0__4_), .Q(word2_reg_4_));
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf66), .D(_0word2_reg_31_0__5_), .Q(word2_reg_5_));
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf65), .D(_0word2_reg_31_0__6_), .Q(word2_reg_6_));
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf64), .D(_0word2_reg_31_0__7_), .Q(word2_reg_7_));
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf63), .D(_0word2_reg_31_0__8_), .Q(word2_reg_8_));
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf62), .D(_0word2_reg_31_0__9_), .Q(word2_reg_9_));
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf61), .D(_0word2_reg_31_0__10_), .Q(word2_reg_10_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf57), .D(_0key0_reg_31_0__15_), .Q(core_key_15_));
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf60), .D(_0word2_reg_31_0__11_), .Q(word2_reg_11_));
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf59), .D(_0word2_reg_31_0__12_), .Q(word2_reg_12_));
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf58), .D(_0word2_reg_31_0__13_), .Q(word2_reg_13_));
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf57), .D(_0word2_reg_31_0__14_), .Q(word2_reg_14_));
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf56), .D(_0word2_reg_31_0__15_), .Q(word2_reg_15_));
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf55), .D(_0word2_reg_31_0__16_), .Q(word2_reg_16_));
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf54), .D(_0word2_reg_31_0__17_), .Q(word2_reg_17_));
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf53), .D(_0word2_reg_31_0__18_), .Q(word2_reg_18_));
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf52), .D(_0word2_reg_31_0__19_), .Q(word2_reg_19_));
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf51), .D(_0word2_reg_31_0__20_), .Q(word2_reg_20_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf56), .D(_0key0_reg_31_0__16_), .Q(core_key_16_));
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf50), .D(_0word2_reg_31_0__21_), .Q(word2_reg_21_));
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf49), .D(_0word2_reg_31_0__22_), .Q(word2_reg_22_));
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf48), .D(_0word2_reg_31_0__23_), .Q(word2_reg_23_));
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf47), .D(_0word2_reg_31_0__24_), .Q(word2_reg_24_));
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf46), .D(_0word2_reg_31_0__25_), .Q(word2_reg_25_));
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf45), .D(_0word2_reg_31_0__26_), .Q(word2_reg_26_));
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf44), .D(_0word2_reg_31_0__27_), .Q(word2_reg_27_));
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf43), .D(_0word2_reg_31_0__28_), .Q(word2_reg_28_));
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf42), .D(_0word2_reg_31_0__29_), .Q(word2_reg_29_));
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf41), .D(_0word2_reg_31_0__30_), .Q(word2_reg_30_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf82), .D(_0ctrl_reg_2_0__2_), .Q(core_finalize));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf55), .D(_0key0_reg_31_0__17_), .Q(core_key_17_));
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf40), .D(_0word2_reg_31_0__31_), .Q(word2_reg_31_));
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf39), .D(_0word3_reg_31_0__0_), .Q(word3_reg_0_));
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf38), .D(_0word3_reg_31_0__1_), .Q(word3_reg_1_));
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf37), .D(_0word3_reg_31_0__2_), .Q(word3_reg_2_));
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf36), .D(_0word3_reg_31_0__3_), .Q(word3_reg_3_));
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf35), .D(_0word3_reg_31_0__4_), .Q(word3_reg_4_));
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf34), .D(_0word3_reg_31_0__5_), .Q(word3_reg_5_));
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf33), .D(_0word3_reg_31_0__6_), .Q(word3_reg_6_));
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf32), .D(_0word3_reg_31_0__7_), .Q(word3_reg_7_));
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf31), .D(_0word3_reg_31_0__8_), .Q(word3_reg_8_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf54), .D(_0key0_reg_31_0__18_), .Q(core_key_18_));
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf30), .D(_0word3_reg_31_0__9_), .Q(word3_reg_9_));
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf29), .D(_0word3_reg_31_0__10_), .Q(word3_reg_10_));
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf28), .D(_0word3_reg_31_0__11_), .Q(word3_reg_11_));
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf27), .D(_0word3_reg_31_0__12_), .Q(word3_reg_12_));
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf26), .D(_0word3_reg_31_0__13_), .Q(word3_reg_13_));
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf25), .D(_0word3_reg_31_0__14_), .Q(word3_reg_14_));
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf24), .D(_0word3_reg_31_0__15_), .Q(word3_reg_15_));
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf23), .D(_0word3_reg_31_0__16_), .Q(word3_reg_16_));
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf22), .D(_0word3_reg_31_0__17_), .Q(word3_reg_17_));
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf21), .D(_0word3_reg_31_0__18_), .Q(word3_reg_18_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf53), .D(_0key0_reg_31_0__19_), .Q(core_key_19_));
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf20), .D(_0word3_reg_31_0__19_), .Q(word3_reg_19_));
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf19), .D(_0word3_reg_31_0__20_), .Q(word3_reg_20_));
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf18), .D(_0word3_reg_31_0__21_), .Q(word3_reg_21_));
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf17), .D(_0word3_reg_31_0__22_), .Q(word3_reg_22_));
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf16), .D(_0word3_reg_31_0__23_), .Q(word3_reg_23_));
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf15), .D(_0word3_reg_31_0__24_), .Q(word3_reg_24_));
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf14), .D(_0word3_reg_31_0__25_), .Q(word3_reg_25_));
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf13), .D(_0word3_reg_31_0__26_), .Q(word3_reg_26_));
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf12), .D(_0word3_reg_31_0__27_), .Q(word3_reg_27_));
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf11), .D(_0word3_reg_31_0__28_), .Q(word3_reg_28_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf52), .D(_0key0_reg_31_0__20_), .Q(core_key_20_));
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf10), .D(_0word3_reg_31_0__29_), .Q(word3_reg_29_));
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf9), .D(_0word3_reg_31_0__30_), .Q(word3_reg_30_));
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf8), .D(_0word3_reg_31_0__31_), .Q(word3_reg_31_));
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf7), .D(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_0_), .Q(core_siphash_ctrl_reg_0_));
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf6), .D(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1470), .Q(core_siphash_ctrl_reg_1_));
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf5), .D(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1474), .Q(core_siphash_ctrl_reg_2_));
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf4), .D(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_3_), .Q(core_siphash_ctrl_reg_3_));
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf3), .D(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_4_), .Q(core_siphash_ctrl_reg_4_));
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf2), .D(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1496), .Q(core_siphash_ctrl_reg_5_));
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf1), .D(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_6_), .Q(core_siphash_ctrl_reg_6_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf51), .D(_0key0_reg_31_0__21_), .Q(core_key_21_));
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf0), .D(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1509), .Q(core_siphash_word1_we));
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf84), .D(core__0v0_reg_63_0__0_), .Q(core_v0_reg_0_));
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf83), .D(core__0v0_reg_63_0__1_), .Q(core_v0_reg_1_));
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf82), .D(core__0v0_reg_63_0__2_), .Q(core_v0_reg_2_));
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf81), .D(core__0v0_reg_63_0__3_), .Q(core_v0_reg_3_));
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf80), .D(core__0v0_reg_63_0__4_), .Q(core_v0_reg_4_));
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf79), .D(core__0v0_reg_63_0__5_), .Q(core_v0_reg_5_));
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf78), .D(core__0v0_reg_63_0__6_), .Q(core_v0_reg_6_));
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf77), .D(core__0v0_reg_63_0__7_), .Q(core_v0_reg_7_));
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf76), .D(core__0v0_reg_63_0__8_), .Q(core_v0_reg_8_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf50), .D(_0key0_reg_31_0__22_), .Q(core_key_22_));
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf75), .D(core__0v0_reg_63_0__9_), .Q(core_v0_reg_9_));
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf74), .D(core__0v0_reg_63_0__10_), .Q(core_v0_reg_10_));
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf73), .D(core__0v0_reg_63_0__11_), .Q(core_v0_reg_11_));
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf72), .D(core__0v0_reg_63_0__12_), .Q(core_v0_reg_12_));
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf71), .D(core__0v0_reg_63_0__13_), .Q(core_v0_reg_13_));
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf70), .D(core__0v0_reg_63_0__14_), .Q(core_v0_reg_14_));
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf69), .D(core__0v0_reg_63_0__15_), .Q(core_v0_reg_15_));
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf68), .D(core__0v0_reg_63_0__16_), .Q(core_v0_reg_16_));
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf67), .D(core__0v0_reg_63_0__17_), .Q(core_v0_reg_17_));
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf66), .D(core__0v0_reg_63_0__18_), .Q(core_v0_reg_18_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf49), .D(_0key0_reg_31_0__23_), .Q(core_key_23_));
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf65), .D(core__0v0_reg_63_0__19_), .Q(core_v0_reg_19_));
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf64), .D(core__0v0_reg_63_0__20_), .Q(core_v0_reg_20_));
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf63), .D(core__0v0_reg_63_0__21_), .Q(core_v0_reg_21_));
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf62), .D(core__0v0_reg_63_0__22_), .Q(core_v0_reg_22_));
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf61), .D(core__0v0_reg_63_0__23_), .Q(core_v0_reg_23_));
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf60), .D(core__0v0_reg_63_0__24_), .Q(core_v0_reg_24_));
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf59), .D(core__0v0_reg_63_0__25_), .Q(core_v0_reg_25_));
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf58), .D(core__0v0_reg_63_0__26_), .Q(core_v0_reg_26_));
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf57), .D(core__0v0_reg_63_0__27_), .Q(core_v0_reg_27_));
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf56), .D(core__0v0_reg_63_0__28_), .Q(core_v0_reg_28_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf48), .D(_0key0_reg_31_0__24_), .Q(core_key_24_));
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf55), .D(core__0v0_reg_63_0__29_), .Q(core_v0_reg_29_));
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf54), .D(core__0v0_reg_63_0__30_), .Q(core_v0_reg_30_));
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf53), .D(core__0v0_reg_63_0__31_), .Q(core_v0_reg_31_));
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf52), .D(core__0v0_reg_63_0__32_), .Q(core_v0_reg_32_));
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf51), .D(core__0v0_reg_63_0__33_), .Q(core_v0_reg_33_));
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf50), .D(core__0v0_reg_63_0__34_), .Q(core_v0_reg_34_));
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf49), .D(core__0v0_reg_63_0__35_), .Q(core_v0_reg_35_));
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf48), .D(core__0v0_reg_63_0__36_), .Q(core_v0_reg_36_));
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf47), .D(core__0v0_reg_63_0__37_), .Q(core_v0_reg_37_));
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf46), .D(core__0v0_reg_63_0__38_), .Q(core_v0_reg_38_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf47), .D(_0key0_reg_31_0__25_), .Q(core_key_25_));
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf45), .D(core__0v0_reg_63_0__39_), .Q(core_v0_reg_39_));
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf44), .D(core__0v0_reg_63_0__40_), .Q(core_v0_reg_40_));
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf43), .D(core__0v0_reg_63_0__41_), .Q(core_v0_reg_41_));
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf42), .D(core__0v0_reg_63_0__42_), .Q(core_v0_reg_42_));
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf41), .D(core__0v0_reg_63_0__43_), .Q(core_v0_reg_43_));
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf40), .D(core__0v0_reg_63_0__44_), .Q(core_v0_reg_44_));
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf39), .D(core__0v0_reg_63_0__45_), .Q(core_v0_reg_45_));
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf38), .D(core__0v0_reg_63_0__46_), .Q(core_v0_reg_46_));
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf37), .D(core__0v0_reg_63_0__47_), .Q(core_v0_reg_47_));
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf36), .D(core__0v0_reg_63_0__48_), .Q(core_v0_reg_48_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf46), .D(_0key0_reg_31_0__26_), .Q(core_key_26_));
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf35), .D(core__0v0_reg_63_0__49_), .Q(core_v0_reg_49_));
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf34), .D(core__0v0_reg_63_0__50_), .Q(core_v0_reg_50_));
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf33), .D(core__0v0_reg_63_0__51_), .Q(core_v0_reg_51_));
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf32), .D(core__0v0_reg_63_0__52_), .Q(core_v0_reg_52_));
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf31), .D(core__0v0_reg_63_0__53_), .Q(core_v0_reg_53_));
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf30), .D(core__0v0_reg_63_0__54_), .Q(core_v0_reg_54_));
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf29), .D(core__0v0_reg_63_0__55_), .Q(core_v0_reg_55_));
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf28), .D(core__0v0_reg_63_0__56_), .Q(core_v0_reg_56_));
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf27), .D(core__0v0_reg_63_0__57_), .Q(core_v0_reg_57_));
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf26), .D(core__0v0_reg_63_0__58_), .Q(core_v0_reg_58_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf81), .D(_0long_reg_0_0_), .Q(core_long));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf45), .D(_0key0_reg_31_0__27_), .Q(core_key_27_));
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf25), .D(core__0v0_reg_63_0__59_), .Q(core_v0_reg_59_));
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf24), .D(core__0v0_reg_63_0__60_), .Q(core_v0_reg_60_));
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf23), .D(core__0v0_reg_63_0__61_), .Q(core_v0_reg_61_));
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf22), .D(core__0v0_reg_63_0__62_), .Q(core_v0_reg_62_));
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf21), .D(core__0v0_reg_63_0__63_), .Q(core_v0_reg_63_));
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf20), .D(core__0v1_reg_63_0__0_), .Q(core_v1_reg_0_));
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf19), .D(core__0v1_reg_63_0__1_), .Q(core_v1_reg_1_));
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf18), .D(core__0v1_reg_63_0__2_), .Q(core_v1_reg_2_));
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf17), .D(core__0v1_reg_63_0__3_), .Q(core_v1_reg_3_));
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf16), .D(core__0v1_reg_63_0__4_), .Q(core_v1_reg_4_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf44), .D(_0key0_reg_31_0__28_), .Q(core_key_28_));
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf15), .D(core__0v1_reg_63_0__5_), .Q(core_v1_reg_5_));
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf14), .D(core__0v1_reg_63_0__6_), .Q(core_v1_reg_6_));
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf13), .D(core__0v1_reg_63_0__7_), .Q(core_v1_reg_7_));
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf12), .D(core__0v1_reg_63_0__8_), .Q(core_v1_reg_8_));
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf11), .D(core__0v1_reg_63_0__9_), .Q(core_v1_reg_9_));
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf10), .D(core__0v1_reg_63_0__10_), .Q(core_v1_reg_10_));
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf9), .D(core__0v1_reg_63_0__11_), .Q(core_v1_reg_11_));
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf8), .D(core__0v1_reg_63_0__12_), .Q(core_v1_reg_12_));
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf7), .D(core__0v1_reg_63_0__13_), .Q(core_v1_reg_13_));
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf6), .D(core__0v1_reg_63_0__14_), .Q(core_v1_reg_14_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf43), .D(_0key0_reg_31_0__29_), .Q(core_key_29_));
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf5), .D(core__0v1_reg_63_0__15_), .Q(core_v1_reg_15_));
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf4), .D(core__0v1_reg_63_0__16_), .Q(core_v1_reg_16_));
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf3), .D(core__0v1_reg_63_0__17_), .Q(core_v1_reg_17_));
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf2), .D(core__0v1_reg_63_0__18_), .Q(core_v1_reg_18_));
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf1), .D(core__0v1_reg_63_0__19_), .Q(core_v1_reg_19_));
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf0), .D(core__0v1_reg_63_0__20_), .Q(core_v1_reg_20_));
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf84), .D(core__0v1_reg_63_0__21_), .Q(core_v1_reg_21_));
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf83), .D(core__0v1_reg_63_0__22_), .Q(core_v1_reg_22_));
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf82), .D(core__0v1_reg_63_0__23_), .Q(core_v1_reg_23_));
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf81), .D(core__0v1_reg_63_0__24_), .Q(core_v1_reg_24_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf42), .D(_0key0_reg_31_0__30_), .Q(core_key_30_));
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf80), .D(core__0v1_reg_63_0__25_), .Q(core_v1_reg_25_));
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf79), .D(core__0v1_reg_63_0__26_), .Q(core_v1_reg_26_));
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf78), .D(core__0v1_reg_63_0__27_), .Q(core_v1_reg_27_));
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf77), .D(core__0v1_reg_63_0__28_), .Q(core_v1_reg_28_));
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf76), .D(core__0v1_reg_63_0__29_), .Q(core_v1_reg_29_));
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf75), .D(core__0v1_reg_63_0__30_), .Q(core_v1_reg_30_));
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf74), .D(core__0v1_reg_63_0__31_), .Q(core_v1_reg_31_));
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf73), .D(core__0v1_reg_63_0__32_), .Q(core_v1_reg_32_));
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf72), .D(core__0v1_reg_63_0__33_), .Q(core_v1_reg_33_));
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf71), .D(core__0v1_reg_63_0__34_), .Q(core_v1_reg_34_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf41), .D(_0key0_reg_31_0__31_), .Q(core_key_31_));
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf70), .D(core__0v1_reg_63_0__35_), .Q(core_v1_reg_35_));
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf69), .D(core__0v1_reg_63_0__36_), .Q(core_v1_reg_36_));
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf68), .D(core__0v1_reg_63_0__37_), .Q(core_v1_reg_37_));
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf67), .D(core__0v1_reg_63_0__38_), .Q(core_v1_reg_38_));
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf66), .D(core__0v1_reg_63_0__39_), .Q(core_v1_reg_39_));
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf65), .D(core__0v1_reg_63_0__40_), .Q(core_v1_reg_40_));
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf64), .D(core__0v1_reg_63_0__41_), .Q(core_v1_reg_41_));
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf63), .D(core__0v1_reg_63_0__42_), .Q(core_v1_reg_42_));
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf62), .D(core__0v1_reg_63_0__43_), .Q(core_v1_reg_43_));
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf61), .D(core__0v1_reg_63_0__44_), .Q(core_v1_reg_44_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf40), .D(_0key1_reg_31_0__0_), .Q(core_key_32_));
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf60), .D(core__0v1_reg_63_0__45_), .Q(core_v1_reg_45_));
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf59), .D(core__0v1_reg_63_0__46_), .Q(core_v1_reg_46_));
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf58), .D(core__0v1_reg_63_0__47_), .Q(core_v1_reg_47_));
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf57), .D(core__0v1_reg_63_0__48_), .Q(core_v1_reg_48_));
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf56), .D(core__0v1_reg_63_0__49_), .Q(core_v1_reg_49_));
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf55), .D(core__0v1_reg_63_0__50_), .Q(core_v1_reg_50_));
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf54), .D(core__0v1_reg_63_0__51_), .Q(core_v1_reg_51_));
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf53), .D(core__0v1_reg_63_0__52_), .Q(core_v1_reg_52_));
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf52), .D(core__0v1_reg_63_0__53_), .Q(core_v1_reg_53_));
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf51), .D(core__0v1_reg_63_0__54_), .Q(core_v1_reg_54_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf39), .D(_0key1_reg_31_0__1_), .Q(core_key_33_));
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf50), .D(core__0v1_reg_63_0__55_), .Q(core_v1_reg_55_));
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf49), .D(core__0v1_reg_63_0__56_), .Q(core_v1_reg_56_));
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf48), .D(core__0v1_reg_63_0__57_), .Q(core_v1_reg_57_));
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf47), .D(core__0v1_reg_63_0__58_), .Q(core_v1_reg_58_));
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf46), .D(core__0v1_reg_63_0__59_), .Q(core_v1_reg_59_));
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf45), .D(core__0v1_reg_63_0__60_), .Q(core_v1_reg_60_));
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf44), .D(core__0v1_reg_63_0__61_), .Q(core_v1_reg_61_));
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf43), .D(core__0v1_reg_63_0__62_), .Q(core_v1_reg_62_));
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf42), .D(core__0v1_reg_63_0__63_), .Q(core_v1_reg_63_));
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf41), .D(core__0v2_reg_63_0__0_), .Q(core_v2_reg_0_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf38), .D(_0key1_reg_31_0__2_), .Q(core_key_34_));
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf40), .D(core__0v2_reg_63_0__1_), .Q(core_v2_reg_1_));
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf39), .D(core__0v2_reg_63_0__2_), .Q(core_v2_reg_2_));
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf38), .D(core__0v2_reg_63_0__3_), .Q(core_v2_reg_3_));
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf37), .D(core__0v2_reg_63_0__4_), .Q(core_v2_reg_4_));
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf36), .D(core__0v2_reg_63_0__5_), .Q(core_v2_reg_5_));
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf35), .D(core__0v2_reg_63_0__6_), .Q(core_v2_reg_6_));
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf34), .D(core__0v2_reg_63_0__7_), .Q(core_v2_reg_7_));
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf33), .D(core__0v2_reg_63_0__8_), .Q(core_v2_reg_8_));
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf32), .D(core__0v2_reg_63_0__9_), .Q(core_v2_reg_9_));
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf31), .D(core__0v2_reg_63_0__10_), .Q(core_v2_reg_10_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf37), .D(_0key1_reg_31_0__3_), .Q(core_key_35_));
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf30), .D(core__0v2_reg_63_0__11_), .Q(core_v2_reg_11_));
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf29), .D(core__0v2_reg_63_0__12_), .Q(core_v2_reg_12_));
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf28), .D(core__0v2_reg_63_0__13_), .Q(core_v2_reg_13_));
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf27), .D(core__0v2_reg_63_0__14_), .Q(core_v2_reg_14_));
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf26), .D(core__0v2_reg_63_0__15_), .Q(core_v2_reg_15_));
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf25), .D(core__0v2_reg_63_0__16_), .Q(core_v2_reg_16_));
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf24), .D(core__0v2_reg_63_0__17_), .Q(core_v2_reg_17_));
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf23), .D(core__0v2_reg_63_0__18_), .Q(core_v2_reg_18_));
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf22), .D(core__0v2_reg_63_0__19_), .Q(core_v2_reg_19_));
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf21), .D(core__0v2_reg_63_0__20_), .Q(core_v2_reg_20_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf36), .D(_0key1_reg_31_0__4_), .Q(core_key_36_));
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf20), .D(core__0v2_reg_63_0__21_), .Q(core_v2_reg_21_));
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf19), .D(core__0v2_reg_63_0__22_), .Q(core_v2_reg_22_));
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf18), .D(core__0v2_reg_63_0__23_), .Q(core_v2_reg_23_));
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf17), .D(core__0v2_reg_63_0__24_), .Q(core_v2_reg_24_));
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf16), .D(core__0v2_reg_63_0__25_), .Q(core_v2_reg_25_));
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf15), .D(core__0v2_reg_63_0__26_), .Q(core_v2_reg_26_));
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf14), .D(core__0v2_reg_63_0__27_), .Q(core_v2_reg_27_));
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf13), .D(core__0v2_reg_63_0__28_), .Q(core_v2_reg_28_));
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf12), .D(core__0v2_reg_63_0__29_), .Q(core_v2_reg_29_));
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf11), .D(core__0v2_reg_63_0__30_), .Q(core_v2_reg_30_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf80), .D(_0param_reg_7_0__0_), .Q(core_compression_rounds_0_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf35), .D(_0key1_reg_31_0__5_), .Q(core_key_37_));
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf10), .D(core__0v2_reg_63_0__31_), .Q(core_v2_reg_31_));
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf9), .D(core__0v2_reg_63_0__32_), .Q(core_v2_reg_32_));
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf8), .D(core__0v2_reg_63_0__33_), .Q(core_v2_reg_33_));
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf7), .D(core__0v2_reg_63_0__34_), .Q(core_v2_reg_34_));
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf6), .D(core__0v2_reg_63_0__35_), .Q(core_v2_reg_35_));
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf5), .D(core__0v2_reg_63_0__36_), .Q(core_v2_reg_36_));
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf4), .D(core__0v2_reg_63_0__37_), .Q(core_v2_reg_37_));
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf3), .D(core__0v2_reg_63_0__38_), .Q(core_v2_reg_38_));
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf2), .D(core__0v2_reg_63_0__39_), .Q(core_v2_reg_39_));
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf1), .D(core__0v2_reg_63_0__40_), .Q(core_v2_reg_40_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf34), .D(_0key1_reg_31_0__6_), .Q(core_key_38_));
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf0), .D(core__0v2_reg_63_0__41_), .Q(core_v2_reg_41_));
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf84), .D(core__0v2_reg_63_0__42_), .Q(core_v2_reg_42_));
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf83), .D(core__0v2_reg_63_0__43_), .Q(core_v2_reg_43_));
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf82), .D(core__0v2_reg_63_0__44_), .Q(core_v2_reg_44_));
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf81), .D(core__0v2_reg_63_0__45_), .Q(core_v2_reg_45_));
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf80), .D(core__0v2_reg_63_0__46_), .Q(core_v2_reg_46_));
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf79), .D(core__0v2_reg_63_0__47_), .Q(core_v2_reg_47_));
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf78), .D(core__0v2_reg_63_0__48_), .Q(core_v2_reg_48_));
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf77), .D(core__0v2_reg_63_0__49_), .Q(core_v2_reg_49_));
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf76), .D(core__0v2_reg_63_0__50_), .Q(core_v2_reg_50_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf33), .D(_0key1_reg_31_0__7_), .Q(core_key_39_));
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf75), .D(core__0v2_reg_63_0__51_), .Q(core_v2_reg_51_));
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf74), .D(core__0v2_reg_63_0__52_), .Q(core_v2_reg_52_));
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf73), .D(core__0v2_reg_63_0__53_), .Q(core_v2_reg_53_));
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf72), .D(core__0v2_reg_63_0__54_), .Q(core_v2_reg_54_));
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf71), .D(core__0v2_reg_63_0__55_), .Q(core_v2_reg_55_));
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf70), .D(core__0v2_reg_63_0__56_), .Q(core_v2_reg_56_));
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf69), .D(core__0v2_reg_63_0__57_), .Q(core_v2_reg_57_));
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf68), .D(core__0v2_reg_63_0__58_), .Q(core_v2_reg_58_));
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf67), .D(core__0v2_reg_63_0__59_), .Q(core_v2_reg_59_));
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf66), .D(core__0v2_reg_63_0__60_), .Q(core_v2_reg_60_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf32), .D(_0key1_reg_31_0__8_), .Q(core_key_40_));
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf65), .D(core__0v2_reg_63_0__61_), .Q(core_v2_reg_61_));
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf64), .D(core__0v2_reg_63_0__62_), .Q(core_v2_reg_62_));
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf63), .D(core__0v2_reg_63_0__63_), .Q(core_v2_reg_63_));
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf62), .D(core__0v3_reg_63_0__0_), .Q(core_v3_reg_0_));
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf61), .D(core__0v3_reg_63_0__1_), .Q(core_v3_reg_1_));
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf60), .D(core__0v3_reg_63_0__2_), .Q(core_v3_reg_2_));
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf59), .D(core__0v3_reg_63_0__3_), .Q(core_v3_reg_3_));
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf58), .D(core__0v3_reg_63_0__4_), .Q(core_v3_reg_4_));
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf57), .D(core__0v3_reg_63_0__5_), .Q(core_v3_reg_5_));
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf56), .D(core__0v3_reg_63_0__6_), .Q(core_v3_reg_6_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf31), .D(_0key1_reg_31_0__9_), .Q(core_key_41_));
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf55), .D(core__0v3_reg_63_0__7_), .Q(core_v3_reg_7_));
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf54), .D(core__0v3_reg_63_0__8_), .Q(core_v3_reg_8_));
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf53), .D(core__0v3_reg_63_0__9_), .Q(core_v3_reg_9_));
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf52), .D(core__0v3_reg_63_0__10_), .Q(core_v3_reg_10_));
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf51), .D(core__0v3_reg_63_0__11_), .Q(core_v3_reg_11_));
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf50), .D(core__0v3_reg_63_0__12_), .Q(core_v3_reg_12_));
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf49), .D(core__0v3_reg_63_0__13_), .Q(core_v3_reg_13_));
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf48), .D(core__0v3_reg_63_0__14_), .Q(core_v3_reg_14_));
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf47), .D(core__0v3_reg_63_0__15_), .Q(core_v3_reg_15_));
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf46), .D(core__0v3_reg_63_0__16_), .Q(core_v3_reg_16_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf30), .D(_0key1_reg_31_0__10_), .Q(core_key_42_));
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf45), .D(core__0v3_reg_63_0__17_), .Q(core_v3_reg_17_));
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf44), .D(core__0v3_reg_63_0__18_), .Q(core_v3_reg_18_));
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf43), .D(core__0v3_reg_63_0__19_), .Q(core_v3_reg_19_));
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf42), .D(core__0v3_reg_63_0__20_), .Q(core_v3_reg_20_));
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf41), .D(core__0v3_reg_63_0__21_), .Q(core_v3_reg_21_));
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf40), .D(core__0v3_reg_63_0__22_), .Q(core_v3_reg_22_));
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf39), .D(core__0v3_reg_63_0__23_), .Q(core_v3_reg_23_));
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf38), .D(core__0v3_reg_63_0__24_), .Q(core_v3_reg_24_));
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf37), .D(core__0v3_reg_63_0__25_), .Q(core_v3_reg_25_));
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf36), .D(core__0v3_reg_63_0__26_), .Q(core_v3_reg_26_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf29), .D(_0key1_reg_31_0__11_), .Q(core_key_43_));
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf35), .D(core__0v3_reg_63_0__27_), .Q(core_v3_reg_27_));
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf34), .D(core__0v3_reg_63_0__28_), .Q(core_v3_reg_28_));
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf33), .D(core__0v3_reg_63_0__29_), .Q(core_v3_reg_29_));
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf32), .D(core__0v3_reg_63_0__30_), .Q(core_v3_reg_30_));
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf31), .D(core__0v3_reg_63_0__31_), .Q(core_v3_reg_31_));
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf30), .D(core__0v3_reg_63_0__32_), .Q(core_v3_reg_32_));
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf29), .D(core__0v3_reg_63_0__33_), .Q(core_v3_reg_33_));
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf28), .D(core__0v3_reg_63_0__34_), .Q(core_v3_reg_34_));
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf27), .D(core__0v3_reg_63_0__35_), .Q(core_v3_reg_35_));
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf26), .D(core__0v3_reg_63_0__36_), .Q(core_v3_reg_36_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf28), .D(_0key1_reg_31_0__12_), .Q(core_key_44_));
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf25), .D(core__0v3_reg_63_0__37_), .Q(core_v3_reg_37_));
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf24), .D(core__0v3_reg_63_0__38_), .Q(core_v3_reg_38_));
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf23), .D(core__0v3_reg_63_0__39_), .Q(core_v3_reg_39_));
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf22), .D(core__0v3_reg_63_0__40_), .Q(core_v3_reg_40_));
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf21), .D(core__0v3_reg_63_0__41_), .Q(core_v3_reg_41_));
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf20), .D(core__0v3_reg_63_0__42_), .Q(core_v3_reg_42_));
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf19), .D(core__0v3_reg_63_0__43_), .Q(core_v3_reg_43_));
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf18), .D(core__0v3_reg_63_0__44_), .Q(core_v3_reg_44_));
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf17), .D(core__0v3_reg_63_0__45_), .Q(core_v3_reg_45_));
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf16), .D(core__0v3_reg_63_0__46_), .Q(core_v3_reg_46_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf27), .D(_0key1_reg_31_0__13_), .Q(core_key_45_));
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf15), .D(core__0v3_reg_63_0__47_), .Q(core_v3_reg_47_));
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf14), .D(core__0v3_reg_63_0__48_), .Q(core_v3_reg_48_));
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf13), .D(core__0v3_reg_63_0__49_), .Q(core_v3_reg_49_));
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf12), .D(core__0v3_reg_63_0__50_), .Q(core_v3_reg_50_));
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf11), .D(core__0v3_reg_63_0__51_), .Q(core_v3_reg_51_));
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf10), .D(core__0v3_reg_63_0__52_), .Q(core_v3_reg_52_));
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf9), .D(core__0v3_reg_63_0__53_), .Q(core_v3_reg_53_));
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf8), .D(core__0v3_reg_63_0__54_), .Q(core_v3_reg_54_));
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf7), .D(core__0v3_reg_63_0__55_), .Q(core_v3_reg_55_));
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf6), .D(core__0v3_reg_63_0__56_), .Q(core_v3_reg_56_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf26), .D(_0key1_reg_31_0__14_), .Q(core_key_46_));
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf5), .D(core__0v3_reg_63_0__57_), .Q(core_v3_reg_57_));
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf4), .D(core__0v3_reg_63_0__58_), .Q(core_v3_reg_58_));
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf3), .D(core__0v3_reg_63_0__59_), .Q(core_v3_reg_59_));
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf2), .D(core__0v3_reg_63_0__60_), .Q(core_v3_reg_60_));
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf1), .D(core__0v3_reg_63_0__61_), .Q(core_v3_reg_61_));
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf0), .D(core__0v3_reg_63_0__62_), .Q(core_v3_reg_62_));
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf84), .D(core__0v3_reg_63_0__63_), .Q(core_v3_reg_63_));
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf83), .D(core__0mi_reg_63_0__0_), .Q(core_mi_reg_0_));
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf82), .D(core__0mi_reg_63_0__1_), .Q(core_mi_reg_1_));
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf81), .D(core__0mi_reg_63_0__2_), .Q(core_mi_reg_2_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf79), .D(_0param_reg_7_0__1_), .Q(core_compression_rounds_1_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf25), .D(_0key1_reg_31_0__15_), .Q(core_key_47_));
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf80), .D(core__0mi_reg_63_0__3_), .Q(core_mi_reg_3_));
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf79), .D(core__0mi_reg_63_0__4_), .Q(core_mi_reg_4_));
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf78), .D(core__0mi_reg_63_0__5_), .Q(core_mi_reg_5_));
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf77), .D(core__0mi_reg_63_0__6_), .Q(core_mi_reg_6_));
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf76), .D(core__0mi_reg_63_0__7_), .Q(core_mi_reg_7_));
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf75), .D(core__0mi_reg_63_0__8_), .Q(core_mi_reg_8_));
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf74), .D(core__0mi_reg_63_0__9_), .Q(core_mi_reg_9_));
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf73), .D(core__0mi_reg_63_0__10_), .Q(core_mi_reg_10_));
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf72), .D(core__0mi_reg_63_0__11_), .Q(core_mi_reg_11_));
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf71), .D(core__0mi_reg_63_0__12_), .Q(core_mi_reg_12_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf24), .D(_0key1_reg_31_0__16_), .Q(core_key_48_));
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf70), .D(core__0mi_reg_63_0__13_), .Q(core_mi_reg_13_));
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf69), .D(core__0mi_reg_63_0__14_), .Q(core_mi_reg_14_));
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf68), .D(core__0mi_reg_63_0__15_), .Q(core_mi_reg_15_));
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf67), .D(core__0mi_reg_63_0__16_), .Q(core_mi_reg_16_));
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf66), .D(core__0mi_reg_63_0__17_), .Q(core_mi_reg_17_));
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf65), .D(core__0mi_reg_63_0__18_), .Q(core_mi_reg_18_));
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf64), .D(core__0mi_reg_63_0__19_), .Q(core_mi_reg_19_));
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf63), .D(core__0mi_reg_63_0__20_), .Q(core_mi_reg_20_));
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf62), .D(core__0mi_reg_63_0__21_), .Q(core_mi_reg_21_));
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf61), .D(core__0mi_reg_63_0__22_), .Q(core_mi_reg_22_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf23), .D(_0key1_reg_31_0__17_), .Q(core_key_49_));
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf60), .D(core__0mi_reg_63_0__23_), .Q(core_mi_reg_23_));
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf59), .D(core__0mi_reg_63_0__24_), .Q(core_mi_reg_24_));
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf58), .D(core__0mi_reg_63_0__25_), .Q(core_mi_reg_25_));
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf57), .D(core__0mi_reg_63_0__26_), .Q(core_mi_reg_26_));
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf56), .D(core__0mi_reg_63_0__27_), .Q(core_mi_reg_27_));
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf55), .D(core__0mi_reg_63_0__28_), .Q(core_mi_reg_28_));
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf54), .D(core__0mi_reg_63_0__29_), .Q(core_mi_reg_29_));
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf53), .D(core__0mi_reg_63_0__30_), .Q(core_mi_reg_30_));
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf52), .D(core__0mi_reg_63_0__31_), .Q(core_mi_reg_31_));
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf51), .D(core__0mi_reg_63_0__32_), .Q(core_mi_reg_32_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf22), .D(_0key1_reg_31_0__18_), .Q(core_key_50_));
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf50), .D(core__0mi_reg_63_0__33_), .Q(core_mi_reg_33_));
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf49), .D(core__0mi_reg_63_0__34_), .Q(core_mi_reg_34_));
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf48), .D(core__0mi_reg_63_0__35_), .Q(core_mi_reg_35_));
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf47), .D(core__0mi_reg_63_0__36_), .Q(core_mi_reg_36_));
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf46), .D(core__0mi_reg_63_0__37_), .Q(core_mi_reg_37_));
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf45), .D(core__0mi_reg_63_0__38_), .Q(core_mi_reg_38_));
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf44), .D(core__0mi_reg_63_0__39_), .Q(core_mi_reg_39_));
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf43), .D(core__0mi_reg_63_0__40_), .Q(core_mi_reg_40_));
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf42), .D(core__0mi_reg_63_0__41_), .Q(core_mi_reg_41_));
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf41), .D(core__0mi_reg_63_0__42_), .Q(core_mi_reg_42_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf21), .D(_0key1_reg_31_0__19_), .Q(core_key_51_));
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf40), .D(core__0mi_reg_63_0__43_), .Q(core_mi_reg_43_));
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf39), .D(core__0mi_reg_63_0__44_), .Q(core_mi_reg_44_));
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf38), .D(core__0mi_reg_63_0__45_), .Q(core_mi_reg_45_));
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf37), .D(core__0mi_reg_63_0__46_), .Q(core_mi_reg_46_));
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf36), .D(core__0mi_reg_63_0__47_), .Q(core_mi_reg_47_));
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf35), .D(core__0mi_reg_63_0__48_), .Q(core_mi_reg_48_));
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf34), .D(core__0mi_reg_63_0__49_), .Q(core_mi_reg_49_));
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf33), .D(core__0mi_reg_63_0__50_), .Q(core_mi_reg_50_));
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf32), .D(core__0mi_reg_63_0__51_), .Q(core_mi_reg_51_));
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf31), .D(core__0mi_reg_63_0__52_), .Q(core_mi_reg_52_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf20), .D(_0key1_reg_31_0__20_), .Q(core_key_52_));
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf30), .D(core__0mi_reg_63_0__53_), .Q(core_mi_reg_53_));
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf29), .D(core__0mi_reg_63_0__54_), .Q(core_mi_reg_54_));
DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf28), .D(core__0mi_reg_63_0__55_), .Q(core_mi_reg_55_));
DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf27), .D(core__0mi_reg_63_0__56_), .Q(core_mi_reg_56_));
DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf26), .D(core__0mi_reg_63_0__57_), .Q(core_mi_reg_57_));
DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf25), .D(core__0mi_reg_63_0__58_), .Q(core_mi_reg_58_));
DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf24), .D(core__0mi_reg_63_0__59_), .Q(core_mi_reg_59_));
DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf23), .D(core__0mi_reg_63_0__60_), .Q(core_mi_reg_60_));
DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf22), .D(core__0mi_reg_63_0__61_), .Q(core_mi_reg_61_));
DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf21), .D(core__0mi_reg_63_0__62_), .Q(core_mi_reg_62_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf19), .D(_0key1_reg_31_0__21_), .Q(core_key_53_));
DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf20), .D(core__0mi_reg_63_0__63_), .Q(core_mi_reg_63_));
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf19), .D(core__0loop_ctr_reg_3_0__0_), .Q(core_loop_ctr_reg_0_));
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf18), .D(core__0loop_ctr_reg_3_0__1_), .Q(core_loop_ctr_reg_1_));
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf17), .D(core__0loop_ctr_reg_3_0__2_), .Q(core_loop_ctr_reg_2_));
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf16), .D(core__0loop_ctr_reg_3_0__3_), .Q(core_loop_ctr_reg_3_));
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf15), .D(core__0ready_reg_0_0_), .Q(core_ready));
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf14), .D(core__0siphash_word0_reg_63_0__0_), .Q(core_siphash_word_0_));
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf13), .D(core__0siphash_word0_reg_63_0__1_), .Q(core_siphash_word_1_));
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf12), .D(core__0siphash_word0_reg_63_0__2_), .Q(core_siphash_word_2_));
DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf11), .D(core__0siphash_word0_reg_63_0__3_), .Q(core_siphash_word_3_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf18), .D(_0key1_reg_31_0__22_), .Q(core_key_54_));
DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf10), .D(core__0siphash_word0_reg_63_0__4_), .Q(core_siphash_word_4_));
DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf9), .D(core__0siphash_word0_reg_63_0__5_), .Q(core_siphash_word_5_));
DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf8), .D(core__0siphash_word0_reg_63_0__6_), .Q(core_siphash_word_6_));
DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf7), .D(core__0siphash_word0_reg_63_0__7_), .Q(core_siphash_word_7_));
DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf6), .D(core__0siphash_word0_reg_63_0__8_), .Q(core_siphash_word_8_));
DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf5), .D(core__0siphash_word0_reg_63_0__9_), .Q(core_siphash_word_9_));
DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf4), .D(core__0siphash_word0_reg_63_0__10_), .Q(core_siphash_word_10_));
DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf3), .D(core__0siphash_word0_reg_63_0__11_), .Q(core_siphash_word_11_));
DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf2), .D(core__0siphash_word0_reg_63_0__12_), .Q(core_siphash_word_12_));
DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf1), .D(core__0siphash_word0_reg_63_0__13_), .Q(core_siphash_word_13_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf17), .D(_0key1_reg_31_0__23_), .Q(core_key_55_));
DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf0), .D(core__0siphash_word0_reg_63_0__14_), .Q(core_siphash_word_14_));
DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_bF_buf84), .D(core__0siphash_word0_reg_63_0__15_), .Q(core_siphash_word_15_));
DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_bF_buf83), .D(core__0siphash_word0_reg_63_0__16_), .Q(core_siphash_word_16_));
DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_bF_buf82), .D(core__0siphash_word0_reg_63_0__17_), .Q(core_siphash_word_17_));
DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_bF_buf81), .D(core__0siphash_word0_reg_63_0__18_), .Q(core_siphash_word_18_));
DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_bF_buf80), .D(core__0siphash_word0_reg_63_0__19_), .Q(core_siphash_word_19_));
DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_bF_buf79), .D(core__0siphash_word0_reg_63_0__20_), .Q(core_siphash_word_20_));
DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_bF_buf78), .D(core__0siphash_word0_reg_63_0__21_), .Q(core_siphash_word_21_));
DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_bF_buf77), .D(core__0siphash_word0_reg_63_0__22_), .Q(core_siphash_word_22_));
DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_bF_buf76), .D(core__0siphash_word0_reg_63_0__23_), .Q(core_siphash_word_23_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf16), .D(_0key1_reg_31_0__24_), .Q(core_key_56_));
DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_bF_buf75), .D(core__0siphash_word0_reg_63_0__24_), .Q(core_siphash_word_24_));
DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_bF_buf74), .D(core__0siphash_word0_reg_63_0__25_), .Q(core_siphash_word_25_));
DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_bF_buf73), .D(core__0siphash_word0_reg_63_0__26_), .Q(core_siphash_word_26_));
DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_bF_buf72), .D(core__0siphash_word0_reg_63_0__27_), .Q(core_siphash_word_27_));
DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_bF_buf71), .D(core__0siphash_word0_reg_63_0__28_), .Q(core_siphash_word_28_));
DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_bF_buf70), .D(core__0siphash_word0_reg_63_0__29_), .Q(core_siphash_word_29_));
DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_bF_buf69), .D(core__0siphash_word0_reg_63_0__30_), .Q(core_siphash_word_30_));
DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_bF_buf68), .D(core__0siphash_word0_reg_63_0__31_), .Q(core_siphash_word_31_));
DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_bF_buf67), .D(core__0siphash_word0_reg_63_0__32_), .Q(core_siphash_word_32_));
DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_bF_buf66), .D(core__0siphash_word0_reg_63_0__33_), .Q(core_siphash_word_33_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf78), .D(_0param_reg_7_0__2_), .Q(core_compression_rounds_2_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf15), .D(_0key1_reg_31_0__25_), .Q(core_key_57_));
DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_bF_buf65), .D(core__0siphash_word0_reg_63_0__34_), .Q(core_siphash_word_34_));
DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_bF_buf64), .D(core__0siphash_word0_reg_63_0__35_), .Q(core_siphash_word_35_));
DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_bF_buf63), .D(core__0siphash_word0_reg_63_0__36_), .Q(core_siphash_word_36_));
DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_bF_buf62), .D(core__0siphash_word0_reg_63_0__37_), .Q(core_siphash_word_37_));
DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_bF_buf61), .D(core__0siphash_word0_reg_63_0__38_), .Q(core_siphash_word_38_));
DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_bF_buf60), .D(core__0siphash_word0_reg_63_0__39_), .Q(core_siphash_word_39_));
DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_bF_buf59), .D(core__0siphash_word0_reg_63_0__40_), .Q(core_siphash_word_40_));
DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_bF_buf58), .D(core__0siphash_word0_reg_63_0__41_), .Q(core_siphash_word_41_));
DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_bF_buf57), .D(core__0siphash_word0_reg_63_0__42_), .Q(core_siphash_word_42_));
DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_bF_buf56), .D(core__0siphash_word0_reg_63_0__43_), .Q(core_siphash_word_43_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf14), .D(_0key1_reg_31_0__26_), .Q(core_key_58_));
DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_bF_buf55), .D(core__0siphash_word0_reg_63_0__44_), .Q(core_siphash_word_44_));
DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_bF_buf54), .D(core__0siphash_word0_reg_63_0__45_), .Q(core_siphash_word_45_));
DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_bF_buf53), .D(core__0siphash_word0_reg_63_0__46_), .Q(core_siphash_word_46_));
DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_bF_buf52), .D(core__0siphash_word0_reg_63_0__47_), .Q(core_siphash_word_47_));
DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_bF_buf51), .D(core__0siphash_word0_reg_63_0__48_), .Q(core_siphash_word_48_));
DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_bF_buf50), .D(core__0siphash_word0_reg_63_0__49_), .Q(core_siphash_word_49_));
DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_bF_buf49), .D(core__0siphash_word0_reg_63_0__50_), .Q(core_siphash_word_50_));
DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_bF_buf48), .D(core__0siphash_word0_reg_63_0__51_), .Q(core_siphash_word_51_));
DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_bF_buf47), .D(core__0siphash_word0_reg_63_0__52_), .Q(core_siphash_word_52_));
DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_bF_buf46), .D(core__0siphash_word0_reg_63_0__53_), .Q(core_siphash_word_53_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf13), .D(_0key1_reg_31_0__27_), .Q(core_key_59_));
DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_bF_buf45), .D(core__0siphash_word0_reg_63_0__54_), .Q(core_siphash_word_54_));
DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_bF_buf44), .D(core__0siphash_word0_reg_63_0__55_), .Q(core_siphash_word_55_));
DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_bF_buf43), .D(core__0siphash_word0_reg_63_0__56_), .Q(core_siphash_word_56_));
DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_bF_buf42), .D(core__0siphash_word0_reg_63_0__57_), .Q(core_siphash_word_57_));
DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_bF_buf41), .D(core__0siphash_word0_reg_63_0__58_), .Q(core_siphash_word_58_));
DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_bF_buf40), .D(core__0siphash_word0_reg_63_0__59_), .Q(core_siphash_word_59_));
DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_bF_buf39), .D(core__0siphash_word0_reg_63_0__60_), .Q(core_siphash_word_60_));
DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_bF_buf38), .D(core__0siphash_word0_reg_63_0__61_), .Q(core_siphash_word_61_));
DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_bF_buf37), .D(core__0siphash_word0_reg_63_0__62_), .Q(core_siphash_word_62_));
DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_bF_buf36), .D(core__0siphash_word0_reg_63_0__63_), .Q(core_siphash_word_63_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf12), .D(_0key1_reg_31_0__28_), .Q(core_key_60_));
DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_bF_buf35), .D(core__0siphash_word1_reg_63_0__0_), .Q(core_siphash_word_64_));
DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_bF_buf34), .D(core__0siphash_word1_reg_63_0__1_), .Q(core_siphash_word_65_));
DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_bF_buf33), .D(core__0siphash_word1_reg_63_0__2_), .Q(core_siphash_word_66_));
DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_bF_buf32), .D(core__0siphash_word1_reg_63_0__3_), .Q(core_siphash_word_67_));
DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_bF_buf31), .D(core__0siphash_word1_reg_63_0__4_), .Q(core_siphash_word_68_));
DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_bF_buf30), .D(core__0siphash_word1_reg_63_0__5_), .Q(core_siphash_word_69_));
DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_bF_buf29), .D(core__0siphash_word1_reg_63_0__6_), .Q(core_siphash_word_70_));
DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_bF_buf28), .D(core__0siphash_word1_reg_63_0__7_), .Q(core_siphash_word_71_));
DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_bF_buf27), .D(core__0siphash_word1_reg_63_0__8_), .Q(core_siphash_word_72_));
DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_bF_buf26), .D(core__0siphash_word1_reg_63_0__9_), .Q(core_siphash_word_73_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf11), .D(_0key1_reg_31_0__29_), .Q(core_key_61_));
DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_bF_buf25), .D(core__0siphash_word1_reg_63_0__10_), .Q(core_siphash_word_74_));
DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_bF_buf24), .D(core__0siphash_word1_reg_63_0__11_), .Q(core_siphash_word_75_));
DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_bF_buf23), .D(core__0siphash_word1_reg_63_0__12_), .Q(core_siphash_word_76_));
DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_bF_buf22), .D(core__0siphash_word1_reg_63_0__13_), .Q(core_siphash_word_77_));
DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_bF_buf21), .D(core__0siphash_word1_reg_63_0__14_), .Q(core_siphash_word_78_));
DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_bF_buf20), .D(core__0siphash_word1_reg_63_0__15_), .Q(core_siphash_word_79_));
DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_bF_buf19), .D(core__0siphash_word1_reg_63_0__16_), .Q(core_siphash_word_80_));
DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_bF_buf18), .D(core__0siphash_word1_reg_63_0__17_), .Q(core_siphash_word_81_));
DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_bF_buf17), .D(core__0siphash_word1_reg_63_0__18_), .Q(core_siphash_word_82_));
DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_bF_buf16), .D(core__0siphash_word1_reg_63_0__19_), .Q(core_siphash_word_83_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf10), .D(_0key1_reg_31_0__30_), .Q(core_key_62_));
DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_bF_buf15), .D(core__0siphash_word1_reg_63_0__20_), .Q(core_siphash_word_84_));
DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_bF_buf14), .D(core__0siphash_word1_reg_63_0__21_), .Q(core_siphash_word_85_));
DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_bF_buf13), .D(core__0siphash_word1_reg_63_0__22_), .Q(core_siphash_word_86_));
DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_bF_buf12), .D(core__0siphash_word1_reg_63_0__23_), .Q(core_siphash_word_87_));
DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_bF_buf11), .D(core__0siphash_word1_reg_63_0__24_), .Q(core_siphash_word_88_));
DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_bF_buf10), .D(core__0siphash_word1_reg_63_0__25_), .Q(core_siphash_word_89_));
DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_bF_buf9), .D(core__0siphash_word1_reg_63_0__26_), .Q(core_siphash_word_90_));
DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_bF_buf8), .D(core__0siphash_word1_reg_63_0__27_), .Q(core_siphash_word_91_));
DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_bF_buf7), .D(core__0siphash_word1_reg_63_0__28_), .Q(core_siphash_word_92_));
DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_bF_buf6), .D(core__0siphash_word1_reg_63_0__29_), .Q(core_siphash_word_93_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf9), .D(_0key1_reg_31_0__31_), .Q(core_key_63_));
DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_bF_buf5), .D(core__0siphash_word1_reg_63_0__30_), .Q(core_siphash_word_94_));
DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_bF_buf4), .D(core__0siphash_word1_reg_63_0__31_), .Q(core_siphash_word_95_));
DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_bF_buf3), .D(core__0siphash_word1_reg_63_0__32_), .Q(core_siphash_word_96_));
DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_bF_buf2), .D(core__0siphash_word1_reg_63_0__33_), .Q(core_siphash_word_97_));
DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_bF_buf1), .D(core__0siphash_word1_reg_63_0__34_), .Q(core_siphash_word_98_));
DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_bF_buf0), .D(core__0siphash_word1_reg_63_0__35_), .Q(core_siphash_word_99_));
DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_bF_buf84), .D(core__0siphash_word1_reg_63_0__36_), .Q(core_siphash_word_100_));
DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_bF_buf83), .D(core__0siphash_word1_reg_63_0__37_), .Q(core_siphash_word_101_));
DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_bF_buf82), .D(core__0siphash_word1_reg_63_0__38_), .Q(core_siphash_word_102_));
DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_bF_buf81), .D(core__0siphash_word1_reg_63_0__39_), .Q(core_siphash_word_103_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf8), .D(_0key2_reg_31_0__0_), .Q(core_key_64_));
DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_bF_buf80), .D(core__0siphash_word1_reg_63_0__40_), .Q(core_siphash_word_104_));
DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_bF_buf79), .D(core__0siphash_word1_reg_63_0__41_), .Q(core_siphash_word_105_));
DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_bF_buf78), .D(core__0siphash_word1_reg_63_0__42_), .Q(core_siphash_word_106_));
DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_bF_buf77), .D(core__0siphash_word1_reg_63_0__43_), .Q(core_siphash_word_107_));
DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_bF_buf76), .D(core__0siphash_word1_reg_63_0__44_), .Q(core_siphash_word_108_));
DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_bF_buf75), .D(core__0siphash_word1_reg_63_0__45_), .Q(core_siphash_word_109_));
DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_bF_buf74), .D(core__0siphash_word1_reg_63_0__46_), .Q(core_siphash_word_110_));
DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_bF_buf73), .D(core__0siphash_word1_reg_63_0__47_), .Q(core_siphash_word_111_));
DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_bF_buf72), .D(core__0siphash_word1_reg_63_0__48_), .Q(core_siphash_word_112_));
DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_bF_buf71), .D(core__0siphash_word1_reg_63_0__49_), .Q(core_siphash_word_113_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf7), .D(_0key2_reg_31_0__1_), .Q(core_key_65_));
DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_bF_buf70), .D(core__0siphash_word1_reg_63_0__50_), .Q(core_siphash_word_114_));
DFFPOSX1 DFFPOSX1_781 ( .CLK(clk_bF_buf69), .D(core__0siphash_word1_reg_63_0__51_), .Q(core_siphash_word_115_));
DFFPOSX1 DFFPOSX1_782 ( .CLK(clk_bF_buf68), .D(core__0siphash_word1_reg_63_0__52_), .Q(core_siphash_word_116_));
DFFPOSX1 DFFPOSX1_783 ( .CLK(clk_bF_buf67), .D(core__0siphash_word1_reg_63_0__53_), .Q(core_siphash_word_117_));
DFFPOSX1 DFFPOSX1_784 ( .CLK(clk_bF_buf66), .D(core__0siphash_word1_reg_63_0__54_), .Q(core_siphash_word_118_));
DFFPOSX1 DFFPOSX1_785 ( .CLK(clk_bF_buf65), .D(core__0siphash_word1_reg_63_0__55_), .Q(core_siphash_word_119_));
DFFPOSX1 DFFPOSX1_786 ( .CLK(clk_bF_buf64), .D(core__0siphash_word1_reg_63_0__56_), .Q(core_siphash_word_120_));
DFFPOSX1 DFFPOSX1_787 ( .CLK(clk_bF_buf63), .D(core__0siphash_word1_reg_63_0__57_), .Q(core_siphash_word_121_));
DFFPOSX1 DFFPOSX1_788 ( .CLK(clk_bF_buf62), .D(core__0siphash_word1_reg_63_0__58_), .Q(core_siphash_word_122_));
DFFPOSX1 DFFPOSX1_789 ( .CLK(clk_bF_buf61), .D(core__0siphash_word1_reg_63_0__59_), .Q(core_siphash_word_123_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf6), .D(_0key2_reg_31_0__2_), .Q(core_key_66_));
DFFPOSX1 DFFPOSX1_790 ( .CLK(clk_bF_buf60), .D(core__0siphash_word1_reg_63_0__60_), .Q(core_siphash_word_124_));
DFFPOSX1 DFFPOSX1_791 ( .CLK(clk_bF_buf59), .D(core__0siphash_word1_reg_63_0__61_), .Q(core_siphash_word_125_));
DFFPOSX1 DFFPOSX1_792 ( .CLK(clk_bF_buf58), .D(core__0siphash_word1_reg_63_0__62_), .Q(core_siphash_word_126_));
DFFPOSX1 DFFPOSX1_793 ( .CLK(clk_bF_buf57), .D(core__0siphash_word1_reg_63_0__63_), .Q(core_siphash_word_127_));
DFFPOSX1 DFFPOSX1_794 ( .CLK(clk_bF_buf56), .D(core__0siphash_valid_reg_0_0_), .Q(core_siphash_valid_reg));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf77), .D(_0param_reg_7_0__3_), .Q(core_compression_rounds_3_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf5), .D(_0key2_reg_31_0__3_), .Q(core_key_67_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf4), .D(_0key2_reg_31_0__4_), .Q(core_key_68_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf3), .D(_0key2_reg_31_0__5_), .Q(core_key_69_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf2), .D(_0key2_reg_31_0__6_), .Q(core_key_70_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf1), .D(_0key2_reg_31_0__7_), .Q(core_key_71_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf0), .D(_0key2_reg_31_0__8_), .Q(core_key_72_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf84), .D(_0key2_reg_31_0__9_), .Q(core_key_73_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf83), .D(_0key2_reg_31_0__10_), .Q(core_key_74_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf82), .D(_0key2_reg_31_0__11_), .Q(core_key_75_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf81), .D(_0key2_reg_31_0__12_), .Q(core_key_76_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf76), .D(_0param_reg_7_0__4_), .Q(core_final_rounds_0_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf80), .D(_0key2_reg_31_0__13_), .Q(core_key_77_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf79), .D(_0key2_reg_31_0__14_), .Q(core_key_78_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf78), .D(_0key2_reg_31_0__15_), .Q(core_key_79_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf77), .D(_0key2_reg_31_0__16_), .Q(core_key_80_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf76), .D(_0key2_reg_31_0__17_), .Q(core_key_81_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf75), .D(_0key2_reg_31_0__18_), .Q(core_key_82_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf74), .D(_0key2_reg_31_0__19_), .Q(core_key_83_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf73), .D(_0key2_reg_31_0__20_), .Q(core_key_84_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf72), .D(_0key2_reg_31_0__21_), .Q(core_key_85_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf71), .D(_0key2_reg_31_0__22_), .Q(core_key_86_));
INVX1 INVX1_1 ( .A(core_initalize), .Y(_abc_19873_new_n870_));
INVX1 INVX1_10 ( .A(core_key_96_), .Y(_abc_19873_new_n910_));
INVX1 INVX1_100 ( .A(word0_reg_11_), .Y(_abc_19873_new_n1150_));
INVX1 INVX1_1000 ( .A(core__abc_21302_new_n5089_), .Y(core__abc_21302_new_n5107_));
INVX1 INVX1_1001 ( .A(core__abc_21302_new_n5109_), .Y(core__abc_21302_new_n5110_));
INVX1 INVX1_1002 ( .A(core__abc_21302_new_n5111_), .Y(core__abc_21302_new_n5112_));
INVX1 INVX1_1003 ( .A(core_v1_reg_21_), .Y(core__abc_21302_new_n5113_));
INVX1 INVX1_1004 ( .A(core__abc_21302_new_n5114_), .Y(core__abc_21302_new_n5115_));
INVX1 INVX1_1005 ( .A(core__abc_21302_new_n5116_), .Y(core__abc_21302_new_n5118_));
INVX1 INVX1_1006 ( .A(core_key_3_), .Y(core__abc_21302_new_n5131_));
INVX1 INVX1_1007 ( .A(core_v1_reg_22_), .Y(core__abc_21302_new_n5136_));
INVX1 INVX1_1008 ( .A(core__abc_21302_new_n5135_), .Y(core__abc_21302_new_n5140_));
INVX1 INVX1_1009 ( .A(core__abc_21302_new_n5137_), .Y(core__abc_21302_new_n5141_));
INVX1 INVX1_101 ( .A(core_mi_43_), .Y(_abc_19873_new_n1151_));
INVX1 INVX1_1010 ( .A(core__abc_21302_new_n5138_), .Y(core__abc_21302_new_n5142_));
INVX1 INVX1_1011 ( .A(core__abc_21302_new_n5159_), .Y(core__abc_21302_new_n5160_));
INVX1 INVX1_1012 ( .A(core__abc_21302_new_n5154_), .Y(core__abc_21302_new_n5164_));
INVX1 INVX1_1013 ( .A(core__abc_21302_new_n5161_), .Y(core__abc_21302_new_n5165_));
INVX1 INVX1_1014 ( .A(core__abc_21302_new_n5166_), .Y(core__abc_21302_new_n5174_));
INVX1 INVX1_1015 ( .A(core__abc_21302_new_n5188_), .Y(core__abc_21302_new_n5190_));
INVX1 INVX1_1016 ( .A(core__abc_21302_new_n5196_), .Y(core__abc_21302_new_n5197_));
INVX1 INVX1_1017 ( .A(core__abc_21302_new_n5191_), .Y(core__abc_21302_new_n5205_));
INVX1 INVX1_1018 ( .A(core__abc_21302_new_n5207_), .Y(core__abc_21302_new_n5208_));
INVX1 INVX1_1019 ( .A(core_v1_reg_26_), .Y(core__abc_21302_new_n5210_));
INVX1 INVX1_102 ( .A(core_mi_12_), .Y(_abc_19873_new_n1155_));
INVX1 INVX1_1020 ( .A(core__abc_21302_new_n5216_), .Y(core__abc_21302_new_n5218_));
INVX1 INVX1_1021 ( .A(core_key_7_), .Y(core__abc_21302_new_n5221_));
INVX1 INVX1_1022 ( .A(core__abc_21302_new_n5227_), .Y(core__abc_21302_new_n5228_));
INVX1 INVX1_1023 ( .A(core__abc_21302_new_n4175_), .Y(core__abc_21302_new_n5236_));
INVX1 INVX1_1024 ( .A(core__abc_21302_new_n5239_), .Y(core__abc_21302_new_n5240_));
INVX1 INVX1_1025 ( .A(core_v1_reg_28_), .Y(core__abc_21302_new_n5248_));
INVX1 INVX1_1026 ( .A(core__abc_21302_new_n5251_), .Y(core__abc_21302_new_n5264_));
INVX1 INVX1_1027 ( .A(core__abc_21302_new_n5265_), .Y(core__abc_21302_new_n5266_));
INVX1 INVX1_1028 ( .A(core_v1_reg_29_), .Y(core__abc_21302_new_n5268_));
INVX1 INVX1_1029 ( .A(core__abc_21302_new_n5278_), .Y(core__abc_21302_new_n5279_));
INVX1 INVX1_103 ( .A(core_key_108_), .Y(_abc_19873_new_n1156_));
INVX1 INVX1_1030 ( .A(core__abc_21302_new_n5286_), .Y(core__abc_21302_new_n5287_));
INVX1 INVX1_1031 ( .A(core__abc_21302_new_n4255_), .Y(core__abc_21302_new_n5290_));
INVX1 INVX1_1032 ( .A(core__abc_21302_new_n5288_), .Y(core__abc_21302_new_n5291_));
INVX1 INVX1_1033 ( .A(core_key_11_), .Y(core__abc_21302_new_n5297_));
INVX1 INVX1_1034 ( .A(core__abc_21302_new_n5272_), .Y(core__abc_21302_new_n5304_));
INVX1 INVX1_1035 ( .A(core__abc_21302_new_n5307_), .Y(core__abc_21302_new_n5308_));
INVX1 INVX1_1036 ( .A(core_v1_reg_31_), .Y(core__abc_21302_new_n5311_));
INVX1 INVX1_1037 ( .A(core__abc_21302_new_n5315_), .Y(core__abc_21302_new_n5322_));
INVX1 INVX1_1038 ( .A(core_v1_reg_32_), .Y(core__abc_21302_new_n5325_));
INVX1 INVX1_1039 ( .A(core__abc_21302_new_n5328_), .Y(core__abc_21302_new_n5330_));
INVX1 INVX1_104 ( .A(core_key_76_), .Y(_abc_19873_new_n1158_));
INVX1 INVX1_1040 ( .A(core__abc_21302_new_n5332_), .Y(core__abc_21302_new_n5333_));
INVX1 INVX1_1041 ( .A(core__abc_21302_new_n5343_), .Y(core__abc_21302_new_n5344_));
INVX1 INVX1_1042 ( .A(core__abc_21302_new_n5346_), .Y(core__abc_21302_new_n5347_));
INVX1 INVX1_1043 ( .A(core__abc_21302_new_n5351_), .Y(core__abc_21302_new_n5354_));
INVX1 INVX1_1044 ( .A(core__abc_21302_new_n5345_), .Y(core__abc_21302_new_n5358_));
INVX1 INVX1_1045 ( .A(core__abc_21302_new_n5368_), .Y(core__abc_21302_new_n5372_));
INVX1 INVX1_1046 ( .A(core__abc_21302_new_n5375_), .Y(core__abc_21302_new_n5376_));
INVX1 INVX1_1047 ( .A(core__abc_21302_new_n5355_), .Y(core__abc_21302_new_n5378_));
INVX1 INVX1_1048 ( .A(core_key_15_), .Y(core__abc_21302_new_n5382_));
INVX1 INVX1_1049 ( .A(core__abc_21302_new_n5391_), .Y(core__abc_21302_new_n5392_));
INVX1 INVX1_105 ( .A(core_key_12_), .Y(_abc_19873_new_n1166_));
INVX1 INVX1_1050 ( .A(core__abc_21302_new_n5404_), .Y(core__abc_21302_new_n5405_));
INVX1 INVX1_1051 ( .A(core__abc_21302_new_n5408_), .Y(core__abc_21302_new_n5419_));
INVX1 INVX1_1052 ( .A(core_v1_reg_36_), .Y(core__abc_21302_new_n5422_));
INVX1 INVX1_1053 ( .A(core__abc_21302_new_n5435_), .Y(core__abc_21302_new_n5436_));
INVX1 INVX1_1054 ( .A(core__abc_21302_new_n5439_), .Y(core__abc_21302_new_n5440_));
INVX1 INVX1_1055 ( .A(core__abc_21302_new_n5447_), .Y(core__abc_21302_new_n5448_));
INVX1 INVX1_1056 ( .A(core_key_19_), .Y(core__abc_21302_new_n5460_));
INVX1 INVX1_1057 ( .A(core__abc_21302_new_n5455_), .Y(core__abc_21302_new_n5466_));
INVX1 INVX1_1058 ( .A(core__abc_21302_new_n5443_), .Y(core__abc_21302_new_n5473_));
INVX1 INVX1_1059 ( .A(core__abc_21302_new_n5474_), .Y(core__abc_21302_new_n5475_));
INVX1 INVX1_106 ( .A(word0_reg_12_), .Y(_abc_19873_new_n1169_));
INVX1 INVX1_1060 ( .A(core_v1_reg_39_), .Y(core__abc_21302_new_n5478_));
INVX1 INVX1_1061 ( .A(core__abc_21302_new_n5479_), .Y(core__abc_21302_new_n5480_));
INVX1 INVX1_1062 ( .A(core__abc_21302_new_n5481_), .Y(core__abc_21302_new_n5482_));
INVX1 INVX1_1063 ( .A(core__abc_21302_new_n5492_), .Y(core__abc_21302_new_n5498_));
INVX1 INVX1_1064 ( .A(core__abc_21302_new_n5496_), .Y(core__abc_21302_new_n5499_));
INVX1 INVX1_1065 ( .A(core_v1_reg_41_), .Y(core__abc_21302_new_n5507_));
INVX1 INVX1_1066 ( .A(core__abc_21302_new_n5509_), .Y(core__abc_21302_new_n5511_));
INVX1 INVX1_1067 ( .A(core__abc_21302_new_n5514_), .Y(core__abc_21302_new_n5515_));
INVX1 INVX1_1068 ( .A(core__abc_21302_new_n5517_), .Y(core__abc_21302_new_n5518_));
INVX1 INVX1_1069 ( .A(core__abc_21302_new_n5519_), .Y(core__abc_21302_new_n5520_));
INVX1 INVX1_107 ( .A(core_mi_44_), .Y(_abc_19873_new_n1170_));
INVX1 INVX1_1070 ( .A(core_v1_reg_42_), .Y(core__abc_21302_new_n5528_));
INVX1 INVX1_1071 ( .A(core__abc_21302_new_n5510_), .Y(core__abc_21302_new_n5536_));
INVX1 INVX1_1072 ( .A(core__abc_21302_new_n5534_), .Y(core__abc_21302_new_n5537_));
INVX1 INVX1_1073 ( .A(core_key_23_), .Y(core__abc_21302_new_n5540_));
INVX1 INVX1_1074 ( .A(core__abc_21302_new_n5531_), .Y(core__abc_21302_new_n5548_));
INVX1 INVX1_1075 ( .A(core__abc_21302_new_n5555_), .Y(core__abc_21302_new_n5556_));
INVX1 INVX1_1076 ( .A(core__abc_21302_new_n5558_), .Y(core__abc_21302_new_n5559_));
INVX1 INVX1_1077 ( .A(core__abc_21302_new_n5560_), .Y(core__abc_21302_new_n5570_));
INVX1 INVX1_1078 ( .A(core__abc_21302_new_n5588_), .Y(core__abc_21302_new_n5589_));
INVX1 INVX1_1079 ( .A(core__abc_21302_new_n5592_), .Y(core__abc_21302_new_n5593_));
INVX1 INVX1_108 ( .A(core_key_45_), .Y(_abc_19873_new_n1174_));
INVX1 INVX1_1080 ( .A(core_v1_reg_46_), .Y(core__abc_21302_new_n5601_));
INVX1 INVX1_1081 ( .A(core__abc_21302_new_n5603_), .Y(core__abc_21302_new_n5605_));
INVX1 INVX1_1082 ( .A(core__abc_21302_new_n5585_), .Y(core__abc_21302_new_n5609_));
INVX1 INVX1_1083 ( .A(core__abc_21302_new_n5607_), .Y(core__abc_21302_new_n5610_));
INVX1 INVX1_1084 ( .A(core__abc_21302_new_n5618_), .Y(core__abc_21302_new_n5619_));
INVX1 INVX1_1085 ( .A(core__abc_21302_new_n5617_), .Y(core__abc_21302_new_n5621_));
INVX1 INVX1_1086 ( .A(core__abc_21302_new_n5625_), .Y(core__abc_21302_new_n5626_));
INVX1 INVX1_1087 ( .A(core__abc_21302_new_n5552_), .Y(core__abc_21302_new_n5632_));
INVX1 INVX1_1088 ( .A(core__abc_21302_new_n5629_), .Y(core__abc_21302_new_n5636_));
INVX1 INVX1_1089 ( .A(core_v1_reg_48_), .Y(core__abc_21302_new_n5646_));
INVX1 INVX1_109 ( .A(core_key_13_), .Y(_abc_19873_new_n1175_));
INVX1 INVX1_1090 ( .A(core__abc_21302_new_n5627_), .Y(core__abc_21302_new_n5651_));
INVX1 INVX1_1091 ( .A(core__abc_21302_new_n5665_), .Y(core__abc_21302_new_n5666_));
INVX1 INVX1_1092 ( .A(core__abc_21302_new_n5673_), .Y(core__abc_21302_new_n5674_));
INVX1 INVX1_1093 ( .A(core__abc_21302_new_n5683_), .Y(core__abc_21302_new_n5684_));
INVX1 INVX1_1094 ( .A(core_v1_reg_50_), .Y(core__abc_21302_new_n5685_));
INVX1 INVX1_1095 ( .A(core__abc_21302_new_n5688_), .Y(core__abc_21302_new_n5689_));
INVX1 INVX1_1096 ( .A(core_key_31_), .Y(core__abc_21302_new_n5694_));
INVX1 INVX1_1097 ( .A(core__abc_21302_new_n5700_), .Y(core__abc_21302_new_n5701_));
INVX1 INVX1_1098 ( .A(core__abc_21302_new_n5045_), .Y(core__abc_21302_new_n5708_));
INVX1 INVX1_1099 ( .A(core_key_35_), .Y(core__abc_21302_new_n5723_));
INVX1 INVX1_11 ( .A(core_compression_rounds_0_), .Y(_abc_19873_new_n916_));
INVX1 INVX1_110 ( .A(word2_reg_13_), .Y(_abc_19873_new_n1177_));
INVX1 INVX1_1100 ( .A(core_v2_reg_36_), .Y(core__abc_21302_new_n5728_));
INVX1 INVX1_1101 ( .A(core__abc_21302_new_n5729_), .Y(core__abc_21302_new_n5730_));
INVX1 INVX1_1102 ( .A(core__abc_21302_new_n5026_), .Y(core__abc_21302_new_n5753_));
INVX1 INVX1_1103 ( .A(core__abc_21302_new_n5028_), .Y(core__abc_21302_new_n5754_));
INVX1 INVX1_1104 ( .A(core_key_39_), .Y(core__abc_21302_new_n5758_));
INVX1 INVX1_1105 ( .A(core_v2_reg_40_), .Y(core__abc_21302_new_n5766_));
INVX1 INVX1_1106 ( .A(core__abc_21302_new_n5775_), .Y(core__abc_21302_new_n5776_));
INVX1 INVX1_1107 ( .A(core__abc_21302_new_n4992_), .Y(core__abc_21302_new_n5797_));
INVX1 INVX1_1108 ( .A(core__abc_21302_new_n5006_), .Y(core__abc_21302_new_n5798_));
INVX1 INVX1_1109 ( .A(core__abc_21302_new_n5801_), .Y(core__abc_21302_new_n5802_));
INVX1 INVX1_111 ( .A(core_key_109_), .Y(_abc_19873_new_n1179_));
INVX1 INVX1_1110 ( .A(core_v2_reg_47_), .Y(core__abc_21302_new_n5828_));
INVX1 INVX1_1111 ( .A(core__abc_21302_new_n4974_), .Y(core__abc_21302_new_n5830_));
INVX1 INVX1_1112 ( .A(core__abc_21302_new_n4987_), .Y(core__abc_21302_new_n5838_));
INVX1 INVX1_1113 ( .A(core__abc_21302_new_n5841_), .Y(core__abc_21302_new_n5849_));
INVX1 INVX1_1114 ( .A(core__abc_21302_new_n5860_), .Y(core__abc_21302_new_n5861_));
INVX1 INVX1_1115 ( .A(core_key_50_), .Y(core__abc_21302_new_n5865_));
INVX1 INVX1_1116 ( .A(core__abc_21302_new_n5879_), .Y(core__abc_21302_new_n5880_));
INVX1 INVX1_1117 ( .A(core__abc_21302_new_n5892_), .Y(core__abc_21302_new_n5893_));
INVX1 INVX1_1118 ( .A(core__abc_21302_new_n4915_), .Y(core__abc_21302_new_n5899_));
INVX1 INVX1_1119 ( .A(core__abc_21302_new_n5909_), .Y(core__abc_21302_new_n5910_));
INVX1 INVX1_112 ( .A(core_key_77_), .Y(_abc_19873_new_n1180_));
INVX1 INVX1_1120 ( .A(core_key_55_), .Y(core__abc_21302_new_n5915_));
INVX1 INVX1_1121 ( .A(core__abc_21302_new_n5923_), .Y(core__abc_21302_new_n5924_));
INVX1 INVX1_1122 ( .A(core__abc_21302_new_n5955_), .Y(core__abc_21302_new_n5956_));
INVX1 INVX1_1123 ( .A(core__abc_21302_new_n5957_), .Y(core__abc_21302_new_n5958_));
INVX1 INVX1_1124 ( .A(core__abc_21302_new_n5965_), .Y(core__abc_21302_new_n5967_));
INVX1 INVX1_1125 ( .A(core__abc_21302_new_n5954_), .Y(core__abc_21302_new_n5968_));
INVX1 INVX1_1126 ( .A(core_key_63_), .Y(core__abc_21302_new_n5985_));
INVX1 INVX1_1127 ( .A(core__abc_21302_new_n2641_), .Y(core__abc_21302_new_n5997_));
INVX1 INVX1_1128 ( .A(core__abc_21302_new_n5702_), .Y(core__abc_21302_new_n6001_));
INVX1 INVX1_1129 ( .A(core__abc_21302_new_n5721_), .Y(core__abc_21302_new_n6023_));
INVX1 INVX1_113 ( .A(core_mi_45_), .Y(_abc_19873_new_n1183_));
INVX1 INVX1_1130 ( .A(core__abc_21302_new_n5739_), .Y(core__abc_21302_new_n6038_));
INVX1 INVX1_1131 ( .A(core__abc_21302_new_n5584_), .Y(core__abc_21302_new_n6081_));
INVX1 INVX1_1132 ( .A(core__abc_21302_new_n5647_), .Y(core__abc_21302_new_n6100_));
INVX1 INVX1_1133 ( .A(core__abc_21302_new_n5041_), .Y(core__abc_21302_new_n6132_));
INVX1 INVX1_1134 ( .A(core_v1_reg_20_), .Y(core__abc_21302_new_n6142_));
INVX1 INVX1_1135 ( .A(core_v1_reg_23_), .Y(core__abc_21302_new_n6162_));
INVX1 INVX1_1136 ( .A(core_v1_reg_25_), .Y(core__abc_21302_new_n6176_));
INVX1 INVX1_1137 ( .A(core_v1_reg_30_), .Y(core__abc_21302_new_n6207_));
INVX1 INVX1_1138 ( .A(core__abc_21302_new_n4950_), .Y(core__abc_21302_new_n6245_));
INVX1 INVX1_1139 ( .A(core__abc_21302_new_n4872_), .Y(core__abc_21302_new_n6282_));
INVX1 INVX1_114 ( .A(core_mi_13_), .Y(_abc_19873_new_n1184_));
INVX1 INVX1_1140 ( .A(core_v1_reg_44_), .Y(core__abc_21302_new_n6304_));
INVX1 INVX1_1141 ( .A(core__abc_21302_new_n6316_), .Y(core__abc_21302_new_n6317_));
INVX1 INVX1_1142 ( .A(core__abc_21302_new_n6330_), .Y(core__abc_21302_new_n6331_));
INVX1 INVX1_1143 ( .A(core__abc_21302_new_n5074_), .Y(core__abc_21302_new_n6337_));
INVX1 INVX1_1144 ( .A(core__abc_21302_new_n5446_), .Y(core__abc_21302_new_n6345_));
INVX1 INVX1_1145 ( .A(core_v1_reg_51_), .Y(core__abc_21302_new_n6354_));
INVX1 INVX1_1146 ( .A(core__abc_21302_new_n5237_), .Y(core__abc_21302_new_n6393_));
INVX1 INVX1_1147 ( .A(core__abc_21302_new_n5271_), .Y(core__abc_21302_new_n6411_));
INVX1 INVX1_1148 ( .A(core__abc_21302_new_n6418_), .Y(core__abc_21302_new_n6419_));
INVX1 INVX1_1149 ( .A(core_key_124_), .Y(core__abc_21302_new_n6422_));
INVX1 INVX1_115 ( .A(core_mi_14_), .Y(_abc_19873_new_n1192_));
INVX1 INVX1_1150 ( .A(core__abc_21302_new_n6464_), .Y(core__abc_21302_new_n6465_));
INVX1 INVX1_1151 ( .A(core__abc_21302_new_n2863_), .Y(core__abc_21302_new_n6492_));
INVX1 INVX1_1152 ( .A(core_key_9_), .Y(core__abc_21302_new_n6514_));
INVX1 INVX1_1153 ( .A(core_key_12_), .Y(core__abc_21302_new_n6536_));
INVX1 INVX1_1154 ( .A(core_key_18_), .Y(core__abc_21302_new_n6579_));
INVX1 INVX1_1155 ( .A(core__abc_21302_new_n3646_), .Y(core__abc_21302_new_n6623_));
INVX1 INVX1_1156 ( .A(core_key_25_), .Y(core__abc_21302_new_n6629_));
INVX1 INVX1_1157 ( .A(core_key_26_), .Y(core__abc_21302_new_n6637_));
INVX1 INVX1_1158 ( .A(core_key_27_), .Y(core__abc_21302_new_n6645_));
INVX1 INVX1_1159 ( .A(core_key_41_), .Y(core__abc_21302_new_n6740_));
INVX1 INVX1_116 ( .A(core_key_110_), .Y(_abc_19873_new_n1193_));
INVX1 INVX1_1160 ( .A(core_key_52_), .Y(core__abc_21302_new_n6817_));
INVX1 INVX1_1161 ( .A(core_key_58_), .Y(core__abc_21302_new_n6861_));
INVX1 INVX1_1162 ( .A(core_key_59_), .Y(core__abc_21302_new_n6869_));
INVX1 INVX1_1163 ( .A(core_long), .Y(core__abc_21302_new_n6909_));
INVX1 INVX1_117 ( .A(core_key_78_), .Y(_abc_19873_new_n1195_));
INVX1 INVX1_118 ( .A(word0_reg_14_), .Y(_abc_19873_new_n1198_));
INVX1 INVX1_119 ( .A(core_key_46_), .Y(_abc_19873_new_n1205_));
INVX1 INVX1_12 ( .A(word3_reg_0_), .Y(_abc_19873_new_n921_));
INVX1 INVX1_120 ( .A(core_key_14_), .Y(_abc_19873_new_n1206_));
INVX1 INVX1_121 ( .A(word3_reg_15_), .Y(_abc_19873_new_n1210_));
INVX1 INVX1_122 ( .A(core_key_111_), .Y(_abc_19873_new_n1212_));
INVX1 INVX1_123 ( .A(core_key_79_), .Y(_abc_19873_new_n1213_));
INVX1 INVX1_124 ( .A(word1_reg_15_), .Y(_abc_19873_new_n1215_));
INVX1 INVX1_125 ( .A(word0_reg_15_), .Y(_abc_19873_new_n1216_));
INVX1 INVX1_126 ( .A(word2_reg_15_), .Y(_abc_19873_new_n1219_));
INVX1 INVX1_127 ( .A(core_key_47_), .Y(_abc_19873_new_n1221_));
INVX1 INVX1_128 ( .A(core_key_15_), .Y(_abc_19873_new_n1222_));
INVX1 INVX1_129 ( .A(core_mi_47_), .Y(_abc_19873_new_n1224_));
INVX1 INVX1_13 ( .A(word1_reg_0_), .Y(_abc_19873_new_n922_));
INVX1 INVX1_130 ( .A(core_mi_15_), .Y(_abc_19873_new_n1225_));
INVX1 INVX1_131 ( .A(core_mi_16_), .Y(_abc_19873_new_n1229_));
INVX1 INVX1_132 ( .A(core_key_112_), .Y(_abc_19873_new_n1230_));
INVX1 INVX1_133 ( .A(core_key_80_), .Y(_abc_19873_new_n1232_));
INVX1 INVX1_134 ( .A(word0_reg_16_), .Y(_abc_19873_new_n1235_));
INVX1 INVX1_135 ( .A(core_key_48_), .Y(_abc_19873_new_n1242_));
INVX1 INVX1_136 ( .A(core_key_16_), .Y(_abc_19873_new_n1243_));
INVX1 INVX1_137 ( .A(core_key_17_), .Y(_abc_19873_new_n1247_));
INVX1 INVX1_138 ( .A(word0_reg_17_), .Y(_abc_19873_new_n1250_));
INVX1 INVX1_139 ( .A(core_mi_49_), .Y(_abc_19873_new_n1251_));
INVX1 INVX1_14 ( .A(we), .Y(_abc_19873_new_n927_));
INVX1 INVX1_140 ( .A(core_key_81_), .Y(_abc_19873_new_n1254_));
INVX1 INVX1_141 ( .A(core_key_49_), .Y(_abc_19873_new_n1255_));
INVX1 INVX1_142 ( .A(core_key_113_), .Y(_abc_19873_new_n1261_));
INVX1 INVX1_143 ( .A(core_mi_18_), .Y(_abc_19873_new_n1266_));
INVX1 INVX1_144 ( .A(core_key_114_), .Y(_abc_19873_new_n1267_));
INVX1 INVX1_145 ( .A(core_key_82_), .Y(_abc_19873_new_n1269_));
INVX1 INVX1_146 ( .A(core_key_18_), .Y(_abc_19873_new_n1276_));
INVX1 INVX1_147 ( .A(word0_reg_18_), .Y(_abc_19873_new_n1279_));
INVX1 INVX1_148 ( .A(core_mi_50_), .Y(_abc_19873_new_n1280_));
INVX1 INVX1_149 ( .A(core_mi_19_), .Y(_abc_19873_new_n1284_));
INVX1 INVX1_15 ( .A(core_compress), .Y(_abc_19873_new_n930_));
INVX1 INVX1_150 ( .A(core_key_115_), .Y(_abc_19873_new_n1285_));
INVX1 INVX1_151 ( .A(core_key_83_), .Y(_abc_19873_new_n1287_));
INVX1 INVX1_152 ( .A(word0_reg_19_), .Y(_abc_19873_new_n1290_));
INVX1 INVX1_153 ( .A(core_key_51_), .Y(_abc_19873_new_n1297_));
INVX1 INVX1_154 ( .A(core_key_19_), .Y(_abc_19873_new_n1298_));
INVX1 INVX1_155 ( .A(core_mi_20_), .Y(_abc_19873_new_n1302_));
INVX1 INVX1_156 ( .A(core_key_116_), .Y(_abc_19873_new_n1303_));
INVX1 INVX1_157 ( .A(core_key_84_), .Y(_abc_19873_new_n1305_));
INVX1 INVX1_158 ( .A(core_key_20_), .Y(_abc_19873_new_n1312_));
INVX1 INVX1_159 ( .A(word0_reg_20_), .Y(_abc_19873_new_n1315_));
INVX1 INVX1_16 ( .A(core_key_65_), .Y(_abc_19873_new_n933_));
INVX1 INVX1_160 ( .A(core_mi_52_), .Y(_abc_19873_new_n1316_));
INVX1 INVX1_161 ( .A(word2_reg_21_), .Y(_abc_19873_new_n1320_));
INVX1 INVX1_162 ( .A(core_key_53_), .Y(_abc_19873_new_n1322_));
INVX1 INVX1_163 ( .A(core_key_21_), .Y(_abc_19873_new_n1323_));
INVX1 INVX1_164 ( .A(core_key_117_), .Y(_abc_19873_new_n1325_));
INVX1 INVX1_165 ( .A(core_key_85_), .Y(_abc_19873_new_n1326_));
INVX1 INVX1_166 ( .A(core_mi_53_), .Y(_abc_19873_new_n1329_));
INVX1 INVX1_167 ( .A(core_mi_21_), .Y(_abc_19873_new_n1330_));
INVX1 INVX1_168 ( .A(core_mi_22_), .Y(_abc_19873_new_n1338_));
INVX1 INVX1_169 ( .A(core_key_118_), .Y(_abc_19873_new_n1339_));
INVX1 INVX1_17 ( .A(core_key_33_), .Y(_abc_19873_new_n934_));
INVX1 INVX1_170 ( .A(core_key_86_), .Y(_abc_19873_new_n1341_));
INVX1 INVX1_171 ( .A(word0_reg_22_), .Y(_abc_19873_new_n1344_));
INVX1 INVX1_172 ( .A(core_key_54_), .Y(_abc_19873_new_n1351_));
INVX1 INVX1_173 ( .A(core_key_22_), .Y(_abc_19873_new_n1352_));
INVX1 INVX1_174 ( .A(word2_reg_23_), .Y(_abc_19873_new_n1356_));
INVX1 INVX1_175 ( .A(core_key_119_), .Y(_abc_19873_new_n1358_));
INVX1 INVX1_176 ( .A(core_key_87_), .Y(_abc_19873_new_n1359_));
INVX1 INVX1_177 ( .A(word1_reg_23_), .Y(_abc_19873_new_n1361_));
INVX1 INVX1_178 ( .A(word0_reg_23_), .Y(_abc_19873_new_n1362_));
INVX1 INVX1_179 ( .A(word3_reg_23_), .Y(_abc_19873_new_n1365_));
INVX1 INVX1_18 ( .A(core_mi_1_), .Y(_abc_19873_new_n941_));
INVX1 INVX1_180 ( .A(core_key_55_), .Y(_abc_19873_new_n1367_));
INVX1 INVX1_181 ( .A(core_key_23_), .Y(_abc_19873_new_n1368_));
INVX1 INVX1_182 ( .A(core_mi_55_), .Y(_abc_19873_new_n1370_));
INVX1 INVX1_183 ( .A(core_mi_23_), .Y(_abc_19873_new_n1371_));
INVX1 INVX1_184 ( .A(core_mi_24_), .Y(_abc_19873_new_n1375_));
INVX1 INVX1_185 ( .A(core_key_120_), .Y(_abc_19873_new_n1376_));
INVX1 INVX1_186 ( .A(core_key_88_), .Y(_abc_19873_new_n1378_));
INVX1 INVX1_187 ( .A(word0_reg_24_), .Y(_abc_19873_new_n1381_));
INVX1 INVX1_188 ( .A(core_key_56_), .Y(_abc_19873_new_n1388_));
INVX1 INVX1_189 ( .A(core_key_24_), .Y(_abc_19873_new_n1389_));
INVX1 INVX1_19 ( .A(core_key_97_), .Y(_abc_19873_new_n942_));
INVX1 INVX1_190 ( .A(core_mi_25_), .Y(_abc_19873_new_n1393_));
INVX1 INVX1_191 ( .A(core_key_121_), .Y(_abc_19873_new_n1394_));
INVX1 INVX1_192 ( .A(core_key_89_), .Y(_abc_19873_new_n1396_));
INVX1 INVX1_193 ( .A(word0_reg_25_), .Y(_abc_19873_new_n1399_));
INVX1 INVX1_194 ( .A(core_key_57_), .Y(_abc_19873_new_n1406_));
INVX1 INVX1_195 ( .A(core_key_25_), .Y(_abc_19873_new_n1407_));
INVX1 INVX1_196 ( .A(word2_reg_26_), .Y(_abc_19873_new_n1411_));
INVX1 INVX1_197 ( .A(core_key_122_), .Y(_abc_19873_new_n1413_));
INVX1 INVX1_198 ( .A(core_key_90_), .Y(_abc_19873_new_n1414_));
INVX1 INVX1_199 ( .A(word1_reg_26_), .Y(_abc_19873_new_n1416_));
INVX1 INVX1_2 ( .A(\addr[2] ), .Y(_abc_19873_new_n872_));
INVX1 INVX1_20 ( .A(core_compression_rounds_1_), .Y(_abc_19873_new_n944_));
INVX1 INVX1_200 ( .A(word0_reg_26_), .Y(_abc_19873_new_n1417_));
INVX1 INVX1_201 ( .A(word3_reg_26_), .Y(_abc_19873_new_n1420_));
INVX1 INVX1_202 ( .A(core_key_58_), .Y(_abc_19873_new_n1422_));
INVX1 INVX1_203 ( .A(core_key_26_), .Y(_abc_19873_new_n1423_));
INVX1 INVX1_204 ( .A(core_mi_58_), .Y(_abc_19873_new_n1425_));
INVX1 INVX1_205 ( .A(core_mi_26_), .Y(_abc_19873_new_n1426_));
INVX1 INVX1_206 ( .A(word3_reg_27_), .Y(_abc_19873_new_n1430_));
INVX1 INVX1_207 ( .A(core_key_123_), .Y(_abc_19873_new_n1432_));
INVX1 INVX1_208 ( .A(core_key_91_), .Y(_abc_19873_new_n1433_));
INVX1 INVX1_209 ( .A(word1_reg_27_), .Y(_abc_19873_new_n1435_));
INVX1 INVX1_21 ( .A(word3_reg_1_), .Y(_abc_19873_new_n947_));
INVX1 INVX1_210 ( .A(word0_reg_27_), .Y(_abc_19873_new_n1436_));
INVX1 INVX1_211 ( .A(word2_reg_27_), .Y(_abc_19873_new_n1439_));
INVX1 INVX1_212 ( .A(core_key_59_), .Y(_abc_19873_new_n1441_));
INVX1 INVX1_213 ( .A(core_key_27_), .Y(_abc_19873_new_n1442_));
INVX1 INVX1_214 ( .A(core_mi_59_), .Y(_abc_19873_new_n1444_));
INVX1 INVX1_215 ( .A(core_mi_27_), .Y(_abc_19873_new_n1445_));
INVX1 INVX1_216 ( .A(core_mi_28_), .Y(_abc_19873_new_n1449_));
INVX1 INVX1_217 ( .A(core_key_124_), .Y(_abc_19873_new_n1450_));
INVX1 INVX1_218 ( .A(core_key_92_), .Y(_abc_19873_new_n1452_));
INVX1 INVX1_219 ( .A(word0_reg_28_), .Y(_abc_19873_new_n1455_));
INVX1 INVX1_22 ( .A(word1_reg_1_), .Y(_abc_19873_new_n948_));
INVX1 INVX1_220 ( .A(core_key_60_), .Y(_abc_19873_new_n1462_));
INVX1 INVX1_221 ( .A(core_key_28_), .Y(_abc_19873_new_n1463_));
INVX1 INVX1_222 ( .A(word1_reg_29_), .Y(_abc_19873_new_n1467_));
INVX1 INVX1_223 ( .A(word0_reg_29_), .Y(_abc_19873_new_n1468_));
INVX1 INVX1_224 ( .A(word3_reg_29_), .Y(_abc_19873_new_n1470_));
INVX1 INVX1_225 ( .A(word2_reg_29_), .Y(_abc_19873_new_n1471_));
INVX1 INVX1_226 ( .A(core_key_93_), .Y(_abc_19873_new_n1477_));
INVX1 INVX1_227 ( .A(core_key_61_), .Y(_abc_19873_new_n1478_));
INVX1 INVX1_228 ( .A(core_mi_30_), .Y(_abc_19873_new_n1487_));
INVX1 INVX1_229 ( .A(core_key_126_), .Y(_abc_19873_new_n1488_));
INVX1 INVX1_23 ( .A(word2_reg_2_), .Y(_abc_19873_new_n952_));
INVX1 INVX1_230 ( .A(core_key_94_), .Y(_abc_19873_new_n1490_));
INVX1 INVX1_231 ( .A(word0_reg_30_), .Y(_abc_19873_new_n1493_));
INVX1 INVX1_232 ( .A(core_key_62_), .Y(_abc_19873_new_n1500_));
INVX1 INVX1_233 ( .A(core_key_30_), .Y(_abc_19873_new_n1501_));
INVX1 INVX1_234 ( .A(word3_reg_31_), .Y(_abc_19873_new_n1505_));
INVX1 INVX1_235 ( .A(core_key_127_), .Y(_abc_19873_new_n1507_));
INVX1 INVX1_236 ( .A(core_key_95_), .Y(_abc_19873_new_n1508_));
INVX1 INVX1_237 ( .A(word1_reg_31_), .Y(_abc_19873_new_n1510_));
INVX1 INVX1_238 ( .A(word0_reg_31_), .Y(_abc_19873_new_n1511_));
INVX1 INVX1_239 ( .A(word2_reg_31_), .Y(_abc_19873_new_n1514_));
INVX1 INVX1_24 ( .A(core_key_98_), .Y(_abc_19873_new_n955_));
INVX1 INVX1_240 ( .A(core_key_63_), .Y(_abc_19873_new_n1516_));
INVX1 INVX1_241 ( .A(core_key_31_), .Y(_abc_19873_new_n1517_));
INVX1 INVX1_242 ( .A(core_mi_63_), .Y(_abc_19873_new_n1519_));
INVX1 INVX1_243 ( .A(core_mi_31_), .Y(_abc_19873_new_n1520_));
INVX1 INVX1_244 ( .A(word3_reg_2_), .Y(_abc_19873_new_n1529_));
INVX1 INVX1_245 ( .A(word3_reg_7_), .Y(_abc_19873_new_n1540_));
INVX1 INVX1_246 ( .A(word3_reg_11_), .Y(_abc_19873_new_n1549_));
INVX1 INVX1_247 ( .A(word3_reg_12_), .Y(_abc_19873_new_n1552_));
INVX1 INVX1_248 ( .A(word3_reg_13_), .Y(_abc_19873_new_n1555_));
INVX1 INVX1_249 ( .A(word3_reg_14_), .Y(_abc_19873_new_n1558_));
INVX1 INVX1_25 ( .A(core_key_66_), .Y(_abc_19873_new_n956_));
INVX1 INVX1_250 ( .A(word3_reg_16_), .Y(_abc_19873_new_n1563_));
INVX1 INVX1_251 ( .A(word3_reg_17_), .Y(_abc_19873_new_n1566_));
INVX1 INVX1_252 ( .A(word3_reg_18_), .Y(_abc_19873_new_n1569_));
INVX1 INVX1_253 ( .A(word3_reg_19_), .Y(_abc_19873_new_n1572_));
INVX1 INVX1_254 ( .A(word3_reg_20_), .Y(_abc_19873_new_n1575_));
INVX1 INVX1_255 ( .A(word3_reg_21_), .Y(_abc_19873_new_n1578_));
INVX1 INVX1_256 ( .A(word3_reg_22_), .Y(_abc_19873_new_n1581_));
INVX1 INVX1_257 ( .A(word3_reg_24_), .Y(_abc_19873_new_n1586_));
INVX1 INVX1_258 ( .A(word3_reg_25_), .Y(_abc_19873_new_n1589_));
INVX1 INVX1_259 ( .A(word3_reg_28_), .Y(_abc_19873_new_n1596_));
INVX1 INVX1_26 ( .A(core_key_34_), .Y(_abc_19873_new_n958_));
INVX1 INVX1_260 ( .A(word3_reg_30_), .Y(_abc_19873_new_n1601_));
INVX1 INVX1_261 ( .A(word2_reg_0_), .Y(_abc_19873_new_n1606_));
INVX1 INVX1_262 ( .A(word2_reg_1_), .Y(_abc_19873_new_n1609_));
INVX1 INVX1_263 ( .A(word2_reg_3_), .Y(_abc_19873_new_n1614_));
INVX1 INVX1_264 ( .A(word2_reg_4_), .Y(_abc_19873_new_n1617_));
INVX1 INVX1_265 ( .A(word2_reg_5_), .Y(_abc_19873_new_n1620_));
INVX1 INVX1_266 ( .A(word2_reg_6_), .Y(_abc_19873_new_n1623_));
INVX1 INVX1_267 ( .A(word2_reg_7_), .Y(_abc_19873_new_n1626_));
INVX1 INVX1_268 ( .A(word2_reg_11_), .Y(_abc_19873_new_n1635_));
INVX1 INVX1_269 ( .A(word2_reg_12_), .Y(_abc_19873_new_n1638_));
INVX1 INVX1_27 ( .A(core_key_2_), .Y(_abc_19873_new_n959_));
INVX1 INVX1_270 ( .A(word2_reg_14_), .Y(_abc_19873_new_n1643_));
INVX1 INVX1_271 ( .A(word2_reg_16_), .Y(_abc_19873_new_n1648_));
INVX1 INVX1_272 ( .A(word2_reg_17_), .Y(_abc_19873_new_n1651_));
INVX1 INVX1_273 ( .A(word2_reg_18_), .Y(_abc_19873_new_n1654_));
INVX1 INVX1_274 ( .A(word2_reg_19_), .Y(_abc_19873_new_n1657_));
INVX1 INVX1_275 ( .A(word2_reg_20_), .Y(_abc_19873_new_n1660_));
INVX1 INVX1_276 ( .A(word2_reg_22_), .Y(_abc_19873_new_n1665_));
INVX1 INVX1_277 ( .A(word2_reg_24_), .Y(_abc_19873_new_n1670_));
INVX1 INVX1_278 ( .A(word2_reg_25_), .Y(_abc_19873_new_n1673_));
INVX1 INVX1_279 ( .A(word2_reg_28_), .Y(_abc_19873_new_n1680_));
INVX1 INVX1_28 ( .A(core_mi_34_), .Y(_abc_19873_new_n967_));
INVX1 INVX1_280 ( .A(word2_reg_30_), .Y(_abc_19873_new_n1685_));
INVX1 INVX1_281 ( .A(word1_reg_2_), .Y(_abc_19873_new_n1694_));
INVX1 INVX1_282 ( .A(word1_reg_3_), .Y(_abc_19873_new_n1697_));
INVX1 INVX1_283 ( .A(word1_reg_4_), .Y(_abc_19873_new_n1700_));
INVX1 INVX1_284 ( .A(word1_reg_6_), .Y(_abc_19873_new_n1705_));
INVX1 INVX1_285 ( .A(word1_reg_7_), .Y(_abc_19873_new_n1708_));
INVX1 INVX1_286 ( .A(word1_reg_11_), .Y(_abc_19873_new_n1717_));
INVX1 INVX1_287 ( .A(word1_reg_12_), .Y(_abc_19873_new_n1720_));
INVX1 INVX1_288 ( .A(word1_reg_13_), .Y(_abc_19873_new_n1723_));
INVX1 INVX1_289 ( .A(word1_reg_14_), .Y(_abc_19873_new_n1726_));
INVX1 INVX1_29 ( .A(core_mi_2_), .Y(_abc_19873_new_n968_));
INVX1 INVX1_290 ( .A(word1_reg_16_), .Y(_abc_19873_new_n1731_));
INVX1 INVX1_291 ( .A(word1_reg_17_), .Y(_abc_19873_new_n1734_));
INVX1 INVX1_292 ( .A(word1_reg_18_), .Y(_abc_19873_new_n1737_));
INVX1 INVX1_293 ( .A(word1_reg_19_), .Y(_abc_19873_new_n1740_));
INVX1 INVX1_294 ( .A(word1_reg_20_), .Y(_abc_19873_new_n1743_));
INVX1 INVX1_295 ( .A(word1_reg_21_), .Y(_abc_19873_new_n1746_));
INVX1 INVX1_296 ( .A(word1_reg_22_), .Y(_abc_19873_new_n1749_));
INVX1 INVX1_297 ( .A(word1_reg_24_), .Y(_abc_19873_new_n1754_));
INVX1 INVX1_298 ( .A(word1_reg_25_), .Y(_abc_19873_new_n1757_));
INVX1 INVX1_299 ( .A(word1_reg_28_), .Y(_abc_19873_new_n1764_));
INVX1 INVX1_3 ( .A(\addr[1] ), .Y(_abc_19873_new_n879_));
INVX1 INVX1_30 ( .A(core_compression_rounds_2_), .Y(_abc_19873_new_n971_));
INVX1 INVX1_300 ( .A(word1_reg_30_), .Y(_abc_19873_new_n1769_));
INVX1 INVX1_301 ( .A(word0_reg_0_), .Y(_abc_19873_new_n1774_));
INVX1 INVX1_302 ( .A(word0_reg_1_), .Y(_abc_19873_new_n1777_));
INVX1 INVX1_303 ( .A(word0_reg_2_), .Y(_abc_19873_new_n1780_));
INVX1 INVX1_304 ( .A(word0_reg_3_), .Y(_abc_19873_new_n1783_));
INVX1 INVX1_305 ( .A(word0_reg_4_), .Y(_abc_19873_new_n1786_));
INVX1 INVX1_306 ( .A(word0_reg_5_), .Y(_abc_19873_new_n1789_));
INVX1 INVX1_307 ( .A(word0_reg_6_), .Y(_abc_19873_new_n1792_));
INVX1 INVX1_308 ( .A(word0_reg_13_), .Y(_abc_19873_new_n1807_));
INVX1 INVX1_309 ( .A(word0_reg_21_), .Y(_abc_19873_new_n1824_));
INVX1 INVX1_31 ( .A(word3_reg_3_), .Y(_abc_19873_new_n976_));
INVX1 INVX1_310 ( .A(core_mi_32_), .Y(_abc_19873_new_n1847_));
INVX1 INVX1_311 ( .A(core_mi_33_), .Y(_abc_19873_new_n1852_));
INVX1 INVX1_312 ( .A(core_mi_37_), .Y(_abc_19873_new_n1861_));
INVX1 INVX1_313 ( .A(core_mi_46_), .Y(_abc_19873_new_n1880_));
INVX1 INVX1_314 ( .A(core_mi_48_), .Y(_abc_19873_new_n1885_));
INVX1 INVX1_315 ( .A(core_mi_51_), .Y(_abc_19873_new_n1892_));
INVX1 INVX1_316 ( .A(core_mi_54_), .Y(_abc_19873_new_n1899_));
INVX1 INVX1_317 ( .A(core_mi_56_), .Y(_abc_19873_new_n1904_));
INVX1 INVX1_318 ( .A(core_mi_57_), .Y(_abc_19873_new_n1907_));
INVX1 INVX1_319 ( .A(core_mi_60_), .Y(_abc_19873_new_n1914_));
INVX1 INVX1_32 ( .A(core_mi_35_), .Y(_abc_19873_new_n978_));
INVX1 INVX1_320 ( .A(core_mi_61_), .Y(_abc_19873_new_n1917_));
INVX1 INVX1_321 ( .A(core_mi_62_), .Y(_abc_19873_new_n1920_));
INVX1 INVX1_322 ( .A(core_mi_17_), .Y(_abc_19873_new_n1960_));
INVX1 INVX1_323 ( .A(core_mi_29_), .Y(_abc_19873_new_n1985_));
INVX1 INVX1_324 ( .A(core_key_125_), .Y(_abc_19873_new_n2051_));
INVX1 INVX1_325 ( .A(core_key_70_), .Y(_abc_19873_new_n2071_));
INVX1 INVX1_326 ( .A(core_key_71_), .Y(_abc_19873_new_n2074_));
INVX1 INVX1_327 ( .A(core_key_35_), .Y(_abc_19873_new_n2132_));
INVX1 INVX1_328 ( .A(core_key_36_), .Y(_abc_19873_new_n2135_));
INVX1 INVX1_329 ( .A(core_key_37_), .Y(_abc_19873_new_n2138_));
INVX1 INVX1_33 ( .A(core_mi_3_), .Y(_abc_19873_new_n979_));
INVX1 INVX1_330 ( .A(core_key_43_), .Y(_abc_19873_new_n2151_));
INVX1 INVX1_331 ( .A(core_key_44_), .Y(_abc_19873_new_n2154_));
INVX1 INVX1_332 ( .A(core_key_50_), .Y(_abc_19873_new_n2167_));
INVX1 INVX1_333 ( .A(core_key_52_), .Y(_abc_19873_new_n2172_));
INVX1 INVX1_334 ( .A(core_key_0_), .Y(_abc_19873_new_n2197_));
INVX1 INVX1_335 ( .A(core_key_1_), .Y(_abc_19873_new_n2201_));
INVX1 INVX1_336 ( .A(core_key_29_), .Y(_abc_19873_new_n2258_));
INVX1 INVX1_337 ( .A(reset_n_bF_buf28), .Y(_abc_19873_new_n2269_));
INVX1 INVX1_338 ( .A(_abc_19873_new_n1848_), .Y(_abc_19873_new_n2284_));
INVX1 INVX1_339 ( .A(_abc_19873_new_n2285_), .Y(_abc_19873_new_n2286_));
INVX1 INVX1_34 ( .A(core_compression_rounds_3_), .Y(_abc_19873_new_n981_));
INVX1 INVX1_340 ( .A(core_long), .Y(_abc_19873_new_n2293_));
INVX1 INVX1_341 ( .A(core__abc_21302_new_n1130_), .Y(core__abc_21302_new_n1131_));
INVX1 INVX1_342 ( .A(core_compression_rounds_3_), .Y(core__abc_21302_new_n1135_));
INVX1 INVX1_343 ( .A(core_loop_ctr_reg_0_), .Y(core__abc_21302_new_n1137_));
INVX1 INVX1_344 ( .A(core_compression_rounds_0_), .Y(core__abc_21302_new_n1138_));
INVX1 INVX1_345 ( .A(core_siphash_ctrl_reg_2_), .Y(core__abc_21302_new_n1149_));
INVX1 INVX1_346 ( .A(core__abc_21302_new_n1152_), .Y(core__abc_21302_new_n1153_));
INVX1 INVX1_347 ( .A(core__abc_21302_new_n1156_), .Y(core__abc_21302_new_n1157_));
INVX1 INVX1_348 ( .A(core__abc_21302_new_n1158_), .Y(core__abc_21302_new_n1159_));
INVX1 INVX1_349 ( .A(core_final_rounds_2_), .Y(core__abc_21302_new_n1160_));
INVX1 INVX1_35 ( .A(core_key_3_), .Y(_abc_19873_new_n989_));
INVX1 INVX1_350 ( .A(core__abc_21302_new_n1164_), .Y(core__abc_21302_new_n1165_));
INVX1 INVX1_351 ( .A(core_final_rounds_0_), .Y(core__abc_21302_new_n1171_));
INVX1 INVX1_352 ( .A(core__abc_21302_new_n1176_), .Y(core__abc_21302_new_n1177_));
INVX1 INVX1_353 ( .A(core__abc_21302_new_n1179_), .Y(core__abc_21302_new_n1180_));
INVX1 INVX1_354 ( .A(core__abc_21302_new_n1182_), .Y(core__abc_21302_new_n1183_));
INVX1 INVX1_355 ( .A(core_siphash_ctrl_reg_0_), .Y(core__abc_21302_new_n1184_));
INVX1 INVX1_356 ( .A(core_siphash_ctrl_reg_4_), .Y(core__abc_21302_new_n1188_));
INVX1 INVX1_357 ( .A(core_siphash_ctrl_reg_5_), .Y(core__abc_21302_new_n1194_));
INVX1 INVX1_358 ( .A(core_siphash_ctrl_reg_3_), .Y(core__abc_21302_new_n1195_));
INVX1 INVX1_359 ( .A(core_compress), .Y(core__abc_21302_new_n1198_));
INVX1 INVX1_36 ( .A(core_key_99_), .Y(_abc_19873_new_n992_));
INVX1 INVX1_360 ( .A(core__abc_21302_new_n1199_), .Y(core__abc_21302_new_n1200_));
INVX1 INVX1_361 ( .A(core_siphash_ctrl_reg_6_), .Y(core__abc_21302_new_n1203_));
INVX1 INVX1_362 ( .A(core__abc_21302_new_n1209_), .Y(core__abc_21302_new_n1210_));
INVX1 INVX1_363 ( .A(core__abc_21302_new_n1213_), .Y(core__abc_21302_new_n1214_));
INVX1 INVX1_364 ( .A(core__abc_21302_new_n1216_), .Y(core__abc_21302_new_n1217_));
INVX1 INVX1_365 ( .A(core__abc_21302_new_n1221_), .Y(core__abc_21302_new_n1222_));
INVX1 INVX1_366 ( .A(core__abc_21302_new_n1224_), .Y(core__abc_21302_new_n1225_));
INVX1 INVX1_367 ( .A(core__abc_21302_new_n1228_), .Y(core__abc_21302_new_n1229_));
INVX1 INVX1_368 ( .A(core__abc_21302_new_n1247_), .Y(core__abc_21302_new_n1248_));
INVX1 INVX1_369 ( .A(core__abc_21302_new_n1257_), .Y(core__abc_21302_new_n1258_));
INVX1 INVX1_37 ( .A(core_key_67_), .Y(_abc_19873_new_n993_));
INVX1 INVX1_370 ( .A(core_v1_reg_5_), .Y(core__abc_21302_new_n1261_));
INVX1 INVX1_371 ( .A(core_v0_reg_5_), .Y(core__abc_21302_new_n1262_));
INVX1 INVX1_372 ( .A(core__abc_21302_new_n1269_), .Y(core__abc_21302_new_n1270_));
INVX1 INVX1_373 ( .A(core__abc_21302_new_n1279_), .Y(core__abc_21302_new_n1280_));
INVX1 INVX1_374 ( .A(core__abc_21302_new_n1289_), .Y(core__abc_21302_new_n1290_));
INVX1 INVX1_375 ( .A(core__abc_21302_new_n1297_), .Y(core__abc_21302_new_n1298_));
INVX1 INVX1_376 ( .A(core__abc_21302_new_n1305_), .Y(core__abc_21302_new_n1306_));
INVX1 INVX1_377 ( .A(core__abc_21302_new_n1308_), .Y(core__abc_21302_new_n1309_));
INVX1 INVX1_378 ( .A(core_v2_reg_10_), .Y(core__abc_21302_new_n1316_));
INVX1 INVX1_379 ( .A(core_v3_reg_10_), .Y(core__abc_21302_new_n1317_));
INVX1 INVX1_38 ( .A(word3_reg_4_), .Y(_abc_19873_new_n997_));
INVX1 INVX1_380 ( .A(core__abc_21302_new_n1320_), .Y(core__abc_21302_new_n1321_));
INVX1 INVX1_381 ( .A(core_v2_reg_11_), .Y(core__abc_21302_new_n1328_));
INVX1 INVX1_382 ( .A(core_v3_reg_11_), .Y(core__abc_21302_new_n1329_));
INVX1 INVX1_383 ( .A(core__abc_21302_new_n1332_), .Y(core__abc_21302_new_n1333_));
INVX1 INVX1_384 ( .A(core_v2_reg_12_), .Y(core__abc_21302_new_n1338_));
INVX1 INVX1_385 ( .A(core__abc_21302_new_n1342_), .Y(core__abc_21302_new_n1343_));
INVX1 INVX1_386 ( .A(core_v2_reg_13_), .Y(core__abc_21302_new_n1350_));
INVX1 INVX1_387 ( .A(core_v3_reg_13_), .Y(core__abc_21302_new_n1351_));
INVX1 INVX1_388 ( .A(core__abc_21302_new_n1354_), .Y(core__abc_21302_new_n1355_));
INVX1 INVX1_389 ( .A(core_v2_reg_14_), .Y(core__abc_21302_new_n1362_));
INVX1 INVX1_39 ( .A(core_mi_36_), .Y(_abc_19873_new_n999_));
INVX1 INVX1_390 ( .A(core_v3_reg_14_), .Y(core__abc_21302_new_n1363_));
INVX1 INVX1_391 ( .A(core__abc_21302_new_n1366_), .Y(core__abc_21302_new_n1367_));
INVX1 INVX1_392 ( .A(core_v2_reg_15_), .Y(core__abc_21302_new_n1373_));
INVX1 INVX1_393 ( .A(core_v3_reg_15_), .Y(core__abc_21302_new_n1374_));
INVX1 INVX1_394 ( .A(core__abc_21302_new_n1378_), .Y(core__abc_21302_new_n1379_));
INVX1 INVX1_395 ( .A(core__abc_21302_new_n1385_), .Y(core__abc_21302_new_n1386_));
INVX1 INVX1_396 ( .A(core__abc_21302_new_n1389_), .Y(core__abc_21302_new_n1390_));
INVX1 INVX1_397 ( .A(core_v2_reg_17_), .Y(core__abc_21302_new_n1397_));
INVX1 INVX1_398 ( .A(core_v3_reg_17_), .Y(core__abc_21302_new_n1398_));
INVX1 INVX1_399 ( .A(core__abc_21302_new_n1401_), .Y(core__abc_21302_new_n1402_));
INVX1 INVX1_4 ( .A(core_key_64_), .Y(_abc_19873_new_n884_));
INVX1 INVX1_40 ( .A(core_mi_4_), .Y(_abc_19873_new_n1000_));
INVX1 INVX1_400 ( .A(core_v2_reg_18_), .Y(core__abc_21302_new_n1409_));
INVX1 INVX1_401 ( .A(core_v3_reg_18_), .Y(core__abc_21302_new_n1410_));
INVX1 INVX1_402 ( .A(core__abc_21302_new_n1413_), .Y(core__abc_21302_new_n1414_));
INVX1 INVX1_403 ( .A(core_v2_reg_19_), .Y(core__abc_21302_new_n1421_));
INVX1 INVX1_404 ( .A(core_v3_reg_19_), .Y(core__abc_21302_new_n1422_));
INVX1 INVX1_405 ( .A(core__abc_21302_new_n1425_), .Y(core__abc_21302_new_n1426_));
INVX1 INVX1_406 ( .A(core_v2_reg_20_), .Y(core__abc_21302_new_n1433_));
INVX1 INVX1_407 ( .A(core_v3_reg_20_), .Y(core__abc_21302_new_n1434_));
INVX1 INVX1_408 ( .A(core__abc_21302_new_n1437_), .Y(core__abc_21302_new_n1438_));
INVX1 INVX1_409 ( .A(core_v2_reg_21_), .Y(core__abc_21302_new_n1445_));
INVX1 INVX1_41 ( .A(core_final_rounds_0_), .Y(_abc_19873_new_n1002_));
INVX1 INVX1_410 ( .A(core_v3_reg_21_), .Y(core__abc_21302_new_n1446_));
INVX1 INVX1_411 ( .A(core__abc_21302_new_n1449_), .Y(core__abc_21302_new_n1450_));
INVX1 INVX1_412 ( .A(core_v2_reg_22_), .Y(core__abc_21302_new_n1457_));
INVX1 INVX1_413 ( .A(core_v3_reg_22_), .Y(core__abc_21302_new_n1458_));
INVX1 INVX1_414 ( .A(core__abc_21302_new_n1461_), .Y(core__abc_21302_new_n1462_));
INVX1 INVX1_415 ( .A(core__abc_21302_new_n1469_), .Y(core__abc_21302_new_n1470_));
INVX1 INVX1_416 ( .A(core_v2_reg_24_), .Y(core__abc_21302_new_n1476_));
INVX1 INVX1_417 ( .A(core_v3_reg_24_), .Y(core__abc_21302_new_n1477_));
INVX1 INVX1_418 ( .A(core__abc_21302_new_n1481_), .Y(core__abc_21302_new_n1482_));
INVX1 INVX1_419 ( .A(core_v2_reg_25_), .Y(core__abc_21302_new_n1487_));
INVX1 INVX1_42 ( .A(core_key_4_), .Y(_abc_19873_new_n1010_));
INVX1 INVX1_420 ( .A(core_v3_reg_25_), .Y(core__abc_21302_new_n1488_));
INVX1 INVX1_421 ( .A(core__abc_21302_new_n1491_), .Y(core__abc_21302_new_n1492_));
INVX1 INVX1_422 ( .A(core_v2_reg_26_), .Y(core__abc_21302_new_n1499_));
INVX1 INVX1_423 ( .A(core_v3_reg_26_), .Y(core__abc_21302_new_n1500_));
INVX1 INVX1_424 ( .A(core__abc_21302_new_n1503_), .Y(core__abc_21302_new_n1504_));
INVX1 INVX1_425 ( .A(core_v2_reg_27_), .Y(core__abc_21302_new_n1511_));
INVX1 INVX1_426 ( .A(core_v3_reg_27_), .Y(core__abc_21302_new_n1512_));
INVX1 INVX1_427 ( .A(core__abc_21302_new_n1515_), .Y(core__abc_21302_new_n1516_));
INVX1 INVX1_428 ( .A(core_v2_reg_28_), .Y(core__abc_21302_new_n1523_));
INVX1 INVX1_429 ( .A(core_v3_reg_28_), .Y(core__abc_21302_new_n1524_));
INVX1 INVX1_43 ( .A(core_key_100_), .Y(_abc_19873_new_n1013_));
INVX1 INVX1_430 ( .A(core__abc_21302_new_n1527_), .Y(core__abc_21302_new_n1528_));
INVX1 INVX1_431 ( .A(core__abc_21302_new_n1532_), .Y(core__abc_21302_new_n1533_));
INVX1 INVX1_432 ( .A(core_v2_reg_29_), .Y(core__abc_21302_new_n1536_));
INVX1 INVX1_433 ( .A(core_v3_reg_29_), .Y(core__abc_21302_new_n1537_));
INVX1 INVX1_434 ( .A(core__abc_21302_new_n1540_), .Y(core__abc_21302_new_n1541_));
INVX1 INVX1_435 ( .A(core_v2_reg_30_), .Y(core__abc_21302_new_n1548_));
INVX1 INVX1_436 ( .A(core_v3_reg_30_), .Y(core__abc_21302_new_n1549_));
INVX1 INVX1_437 ( .A(core__abc_21302_new_n1552_), .Y(core__abc_21302_new_n1553_));
INVX1 INVX1_438 ( .A(core__abc_21302_new_n1560_), .Y(core__abc_21302_new_n1561_));
INVX1 INVX1_439 ( .A(core__abc_21302_new_n1565_), .Y(core__abc_21302_new_n1566_));
INVX1 INVX1_44 ( .A(core_key_68_), .Y(_abc_19873_new_n1014_));
INVX1 INVX1_440 ( .A(core__abc_21302_new_n1568_), .Y(core__abc_21302_new_n1569_));
INVX1 INVX1_441 ( .A(core__abc_21302_new_n1572_), .Y(core__abc_21302_new_n1573_));
INVX1 INVX1_442 ( .A(core_v1_reg_33_), .Y(core__abc_21302_new_n1576_));
INVX1 INVX1_443 ( .A(core_v0_reg_33_), .Y(core__abc_21302_new_n1577_));
INVX1 INVX1_444 ( .A(core__abc_21302_new_n1584_), .Y(core__abc_21302_new_n1585_));
INVX1 INVX1_445 ( .A(core_v1_reg_34_), .Y(core__abc_21302_new_n1588_));
INVX1 INVX1_446 ( .A(core_v0_reg_34_), .Y(core__abc_21302_new_n1589_));
INVX1 INVX1_447 ( .A(core_v2_reg_34_), .Y(core__abc_21302_new_n1593_));
INVX1 INVX1_448 ( .A(core_v3_reg_34_), .Y(core__abc_21302_new_n1594_));
INVX1 INVX1_449 ( .A(core__abc_21302_new_n1598_), .Y(core__abc_21302_new_n1599_));
INVX1 INVX1_45 ( .A(core_key_69_), .Y(_abc_19873_new_n1020_));
INVX1 INVX1_450 ( .A(core_v2_reg_35_), .Y(core__abc_21302_new_n1606_));
INVX1 INVX1_451 ( .A(core_v3_reg_35_), .Y(core__abc_21302_new_n1607_));
INVX1 INVX1_452 ( .A(core__abc_21302_new_n1610_), .Y(core__abc_21302_new_n1611_));
INVX1 INVX1_453 ( .A(core__abc_21302_new_n1618_), .Y(core__abc_21302_new_n1619_));
INVX1 INVX1_454 ( .A(core__abc_21302_new_n1621_), .Y(core__abc_21302_new_n1622_));
INVX1 INVX1_455 ( .A(core_v0_reg_37_), .Y(core__abc_21302_new_n1626_));
INVX1 INVX1_456 ( .A(core__abc_21302_new_n1630_), .Y(core__abc_21302_new_n1631_));
INVX1 INVX1_457 ( .A(core__abc_21302_new_n1634_), .Y(core__abc_21302_new_n1635_));
INVX1 INVX1_458 ( .A(core__abc_21302_new_n1640_), .Y(core__abc_21302_new_n1641_));
INVX1 INVX1_459 ( .A(core__abc_21302_new_n1643_), .Y(core__abc_21302_new_n1644_));
INVX1 INVX1_46 ( .A(core_final_rounds_1_), .Y(_abc_19873_new_n1021_));
INVX1 INVX1_460 ( .A(core__abc_21302_new_n1650_), .Y(core__abc_21302_new_n1651_));
INVX1 INVX1_461 ( .A(core__abc_21302_new_n1654_), .Y(core__abc_21302_new_n1655_));
INVX1 INVX1_462 ( .A(core__abc_21302_new_n1661_), .Y(core__abc_21302_new_n1662_));
INVX1 INVX1_463 ( .A(core__abc_21302_new_n1665_), .Y(core__abc_21302_new_n1666_));
INVX1 INVX1_464 ( .A(core__abc_21302_new_n1672_), .Y(core__abc_21302_new_n1673_));
INVX1 INVX1_465 ( .A(core__abc_21302_new_n1676_), .Y(core__abc_21302_new_n1677_));
INVX1 INVX1_466 ( .A(core__abc_21302_new_n1687_), .Y(core__abc_21302_new_n1688_));
INVX1 INVX1_467 ( .A(core__abc_21302_new_n1695_), .Y(core__abc_21302_new_n1696_));
INVX1 INVX1_468 ( .A(core__abc_21302_new_n1698_), .Y(core__abc_21302_new_n1699_));
INVX1 INVX1_469 ( .A(core__abc_21302_new_n1707_), .Y(core__abc_21302_new_n1708_));
INVX1 INVX1_47 ( .A(core_key_5_), .Y(_abc_19873_new_n1028_));
INVX1 INVX1_470 ( .A(core__abc_21302_new_n1710_), .Y(core__abc_21302_new_n1711_));
INVX1 INVX1_471 ( .A(core__abc_21302_new_n1718_), .Y(core__abc_21302_new_n1719_));
INVX1 INVX1_472 ( .A(core__abc_21302_new_n1721_), .Y(core__abc_21302_new_n1722_));
INVX1 INVX1_473 ( .A(core__abc_21302_new_n1726_), .Y(core__abc_21302_new_n1727_));
INVX1 INVX1_474 ( .A(core__abc_21302_new_n1730_), .Y(core__abc_21302_new_n1731_));
INVX1 INVX1_475 ( .A(core__abc_21302_new_n1733_), .Y(core__abc_21302_new_n1734_));
INVX1 INVX1_476 ( .A(core__abc_21302_new_n1741_), .Y(core__abc_21302_new_n1742_));
INVX1 INVX1_477 ( .A(core__abc_21302_new_n1744_), .Y(core__abc_21302_new_n1745_));
INVX1 INVX1_478 ( .A(core__abc_21302_new_n1749_), .Y(core__abc_21302_new_n1750_));
INVX1 INVX1_479 ( .A(core_v2_reg_48_), .Y(core__abc_21302_new_n1753_));
INVX1 INVX1_48 ( .A(core_mi_5_), .Y(_abc_19873_new_n1031_));
INVX1 INVX1_480 ( .A(core_v3_reg_48_), .Y(core__abc_21302_new_n1754_));
INVX1 INVX1_481 ( .A(core__abc_21302_new_n1757_), .Y(core__abc_21302_new_n1758_));
INVX1 INVX1_482 ( .A(core_v2_reg_49_), .Y(core__abc_21302_new_n1763_));
INVX1 INVX1_483 ( .A(core_v3_reg_49_), .Y(core__abc_21302_new_n1764_));
INVX1 INVX1_484 ( .A(core__abc_21302_new_n1775_), .Y(core__abc_21302_new_n1776_));
INVX1 INVX1_485 ( .A(core__abc_21302_new_n1778_), .Y(core__abc_21302_new_n1779_));
INVX1 INVX1_486 ( .A(core__abc_21302_new_n1783_), .Y(core__abc_21302_new_n1784_));
INVX1 INVX1_487 ( .A(core__abc_21302_new_n1789_), .Y(core__abc_21302_new_n1790_));
INVX1 INVX1_488 ( .A(core_v1_reg_52_), .Y(core__abc_21302_new_n1794_));
INVX1 INVX1_489 ( .A(core_v0_reg_52_), .Y(core__abc_21302_new_n1795_));
INVX1 INVX1_49 ( .A(core_key_101_), .Y(_abc_19873_new_n1032_));
INVX1 INVX1_490 ( .A(core_v2_reg_52_), .Y(core__abc_21302_new_n1799_));
INVX1 INVX1_491 ( .A(core_v3_reg_52_), .Y(core__abc_21302_new_n1800_));
INVX1 INVX1_492 ( .A(core__abc_21302_new_n1803_), .Y(core__abc_21302_new_n1804_));
INVX1 INVX1_493 ( .A(core_v0_reg_53_), .Y(core__abc_21302_new_n1808_));
INVX1 INVX1_494 ( .A(core__abc_21302_new_n1819_), .Y(core__abc_21302_new_n1820_));
INVX1 INVX1_495 ( .A(core_v2_reg_54_), .Y(core__abc_21302_new_n1823_));
INVX1 INVX1_496 ( .A(core_v3_reg_54_), .Y(core__abc_21302_new_n1824_));
INVX1 INVX1_497 ( .A(core__abc_21302_new_n1827_), .Y(core__abc_21302_new_n1828_));
INVX1 INVX1_498 ( .A(core__abc_21302_new_n1832_), .Y(core__abc_21302_new_n1833_));
INVX1 INVX1_499 ( .A(core_v2_reg_55_), .Y(core__abc_21302_new_n1836_));
INVX1 INVX1_5 ( .A(core_key_32_), .Y(_abc_19873_new_n885_));
INVX1 INVX1_50 ( .A(word3_reg_5_), .Y(_abc_19873_new_n1034_));
INVX1 INVX1_500 ( .A(core_v3_reg_55_), .Y(core__abc_21302_new_n1837_));
INVX1 INVX1_501 ( .A(core__abc_21302_new_n1840_), .Y(core__abc_21302_new_n1841_));
INVX1 INVX1_502 ( .A(core_v0_reg_56_), .Y(core__abc_21302_new_n1846_));
INVX1 INVX1_503 ( .A(core_v2_reg_56_), .Y(core__abc_21302_new_n1850_));
INVX1 INVX1_504 ( .A(core_v3_reg_56_), .Y(core__abc_21302_new_n1851_));
INVX1 INVX1_505 ( .A(core__abc_21302_new_n1854_), .Y(core__abc_21302_new_n1855_));
INVX1 INVX1_506 ( .A(core__abc_21302_new_n1859_), .Y(core__abc_21302_new_n1860_));
INVX1 INVX1_507 ( .A(core__abc_21302_new_n1863_), .Y(core__abc_21302_new_n1864_));
INVX1 INVX1_508 ( .A(core__abc_21302_new_n1866_), .Y(core__abc_21302_new_n1867_));
INVX1 INVX1_509 ( .A(core_v1_reg_58_), .Y(core__abc_21302_new_n1871_));
INVX1 INVX1_51 ( .A(word1_reg_5_), .Y(_abc_19873_new_n1035_));
INVX1 INVX1_510 ( .A(core_v0_reg_58_), .Y(core__abc_21302_new_n1872_));
INVX1 INVX1_511 ( .A(core_v2_reg_58_), .Y(core__abc_21302_new_n1876_));
INVX1 INVX1_512 ( .A(core_v3_reg_58_), .Y(core__abc_21302_new_n1877_));
INVX1 INVX1_513 ( .A(core__abc_21302_new_n1880_), .Y(core__abc_21302_new_n1881_));
INVX1 INVX1_514 ( .A(core__abc_21302_new_n1885_), .Y(core__abc_21302_new_n1886_));
INVX1 INVX1_515 ( .A(core__abc_21302_new_n1889_), .Y(core__abc_21302_new_n1890_));
INVX1 INVX1_516 ( .A(core__abc_21302_new_n1892_), .Y(core__abc_21302_new_n1893_));
INVX1 INVX1_517 ( .A(core_v1_reg_60_), .Y(core__abc_21302_new_n1897_));
INVX1 INVX1_518 ( .A(core_v0_reg_60_), .Y(core__abc_21302_new_n1898_));
INVX1 INVX1_519 ( .A(core_v2_reg_60_), .Y(core__abc_21302_new_n1902_));
INVX1 INVX1_52 ( .A(word3_reg_6_), .Y(_abc_19873_new_n1039_));
INVX1 INVX1_520 ( .A(core_v3_reg_60_), .Y(core__abc_21302_new_n1903_));
INVX1 INVX1_521 ( .A(core__abc_21302_new_n1906_), .Y(core__abc_21302_new_n1907_));
INVX1 INVX1_522 ( .A(core_v0_reg_61_), .Y(core__abc_21302_new_n1912_));
INVX1 INVX1_523 ( .A(core_v2_reg_61_), .Y(core__abc_21302_new_n1916_));
INVX1 INVX1_524 ( .A(core_v3_reg_61_), .Y(core__abc_21302_new_n1917_));
INVX1 INVX1_525 ( .A(core__abc_21302_new_n1920_), .Y(core__abc_21302_new_n1921_));
INVX1 INVX1_526 ( .A(core__abc_21302_new_n1925_), .Y(core__abc_21302_new_n1926_));
INVX1 INVX1_527 ( .A(core_v2_reg_62_), .Y(core__abc_21302_new_n1929_));
INVX1 INVX1_528 ( .A(core_v3_reg_62_), .Y(core__abc_21302_new_n1930_));
INVX1 INVX1_529 ( .A(core__abc_21302_new_n1933_), .Y(core__abc_21302_new_n1934_));
INVX1 INVX1_53 ( .A(core_mi_38_), .Y(_abc_19873_new_n1041_));
INVX1 INVX1_530 ( .A(core__abc_21302_new_n1939_), .Y(core__abc_21302_new_n1940_));
INVX1 INVX1_531 ( .A(core__abc_21302_new_n2138_), .Y(core__abc_21302_new_n2139_));
INVX1 INVX1_532 ( .A(core__abc_21302_new_n2142_), .Y(core__abc_21302_new_n2143_));
INVX1 INVX1_533 ( .A(core__abc_21302_new_n2145_), .Y(core__abc_21302_new_n2149_));
INVX1 INVX1_534 ( .A(core__abc_21302_new_n2150_), .Y(core__abc_21302_new_n2154_));
INVX1 INVX1_535 ( .A(core__abc_21302_new_n2158_), .Y(core__abc_21302_new_n2161_));
INVX1 INVX1_536 ( .A(core_mi_reg_0_), .Y(core__abc_21302_new_n2164_));
INVX1 INVX1_537 ( .A(core__abc_21302_new_n2165_), .Y(core__abc_21302_new_n2166_));
INVX1 INVX1_538 ( .A(core_mi_reg_1_), .Y(core__abc_21302_new_n2171_));
INVX1 INVX1_539 ( .A(core_mi_reg_2_), .Y(core__abc_21302_new_n2174_));
INVX1 INVX1_54 ( .A(core_mi_6_), .Y(_abc_19873_new_n1042_));
INVX1 INVX1_540 ( .A(core_mi_reg_3_), .Y(core__abc_21302_new_n2177_));
INVX1 INVX1_541 ( .A(core_mi_reg_4_), .Y(core__abc_21302_new_n2180_));
INVX1 INVX1_542 ( .A(core_mi_reg_5_), .Y(core__abc_21302_new_n2183_));
INVX1 INVX1_543 ( .A(core_mi_reg_6_), .Y(core__abc_21302_new_n2186_));
INVX1 INVX1_544 ( .A(core_mi_reg_7_), .Y(core__abc_21302_new_n2189_));
INVX1 INVX1_545 ( .A(core_mi_reg_8_), .Y(core__abc_21302_new_n2192_));
INVX1 INVX1_546 ( .A(core_mi_reg_9_), .Y(core__abc_21302_new_n2195_));
INVX1 INVX1_547 ( .A(core_mi_reg_10_), .Y(core__abc_21302_new_n2198_));
INVX1 INVX1_548 ( .A(core_mi_reg_11_), .Y(core__abc_21302_new_n2201_));
INVX1 INVX1_549 ( .A(core_mi_reg_12_), .Y(core__abc_21302_new_n2204_));
INVX1 INVX1_55 ( .A(core_key_6_), .Y(_abc_19873_new_n1044_));
INVX1 INVX1_550 ( .A(core_mi_reg_13_), .Y(core__abc_21302_new_n2207_));
INVX1 INVX1_551 ( .A(core_mi_reg_14_), .Y(core__abc_21302_new_n2210_));
INVX1 INVX1_552 ( .A(core_mi_reg_15_), .Y(core__abc_21302_new_n2213_));
INVX1 INVX1_553 ( .A(core_mi_reg_16_), .Y(core__abc_21302_new_n2216_));
INVX1 INVX1_554 ( .A(core_mi_reg_17_), .Y(core__abc_21302_new_n2219_));
INVX1 INVX1_555 ( .A(core_mi_reg_18_), .Y(core__abc_21302_new_n2222_));
INVX1 INVX1_556 ( .A(core_mi_reg_19_), .Y(core__abc_21302_new_n2225_));
INVX1 INVX1_557 ( .A(core_mi_reg_20_), .Y(core__abc_21302_new_n2228_));
INVX1 INVX1_558 ( .A(core_mi_reg_21_), .Y(core__abc_21302_new_n2231_));
INVX1 INVX1_559 ( .A(core_mi_reg_22_), .Y(core__abc_21302_new_n2234_));
INVX1 INVX1_56 ( .A(core_final_rounds_2_), .Y(_abc_19873_new_n1045_));
INVX1 INVX1_560 ( .A(core_mi_reg_23_), .Y(core__abc_21302_new_n2237_));
INVX1 INVX1_561 ( .A(core_mi_reg_24_), .Y(core__abc_21302_new_n2240_));
INVX1 INVX1_562 ( .A(core_mi_reg_25_), .Y(core__abc_21302_new_n2243_));
INVX1 INVX1_563 ( .A(core_mi_reg_26_), .Y(core__abc_21302_new_n2246_));
INVX1 INVX1_564 ( .A(core_mi_reg_27_), .Y(core__abc_21302_new_n2249_));
INVX1 INVX1_565 ( .A(core_mi_reg_28_), .Y(core__abc_21302_new_n2252_));
INVX1 INVX1_566 ( .A(core_mi_reg_29_), .Y(core__abc_21302_new_n2255_));
INVX1 INVX1_567 ( .A(core_mi_reg_30_), .Y(core__abc_21302_new_n2258_));
INVX1 INVX1_568 ( .A(core_mi_reg_31_), .Y(core__abc_21302_new_n2261_));
INVX1 INVX1_569 ( .A(core_mi_reg_32_), .Y(core__abc_21302_new_n2264_));
INVX1 INVX1_57 ( .A(core_key_102_), .Y(_abc_19873_new_n1052_));
INVX1 INVX1_570 ( .A(core_mi_reg_33_), .Y(core__abc_21302_new_n2267_));
INVX1 INVX1_571 ( .A(core_mi_reg_34_), .Y(core__abc_21302_new_n2270_));
INVX1 INVX1_572 ( .A(core_mi_reg_35_), .Y(core__abc_21302_new_n2273_));
INVX1 INVX1_573 ( .A(core_mi_reg_36_), .Y(core__abc_21302_new_n2276_));
INVX1 INVX1_574 ( .A(core_mi_reg_37_), .Y(core__abc_21302_new_n2279_));
INVX1 INVX1_575 ( .A(core_mi_reg_38_), .Y(core__abc_21302_new_n2282_));
INVX1 INVX1_576 ( .A(core_mi_reg_39_), .Y(core__abc_21302_new_n2285_));
INVX1 INVX1_577 ( .A(core_mi_reg_40_), .Y(core__abc_21302_new_n2288_));
INVX1 INVX1_578 ( .A(core_mi_reg_41_), .Y(core__abc_21302_new_n2291_));
INVX1 INVX1_579 ( .A(core_mi_reg_42_), .Y(core__abc_21302_new_n2294_));
INVX1 INVX1_58 ( .A(core_key_38_), .Y(_abc_19873_new_n1055_));
INVX1 INVX1_580 ( .A(core_mi_reg_43_), .Y(core__abc_21302_new_n2297_));
INVX1 INVX1_581 ( .A(core_mi_reg_44_), .Y(core__abc_21302_new_n2300_));
INVX1 INVX1_582 ( .A(core_mi_reg_45_), .Y(core__abc_21302_new_n2303_));
INVX1 INVX1_583 ( .A(core_mi_reg_46_), .Y(core__abc_21302_new_n2306_));
INVX1 INVX1_584 ( .A(core_mi_reg_47_), .Y(core__abc_21302_new_n2309_));
INVX1 INVX1_585 ( .A(core_mi_reg_48_), .Y(core__abc_21302_new_n2312_));
INVX1 INVX1_586 ( .A(core_mi_reg_49_), .Y(core__abc_21302_new_n2315_));
INVX1 INVX1_587 ( .A(core_mi_reg_50_), .Y(core__abc_21302_new_n2318_));
INVX1 INVX1_588 ( .A(core_mi_reg_51_), .Y(core__abc_21302_new_n2321_));
INVX1 INVX1_589 ( .A(core_mi_reg_52_), .Y(core__abc_21302_new_n2324_));
INVX1 INVX1_59 ( .A(core_key_7_), .Y(_abc_19873_new_n1059_));
INVX1 INVX1_590 ( .A(core_mi_reg_53_), .Y(core__abc_21302_new_n2327_));
INVX1 INVX1_591 ( .A(core_mi_reg_54_), .Y(core__abc_21302_new_n2330_));
INVX1 INVX1_592 ( .A(core_mi_reg_55_), .Y(core__abc_21302_new_n2333_));
INVX1 INVX1_593 ( .A(core_mi_reg_56_), .Y(core__abc_21302_new_n2336_));
INVX1 INVX1_594 ( .A(core_mi_reg_57_), .Y(core__abc_21302_new_n2339_));
INVX1 INVX1_595 ( .A(core_mi_reg_58_), .Y(core__abc_21302_new_n2342_));
INVX1 INVX1_596 ( .A(core_mi_reg_59_), .Y(core__abc_21302_new_n2345_));
INVX1 INVX1_597 ( .A(core_mi_reg_60_), .Y(core__abc_21302_new_n2348_));
INVX1 INVX1_598 ( .A(core_mi_reg_61_), .Y(core__abc_21302_new_n2351_));
INVX1 INVX1_599 ( .A(core_mi_reg_62_), .Y(core__abc_21302_new_n2354_));
INVX1 INVX1_6 ( .A(\addr[5] ), .Y(_abc_19873_new_n887_));
INVX1 INVX1_60 ( .A(core_key_39_), .Y(_abc_19873_new_n1060_));
INVX1 INVX1_600 ( .A(core_mi_reg_63_), .Y(core__abc_21302_new_n2357_));
INVX1 INVX1_601 ( .A(core_v3_reg_0_), .Y(core__abc_21302_new_n2360_));
INVX1 INVX1_602 ( .A(core__abc_21302_new_n1567_), .Y(core__abc_21302_new_n2371_));
INVX1 INVX1_603 ( .A(core__abc_21302_new_n2392_), .Y(core__abc_21302_new_n2393_));
INVX1 INVX1_604 ( .A(core__abc_21302_new_n2394_), .Y(core__abc_21302_new_n2395_));
INVX1 INVX1_605 ( .A(core_v1_reg_8_), .Y(core__abc_21302_new_n2405_));
INVX1 INVX1_606 ( .A(core_v0_reg_8_), .Y(core__abc_21302_new_n2406_));
INVX1 INVX1_607 ( .A(core__abc_21302_new_n1324_), .Y(core__abc_21302_new_n2410_));
INVX1 INVX1_608 ( .A(core_v1_reg_16_), .Y(core__abc_21302_new_n2436_));
INVX1 INVX1_609 ( .A(core_v0_reg_16_), .Y(core__abc_21302_new_n2437_));
INVX1 INVX1_61 ( .A(word0_reg_7_), .Y(_abc_19873_new_n1062_));
INVX1 INVX1_610 ( .A(core__abc_21302_new_n2443_), .Y(core__abc_21302_new_n2444_));
INVX1 INVX1_611 ( .A(core__abc_21302_new_n2448_), .Y(core__abc_21302_new_n2449_));
INVX1 INVX1_612 ( .A(core_v0_reg_24_), .Y(core__abc_21302_new_n2454_));
INVX1 INVX1_613 ( .A(core_v0_reg_2_), .Y(core__abc_21302_new_n2469_));
INVX1 INVX1_614 ( .A(core__abc_21302_new_n2377_), .Y(core__abc_21302_new_n2474_));
INVX1 INVX1_615 ( .A(core__abc_21302_new_n2409_), .Y(core__abc_21302_new_n2487_));
INVX1 INVX1_616 ( .A(core__abc_21302_new_n2418_), .Y(core__abc_21302_new_n2490_));
INVX1 INVX1_617 ( .A(core__abc_21302_new_n2451_), .Y(core__abc_21302_new_n2499_));
INVX1 INVX1_618 ( .A(core__abc_21302_new_n2464_), .Y(core__abc_21302_new_n2502_));
INVX1 INVX1_619 ( .A(core__abc_21302_new_n2507_), .Y(core__abc_21302_new_n2510_));
INVX1 INVX1_62 ( .A(core_mi_39_), .Y(_abc_19873_new_n1063_));
INVX1 INVX1_620 ( .A(core__abc_21302_new_n1697_), .Y(core__abc_21302_new_n2513_));
INVX1 INVX1_621 ( .A(core__abc_21302_new_n1245_), .Y(core__abc_21302_new_n2515_));
INVX1 INVX1_622 ( .A(core__abc_21302_new_n2537_), .Y(core__abc_21302_new_n2538_));
INVX1 INVX1_623 ( .A(core__abc_21302_new_n1468_), .Y(core__abc_21302_new_n2576_));
INVX1 INVX1_624 ( .A(core__abc_21302_new_n2578_), .Y(core__abc_21302_new_n2579_));
INVX1 INVX1_625 ( .A(core__abc_21302_new_n1456_), .Y(core__abc_21302_new_n2580_));
INVX1 INVX1_626 ( .A(core_v2_reg_23_), .Y(core__abc_21302_new_n2581_));
INVX1 INVX1_627 ( .A(core_v3_reg_23_), .Y(core__abc_21302_new_n2582_));
INVX1 INVX1_628 ( .A(core_v2_reg_31_), .Y(core__abc_21302_new_n2587_));
INVX1 INVX1_629 ( .A(core_v3_reg_31_), .Y(core__abc_21302_new_n2588_));
INVX1 INVX1_63 ( .A(core_final_rounds_3_), .Y(_abc_19873_new_n1071_));
INVX1 INVX1_630 ( .A(core__abc_21302_new_n1547_), .Y(core__abc_21302_new_n2589_));
INVX1 INVX1_631 ( .A(core__abc_21302_new_n1653_), .Y(core__abc_21302_new_n2615_));
INVX1 INVX1_632 ( .A(core__abc_21302_new_n2621_), .Y(core__abc_21302_new_n2622_));
INVX1 INVX1_633 ( .A(core__abc_21302_new_n2367_), .Y(core__abc_21302_new_n2637_));
INVX1 INVX1_634 ( .A(core__abc_21302_new_n1580_), .Y(core__abc_21302_new_n2647_));
INVX1 INVX1_635 ( .A(core__abc_21302_new_n2655_), .Y(core__abc_21302_new_n2656_));
INVX1 INVX1_636 ( .A(core__abc_21302_new_n2514_), .Y(core__abc_21302_new_n2659_));
INVX1 INVX1_637 ( .A(core__abc_21302_new_n1592_), .Y(core__abc_21302_new_n2682_));
INVX1 INVX1_638 ( .A(core__abc_21302_new_n2684_), .Y(core__abc_21302_new_n2685_));
INVX1 INVX1_639 ( .A(core__abc_21302_new_n2687_), .Y(core__abc_21302_new_n2688_));
INVX1 INVX1_64 ( .A(core_mi_7_), .Y(_abc_19873_new_n1074_));
INVX1 INVX1_640 ( .A(core__abc_21302_new_n2689_), .Y(core__abc_21302_new_n2695_));
INVX1 INVX1_641 ( .A(core__abc_21302_new_n2697_), .Y(core__abc_21302_new_n2698_));
INVX1 INVX1_642 ( .A(core_v2_reg_44_), .Y(core__abc_21302_new_n2702_));
INVX1 INVX1_643 ( .A(core_v3_reg_44_), .Y(core__abc_21302_new_n2703_));
INVX1 INVX1_644 ( .A(core__abc_21302_new_n2709_), .Y(core__abc_21302_new_n2710_));
INVX1 INVX1_645 ( .A(core_key_66_), .Y(core__abc_21302_new_n2714_));
INVX1 INVX1_646 ( .A(core__abc_21302_new_n2719_), .Y(core__abc_21302_new_n2720_));
INVX1 INVX1_647 ( .A(core__abc_21302_new_n2722_), .Y(core__abc_21302_new_n2723_));
INVX1 INVX1_648 ( .A(core__abc_21302_new_n1732_), .Y(core__abc_21302_new_n2725_));
INVX1 INVX1_649 ( .A(core__abc_21302_new_n2732_), .Y(core__abc_21302_new_n2733_));
INVX1 INVX1_65 ( .A(core_key_103_), .Y(_abc_19873_new_n1075_));
INVX1 INVX1_650 ( .A(core__abc_21302_new_n1591_), .Y(core__abc_21302_new_n2736_));
INVX1 INVX1_651 ( .A(core__abc_21302_new_n1604_), .Y(core__abc_21302_new_n2737_));
INVX1 INVX1_652 ( .A(core_v3_reg_51_), .Y(core__abc_21302_new_n2740_));
INVX1 INVX1_653 ( .A(core_v2_reg_2_), .Y(core__abc_21302_new_n2741_));
INVX1 INVX1_654 ( .A(core_v3_reg_2_), .Y(core__abc_21302_new_n2742_));
INVX1 INVX1_655 ( .A(core__abc_21302_new_n2745_), .Y(core__abc_21302_new_n2746_));
INVX1 INVX1_656 ( .A(core__abc_21302_new_n2748_), .Y(core__abc_21302_new_n2749_));
INVX1 INVX1_657 ( .A(core__abc_21302_new_n2751_), .Y(core__abc_21302_new_n2752_));
INVX1 INVX1_658 ( .A(core_key_67_), .Y(core__abc_21302_new_n2757_));
INVX1 INVX1_659 ( .A(core__abc_21302_new_n2519_), .Y(core__abc_21302_new_n2770_));
INVX1 INVX1_66 ( .A(word2_reg_8_), .Y(_abc_19873_new_n1079_));
INVX1 INVX1_660 ( .A(core__abc_21302_new_n2774_), .Y(core__abc_21302_new_n2775_));
INVX1 INVX1_661 ( .A(core__abc_21302_new_n1743_), .Y(core__abc_21302_new_n2783_));
INVX1 INVX1_662 ( .A(core__abc_21302_new_n2780_), .Y(core__abc_21302_new_n2798_));
INVX1 INVX1_663 ( .A(core__abc_21302_new_n1629_), .Y(core__abc_21302_new_n2800_));
INVX1 INVX1_664 ( .A(core_v3_reg_53_), .Y(core__abc_21302_new_n2804_));
INVX1 INVX1_665 ( .A(core__abc_21302_new_n2807_), .Y(core__abc_21302_new_n2810_));
INVX1 INVX1_666 ( .A(core__abc_21302_new_n1756_), .Y(core__abc_21302_new_n2827_));
INVX1 INVX1_667 ( .A(core__abc_21302_new_n2523_), .Y(core__abc_21302_new_n2846_));
INVX1 INVX1_668 ( .A(core__abc_21302_new_n2851_), .Y(core__abc_21302_new_n2854_));
INVX1 INVX1_669 ( .A(core__abc_21302_new_n2856_), .Y(core__abc_21302_new_n2857_));
INVX1 INVX1_67 ( .A(core_key_104_), .Y(_abc_19873_new_n1081_));
INVX1 INVX1_670 ( .A(core__abc_21302_new_n1755_), .Y(core__abc_21302_new_n2864_));
INVX1 INVX1_671 ( .A(core_v2_reg_6_), .Y(core__abc_21302_new_n2882_));
INVX1 INVX1_672 ( .A(core_v3_reg_6_), .Y(core__abc_21302_new_n2883_));
INVX1 INVX1_673 ( .A(core__abc_21302_new_n2886_), .Y(core__abc_21302_new_n2887_));
INVX1 INVX1_674 ( .A(core__abc_21302_new_n1649_), .Y(core__abc_21302_new_n2889_));
INVX1 INVX1_675 ( .A(core__abc_21302_new_n1766_), .Y(core__abc_21302_new_n2896_));
INVX1 INVX1_676 ( .A(core__abc_21302_new_n1660_), .Y(core__abc_21302_new_n2920_));
INVX1 INVX1_677 ( .A(core__abc_21302_new_n2922_), .Y(core__abc_21302_new_n2931_));
INVX1 INVX1_678 ( .A(core__abc_21302_new_n1296_), .Y(core__abc_21302_new_n2938_));
INVX1 INVX1_679 ( .A(core__abc_21302_new_n2940_), .Y(core__abc_21302_new_n2941_));
INVX1 INVX1_68 ( .A(core_key_72_), .Y(_abc_19873_new_n1082_));
INVX1 INVX1_680 ( .A(core__abc_21302_new_n1788_), .Y(core__abc_21302_new_n2948_));
INVX1 INVX1_681 ( .A(core__abc_21302_new_n2952_), .Y(core__abc_21302_new_n2953_));
INVX1 INVX1_682 ( .A(core__abc_21302_new_n1671_), .Y(core__abc_21302_new_n2966_));
INVX1 INVX1_683 ( .A(core__abc_21302_new_n2971_), .Y(core__abc_21302_new_n2974_));
INVX1 INVX1_684 ( .A(core__abc_21302_new_n2942_), .Y(core__abc_21302_new_n2977_));
INVX1 INVX1_685 ( .A(core_v3_reg_36_), .Y(core__abc_21302_new_n2980_));
INVX1 INVX1_686 ( .A(core__abc_21302_new_n2919_), .Y(core__abc_21302_new_n3001_));
INVX1 INVX1_687 ( .A(core__abc_21302_new_n2972_), .Y(core__abc_21302_new_n3003_));
INVX1 INVX1_688 ( .A(core__abc_21302_new_n1682_), .Y(core__abc_21302_new_n3006_));
INVX1 INVX1_689 ( .A(core__abc_21302_new_n3007_), .Y(core__abc_21302_new_n3008_));
INVX1 INVX1_69 ( .A(word1_reg_8_), .Y(_abc_19873_new_n1084_));
INVX1 INVX1_690 ( .A(core__abc_21302_new_n1669_), .Y(core__abc_21302_new_n3009_));
INVX1 INVX1_691 ( .A(core__abc_21302_new_n3010_), .Y(core__abc_21302_new_n3011_));
INVX1 INVX1_692 ( .A(core__abc_21302_new_n3019_), .Y(core__abc_21302_new_n3022_));
INVX1 INVX1_693 ( .A(core__abc_21302_new_n3029_), .Y(core__abc_21302_new_n3030_));
INVX1 INVX1_694 ( .A(core__abc_21302_new_n3033_), .Y(core__abc_21302_new_n3034_));
INVX1 INVX1_695 ( .A(core__abc_21302_new_n3021_), .Y(core__abc_21302_new_n3042_));
INVX1 INVX1_696 ( .A(core__abc_21302_new_n1693_), .Y(core__abc_21302_new_n3047_));
INVX1 INVX1_697 ( .A(core_v3_reg_38_), .Y(core__abc_21302_new_n3063_));
INVX1 INVX1_698 ( .A(core__abc_21302_new_n3073_), .Y(core__abc_21302_new_n3074_));
INVX1 INVX1_699 ( .A(core__abc_21302_new_n3086_), .Y(core__abc_21302_new_n3087_));
INVX1 INVX1_7 ( .A(\addr[0] ), .Y(_abc_19873_new_n891_));
INVX1 INVX1_70 ( .A(word0_reg_8_), .Y(_abc_19873_new_n1085_));
INVX1 INVX1_700 ( .A(core__abc_21302_new_n3088_), .Y(core__abc_21302_new_n3089_));
INVX1 INVX1_701 ( .A(core__abc_21302_new_n3093_), .Y(core__abc_21302_new_n3094_));
INVX1 INVX1_702 ( .A(core__abc_21302_new_n3095_), .Y(core__abc_21302_new_n3096_));
INVX1 INVX1_703 ( .A(core__abc_21302_new_n2541_), .Y(core__abc_21302_new_n3102_));
INVX1 INVX1_704 ( .A(core__abc_21302_new_n3104_), .Y(core__abc_21302_new_n3105_));
INVX1 INVX1_705 ( .A(core_v3_reg_39_), .Y(core__abc_21302_new_n3111_));
INVX1 INVX1_706 ( .A(core__abc_21302_new_n1825_), .Y(core__abc_21302_new_n3112_));
INVX1 INVX1_707 ( .A(core__abc_21302_new_n1839_), .Y(core__abc_21302_new_n3114_));
INVX1 INVX1_708 ( .A(core__abc_21302_new_n3118_), .Y(core__abc_21302_new_n3119_));
INVX1 INVX1_709 ( .A(core__abc_21302_new_n3120_), .Y(core__abc_21302_new_n3121_));
INVX1 INVX1_71 ( .A(word3_reg_8_), .Y(_abc_19873_new_n1088_));
INVX1 INVX1_710 ( .A(core__abc_21302_new_n1705_), .Y(core__abc_21302_new_n3130_));
INVX1 INVX1_711 ( .A(core__abc_21302_new_n1716_), .Y(core__abc_21302_new_n3134_));
INVX1 INVX1_712 ( .A(core__abc_21302_new_n1353_), .Y(core__abc_21302_new_n3137_));
INVX1 INVX1_713 ( .A(core__abc_21302_new_n3146_), .Y(core__abc_21302_new_n3147_));
INVX1 INVX1_714 ( .A(core__abc_21302_new_n1838_), .Y(core__abc_21302_new_n3156_));
INVX1 INVX1_715 ( .A(core__abc_21302_new_n3065_), .Y(core__abc_21302_new_n3159_));
INVX1 INVX1_716 ( .A(core__abc_21302_new_n1728_), .Y(core__abc_21302_new_n3177_));
INVX1 INVX1_717 ( .A(core__abc_21302_new_n3179_), .Y(core__abc_21302_new_n3180_));
INVX1 INVX1_718 ( .A(core__abc_21302_new_n3178_), .Y(core__abc_21302_new_n3183_));
INVX1 INVX1_719 ( .A(core__abc_21302_new_n1365_), .Y(core__abc_21302_new_n3186_));
INVX1 INVX1_72 ( .A(core_key_40_), .Y(_abc_19873_new_n1090_));
INVX1 INVX1_720 ( .A(core__abc_21302_new_n2543_), .Y(core__abc_21302_new_n3187_));
INVX1 INVX1_721 ( .A(core__abc_21302_new_n3203_), .Y(core__abc_21302_new_n3204_));
INVX1 INVX1_722 ( .A(core_v3_reg_41_), .Y(core__abc_21302_new_n3212_));
INVX1 INVX1_723 ( .A(core_v3_reg_63_), .Y(core__abc_21302_new_n3232_));
INVX1 INVX1_724 ( .A(core__abc_21302_new_n1739_), .Y(core__abc_21302_new_n3237_));
INVX1 INVX1_725 ( .A(core_v3_reg_42_), .Y(core__abc_21302_new_n3246_));
INVX1 INVX1_726 ( .A(core__abc_21302_new_n3255_), .Y(core__abc_21302_new_n3256_));
INVX1 INVX1_727 ( .A(core__abc_21302_new_n3277_), .Y(core__abc_21302_new_n3278_));
INVX1 INVX1_728 ( .A(core__abc_21302_new_n3283_), .Y(core__abc_21302_new_n3284_));
INVX1 INVX1_729 ( .A(core__abc_21302_new_n3288_), .Y(core__abc_21302_new_n3289_));
INVX1 INVX1_73 ( .A(core_key_8_), .Y(_abc_19873_new_n1091_));
INVX1 INVX1_730 ( .A(core__abc_21302_new_n3292_), .Y(core__abc_21302_new_n3293_));
INVX1 INVX1_731 ( .A(core__abc_21302_new_n3300_), .Y(core__abc_21302_new_n3301_));
INVX1 INVX1_732 ( .A(core__abc_21302_new_n3305_), .Y(core__abc_21302_new_n3306_));
INVX1 INVX1_733 ( .A(core__abc_21302_new_n3307_), .Y(core__abc_21302_new_n3308_));
INVX1 INVX1_734 ( .A(core_v3_reg_43_), .Y(core__abc_21302_new_n3311_));
INVX1 INVX1_735 ( .A(core__abc_21302_new_n1878_), .Y(core__abc_21302_new_n3312_));
INVX1 INVX1_736 ( .A(core__abc_21302_new_n1891_), .Y(core__abc_21302_new_n3313_));
INVX1 INVX1_737 ( .A(core__abc_21302_new_n3321_), .Y(core__abc_21302_new_n3322_));
INVX1 INVX1_738 ( .A(core__abc_21302_new_n3341_), .Y(core__abc_21302_new_n3343_));
INVX1 INVX1_739 ( .A(core__abc_21302_new_n3345_), .Y(core__abc_21302_new_n3346_));
INVX1 INVX1_74 ( .A(core_mi_40_), .Y(_abc_19873_new_n1093_));
INVX1 INVX1_740 ( .A(core__abc_21302_new_n3350_), .Y(core__abc_21302_new_n3351_));
INVX1 INVX1_741 ( .A(core__abc_21302_new_n1905_), .Y(core__abc_21302_new_n3357_));
INVX1 INVX1_742 ( .A(core__abc_21302_new_n3304_), .Y(core__abc_21302_new_n3370_));
INVX1 INVX1_743 ( .A(core__abc_21302_new_n3374_), .Y(core__abc_21302_new_n3375_));
INVX1 INVX1_744 ( .A(core__abc_21302_new_n1773_), .Y(core__abc_21302_new_n3377_));
INVX1 INVX1_745 ( .A(core__abc_21302_new_n3335_), .Y(core__abc_21302_new_n3378_));
INVX1 INVX1_746 ( .A(core_v1_reg_49_), .Y(core__abc_21302_new_n3379_));
INVX1 INVX1_747 ( .A(core_v0_reg_49_), .Y(core__abc_21302_new_n3380_));
INVX1 INVX1_748 ( .A(core__abc_21302_new_n2564_), .Y(core__abc_21302_new_n3385_));
INVX1 INVX1_749 ( .A(core__abc_21302_new_n3395_), .Y(core__abc_21302_new_n3396_));
INVX1 INVX1_75 ( .A(core_mi_8_), .Y(_abc_19873_new_n1094_));
INVX1 INVX1_750 ( .A(core__abc_21302_new_n1904_), .Y(core__abc_21302_new_n3398_));
INVX1 INVX1_751 ( .A(core__abc_21302_new_n1919_), .Y(core__abc_21302_new_n3399_));
INVX1 INVX1_752 ( .A(core_v3_reg_45_), .Y(core__abc_21302_new_n3403_));
INVX1 INVX1_753 ( .A(core__abc_21302_new_n3394_), .Y(core__abc_21302_new_n3415_));
INVX1 INVX1_754 ( .A(core__abc_21302_new_n1785_), .Y(core__abc_21302_new_n3418_));
INVX1 INVX1_755 ( .A(core_v3_reg_3_), .Y(core__abc_21302_new_n3424_));
INVX1 INVX1_756 ( .A(core__abc_21302_new_n3434_), .Y(core__abc_21302_new_n3435_));
INVX1 INVX1_757 ( .A(core__abc_21302_new_n1918_), .Y(core__abc_21302_new_n3439_));
INVX1 INVX1_758 ( .A(core__abc_21302_new_n3446_), .Y(core__abc_21302_new_n3447_));
INVX1 INVX1_759 ( .A(core_key_83_), .Y(core__abc_21302_new_n3452_));
INVX1 INVX1_76 ( .A(word3_reg_9_), .Y(_abc_19873_new_n1098_));
INVX1 INVX1_760 ( .A(core__abc_21302_new_n3389_), .Y(core__abc_21302_new_n3461_));
INVX1 INVX1_761 ( .A(core__abc_21302_new_n3466_), .Y(core__abc_21302_new_n3467_));
INVX1 INVX1_762 ( .A(core__abc_21302_new_n3473_), .Y(core__abc_21302_new_n3474_));
INVX1 INVX1_763 ( .A(core__abc_21302_new_n2573_), .Y(core__abc_21302_new_n3477_));
INVX1 INVX1_764 ( .A(core__abc_21302_new_n3485_), .Y(core__abc_21302_new_n3486_));
INVX1 INVX1_765 ( .A(core__abc_21302_new_n3487_), .Y(core__abc_21302_new_n3488_));
INVX1 INVX1_766 ( .A(core__abc_21302_new_n3472_), .Y(core__abc_21302_new_n3500_));
INVX1 INVX1_767 ( .A(core__abc_21302_new_n1796_), .Y(core__abc_21302_new_n3504_));
INVX1 INVX1_768 ( .A(core__abc_21302_new_n1448_), .Y(core__abc_21302_new_n3507_));
INVX1 INVX1_769 ( .A(core__abc_21302_new_n3508_), .Y(core__abc_21302_new_n3509_));
INVX1 INVX1_77 ( .A(core_key_105_), .Y(_abc_19873_new_n1100_));
INVX1 INVX1_770 ( .A(core_v3_reg_5_), .Y(core__abc_21302_new_n3513_));
INVX1 INVX1_771 ( .A(core__abc_21302_new_n3522_), .Y(core__abc_21302_new_n3523_));
INVX1 INVX1_772 ( .A(core__abc_21302_new_n3534_), .Y(core__abc_21302_new_n3535_));
INVX1 INVX1_773 ( .A(core__abc_21302_new_n1821_), .Y(core__abc_21302_new_n3537_));
INVX1 INVX1_774 ( .A(core__abc_21302_new_n1810_), .Y(core__abc_21302_new_n3538_));
INVX1 INVX1_775 ( .A(core__abc_21302_new_n3539_), .Y(core__abc_21302_new_n3540_));
INVX1 INVX1_776 ( .A(core__abc_21302_new_n3544_), .Y(core__abc_21302_new_n3545_));
INVX1 INVX1_777 ( .A(core__abc_21302_new_n2558_), .Y(core__abc_21302_new_n3548_));
INVX1 INVX1_778 ( .A(core__abc_21302_new_n2693_), .Y(core__abc_21302_new_n3573_));
INVX1 INVX1_779 ( .A(core__abc_21302_new_n3561_), .Y(core__abc_21302_new_n3574_));
INVX1 INVX1_78 ( .A(core_key_73_), .Y(_abc_19873_new_n1101_));
INVX1 INVX1_780 ( .A(core__abc_21302_new_n1834_), .Y(core__abc_21302_new_n3576_));
INVX1 INVX1_781 ( .A(core_v3_reg_7_), .Y(core__abc_21302_new_n3583_));
INVX1 INVX1_782 ( .A(core__abc_21302_new_n3587_), .Y(core__abc_21302_new_n3609_));
INVX1 INVX1_783 ( .A(core__abc_21302_new_n1848_), .Y(core__abc_21302_new_n3617_));
INVX1 INVX1_784 ( .A(core__abc_21302_new_n3619_), .Y(core__abc_21302_new_n3620_));
INVX1 INVX1_785 ( .A(core__abc_21302_new_n3621_), .Y(core__abc_21302_new_n3628_));
INVX1 INVX1_786 ( .A(core__abc_21302_new_n2566_), .Y(core__abc_21302_new_n3633_));
INVX1 INVX1_787 ( .A(core__abc_21302_new_n3639_), .Y(core__abc_21302_new_n3640_));
INVX1 INVX1_788 ( .A(core__abc_21302_new_n3644_), .Y(core__abc_21302_new_n3645_));
INVX1 INVX1_789 ( .A(core__abc_21302_new_n1847_), .Y(core__abc_21302_new_n3655_));
INVX1 INVX1_79 ( .A(word1_reg_9_), .Y(_abc_19873_new_n1103_));
INVX1 INVX1_790 ( .A(core__abc_21302_new_n3656_), .Y(core__abc_21302_new_n3657_));
INVX1 INVX1_791 ( .A(core__abc_21302_new_n1490_), .Y(core__abc_21302_new_n3661_));
INVX1 INVX1_792 ( .A(core__abc_21302_new_n1478_), .Y(core__abc_21302_new_n3662_));
INVX1 INVX1_793 ( .A(core__abc_21302_new_n3663_), .Y(core__abc_21302_new_n3664_));
INVX1 INVX1_794 ( .A(core_v3_reg_9_), .Y(core__abc_21302_new_n3669_));
INVX1 INVX1_795 ( .A(core__abc_21302_new_n3671_), .Y(core__abc_21302_new_n3672_));
INVX1 INVX1_796 ( .A(core_key_89_), .Y(core__abc_21302_new_n3682_));
INVX1 INVX1_797 ( .A(core_key_90_), .Y(core__abc_21302_new_n3687_));
INVX1 INVX1_798 ( .A(core__abc_21302_new_n3616_), .Y(core__abc_21302_new_n3689_));
INVX1 INVX1_799 ( .A(core__abc_21302_new_n3690_), .Y(core__abc_21302_new_n3691_));
INVX1 INVX1_8 ( .A(\addr[4] ), .Y(_abc_19873_new_n899_));
INVX1 INVX1_80 ( .A(word0_reg_9_), .Y(_abc_19873_new_n1104_));
INVX1 INVX1_800 ( .A(core__abc_21302_new_n1861_), .Y(core__abc_21302_new_n3694_));
INVX1 INVX1_801 ( .A(core__abc_21302_new_n3695_), .Y(core__abc_21302_new_n3696_));
INVX1 INVX1_802 ( .A(core__abc_21302_new_n3697_), .Y(core__abc_21302_new_n3698_));
INVX1 INVX1_803 ( .A(core__abc_21302_new_n3700_), .Y(core__abc_21302_new_n3701_));
INVX1 INVX1_804 ( .A(core__abc_21302_new_n2595_), .Y(core__abc_21302_new_n3703_));
INVX1 INVX1_805 ( .A(core__abc_21302_new_n3716_), .Y(core__abc_21302_new_n3727_));
INVX1 INVX1_806 ( .A(core__abc_21302_new_n1498_), .Y(core__abc_21302_new_n3736_));
INVX1 INVX1_807 ( .A(core__abc_21302_new_n3731_), .Y(core__abc_21302_new_n3744_));
INVX1 INVX1_808 ( .A(core__abc_21302_new_n3764_), .Y(core__abc_21302_new_n3765_));
INVX1 INVX1_809 ( .A(core__abc_21302_new_n1900_), .Y(core__abc_21302_new_n3768_));
INVX1 INVX1_81 ( .A(word2_reg_9_), .Y(_abc_19873_new_n1107_));
INVX1 INVX1_810 ( .A(core__abc_21302_new_n2555_), .Y(core__abc_21302_new_n3775_));
INVX1 INVX1_811 ( .A(core__abc_21302_new_n3770_), .Y(core__abc_21302_new_n3799_));
INVX1 INVX1_812 ( .A(core__abc_21302_new_n1914_), .Y(core__abc_21302_new_n3801_));
INVX1 INVX1_813 ( .A(core__abc_21302_new_n3802_), .Y(core__abc_21302_new_n3803_));
INVX1 INVX1_814 ( .A(core__abc_21302_new_n1539_), .Y(core__abc_21302_new_n3806_));
INVX1 INVX1_815 ( .A(core__abc_21302_new_n1526_), .Y(core__abc_21302_new_n3807_));
INVX1 INVX1_816 ( .A(core__abc_21302_new_n3818_), .Y(core__abc_21302_new_n3819_));
INVX1 INVX1_817 ( .A(core__abc_21302_new_n1927_), .Y(core__abc_21302_new_n3831_));
INVX1 INVX1_818 ( .A(core__abc_21302_new_n1551_), .Y(core__abc_21302_new_n3841_));
INVX1 INVX1_819 ( .A(core__abc_21302_new_n2550_), .Y(core__abc_21302_new_n3842_));
INVX1 INVX1_82 ( .A(core_key_41_), .Y(_abc_19873_new_n1109_));
INVX1 INVX1_820 ( .A(core__abc_21302_new_n3856_), .Y(core__abc_21302_new_n3857_));
INVX1 INVX1_821 ( .A(core__abc_21302_new_n1899_), .Y(core__abc_21302_new_n3858_));
INVX1 INVX1_822 ( .A(core__abc_21302_new_n3862_), .Y(core__abc_21302_new_n3863_));
INVX1 INVX1_823 ( .A(core__abc_21302_new_n3853_), .Y(core__abc_21302_new_n3877_));
INVX1 INVX1_824 ( .A(core__abc_21302_new_n1937_), .Y(core__abc_21302_new_n3879_));
INVX1 INVX1_825 ( .A(core__abc_21302_new_n1559_), .Y(core__abc_21302_new_n3883_));
INVX1 INVX1_826 ( .A(core__abc_21302_new_n1571_), .Y(core__abc_21302_new_n3923_));
INVX1 INVX1_827 ( .A(core_key_96_), .Y(core__abc_21302_new_n3937_));
INVX1 INVX1_828 ( .A(core__abc_21302_new_n3927_), .Y(core__abc_21302_new_n3943_));
INVX1 INVX1_829 ( .A(core__abc_21302_new_n3947_), .Y(core__abc_21302_new_n3948_));
INVX1 INVX1_83 ( .A(core_key_9_), .Y(_abc_19873_new_n1110_));
INVX1 INVX1_830 ( .A(core__abc_21302_new_n1583_), .Y(core__abc_21302_new_n3949_));
INVX1 INVX1_831 ( .A(core__abc_21302_new_n3959_), .Y(core__abc_21302_new_n3971_));
INVX1 INVX1_832 ( .A(core__abc_21302_new_n3978_), .Y(core__abc_21302_new_n3979_));
INVX1 INVX1_833 ( .A(core__abc_21302_new_n1597_), .Y(core__abc_21302_new_n3980_));
INVX1 INVX1_834 ( .A(core__abc_21302_new_n2606_), .Y(core__abc_21302_new_n3981_));
INVX1 INVX1_835 ( .A(core__abc_21302_new_n2611_), .Y(core__abc_21302_new_n3982_));
INVX1 INVX1_836 ( .A(core__abc_21302_new_n3984_), .Y(core__abc_21302_new_n3985_));
INVX1 INVX1_837 ( .A(core__abc_21302_new_n3986_), .Y(core__abc_21302_new_n3988_));
INVX1 INVX1_838 ( .A(core__abc_21302_new_n1609_), .Y(core__abc_21302_new_n4006_));
INVX1 INVX1_839 ( .A(core__abc_21302_new_n4005_), .Y(core__abc_21302_new_n4016_));
INVX1 INVX1_84 ( .A(core_mi_41_), .Y(_abc_19873_new_n1112_));
INVX1 INVX1_840 ( .A(core_key_99_), .Y(core__abc_21302_new_n4025_));
INVX1 INVX1_841 ( .A(core__abc_21302_new_n3990_), .Y(core__abc_21302_new_n4033_));
INVX1 INVX1_842 ( .A(core__abc_21302_new_n4037_), .Y(core__abc_21302_new_n4038_));
INVX1 INVX1_843 ( .A(core__abc_21302_new_n4043_), .Y(core__abc_21302_new_n4044_));
INVX1 INVX1_844 ( .A(core__abc_21302_new_n1620_), .Y(core__abc_21302_new_n4048_));
INVX1 INVX1_845 ( .A(core__abc_21302_new_n4054_), .Y(core__abc_21302_new_n4055_));
INVX1 INVX1_846 ( .A(core__abc_21302_new_n4064_), .Y(core__abc_21302_new_n4065_));
INVX1 INVX1_847 ( .A(core__abc_21302_new_n1633_), .Y(core__abc_21302_new_n4066_));
INVX1 INVX1_848 ( .A(core__abc_21302_new_n4067_), .Y(core__abc_21302_new_n4069_));
INVX1 INVX1_849 ( .A(core__abc_21302_new_n4075_), .Y(core__abc_21302_new_n4076_));
INVX1 INVX1_85 ( .A(core_mi_9_), .Y(_abc_19873_new_n1113_));
INVX1 INVX1_850 ( .A(core__abc_21302_new_n4092_), .Y(core__abc_21302_new_n4093_));
INVX1 INVX1_851 ( .A(core__abc_21302_new_n4077_), .Y(core__abc_21302_new_n4094_));
INVX1 INVX1_852 ( .A(core__abc_21302_new_n4099_), .Y(core__abc_21302_new_n4108_));
INVX1 INVX1_853 ( .A(core__abc_21302_new_n4112_), .Y(core__abc_21302_new_n4113_));
INVX1 INVX1_854 ( .A(core__abc_21302_new_n4095_), .Y(core__abc_21302_new_n4115_));
INVX1 INVX1_855 ( .A(core__abc_21302_new_n4141_), .Y(core__abc_21302_new_n4142_));
INVX1 INVX1_856 ( .A(core__abc_21302_new_n4140_), .Y(core__abc_21302_new_n4144_));
INVX1 INVX1_857 ( .A(core__abc_21302_new_n4179_), .Y(core__abc_21302_new_n4182_));
INVX1 INVX1_858 ( .A(core__abc_21302_new_n4194_), .Y(core__abc_21302_new_n4195_));
INVX1 INVX1_859 ( .A(core__abc_21302_new_n1664_), .Y(core__abc_21302_new_n4196_));
INVX1 INVX1_86 ( .A(word2_reg_10_), .Y(_abc_19873_new_n1117_));
INVX1 INVX1_860 ( .A(core__abc_21302_new_n1675_), .Y(core__abc_21302_new_n4200_));
INVX1 INVX1_861 ( .A(core__abc_21302_new_n4199_), .Y(core__abc_21302_new_n4204_));
INVX1 INVX1_862 ( .A(core__abc_21302_new_n4202_), .Y(core__abc_21302_new_n4205_));
INVX1 INVX1_863 ( .A(core_key_105_), .Y(core__abc_21302_new_n4212_));
INVX1 INVX1_864 ( .A(core__abc_21302_new_n4219_), .Y(core__abc_21302_new_n4220_));
INVX1 INVX1_865 ( .A(core__abc_21302_new_n1686_), .Y(core__abc_21302_new_n4221_));
INVX1 INVX1_866 ( .A(core__abc_21302_new_n4237_), .Y(core__abc_21302_new_n4238_));
INVX1 INVX1_867 ( .A(core_v0_reg_10_), .Y(core__abc_21302_new_n4249_));
INVX1 INVX1_868 ( .A(core__abc_21302_new_n4259_), .Y(core__abc_21302_new_n4260_));
INVX1 INVX1_869 ( .A(core__abc_21302_new_n4227_), .Y(core__abc_21302_new_n4262_));
INVX1 INVX1_87 ( .A(core_key_106_), .Y(_abc_19873_new_n1119_));
INVX1 INVX1_870 ( .A(core_key_107_), .Y(core__abc_21302_new_n4268_));
INVX1 INVX1_871 ( .A(core__abc_21302_new_n4161_), .Y(core__abc_21302_new_n4278_));
INVX1 INVX1_872 ( .A(core__abc_21302_new_n4171_), .Y(core__abc_21302_new_n4279_));
INVX1 INVX1_873 ( .A(core__abc_21302_new_n4285_), .Y(core__abc_21302_new_n4286_));
INVX1 INVX1_874 ( .A(core__abc_21302_new_n4289_), .Y(core__abc_21302_new_n4290_));
INVX1 INVX1_875 ( .A(core_key_108_), .Y(core__abc_21302_new_n4294_));
INVX1 INVX1_876 ( .A(core__abc_21302_new_n4305_), .Y(core__abc_21302_new_n4307_));
INVX1 INVX1_877 ( .A(core__abc_21302_new_n4309_), .Y(core__abc_21302_new_n4313_));
INVX1 INVX1_878 ( .A(core__abc_21302_new_n4323_), .Y(core__abc_21302_new_n4324_));
INVX1 INVX1_879 ( .A(core__abc_21302_new_n4326_), .Y(core__abc_21302_new_n4327_));
INVX1 INVX1_88 ( .A(core_key_74_), .Y(_abc_19873_new_n1120_));
INVX1 INVX1_880 ( .A(core__abc_21302_new_n4328_), .Y(core__abc_21302_new_n4329_));
INVX1 INVX1_881 ( .A(core__abc_21302_new_n4337_), .Y(core__abc_21302_new_n4339_));
INVX1 INVX1_882 ( .A(core__abc_21302_new_n4277_), .Y(core__abc_21302_new_n4345_));
INVX1 INVX1_883 ( .A(core__abc_21302_new_n4281_), .Y(core__abc_21302_new_n4346_));
INVX1 INVX1_884 ( .A(core_v1_reg_14_), .Y(core__abc_21302_new_n4360_));
INVX1 INVX1_885 ( .A(core_v0_reg_14_), .Y(core__abc_21302_new_n4361_));
INVX1 INVX1_886 ( .A(core__abc_21302_new_n4340_), .Y(core__abc_21302_new_n4369_));
INVX1 INVX1_887 ( .A(core__abc_21302_new_n4367_), .Y(core__abc_21302_new_n4372_));
INVX1 INVX1_888 ( .A(core__abc_21302_new_n1384_), .Y(core__abc_21302_new_n4397_));
INVX1 INVX1_889 ( .A(core__abc_21302_new_n4399_), .Y(core__abc_21302_new_n4400_));
INVX1 INVX1_89 ( .A(word1_reg_10_), .Y(_abc_19873_new_n1122_));
INVX1 INVX1_890 ( .A(core__abc_21302_new_n4402_), .Y(core__abc_21302_new_n4403_));
INVX1 INVX1_891 ( .A(core__abc_21302_new_n1383_), .Y(core__abc_21302_new_n4411_));
INVX1 INVX1_892 ( .A(core__abc_21302_new_n4414_), .Y(core__abc_21302_new_n4415_));
INVX1 INVX1_893 ( .A(core__abc_21302_new_n4417_), .Y(core__abc_21302_new_n4418_));
INVX1 INVX1_894 ( .A(core__abc_21302_new_n4419_), .Y(core__abc_21302_new_n4425_));
INVX1 INVX1_895 ( .A(core_key_113_), .Y(core__abc_21302_new_n4437_));
INVX1 INVX1_896 ( .A(core__abc_21302_new_n2440_), .Y(core__abc_21302_new_n4444_));
INVX1 INVX1_897 ( .A(core__abc_21302_new_n4450_), .Y(core__abc_21302_new_n4451_));
INVX1 INVX1_898 ( .A(core__abc_21302_new_n4453_), .Y(core__abc_21302_new_n4454_));
INVX1 INVX1_899 ( .A(core__abc_21302_new_n4455_), .Y(core__abc_21302_new_n4456_));
INVX1 INVX1_9 ( .A(core_mi_0_), .Y(_abc_19873_new_n909_));
INVX1 INVX1_90 ( .A(word0_reg_10_), .Y(_abc_19873_new_n1123_));
INVX1 INVX1_900 ( .A(core__abc_21302_new_n4431_), .Y(core__abc_21302_new_n4457_));
INVX1 INVX1_901 ( .A(core__abc_21302_new_n4443_), .Y(core__abc_21302_new_n4458_));
INVX1 INVX1_902 ( .A(core__abc_21302_new_n4470_), .Y(core__abc_21302_new_n4471_));
INVX1 INVX1_903 ( .A(core__abc_21302_new_n4475_), .Y(core__abc_21302_new_n4476_));
INVX1 INVX1_904 ( .A(core__abc_21302_new_n4478_), .Y(core__abc_21302_new_n4480_));
INVX1 INVX1_905 ( .A(core_key_115_), .Y(core__abc_21302_new_n4486_));
INVX1 INVX1_906 ( .A(core__abc_21302_new_n4495_), .Y(core__abc_21302_new_n4496_));
INVX1 INVX1_907 ( .A(core__abc_21302_new_n4430_), .Y(core__abc_21302_new_n4497_));
INVX1 INVX1_908 ( .A(core__abc_21302_new_n4507_), .Y(core__abc_21302_new_n4516_));
INVX1 INVX1_909 ( .A(core__abc_21302_new_n4521_), .Y(core__abc_21302_new_n4522_));
INVX1 INVX1_91 ( .A(word3_reg_10_), .Y(_abc_19873_new_n1126_));
INVX1 INVX1_910 ( .A(core__abc_21302_new_n3926_), .Y(core__abc_21302_new_n4530_));
INVX1 INVX1_911 ( .A(core__abc_21302_new_n4542_), .Y(core__abc_21302_new_n4543_));
INVX1 INVX1_912 ( .A(core__abc_21302_new_n4553_), .Y(core__abc_21302_new_n4554_));
INVX1 INVX1_913 ( .A(core__abc_21302_new_n4001_), .Y(core__abc_21302_new_n4564_));
INVX1 INVX1_914 ( .A(core__abc_21302_new_n4551_), .Y(core__abc_21302_new_n4566_));
INVX1 INVX1_915 ( .A(core__abc_21302_new_n3117_), .Y(core__abc_21302_new_n4568_));
INVX1 INVX1_916 ( .A(core__abc_21302_new_n1454_), .Y(core__abc_21302_new_n4569_));
INVX1 INVX1_917 ( .A(core__abc_21302_new_n1467_), .Y(core__abc_21302_new_n4571_));
INVX1 INVX1_918 ( .A(core__abc_21302_new_n4573_), .Y(core__abc_21302_new_n4575_));
INVX1 INVX1_919 ( .A(core__abc_21302_new_n4549_), .Y(core__abc_21302_new_n4579_));
INVX1 INVX1_92 ( .A(core_key_42_), .Y(_abc_19873_new_n1128_));
INVX1 INVX1_920 ( .A(core__abc_21302_new_n4577_), .Y(core__abc_21302_new_n4580_));
INVX1 INVX1_921 ( .A(core__abc_21302_new_n4052_), .Y(core__abc_21302_new_n4617_));
INVX1 INVX1_922 ( .A(core__abc_21302_new_n3167_), .Y(core__abc_21302_new_n4618_));
INVX1 INVX1_923 ( .A(core__abc_21302_new_n4624_), .Y(core__abc_21302_new_n4626_));
INVX1 INVX1_924 ( .A(core__abc_21302_new_n4630_), .Y(core__abc_21302_new_n4631_));
INVX1 INVX1_925 ( .A(core__abc_21302_new_n4629_), .Y(core__abc_21302_new_n4633_));
INVX1 INVX1_926 ( .A(core__abc_21302_new_n4647_), .Y(core__abc_21302_new_n4648_));
INVX1 INVX1_927 ( .A(core__abc_21302_new_n4651_), .Y(core__abc_21302_new_n4652_));
INVX1 INVX1_928 ( .A(core__abc_21302_new_n4657_), .Y(core__abc_21302_new_n4658_));
INVX1 INVX1_929 ( .A(core__abc_21302_new_n4659_), .Y(core__abc_21302_new_n4660_));
INVX1 INVX1_93 ( .A(core_key_10_), .Y(_abc_19873_new_n1129_));
INVX1 INVX1_930 ( .A(core__abc_21302_new_n4642_), .Y(core__abc_21302_new_n4664_));
INVX1 INVX1_931 ( .A(core__abc_21302_new_n4653_), .Y(core__abc_21302_new_n4684_));
INVX1 INVX1_932 ( .A(core__abc_21302_new_n4682_), .Y(core__abc_21302_new_n4685_));
INVX1 INVX1_933 ( .A(core_key_123_), .Y(core__abc_21302_new_n4692_));
INVX1 INVX1_934 ( .A(core__abc_21302_new_n2459_), .Y(core__abc_21302_new_n4706_));
INVX1 INVX1_935 ( .A(core__abc_21302_new_n4709_), .Y(core__abc_21302_new_n4710_));
INVX1 INVX1_936 ( .A(core__abc_21302_new_n4712_), .Y(core__abc_21302_new_n4716_));
INVX1 INVX1_937 ( .A(core__abc_21302_new_n4720_), .Y(core__abc_21302_new_n4721_));
INVX1 INVX1_938 ( .A(core__abc_21302_new_n4176_), .Y(core__abc_21302_new_n4731_));
INVX1 INVX1_939 ( .A(core__abc_21302_new_n4596_), .Y(core__abc_21302_new_n4732_));
INVX1 INVX1_94 ( .A(core_mi_42_), .Y(_abc_19873_new_n1131_));
INVX1 INVX1_940 ( .A(core__abc_21302_new_n1534_), .Y(core__abc_21302_new_n4742_));
INVX1 INVX1_941 ( .A(core__abc_21302_new_n4745_), .Y(core__abc_21302_new_n4746_));
INVX1 INVX1_942 ( .A(core__abc_21302_new_n4713_), .Y(core__abc_21302_new_n4750_));
INVX1 INVX1_943 ( .A(core__abc_21302_new_n4748_), .Y(core__abc_21302_new_n4751_));
INVX1 INVX1_944 ( .A(core__abc_21302_new_n4232_), .Y(core__abc_21302_new_n4763_));
INVX1 INVX1_945 ( .A(core__abc_21302_new_n4766_), .Y(core__abc_21302_new_n4767_));
INVX1 INVX1_946 ( .A(core__abc_21302_new_n4769_), .Y(core__abc_21302_new_n4770_));
INVX1 INVX1_947 ( .A(core__abc_21302_new_n4772_), .Y(core__abc_21302_new_n4773_));
INVX1 INVX1_948 ( .A(core__abc_21302_new_n4774_), .Y(core__abc_21302_new_n4775_));
INVX1 INVX1_949 ( .A(core__abc_21302_new_n3448_), .Y(core__abc_21302_new_n4777_));
INVX1 INVX1_95 ( .A(core_mi_10_), .Y(_abc_19873_new_n1132_));
INVX1 INVX1_950 ( .A(core__abc_21302_new_n4779_), .Y(core__abc_21302_new_n4780_));
INVX1 INVX1_951 ( .A(core__abc_21302_new_n4796_), .Y(core__abc_21302_new_n4797_));
INVX1 INVX1_952 ( .A(core__abc_21302_new_n1545_), .Y(core__abc_21302_new_n4798_));
INVX1 INVX1_953 ( .A(core__abc_21302_new_n4795_), .Y(core__abc_21302_new_n4811_));
INVX1 INVX1_954 ( .A(core_key_127_), .Y(core__abc_21302_new_n4817_));
INVX1 INVX1_955 ( .A(core_v1_reg_18_), .Y(core__abc_21302_new_n4824_));
INVX1 INVX1_956 ( .A(core__abc_21302_new_n4825_), .Y(core__abc_21302_new_n4826_));
INVX1 INVX1_957 ( .A(core__abc_21302_new_n4823_), .Y(core__abc_21302_new_n4830_));
INVX1 INVX1_958 ( .A(core_v1_reg_17_), .Y(core__abc_21302_new_n4833_));
INVX1 INVX1_959 ( .A(core__abc_21302_new_n4840_), .Y(core__abc_21302_new_n4841_));
INVX1 INVX1_96 ( .A(core_mi_11_), .Y(_abc_19873_new_n1136_));
INVX1 INVX1_960 ( .A(core__abc_21302_new_n4839_), .Y(core__abc_21302_new_n4844_));
INVX1 INVX1_961 ( .A(core__abc_21302_new_n4842_), .Y(core__abc_21302_new_n4845_));
INVX1 INVX1_962 ( .A(core_v1_reg_15_), .Y(core__abc_21302_new_n4847_));
INVX1 INVX1_963 ( .A(core__abc_21302_new_n4854_), .Y(core__abc_21302_new_n4859_));
INVX1 INVX1_964 ( .A(core__abc_21302_new_n4862_), .Y(core__abc_21302_new_n4864_));
INVX1 INVX1_965 ( .A(core_v1_reg_12_), .Y(core__abc_21302_new_n4868_));
INVX1 INVX1_966 ( .A(core_v1_reg_11_), .Y(core__abc_21302_new_n4871_));
INVX1 INVX1_967 ( .A(core__abc_21302_new_n4843_), .Y(core__abc_21302_new_n4879_));
INVX1 INVX1_968 ( .A(core__abc_21302_new_n4880_), .Y(core__abc_21302_new_n4881_));
INVX1 INVX1_969 ( .A(core__abc_21302_new_n4883_), .Y(core__abc_21302_new_n4884_));
INVX1 INVX1_97 ( .A(core_key_107_), .Y(_abc_19873_new_n1137_));
INVX1 INVX1_970 ( .A(core__abc_21302_new_n4867_), .Y(core__abc_21302_new_n4889_));
INVX1 INVX1_971 ( .A(core__abc_21302_new_n4895_), .Y(core__abc_21302_new_n4901_));
INVX1 INVX1_972 ( .A(core_v1_reg_9_), .Y(core__abc_21302_new_n4906_));
INVX1 INVX1_973 ( .A(core__abc_21302_new_n4547_), .Y(core__abc_21302_new_n4908_));
INVX1 INVX1_974 ( .A(core__abc_21302_new_n4905_), .Y(core__abc_21302_new_n4911_));
INVX1 INVX1_975 ( .A(core__abc_21302_new_n4917_), .Y(core__abc_21302_new_n4918_));
INVX1 INVX1_976 ( .A(core__abc_21302_new_n3514_), .Y(core__abc_21302_new_n4921_));
INVX1 INVX1_977 ( .A(core__abc_21302_new_n4919_), .Y(core__abc_21302_new_n4922_));
INVX1 INVX1_978 ( .A(core_v1_reg_7_), .Y(core__abc_21302_new_n4924_));
INVX1 INVX1_979 ( .A(core_v1_reg_6_), .Y(core__abc_21302_new_n4933_));
INVX1 INVX1_98 ( .A(core_key_75_), .Y(_abc_19873_new_n1139_));
INVX1 INVX1_980 ( .A(core__abc_21302_new_n4934_), .Y(core__abc_21302_new_n4935_));
INVX1 INVX1_981 ( .A(core__abc_21302_new_n4932_), .Y(core__abc_21302_new_n4938_));
INVX1 INVX1_982 ( .A(core__abc_21302_new_n4936_), .Y(core__abc_21302_new_n4939_));
INVX1 INVX1_983 ( .A(core__abc_21302_new_n4930_), .Y(core__abc_21302_new_n4951_));
INVX1 INVX1_984 ( .A(core__abc_21302_new_n4900_), .Y(core__abc_21302_new_n4959_));
INVX1 INVX1_985 ( .A(core__abc_21302_new_n4910_), .Y(core__abc_21302_new_n4960_));
INVX1 INVX1_986 ( .A(core_v1_reg_1_), .Y(core__abc_21302_new_n4970_));
INVX1 INVX1_987 ( .A(core_v1_reg_63_), .Y(core__abc_21302_new_n4978_));
INVX1 INVX1_988 ( .A(core__abc_21302_new_n4979_), .Y(core__abc_21302_new_n4980_));
INVX1 INVX1_989 ( .A(core__abc_21302_new_n4967_), .Y(core__abc_21302_new_n4984_));
INVX1 INVX1_99 ( .A(core_key_11_), .Y(_abc_19873_new_n1147_));
INVX1 INVX1_990 ( .A(core__abc_21302_new_n3053_), .Y(core__abc_21302_new_n4995_));
INVX1 INVX1_991 ( .A(core_v1_reg_62_), .Y(core__abc_21302_new_n4996_));
INVX1 INVX1_992 ( .A(core__abc_21302_new_n5020_), .Y(core__abc_21302_new_n5021_));
INVX1 INVX1_993 ( .A(core__abc_21302_new_n2885_), .Y(core__abc_21302_new_n5022_));
INVX1 INVX1_994 ( .A(core_v1_reg_57_), .Y(core__abc_21302_new_n5024_));
INVX1 INVX1_995 ( .A(core__abc_21302_new_n5032_), .Y(core__abc_21302_new_n5033_));
INVX1 INVX1_996 ( .A(core_v1_reg_55_), .Y(core__abc_21302_new_n5034_));
INVX1 INVX1_997 ( .A(core__abc_21302_new_n5038_), .Y(core__abc_21302_new_n5039_));
INVX1 INVX1_998 ( .A(core__abc_21302_new_n1215_), .Y(core__abc_21302_new_n5046_));
INVX1 INVX1_999 ( .A(core__abc_21302_new_n5077_), .Y(core__abc_21302_new_n5078_));
INVX2 INVX2_1 ( .A(core_initalize), .Y(core__abc_21302_new_n1147_));
INVX2 INVX2_10 ( .A(core_v1_reg_61_), .Y(core__abc_21302_new_n1911_));
INVX2 INVX2_11 ( .A(core__abc_21302_new_n2369__bF_buf7), .Y(core__abc_21302_new_n2370_));
INVX2 INVX2_12 ( .A(core_v1_reg_24_), .Y(core__abc_21302_new_n2453_));
INVX2 INVX2_13 ( .A(core_v1_reg_2_), .Y(core__abc_21302_new_n2471_));
INVX2 INVX2_14 ( .A(core__abc_21302_new_n1460_), .Y(core__abc_21302_new_n2575_));
INVX2 INVX2_15 ( .A(core__abc_21302_new_n2624_), .Y(core__abc_21302_new_n2626_));
INVX2 INVX2_16 ( .A(core__abc_21302_new_n2652_), .Y(core__abc_21302_new_n2653_));
INVX2 INVX2_17 ( .A(core__abc_21302_new_n2724_), .Y(core__abc_21302_new_n2729_));
INVX2 INVX2_18 ( .A(core__abc_21302_new_n2867_), .Y(core__abc_21302_new_n2868_));
INVX2 INVX2_19 ( .A(core__abc_21302_new_n1777_), .Y(core__abc_21302_new_n2895_));
INVX2 INVX2_2 ( .A(core__abc_21302_new_n1154_), .Y(core__abc_21302_new_n1155_));
INVX2 INVX2_20 ( .A(core__abc_21302_new_n3067_), .Y(core__abc_21302_new_n3068_));
INVX2 INVX2_21 ( .A(core__abc_21302_new_n3192_), .Y(core__abc_21302_new_n3193_));
INVX2 INVX2_22 ( .A(core__abc_21302_new_n1873_), .Y(core__abc_21302_new_n3730_));
INVX2 INVX2_23 ( .A(core_v1_reg_10_), .Y(core__abc_21302_new_n4248_));
INVX2 INVX2_24 ( .A(core__abc_21302_new_n4341_), .Y(core__abc_21302_new_n4342_));
INVX2 INVX2_25 ( .A(core__abc_21302_new_n4545_), .Y(core__abc_21302_new_n4546_));
INVX2 INVX2_26 ( .A(core__abc_21302_new_n4678_), .Y(core__abc_21302_new_n4679_));
INVX2 INVX2_27 ( .A(core__abc_21302_new_n3387_), .Y(core__abc_21302_new_n4929_));
INVX2 INVX2_28 ( .A(core__abc_21302_new_n3340_), .Y(core__abc_21302_new_n4943_));
INVX2 INVX2_29 ( .A(core__abc_21302_new_n5669_), .Y(core__abc_21302_new_n5670_));
INVX2 INVX2_3 ( .A(core_v3_reg_12_), .Y(core__abc_21302_new_n1339_));
INVX2 INVX2_30 ( .A(core__abc_21302_new_n6009__bF_buf3), .Y(core__abc_21302_new_n6068_));
INVX2 INVX2_4 ( .A(core_v1_reg_37_), .Y(core__abc_21302_new_n1625_));
INVX2 INVX2_5 ( .A(core__abc_21302_new_n1683_), .Y(core__abc_21302_new_n1684_));
INVX2 INVX2_6 ( .A(core__abc_21302_new_n1703_), .Y(core__abc_21302_new_n1704_));
INVX2 INVX2_7 ( .A(core__abc_21302_new_n1771_), .Y(core__abc_21302_new_n1772_));
INVX2 INVX2_8 ( .A(core_v1_reg_53_), .Y(core__abc_21302_new_n1807_));
INVX2 INVX2_9 ( .A(core_v1_reg_56_), .Y(core__abc_21302_new_n1845_));
INVX4 INVX4_1 ( .A(_abc_19873_new_n2265_), .Y(_abc_19873_new_n2266_));
INVX8 INVX8_1 ( .A(core_siphash_valid_reg), .Y(_abc_19873_new_n1524_));
INVX8 INVX8_2 ( .A(reset_n_bF_buf20), .Y(core__abc_21302_new_n1185_));
INVX8 INVX8_3 ( .A(core__abc_21302_new_n2167_), .Y(core__abc_21302_new_n2168_));
INVX8 INVX8_4 ( .A(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n2363_));
INVX8 INVX8_5 ( .A(core__abc_21302_new_n2364__bF_buf5), .Y(core__abc_21302_new_n2365_));
INVX8 INVX8_6 ( .A(core__abc_21302_new_n2639__bF_buf6), .Y(core__abc_21302_new_n2640_));
INVX8 INVX8_7 ( .A(core__abc_21302_new_n2634__bF_buf7), .Y(core__abc_21302_new_n2673_));
INVX8 INVX8_8 ( .A(core__abc_21302_new_n5085__bF_buf3), .Y(core__abc_21302_new_n5104_));
INVX8 INVX8_9 ( .A(core__abc_21302_new_n5998__bF_buf3), .Y(core__abc_21302_new_n5999_));
MUX2X1 MUX2X1_1 ( .A(core__abc_21302_new_n1138_), .B(core__abc_21302_new_n1137_), .S(core__abc_21302_new_n1139_), .Y(core__abc_21302_new_n1140_));
MUX2X1 MUX2X1_2 ( .A(core__abc_21302_new_n1171_), .B(core__abc_21302_new_n1137_), .S(core__abc_21302_new_n1172_), .Y(core__abc_21302_new_n1173_));
NAND2X1 NAND2X1_1 ( .A(\addr[3] ), .B(_abc_19873_new_n872_), .Y(_abc_19873_new_n873_));
NAND2X1 NAND2X1_10 ( .A(_abc_19873_new_n912__bF_buf3), .B(_abc_19873_new_n889__bF_buf1), .Y(_abc_19873_new_n913_));
NAND2X1 NAND2X1_100 ( .A(core_v1_reg_29_), .B(core_v0_reg_29_), .Y(core__abc_21302_new_n1532_));
NAND2X1 NAND2X1_1000 ( .A(core__abc_21302_new_n6796_), .B(core__abc_21302_new_n6449__bF_buf5), .Y(core__abc_21302_new_n6797_));
NAND2X1 NAND2X1_1001 ( .A(core_v0_reg_49_), .B(core__abc_21302_new_n6450__bF_buf6), .Y(core__abc_21302_new_n6800_));
NAND2X1 NAND2X1_1002 ( .A(core__abc_21302_new_n6803_), .B(core__abc_21302_new_n6449__bF_buf4), .Y(core__abc_21302_new_n6804_));
NAND2X1 NAND2X1_1003 ( .A(core_v0_reg_50_), .B(core__abc_21302_new_n6450__bF_buf5), .Y(core__abc_21302_new_n6807_));
NAND2X1 NAND2X1_1004 ( .A(core__abc_21302_new_n6810_), .B(core__abc_21302_new_n6449__bF_buf3), .Y(core__abc_21302_new_n6811_));
NAND2X1 NAND2X1_1005 ( .A(core_v0_reg_51_), .B(core__abc_21302_new_n6450__bF_buf4), .Y(core__abc_21302_new_n6814_));
NAND2X1 NAND2X1_1006 ( .A(core__abc_21302_new_n6818_), .B(core__abc_21302_new_n6449__bF_buf2), .Y(core__abc_21302_new_n6819_));
NAND2X1 NAND2X1_1007 ( .A(core_v0_reg_52_), .B(core__abc_21302_new_n6450__bF_buf3), .Y(core__abc_21302_new_n6822_));
NAND2X1 NAND2X1_1008 ( .A(core__abc_21302_new_n6825_), .B(core__abc_21302_new_n6449__bF_buf1), .Y(core__abc_21302_new_n6826_));
NAND2X1 NAND2X1_1009 ( .A(core_v0_reg_53_), .B(core__abc_21302_new_n6450__bF_buf2), .Y(core__abc_21302_new_n6829_));
NAND2X1 NAND2X1_101 ( .A(core_v2_reg_29_), .B(core_v3_reg_29_), .Y(core__abc_21302_new_n1535_));
NAND2X1 NAND2X1_1010 ( .A(core__abc_21302_new_n6832_), .B(core__abc_21302_new_n6449__bF_buf0), .Y(core__abc_21302_new_n6833_));
NAND2X1 NAND2X1_1011 ( .A(core_v0_reg_54_), .B(core__abc_21302_new_n6450__bF_buf1), .Y(core__abc_21302_new_n6836_));
NAND2X1 NAND2X1_1012 ( .A(core__abc_21302_new_n6839_), .B(core__abc_21302_new_n6449__bF_buf7), .Y(core__abc_21302_new_n6840_));
NAND2X1 NAND2X1_1013 ( .A(core_v0_reg_55_), .B(core__abc_21302_new_n6450__bF_buf0), .Y(core__abc_21302_new_n6843_));
NAND2X1 NAND2X1_1014 ( .A(core__abc_21302_new_n6846_), .B(core__abc_21302_new_n6449__bF_buf6), .Y(core__abc_21302_new_n6847_));
NAND2X1 NAND2X1_1015 ( .A(core_v0_reg_56_), .B(core__abc_21302_new_n6450__bF_buf7), .Y(core__abc_21302_new_n6850_));
NAND2X1 NAND2X1_1016 ( .A(core__abc_21302_new_n4630_), .B(core__abc_21302_new_n4633_), .Y(core__abc_21302_new_n6852_));
NAND2X1 NAND2X1_1017 ( .A(core__abc_21302_new_n6854_), .B(core__abc_21302_new_n6449__bF_buf5), .Y(core__abc_21302_new_n6855_));
NAND2X1 NAND2X1_1018 ( .A(core_v0_reg_57_), .B(core__abc_21302_new_n6450__bF_buf6), .Y(core__abc_21302_new_n6858_));
NAND2X1 NAND2X1_1019 ( .A(core__abc_21302_new_n6862_), .B(core__abc_21302_new_n6449__bF_buf4), .Y(core__abc_21302_new_n6863_));
NAND2X1 NAND2X1_102 ( .A(core__abc_21302_new_n1536_), .B(core__abc_21302_new_n1537_), .Y(core__abc_21302_new_n1538_));
NAND2X1 NAND2X1_1020 ( .A(core_v0_reg_58_), .B(core__abc_21302_new_n6450__bF_buf5), .Y(core__abc_21302_new_n6866_));
NAND2X1 NAND2X1_1021 ( .A(core__abc_21302_new_n6870_), .B(core__abc_21302_new_n6449__bF_buf3), .Y(core__abc_21302_new_n6871_));
NAND2X1 NAND2X1_1022 ( .A(core_v0_reg_59_), .B(core__abc_21302_new_n6450__bF_buf4), .Y(core__abc_21302_new_n6874_));
NAND2X1 NAND2X1_1023 ( .A(core__abc_21302_new_n6877_), .B(core__abc_21302_new_n6449__bF_buf2), .Y(core__abc_21302_new_n6878_));
NAND2X1 NAND2X1_1024 ( .A(core_v0_reg_60_), .B(core__abc_21302_new_n6450__bF_buf3), .Y(core__abc_21302_new_n6881_));
NAND2X1 NAND2X1_1025 ( .A(core__abc_21302_new_n6884_), .B(core__abc_21302_new_n6449__bF_buf1), .Y(core__abc_21302_new_n6885_));
NAND2X1 NAND2X1_1026 ( .A(core_v0_reg_61_), .B(core__abc_21302_new_n6450__bF_buf2), .Y(core__abc_21302_new_n6888_));
NAND2X1 NAND2X1_1027 ( .A(core__abc_21302_new_n4785_), .B(core__abc_21302_new_n4781_), .Y(core__abc_21302_new_n6890_));
NAND2X1 NAND2X1_1028 ( .A(core__abc_21302_new_n6892_), .B(core__abc_21302_new_n6449__bF_buf0), .Y(core__abc_21302_new_n6893_));
NAND2X1 NAND2X1_1029 ( .A(core_v0_reg_62_), .B(core__abc_21302_new_n6450__bF_buf1), .Y(core__abc_21302_new_n6896_));
NAND2X1 NAND2X1_103 ( .A(core__abc_21302_new_n1535_), .B(core__abc_21302_new_n1538_), .Y(core__abc_21302_new_n1539_));
NAND2X1 NAND2X1_1030 ( .A(core__abc_21302_new_n6899_), .B(core__abc_21302_new_n6449__bF_buf7), .Y(core__abc_21302_new_n6900_));
NAND2X1 NAND2X1_1031 ( .A(core_v0_reg_63_), .B(core__abc_21302_new_n6450__bF_buf0), .Y(core__abc_21302_new_n6903_));
NAND2X1 NAND2X1_104 ( .A(core_v2_reg_30_), .B(core_v3_reg_30_), .Y(core__abc_21302_new_n1547_));
NAND2X1 NAND2X1_105 ( .A(core__abc_21302_new_n1548_), .B(core__abc_21302_new_n1549_), .Y(core__abc_21302_new_n1550_));
NAND2X1 NAND2X1_106 ( .A(core__abc_21302_new_n1547_), .B(core__abc_21302_new_n1550_), .Y(core__abc_21302_new_n1551_));
NAND2X1 NAND2X1_107 ( .A(core_v1_reg_32_), .B(core_v0_reg_32_), .Y(core__abc_21302_new_n1565_));
NAND2X1 NAND2X1_108 ( .A(core_v2_reg_32_), .B(core_v3_reg_32_), .Y(core__abc_21302_new_n1568_));
NAND2X1 NAND2X1_109 ( .A(core__abc_21302_new_n1576_), .B(core__abc_21302_new_n1577_), .Y(core__abc_21302_new_n1578_));
NAND2X1 NAND2X1_11 ( .A(_abc_19873_new_n889__bF_buf0), .B(_abc_19873_new_n874_), .Y(_abc_19873_new_n914_));
NAND2X1 NAND2X1_110 ( .A(core_v1_reg_33_), .B(core_v0_reg_33_), .Y(core__abc_21302_new_n1579_));
NAND2X1 NAND2X1_111 ( .A(core__abc_21302_new_n1579_), .B(core__abc_21302_new_n1578_), .Y(core__abc_21302_new_n1580_));
NAND2X1 NAND2X1_112 ( .A(core_v2_reg_33_), .B(core_v3_reg_33_), .Y(core__abc_21302_new_n1581_));
NAND2X1 NAND2X1_113 ( .A(core__abc_21302_new_n1581_), .B(core__abc_21302_new_n1582_), .Y(core__abc_21302_new_n1583_));
NAND2X1 NAND2X1_114 ( .A(core__abc_21302_new_n1588_), .B(core__abc_21302_new_n1589_), .Y(core__abc_21302_new_n1590_));
NAND2X1 NAND2X1_115 ( .A(core_v1_reg_34_), .B(core_v0_reg_34_), .Y(core__abc_21302_new_n1591_));
NAND2X1 NAND2X1_116 ( .A(core__abc_21302_new_n1591_), .B(core__abc_21302_new_n1590_), .Y(core__abc_21302_new_n1592_));
NAND2X1 NAND2X1_117 ( .A(core__abc_21302_new_n1593_), .B(core__abc_21302_new_n1594_), .Y(core__abc_21302_new_n1595_));
NAND2X1 NAND2X1_118 ( .A(core_v2_reg_34_), .B(core_v3_reg_34_), .Y(core__abc_21302_new_n1596_));
NAND2X1 NAND2X1_119 ( .A(core__abc_21302_new_n1596_), .B(core__abc_21302_new_n1595_), .Y(core__abc_21302_new_n1597_));
NAND2X1 NAND2X1_12 ( .A(_abc_19873_new_n877_), .B(_abc_19873_new_n917_), .Y(_abc_19873_new_n918_));
NAND2X1 NAND2X1_120 ( .A(core_v2_reg_35_), .B(core_v3_reg_35_), .Y(core__abc_21302_new_n1605_));
NAND2X1 NAND2X1_121 ( .A(core__abc_21302_new_n1606_), .B(core__abc_21302_new_n1607_), .Y(core__abc_21302_new_n1608_));
NAND2X1 NAND2X1_122 ( .A(core__abc_21302_new_n1605_), .B(core__abc_21302_new_n1608_), .Y(core__abc_21302_new_n1609_));
NAND2X1 NAND2X1_123 ( .A(core_v2_reg_36_), .B(core_v3_reg_36_), .Y(core__abc_21302_new_n1618_));
NAND2X1 NAND2X1_124 ( .A(core__abc_21302_new_n1625_), .B(core__abc_21302_new_n1626_), .Y(core__abc_21302_new_n1627_));
NAND2X1 NAND2X1_125 ( .A(core_v1_reg_37_), .B(core_v0_reg_37_), .Y(core__abc_21302_new_n1628_));
NAND2X1 NAND2X1_126 ( .A(core__abc_21302_new_n1628_), .B(core__abc_21302_new_n1627_), .Y(core__abc_21302_new_n1629_));
NAND2X1 NAND2X1_127 ( .A(core_v2_reg_37_), .B(core_v3_reg_37_), .Y(core__abc_21302_new_n1630_));
NAND2X1 NAND2X1_128 ( .A(core_v2_reg_38_), .B(core_v3_reg_38_), .Y(core__abc_21302_new_n1640_));
NAND2X1 NAND2X1_129 ( .A(core_v2_reg_39_), .B(core_v3_reg_39_), .Y(core__abc_21302_new_n1650_));
NAND2X1 NAND2X1_13 ( .A(_abc_19873_new_n895__bF_buf3), .B(_abc_19873_new_n901__bF_buf5), .Y(_abc_19873_new_n923_));
NAND2X1 NAND2X1_130 ( .A(core_v2_reg_40_), .B(core_v3_reg_40_), .Y(core__abc_21302_new_n1661_));
NAND2X1 NAND2X1_131 ( .A(core_v2_reg_41_), .B(core_v3_reg_41_), .Y(core__abc_21302_new_n1672_));
NAND2X1 NAND2X1_132 ( .A(core_v2_reg_42_), .B(core_v3_reg_42_), .Y(core__abc_21302_new_n1683_));
NAND2X1 NAND2X1_133 ( .A(core_v2_reg_43_), .B(core_v3_reg_43_), .Y(core__abc_21302_new_n1695_));
NAND2X1 NAND2X1_134 ( .A(core_v1_reg_44_), .B(core_v0_reg_44_), .Y(core__abc_21302_new_n1703_));
NAND2X1 NAND2X1_135 ( .A(core_v2_reg_44_), .B(core_v3_reg_44_), .Y(core__abc_21302_new_n1707_));
NAND2X1 NAND2X1_136 ( .A(core_v1_reg_45_), .B(core_v0_reg_45_), .Y(core__abc_21302_new_n1715_));
NAND2X1 NAND2X1_137 ( .A(core__abc_21302_new_n1715_), .B(core__abc_21302_new_n1714_), .Y(core__abc_21302_new_n1716_));
NAND2X1 NAND2X1_138 ( .A(core_v2_reg_45_), .B(core_v3_reg_45_), .Y(core__abc_21302_new_n1718_));
NAND2X1 NAND2X1_139 ( .A(core_v1_reg_46_), .B(core_v0_reg_46_), .Y(core__abc_21302_new_n1726_));
NAND2X1 NAND2X1_14 ( .A(_abc_19873_new_n912__bF_buf2), .B(_abc_19873_new_n901__bF_buf4), .Y(_abc_19873_new_n924_));
NAND2X1 NAND2X1_140 ( .A(core_v2_reg_46_), .B(core_v3_reg_46_), .Y(core__abc_21302_new_n1730_));
NAND2X1 NAND2X1_141 ( .A(core_v2_reg_47_), .B(core_v3_reg_47_), .Y(core__abc_21302_new_n1741_));
NAND2X1 NAND2X1_142 ( .A(core_v1_reg_48_), .B(core_v0_reg_48_), .Y(core__abc_21302_new_n1749_));
NAND2X1 NAND2X1_143 ( .A(core_v1_reg_50_), .B(core_v0_reg_50_), .Y(core__abc_21302_new_n1771_));
NAND2X1 NAND2X1_144 ( .A(core_v2_reg_50_), .B(core_v3_reg_50_), .Y(core__abc_21302_new_n1775_));
NAND2X1 NAND2X1_145 ( .A(core_v1_reg_51_), .B(core_v0_reg_51_), .Y(core__abc_21302_new_n1783_));
NAND2X1 NAND2X1_146 ( .A(core_v1_reg_54_), .B(core_v0_reg_54_), .Y(core__abc_21302_new_n1819_));
NAND2X1 NAND2X1_147 ( .A(core_v1_reg_55_), .B(core_v0_reg_55_), .Y(core__abc_21302_new_n1832_));
NAND2X1 NAND2X1_148 ( .A(core_v1_reg_57_), .B(core_v0_reg_57_), .Y(core__abc_21302_new_n1859_));
NAND2X1 NAND2X1_149 ( .A(core_v2_reg_57_), .B(core_v3_reg_57_), .Y(core__abc_21302_new_n1863_));
NAND2X1 NAND2X1_15 ( .A(cs), .B(_abc_19873_new_n927_), .Y(_abc_19873_new_n928_));
NAND2X1 NAND2X1_150 ( .A(core_v1_reg_59_), .B(core_v0_reg_59_), .Y(core__abc_21302_new_n1885_));
NAND2X1 NAND2X1_151 ( .A(core_v2_reg_59_), .B(core_v3_reg_59_), .Y(core__abc_21302_new_n1889_));
NAND2X1 NAND2X1_152 ( .A(core_v1_reg_62_), .B(core_v0_reg_62_), .Y(core__abc_21302_new_n1925_));
NAND2X1 NAND2X1_153 ( .A(core__abc_21302_new_n1184_), .B(core__abc_21302_new_n1943_), .Y(core__abc_21302_new_n1944_));
NAND2X1 NAND2X1_154 ( .A(core__abc_21302_new_n1945__bF_buf10), .B(core__abc_21302_new_n1217_), .Y(core__abc_21302_new_n1946_));
NAND2X1 NAND2X1_155 ( .A(core__abc_21302_new_n1945__bF_buf8), .B(core__abc_21302_new_n1229_), .Y(core__abc_21302_new_n1949_));
NAND2X1 NAND2X1_156 ( .A(core__abc_21302_new_n1238_), .B(core__abc_21302_new_n1945__bF_buf6), .Y(core__abc_21302_new_n1952_));
NAND2X1 NAND2X1_157 ( .A(core__abc_21302_new_n1945__bF_buf4), .B(core__abc_21302_new_n1248_), .Y(core__abc_21302_new_n1955_));
NAND2X1 NAND2X1_158 ( .A(core__abc_21302_new_n1945__bF_buf2), .B(core__abc_21302_new_n1258_), .Y(core__abc_21302_new_n1958_));
NAND2X1 NAND2X1_159 ( .A(core__abc_21302_new_n1945__bF_buf0), .B(core__abc_21302_new_n1270_), .Y(core__abc_21302_new_n1961_));
NAND2X1 NAND2X1_16 ( .A(_abc_19873_new_n901__bF_buf1), .B(_abc_19873_new_n893__bF_buf1), .Y(_abc_19873_new_n953_));
NAND2X1 NAND2X1_160 ( .A(core__abc_21302_new_n1945__bF_buf9), .B(core__abc_21302_new_n1280_), .Y(core__abc_21302_new_n1964_));
NAND2X1 NAND2X1_161 ( .A(core__abc_21302_new_n1945__bF_buf7), .B(core__abc_21302_new_n1290_), .Y(core__abc_21302_new_n1967_));
NAND2X1 NAND2X1_162 ( .A(core__abc_21302_new_n1945__bF_buf5), .B(core__abc_21302_new_n1298_), .Y(core__abc_21302_new_n1970_));
NAND2X1 NAND2X1_163 ( .A(core__abc_21302_new_n1945__bF_buf3), .B(core__abc_21302_new_n1309_), .Y(core__abc_21302_new_n1973_));
NAND2X1 NAND2X1_164 ( .A(core__abc_21302_new_n1945__bF_buf1), .B(core__abc_21302_new_n1321_), .Y(core__abc_21302_new_n1976_));
NAND2X1 NAND2X1_165 ( .A(core__abc_21302_new_n1945__bF_buf10), .B(core__abc_21302_new_n1333_), .Y(core__abc_21302_new_n1979_));
NAND2X1 NAND2X1_166 ( .A(core__abc_21302_new_n1945__bF_buf8), .B(core__abc_21302_new_n1343_), .Y(core__abc_21302_new_n1982_));
NAND2X1 NAND2X1_167 ( .A(core__abc_21302_new_n1945__bF_buf6), .B(core__abc_21302_new_n1355_), .Y(core__abc_21302_new_n1985_));
NAND2X1 NAND2X1_168 ( .A(core__abc_21302_new_n1945__bF_buf4), .B(core__abc_21302_new_n1367_), .Y(core__abc_21302_new_n1988_));
NAND2X1 NAND2X1_169 ( .A(core__abc_21302_new_n1945__bF_buf2), .B(core__abc_21302_new_n1379_), .Y(core__abc_21302_new_n1991_));
NAND2X1 NAND2X1_17 ( .A(_abc_19873_new_n905__bF_buf3), .B(_abc_19873_new_n889__bF_buf1), .Y(_abc_19873_new_n960_));
NAND2X1 NAND2X1_170 ( .A(core__abc_21302_new_n1945__bF_buf0), .B(core__abc_21302_new_n1390_), .Y(core__abc_21302_new_n1994_));
NAND2X1 NAND2X1_171 ( .A(core__abc_21302_new_n1945__bF_buf9), .B(core__abc_21302_new_n1402_), .Y(core__abc_21302_new_n1997_));
NAND2X1 NAND2X1_172 ( .A(core__abc_21302_new_n1945__bF_buf7), .B(core__abc_21302_new_n1414_), .Y(core__abc_21302_new_n2000_));
NAND2X1 NAND2X1_173 ( .A(core__abc_21302_new_n1945__bF_buf5), .B(core__abc_21302_new_n1426_), .Y(core__abc_21302_new_n2003_));
NAND2X1 NAND2X1_174 ( .A(core__abc_21302_new_n1945__bF_buf3), .B(core__abc_21302_new_n1438_), .Y(core__abc_21302_new_n2006_));
NAND2X1 NAND2X1_175 ( .A(core__abc_21302_new_n1945__bF_buf1), .B(core__abc_21302_new_n1450_), .Y(core__abc_21302_new_n2009_));
NAND2X1 NAND2X1_176 ( .A(core__abc_21302_new_n1945__bF_buf10), .B(core__abc_21302_new_n1462_), .Y(core__abc_21302_new_n2012_));
NAND2X1 NAND2X1_177 ( .A(core__abc_21302_new_n1945__bF_buf8), .B(core__abc_21302_new_n1470_), .Y(core__abc_21302_new_n2015_));
NAND2X1 NAND2X1_178 ( .A(core__abc_21302_new_n1945__bF_buf6), .B(core__abc_21302_new_n1482_), .Y(core__abc_21302_new_n2018_));
NAND2X1 NAND2X1_179 ( .A(core__abc_21302_new_n1945__bF_buf4), .B(core__abc_21302_new_n1492_), .Y(core__abc_21302_new_n2021_));
NAND2X1 NAND2X1_18 ( .A(_abc_19873_new_n889__bF_buf0), .B(_abc_19873_new_n881_), .Y(_abc_19873_new_n969_));
NAND2X1 NAND2X1_180 ( .A(core__abc_21302_new_n1945__bF_buf2), .B(core__abc_21302_new_n1504_), .Y(core__abc_21302_new_n2024_));
NAND2X1 NAND2X1_181 ( .A(core__abc_21302_new_n1945__bF_buf0), .B(core__abc_21302_new_n1516_), .Y(core__abc_21302_new_n2027_));
NAND2X1 NAND2X1_182 ( .A(core__abc_21302_new_n1945__bF_buf9), .B(core__abc_21302_new_n1528_), .Y(core__abc_21302_new_n2030_));
NAND2X1 NAND2X1_183 ( .A(core__abc_21302_new_n1945__bF_buf7), .B(core__abc_21302_new_n1541_), .Y(core__abc_21302_new_n2033_));
NAND2X1 NAND2X1_184 ( .A(core__abc_21302_new_n1945__bF_buf5), .B(core__abc_21302_new_n1553_), .Y(core__abc_21302_new_n2036_));
NAND2X1 NAND2X1_185 ( .A(core__abc_21302_new_n1945__bF_buf3), .B(core__abc_21302_new_n1561_), .Y(core__abc_21302_new_n2039_));
NAND2X1 NAND2X1_186 ( .A(core__abc_21302_new_n1945__bF_buf1), .B(core__abc_21302_new_n1573_), .Y(core__abc_21302_new_n2042_));
NAND2X1 NAND2X1_187 ( .A(core__abc_21302_new_n1945__bF_buf10), .B(core__abc_21302_new_n1585_), .Y(core__abc_21302_new_n2045_));
NAND2X1 NAND2X1_188 ( .A(core__abc_21302_new_n1945__bF_buf8), .B(core__abc_21302_new_n1599_), .Y(core__abc_21302_new_n2048_));
NAND2X1 NAND2X1_189 ( .A(core__abc_21302_new_n1945__bF_buf6), .B(core__abc_21302_new_n1611_), .Y(core__abc_21302_new_n2051_));
NAND2X1 NAND2X1_19 ( .A(_abc_19873_new_n877_), .B(_abc_19873_new_n905__bF_buf1), .Y(_abc_19873_new_n982_));
NAND2X1 NAND2X1_190 ( .A(core__abc_21302_new_n1945__bF_buf4), .B(core__abc_21302_new_n1622_), .Y(core__abc_21302_new_n2054_));
NAND2X1 NAND2X1_191 ( .A(core__abc_21302_new_n1945__bF_buf2), .B(core__abc_21302_new_n1635_), .Y(core__abc_21302_new_n2057_));
NAND2X1 NAND2X1_192 ( .A(core__abc_21302_new_n1945__bF_buf0), .B(core__abc_21302_new_n1644_), .Y(core__abc_21302_new_n2060_));
NAND2X1 NAND2X1_193 ( .A(core__abc_21302_new_n1945__bF_buf9), .B(core__abc_21302_new_n1655_), .Y(core__abc_21302_new_n2063_));
NAND2X1 NAND2X1_194 ( .A(core__abc_21302_new_n1945__bF_buf7), .B(core__abc_21302_new_n1666_), .Y(core__abc_21302_new_n2066_));
NAND2X1 NAND2X1_195 ( .A(core__abc_21302_new_n1945__bF_buf5), .B(core__abc_21302_new_n1677_), .Y(core__abc_21302_new_n2069_));
NAND2X1 NAND2X1_196 ( .A(core__abc_21302_new_n1945__bF_buf3), .B(core__abc_21302_new_n1688_), .Y(core__abc_21302_new_n2072_));
NAND2X1 NAND2X1_197 ( .A(core__abc_21302_new_n1945__bF_buf1), .B(core__abc_21302_new_n1699_), .Y(core__abc_21302_new_n2075_));
NAND2X1 NAND2X1_198 ( .A(core__abc_21302_new_n1945__bF_buf10), .B(core__abc_21302_new_n1711_), .Y(core__abc_21302_new_n2078_));
NAND2X1 NAND2X1_199 ( .A(core__abc_21302_new_n1945__bF_buf8), .B(core__abc_21302_new_n1722_), .Y(core__abc_21302_new_n2081_));
NAND2X1 NAND2X1_2 ( .A(_abc_19873_new_n877_), .B(_abc_19873_new_n874_), .Y(_abc_19873_new_n878_));
NAND2X1 NAND2X1_20 ( .A(_abc_19873_new_n877_), .B(_abc_19873_new_n893__bF_buf4), .Y(_abc_19873_new_n1003_));
NAND2X1 NAND2X1_200 ( .A(core__abc_21302_new_n1945__bF_buf6), .B(core__abc_21302_new_n1734_), .Y(core__abc_21302_new_n2084_));
NAND2X1 NAND2X1_201 ( .A(core__abc_21302_new_n1945__bF_buf4), .B(core__abc_21302_new_n1745_), .Y(core__abc_21302_new_n2087_));
NAND2X1 NAND2X1_202 ( .A(core__abc_21302_new_n1945__bF_buf2), .B(core__abc_21302_new_n1758_), .Y(core__abc_21302_new_n2090_));
NAND2X1 NAND2X1_203 ( .A(core__abc_21302_new_n1945__bF_buf0), .B(core__abc_21302_new_n1767_), .Y(core__abc_21302_new_n2093_));
NAND2X1 NAND2X1_204 ( .A(core__abc_21302_new_n1945__bF_buf9), .B(core__abc_21302_new_n1779_), .Y(core__abc_21302_new_n2096_));
NAND2X1 NAND2X1_205 ( .A(core__abc_21302_new_n1945__bF_buf7), .B(core__abc_21302_new_n1790_), .Y(core__abc_21302_new_n2099_));
NAND2X1 NAND2X1_206 ( .A(core__abc_21302_new_n1945__bF_buf5), .B(core__abc_21302_new_n1804_), .Y(core__abc_21302_new_n2102_));
NAND2X1 NAND2X1_207 ( .A(core__abc_21302_new_n1945__bF_buf3), .B(core__abc_21302_new_n1815_), .Y(core__abc_21302_new_n2105_));
NAND2X1 NAND2X1_208 ( .A(core__abc_21302_new_n1945__bF_buf1), .B(core__abc_21302_new_n1828_), .Y(core__abc_21302_new_n2108_));
NAND2X1 NAND2X1_209 ( .A(core__abc_21302_new_n1945__bF_buf10), .B(core__abc_21302_new_n1841_), .Y(core__abc_21302_new_n2111_));
NAND2X1 NAND2X1_21 ( .A(_abc_19873_new_n1003_), .B(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1019_));
NAND2X1 NAND2X1_210 ( .A(core__abc_21302_new_n1945__bF_buf8), .B(core__abc_21302_new_n1855_), .Y(core__abc_21302_new_n2114_));
NAND2X1 NAND2X1_211 ( .A(core__abc_21302_new_n1945__bF_buf6), .B(core__abc_21302_new_n1867_), .Y(core__abc_21302_new_n2117_));
NAND2X1 NAND2X1_212 ( .A(core__abc_21302_new_n1945__bF_buf4), .B(core__abc_21302_new_n1881_), .Y(core__abc_21302_new_n2120_));
NAND2X1 NAND2X1_213 ( .A(core__abc_21302_new_n1945__bF_buf2), .B(core__abc_21302_new_n1893_), .Y(core__abc_21302_new_n2123_));
NAND2X1 NAND2X1_214 ( .A(core__abc_21302_new_n1945__bF_buf0), .B(core__abc_21302_new_n1907_), .Y(core__abc_21302_new_n2126_));
NAND2X1 NAND2X1_215 ( .A(core__abc_21302_new_n1945__bF_buf9), .B(core__abc_21302_new_n1921_), .Y(core__abc_21302_new_n2129_));
NAND2X1 NAND2X1_216 ( .A(core__abc_21302_new_n1945__bF_buf7), .B(core__abc_21302_new_n1934_), .Y(core__abc_21302_new_n2132_));
NAND2X1 NAND2X1_217 ( .A(core__abc_21302_new_n1945__bF_buf5), .B(core__abc_21302_new_n1940_), .Y(core__abc_21302_new_n2135_));
NAND2X1 NAND2X1_218 ( .A(core__abc_21302_new_n1192_), .B(core__abc_21302_new_n2140_), .Y(core__0ready_reg_0_0_));
NAND2X1 NAND2X1_219 ( .A(core__abc_21302_new_n1184_), .B(core__abc_21302_new_n1176_), .Y(core__abc_21302_new_n2142_));
NAND2X1 NAND2X1_22 ( .A(_abc_19873_new_n905__bF_buf3), .B(_abc_19873_new_n901__bF_buf2), .Y(_abc_19873_new_n1064_));
NAND2X1 NAND2X1_220 ( .A(core_loop_ctr_reg_0_), .B(core_loop_ctr_reg_1_), .Y(core__abc_21302_new_n2150_));
NAND2X1 NAND2X1_221 ( .A(core__abc_21302_new_n2150_), .B(core__abc_21302_new_n2143_), .Y(core__abc_21302_new_n2151_));
NAND2X1 NAND2X1_222 ( .A(core_loop_ctr_reg_2_), .B(core__abc_21302_new_n2154_), .Y(core__abc_21302_new_n2156_));
NAND2X1 NAND2X1_223 ( .A(reset_n_bF_buf22), .B(core__abc_21302_new_n2158_), .Y(core__abc_21302_new_n2159_));
NAND2X1 NAND2X1_224 ( .A(core__abc_21302_new_n1205_), .B(core__abc_21302_new_n2165_), .Y(core__abc_21302_new_n2364_));
NAND2X1 NAND2X1_225 ( .A(core__abc_21302_new_n2377_), .B(core__abc_21302_new_n2376_), .Y(core__abc_21302_new_n2378_));
NAND2X1 NAND2X1_226 ( .A(core__abc_21302_new_n2381_), .B(core__abc_21302_new_n2384_), .Y(core__abc_21302_new_n2385_));
NAND2X1 NAND2X1_227 ( .A(core__abc_21302_new_n2389_), .B(core__abc_21302_new_n2386_), .Y(core__abc_21302_new_n2390_));
NAND2X1 NAND2X1_228 ( .A(core__abc_21302_new_n1360_), .B(core__abc_21302_new_n1372_), .Y(core__abc_21302_new_n2398_));
NAND2X1 NAND2X1_229 ( .A(core__abc_21302_new_n1348_), .B(core__abc_21302_new_n1336_), .Y(core__abc_21302_new_n2399_));
NAND2X1 NAND2X1_23 ( .A(_abc_19873_new_n877_), .B(_abc_19873_new_n895__bF_buf3), .Y(_abc_19873_new_n1140_));
NAND2X1 NAND2X1_230 ( .A(core__abc_21302_new_n1303_), .B(core__abc_21302_new_n1293_), .Y(core__abc_21302_new_n2401_));
NAND2X1 NAND2X1_231 ( .A(core__abc_21302_new_n1314_), .B(core__abc_21302_new_n1326_), .Y(core__abc_21302_new_n2402_));
NAND2X1 NAND2X1_232 ( .A(core__abc_21302_new_n2400_), .B(core__abc_21302_new_n2403_), .Y(core__abc_21302_new_n2404_));
NAND2X1 NAND2X1_233 ( .A(core_v1_reg_9_), .B(core_v0_reg_9_), .Y(core__abc_21302_new_n2407_));
NAND2X1 NAND2X1_234 ( .A(core_v1_reg_12_), .B(core_v0_reg_12_), .Y(core__abc_21302_new_n2413_));
NAND2X1 NAND2X1_235 ( .A(core_v1_reg_13_), .B(core_v0_reg_13_), .Y(core__abc_21302_new_n2414_));
NAND2X1 NAND2X1_236 ( .A(core__abc_21302_new_n2416_), .B(core__abc_21302_new_n2417_), .Y(core__abc_21302_new_n2418_));
NAND2X1 NAND2X1_237 ( .A(core__abc_21302_new_n1546_), .B(core__abc_21302_new_n1558_), .Y(core__abc_21302_new_n2421_));
NAND2X1 NAND2X1_238 ( .A(core__abc_21302_new_n1521_), .B(core__abc_21302_new_n1534_), .Y(core__abc_21302_new_n2422_));
NAND2X1 NAND2X1_239 ( .A(core__abc_21302_new_n1475_), .B(core__abc_21302_new_n1485_), .Y(core__abc_21302_new_n2424_));
NAND2X1 NAND2X1_24 ( .A(_abc_19873_new_n1474_), .B(_abc_19873_new_n1475_), .Y(_abc_19873_new_n1476_));
NAND2X1 NAND2X1_240 ( .A(core__abc_21302_new_n1497_), .B(core__abc_21302_new_n1509_), .Y(core__abc_21302_new_n2425_));
NAND2X1 NAND2X1_241 ( .A(core__abc_21302_new_n2426_), .B(core__abc_21302_new_n2423_), .Y(core__abc_21302_new_n2427_));
NAND2X1 NAND2X1_242 ( .A(core__abc_21302_new_n1455_), .B(core__abc_21302_new_n1467_), .Y(core__abc_21302_new_n2428_));
NAND2X1 NAND2X1_243 ( .A(core__abc_21302_new_n1431_), .B(core__abc_21302_new_n1443_), .Y(core__abc_21302_new_n2429_));
NAND2X1 NAND2X1_244 ( .A(core__abc_21302_new_n1407_), .B(core__abc_21302_new_n1419_), .Y(core__abc_21302_new_n2435_));
NAND2X1 NAND2X1_245 ( .A(core_v1_reg_17_), .B(core_v0_reg_17_), .Y(core__abc_21302_new_n2438_));
NAND2X1 NAND2X1_246 ( .A(core_v1_reg_18_), .B(core_v0_reg_18_), .Y(core__abc_21302_new_n2441_));
NAND2X1 NAND2X1_247 ( .A(core_v1_reg_19_), .B(core_v0_reg_19_), .Y(core__abc_21302_new_n2442_));
NAND2X1 NAND2X1_248 ( .A(core_v1_reg_20_), .B(core_v0_reg_20_), .Y(core__abc_21302_new_n2446_));
NAND2X1 NAND2X1_249 ( .A(core_v1_reg_21_), .B(core_v0_reg_21_), .Y(core__abc_21302_new_n2447_));
NAND2X1 NAND2X1_25 ( .A(we), .B(cs), .Y(_abc_19873_new_n1848_));
NAND2X1 NAND2X1_250 ( .A(core_v1_reg_25_), .B(core_v0_reg_25_), .Y(core__abc_21302_new_n2455_));
NAND2X1 NAND2X1_251 ( .A(core_v1_reg_28_), .B(core_v0_reg_28_), .Y(core__abc_21302_new_n2461_));
NAND2X1 NAND2X1_252 ( .A(core__abc_21302_new_n2463_), .B(core__abc_21302_new_n2460_), .Y(core__abc_21302_new_n2464_));
NAND2X1 NAND2X1_253 ( .A(core_v1_reg_2_), .B(core__abc_21302_new_n2469_), .Y(core__abc_21302_new_n2470_));
NAND2X1 NAND2X1_254 ( .A(core_v0_reg_2_), .B(core__abc_21302_new_n2471_), .Y(core__abc_21302_new_n2472_));
NAND2X1 NAND2X1_255 ( .A(core__abc_21302_new_n2476_), .B(core__abc_21302_new_n2477_), .Y(core__abc_21302_new_n2478_));
NAND2X1 NAND2X1_256 ( .A(core__abc_21302_new_n2481_), .B(core__abc_21302_new_n2482_), .Y(core__abc_21302_new_n2483_));
NAND2X1 NAND2X1_257 ( .A(core__abc_21302_new_n2432_), .B(core__abc_21302_new_n2431_), .Y(core__abc_21302_new_n2495_));
NAND2X1 NAND2X1_258 ( .A(core__abc_21302_new_n2493_), .B(core__abc_21302_new_n2496_), .Y(core__abc_21302_new_n2497_));
NAND2X1 NAND2X1_259 ( .A(core__abc_21302_new_n2430_), .B(core__abc_21302_new_n2445_), .Y(core__abc_21302_new_n2498_));
NAND2X1 NAND2X1_26 ( .A(reset_n_bF_buf22), .B(_abc_19873_new_n2284_), .Y(_abc_19873_new_n2285_));
NAND2X1 NAND2X1_260 ( .A(core__abc_21302_new_n2499_), .B(core__abc_21302_new_n2498_), .Y(core__abc_21302_new_n2500_));
NAND2X1 NAND2X1_261 ( .A(core__abc_21302_new_n2459_), .B(core__abc_21302_new_n2423_), .Y(core__abc_21302_new_n2501_));
NAND2X1 NAND2X1_262 ( .A(core__abc_21302_new_n2502_), .B(core__abc_21302_new_n2501_), .Y(core__abc_21302_new_n2503_));
NAND2X1 NAND2X1_263 ( .A(core__abc_21302_new_n2510_), .B(core__abc_21302_new_n2509_), .Y(core__abc_21302_new_n2511_));
NAND2X1 NAND2X1_264 ( .A(core__abc_21302_new_n2508_), .B(core__abc_21302_new_n2511_), .Y(core__abc_21302_new_n2512_));
NAND2X1 NAND2X1_265 ( .A(core__abc_21302_new_n2516_), .B(core__abc_21302_new_n2518_), .Y(core__abc_21302_new_n2519_));
NAND2X1 NAND2X1_266 ( .A(core__abc_21302_new_n1278_), .B(core__abc_21302_new_n1288_), .Y(core__abc_21302_new_n2520_));
NAND2X1 NAND2X1_267 ( .A(core__abc_21302_new_n1256_), .B(core__abc_21302_new_n1268_), .Y(core__abc_21302_new_n2521_));
NAND2X1 NAND2X1_268 ( .A(core__abc_21302_new_n1365_), .B(core__abc_21302_new_n1377_), .Y(core__abc_21302_new_n2527_));
NAND2X1 NAND2X1_269 ( .A(core__abc_21302_new_n1341_), .B(core__abc_21302_new_n1353_), .Y(core__abc_21302_new_n2528_));
NAND2X1 NAND2X1_27 ( .A(\write_data[0] ), .B(_abc_19873_new_n2286_), .Y(_abc_19873_new_n2287_));
NAND2X1 NAND2X1_270 ( .A(core__abc_21302_new_n2529_), .B(core__abc_21302_new_n2532_), .Y(core__abc_21302_new_n2533_));
NAND2X1 NAND2X1_271 ( .A(core__abc_21302_new_n2534_), .B(core__abc_21302_new_n2535_), .Y(core__abc_21302_new_n2536_));
NAND2X1 NAND2X1_272 ( .A(core__abc_21302_new_n2551_), .B(core__abc_21302_new_n2552_), .Y(core__abc_21302_new_n2553_));
NAND2X1 NAND2X1_273 ( .A(core__abc_21302_new_n1490_), .B(core__abc_21302_new_n1480_), .Y(core__abc_21302_new_n2554_));
NAND2X1 NAND2X1_274 ( .A(core__abc_21302_new_n2560_), .B(core__abc_21302_new_n2561_), .Y(core__abc_21302_new_n2562_));
NAND2X1 NAND2X1_275 ( .A(core__abc_21302_new_n1388_), .B(core__abc_21302_new_n2563_), .Y(core__abc_21302_new_n2564_));
NAND2X1 NAND2X1_276 ( .A(core__abc_21302_new_n2559_), .B(core__abc_21302_new_n2565_), .Y(core__abc_21302_new_n2566_));
NAND2X1 NAND2X1_277 ( .A(core__abc_21302_new_n2557_), .B(core__abc_21302_new_n2558_), .Y(core__abc_21302_new_n2569_));
NAND2X1 NAND2X1_278 ( .A(core__abc_21302_new_n2576_), .B(core__abc_21302_new_n2575_), .Y(core__abc_21302_new_n2577_));
NAND2X1 NAND2X1_279 ( .A(core__abc_21302_new_n2549_), .B(core__abc_21302_new_n2550_), .Y(core__abc_21302_new_n2592_));
NAND2X1 NAND2X1_28 ( .A(\write_data[1] ), .B(_abc_19873_new_n2286_), .Y(_abc_19873_new_n2289_));
NAND2X1 NAND2X1_280 ( .A(core__abc_21302_new_n2549_), .B(core__abc_21302_new_n2598_), .Y(core__abc_21302_new_n2599_));
NAND2X1 NAND2X1_281 ( .A(core__abc_21302_new_n2603_), .B(core__abc_21302_new_n2604_), .Y(core__abc_21302_new_n2605_));
NAND2X1 NAND2X1_282 ( .A(core__abc_21302_new_n2607_), .B(core__abc_21302_new_n2606_), .Y(core__abc_21302_new_n2608_));
NAND2X1 NAND2X1_283 ( .A(core__abc_21302_new_n2617_), .B(core__abc_21302_new_n2603_), .Y(core__abc_21302_new_n2618_));
NAND2X1 NAND2X1_284 ( .A(core__abc_21302_new_n2616_), .B(core__abc_21302_new_n2618_), .Y(core__abc_21302_new_n2619_));
NAND2X1 NAND2X1_285 ( .A(core__abc_21302_new_n2367_), .B(core__abc_21302_new_n2366_), .Y(core__abc_21302_new_n2633_));
NAND2X1 NAND2X1_286 ( .A(core__abc_21302_new_n2637_), .B(core__abc_21302_new_n2366_), .Y(core__abc_21302_new_n2638_));
NAND2X1 NAND2X1_287 ( .A(core__abc_21302_new_n1686_), .B(core__abc_21302_new_n1697_), .Y(core__abc_21302_new_n2660_));
NAND2X1 NAND2X1_288 ( .A(core__abc_21302_new_n2667_), .B(core__abc_21302_new_n2666_), .Y(core__abc_21302_new_n2668_));
NAND2X1 NAND2X1_289 ( .A(core_v3_reg_28_), .B(core__abc_21302_new_n2668_), .Y(core__abc_21302_new_n2669_));
NAND2X1 NAND2X1_29 ( .A(\write_data[2] ), .B(_abc_19873_new_n2286_), .Y(_abc_19873_new_n2291_));
NAND2X1 NAND2X1_290 ( .A(core__abc_21302_new_n1524_), .B(core__abc_21302_new_n2670_), .Y(core__abc_21302_new_n2671_));
NAND2X1 NAND2X1_291 ( .A(core__abc_21302_new_n2669_), .B(core__abc_21302_new_n2671_), .Y(core__abc_21302_new_n2672_));
NAND2X1 NAND2X1_292 ( .A(core__abc_21302_new_n1567_), .B(core__abc_21302_new_n2647_), .Y(core__abc_21302_new_n2683_));
NAND2X1 NAND2X1_293 ( .A(core__abc_21302_new_n2682_), .B(core__abc_21302_new_n2686_), .Y(core__abc_21302_new_n2687_));
NAND2X1 NAND2X1_294 ( .A(core__abc_21302_new_n1237_), .B(core__abc_21302_new_n2517_), .Y(core__abc_21302_new_n2690_));
NAND2X1 NAND2X1_295 ( .A(core__abc_21302_new_n2690_), .B(core__abc_21302_new_n2691_), .Y(core__abc_21302_new_n2692_));
NAND2X1 NAND2X1_296 ( .A(core__abc_21302_new_n2687_), .B(core__abc_21302_new_n2695_), .Y(core__abc_21302_new_n2696_));
NAND2X1 NAND2X1_297 ( .A(core__abc_21302_new_n2694_), .B(core__abc_21302_new_n2698_), .Y(core__abc_21302_new_n2699_));
NAND2X1 NAND2X1_298 ( .A(core__abc_21302_new_n1709_), .B(core__abc_21302_new_n1720_), .Y(core__abc_21302_new_n2719_));
NAND2X1 NAND2X1_299 ( .A(core__abc_21302_new_n2728_), .B(core__abc_21302_new_n2731_), .Y(core__abc_21302_new_n2732_));
NAND2X1 NAND2X1_3 ( .A(\addr[0] ), .B(_abc_19873_new_n879_), .Y(_abc_19873_new_n880_));
NAND2X1 NAND2X1_30 ( .A(core_loop_ctr_reg_3_), .B(core__abc_21302_new_n1133_), .Y(core__abc_21302_new_n1134_));
NAND2X1 NAND2X1_300 ( .A(core__abc_21302_new_n2735_), .B(core__abc_21302_new_n2738_), .Y(core__abc_21302_new_n2739_));
NAND2X1 NAND2X1_301 ( .A(core__abc_21302_new_n2749_), .B(core__abc_21302_new_n2747_), .Y(core__abc_21302_new_n2750_));
NAND2X1 NAND2X1_302 ( .A(core__abc_21302_new_n2682_), .B(core__abc_21302_new_n2737_), .Y(core__abc_21302_new_n2765_));
NAND2X1 NAND2X1_303 ( .A(core__abc_21302_new_n1256_), .B(core__abc_21302_new_n2519_), .Y(core__abc_21302_new_n2772_));
NAND2X1 NAND2X1_304 ( .A(core__abc_21302_new_n2772_), .B(core__abc_21302_new_n2771_), .Y(core__abc_21302_new_n2773_));
NAND2X1 NAND2X1_305 ( .A(core__abc_21302_new_n2774_), .B(core__abc_21302_new_n2777_), .Y(core__abc_21302_new_n2778_));
NAND2X1 NAND2X1_306 ( .A(core__abc_21302_new_n2776_), .B(core__abc_21302_new_n2778_), .Y(core__abc_21302_new_n2779_));
NAND2X1 NAND2X1_307 ( .A(core__abc_21302_new_n2800_), .B(core__abc_21302_new_n2801_), .Y(core__abc_21302_new_n2802_));
NAND2X1 NAND2X1_308 ( .A(core__abc_21302_new_n2803_), .B(core__abc_21302_new_n2802_), .Y(core__abc_21302_new_n2809_));
NAND2X1 NAND2X1_309 ( .A(core__abc_21302_new_n2810_), .B(core__abc_21302_new_n2809_), .Y(core__abc_21302_new_n2811_));
NAND2X1 NAND2X1_31 ( .A(core_siphash_ctrl_reg_4_), .B(core__abc_21302_new_n1145_), .Y(core__abc_21302_new_n1146_));
NAND2X1 NAND2X1_310 ( .A(core__abc_21302_new_n2808_), .B(core__abc_21302_new_n2811_), .Y(core__abc_21302_new_n2812_));
NAND2X1 NAND2X1_311 ( .A(core__abc_21302_new_n2814_), .B(core__abc_21302_new_n2720_), .Y(core__abc_21302_new_n2815_));
NAND2X1 NAND2X1_312 ( .A(core__abc_21302_new_n2824_), .B(core__abc_21302_new_n2818_), .Y(core__abc_21302_new_n2825_));
NAND2X1 NAND2X1_313 ( .A(core__abc_21302_new_n2847_), .B(core__abc_21302_new_n2849_), .Y(core__abc_21302_new_n2850_));
NAND2X1 NAND2X1_314 ( .A(core__abc_21302_new_n2854_), .B(core__abc_21302_new_n2853_), .Y(core__abc_21302_new_n2855_));
NAND2X1 NAND2X1_315 ( .A(core__abc_21302_new_n2852_), .B(core__abc_21302_new_n2855_), .Y(core__abc_21302_new_n2856_));
NAND2X1 NAND2X1_316 ( .A(core__abc_21302_new_n2807_), .B(core__abc_21302_new_n2809_), .Y(core__abc_21302_new_n2858_));
NAND2X1 NAND2X1_317 ( .A(core__abc_21302_new_n2887_), .B(core__abc_21302_new_n2881_), .Y(core__abc_21302_new_n2888_));
NAND2X1 NAND2X1_318 ( .A(core__abc_21302_new_n2886_), .B(core__abc_21302_new_n2890_), .Y(core__abc_21302_new_n2891_));
NAND2X1 NAND2X1_319 ( .A(core__abc_21302_new_n2891_), .B(core__abc_21302_new_n2888_), .Y(core__abc_21302_new_n2892_));
NAND2X1 NAND2X1_32 ( .A(core__abc_21302_new_n1149_), .B(core__abc_21302_new_n1150_), .Y(core__abc_21302_new_n1151_));
NAND2X1 NAND2X1_320 ( .A(core_v3_reg_34_), .B(core__abc_21302_new_n2904_), .Y(core__abc_21302_new_n2905_));
NAND2X1 NAND2X1_321 ( .A(core__abc_21302_new_n2903_), .B(core__abc_21302_new_n2905_), .Y(core__abc_21302_new_n2906_));
NAND2X1 NAND2X1_322 ( .A(core__abc_21302_new_n2921_), .B(core__abc_21302_new_n2841_), .Y(core__abc_21302_new_n2922_));
NAND2X1 NAND2X1_323 ( .A(core__abc_21302_new_n2840_), .B(core__abc_21302_new_n2921_), .Y(core__abc_21302_new_n2923_));
NAND2X1 NAND2X1_324 ( .A(core__abc_21302_new_n2923_), .B(core__abc_21302_new_n2924_), .Y(core__abc_21302_new_n2932_));
NAND2X1 NAND2X1_325 ( .A(core__abc_21302_new_n2941_), .B(core__abc_21302_new_n2937_), .Y(core__abc_21302_new_n2942_));
NAND2X1 NAND2X1_326 ( .A(core__abc_21302_new_n2951_), .B(core__abc_21302_new_n2950_), .Y(core__abc_21302_new_n2952_));
NAND2X1 NAND2X1_327 ( .A(core_v3_reg_35_), .B(core__abc_21302_new_n2953_), .Y(core__abc_21302_new_n2954_));
NAND2X1 NAND2X1_328 ( .A(core__abc_21302_new_n1607_), .B(core__abc_21302_new_n2952_), .Y(core__abc_21302_new_n2955_));
NAND2X1 NAND2X1_329 ( .A(core__abc_21302_new_n2955_), .B(core__abc_21302_new_n2954_), .Y(core__abc_21302_new_n2956_));
NAND2X1 NAND2X1_33 ( .A(core__abc_21302_new_n1160_), .B(core__abc_21302_new_n1161_), .Y(core__abc_21302_new_n1162_));
NAND2X1 NAND2X1_330 ( .A(core__abc_21302_new_n1671_), .B(core__abc_21302_new_n2964_), .Y(core__abc_21302_new_n2965_));
NAND2X1 NAND2X1_331 ( .A(core__abc_21302_new_n2967_), .B(core__abc_21302_new_n2965_), .Y(core__abc_21302_new_n2968_));
NAND2X1 NAND2X1_332 ( .A(core__abc_21302_new_n2971_), .B(core__abc_21302_new_n2968_), .Y(core__abc_21302_new_n2972_));
NAND2X1 NAND2X1_333 ( .A(core__abc_21302_new_n2974_), .B(core__abc_21302_new_n2973_), .Y(core__abc_21302_new_n2975_));
NAND2X1 NAND2X1_334 ( .A(core__abc_21302_new_n2972_), .B(core__abc_21302_new_n2975_), .Y(core__abc_21302_new_n2976_));
NAND2X1 NAND2X1_335 ( .A(core__abc_21302_new_n2981_), .B(core__abc_21302_new_n2897_), .Y(core__abc_21302_new_n2982_));
NAND2X1 NAND2X1_336 ( .A(core__abc_21302_new_n2985_), .B(core__abc_21302_new_n2984_), .Y(core__abc_21302_new_n2986_));
NAND2X1 NAND2X1_337 ( .A(core__abc_21302_new_n2989_), .B(core__abc_21302_new_n2988_), .Y(core__abc_21302_new_n2990_));
NAND2X1 NAND2X1_338 ( .A(core__abc_21302_new_n1660_), .B(core__abc_21302_new_n1671_), .Y(core__abc_21302_new_n3007_));
NAND2X1 NAND2X1_339 ( .A(core__abc_21302_new_n2538_), .B(core__abc_21302_new_n3016_), .Y(core__abc_21302_new_n3017_));
NAND2X1 NAND2X1_34 ( .A(core__abc_21302_new_n1166_), .B(core__abc_21302_new_n1162_), .Y(core__abc_21302_new_n1167_));
NAND2X1 NAND2X1_340 ( .A(core__abc_21302_new_n3022_), .B(core__abc_21302_new_n3021_), .Y(core__abc_21302_new_n3023_));
NAND2X1 NAND2X1_341 ( .A(core__abc_21302_new_n1814_), .B(core__abc_21302_new_n3026_), .Y(core__abc_21302_new_n3028_));
NAND2X1 NAND2X1_342 ( .A(core__abc_21302_new_n3028_), .B(core__abc_21302_new_n3027_), .Y(core__abc_21302_new_n3029_));
NAND2X1 NAND2X1_343 ( .A(core_v3_reg_37_), .B(core__abc_21302_new_n3030_), .Y(core__abc_21302_new_n3032_));
NAND2X1 NAND2X1_344 ( .A(core__abc_21302_new_n3032_), .B(core__abc_21302_new_n3031_), .Y(core__abc_21302_new_n3033_));
NAND2X1 NAND2X1_345 ( .A(core__abc_21302_new_n3024_), .B(core__abc_21302_new_n3005_), .Y(core__abc_21302_new_n3043_));
NAND2X1 NAND2X1_346 ( .A(core__abc_21302_new_n1693_), .B(core__abc_21302_new_n3045_), .Y(core__abc_21302_new_n3046_));
NAND2X1 NAND2X1_347 ( .A(core__abc_21302_new_n2534_), .B(core__abc_21302_new_n3017_), .Y(core__abc_21302_new_n3049_));
NAND2X1 NAND2X1_348 ( .A(core__abc_21302_new_n1331_), .B(core__abc_21302_new_n3050_), .Y(core__abc_21302_new_n3052_));
NAND2X1 NAND2X1_349 ( .A(core_v3_reg_59_), .B(core__abc_21302_new_n3053_), .Y(core__abc_21302_new_n3054_));
NAND2X1 NAND2X1_35 ( .A(core__abc_21302_new_n1147_), .B(core__abc_21302_new_n1181_), .Y(core__abc_21302_new_n1182_));
NAND2X1 NAND2X1_350 ( .A(core__abc_21302_new_n3048_), .B(core__abc_21302_new_n3046_), .Y(core__abc_21302_new_n3058_));
NAND2X1 NAND2X1_351 ( .A(core__abc_21302_new_n3054_), .B(core__abc_21302_new_n3055_), .Y(core__abc_21302_new_n3059_));
NAND2X1 NAND2X1_352 ( .A(core__abc_21302_new_n3059_), .B(core__abc_21302_new_n3058_), .Y(core__abc_21302_new_n3060_));
NAND2X1 NAND2X1_353 ( .A(core__abc_21302_new_n3060_), .B(core__abc_21302_new_n3057_), .Y(core__abc_21302_new_n3061_));
NAND2X1 NAND2X1_354 ( .A(core__abc_21302_new_n1814_), .B(core__abc_21302_new_n1802_), .Y(core__abc_21302_new_n3064_));
NAND2X1 NAND2X1_355 ( .A(core__abc_21302_new_n1826_), .B(core__abc_21302_new_n3066_), .Y(core__abc_21302_new_n3067_));
NAND2X1 NAND2X1_356 ( .A(core_v3_reg_38_), .B(core__abc_21302_new_n3071_), .Y(core__abc_21302_new_n3072_));
NAND2X1 NAND2X1_357 ( .A(core__abc_21302_new_n3070_), .B(core__abc_21302_new_n3072_), .Y(core__abc_21302_new_n3073_));
NAND2X1 NAND2X1_358 ( .A(core__abc_21302_new_n3057_), .B(core__abc_21302_new_n3084_), .Y(core__abc_21302_new_n3085_));
NAND2X1 NAND2X1_359 ( .A(core__abc_21302_new_n1682_), .B(core__abc_21302_new_n1693_), .Y(core__abc_21302_new_n3091_));
NAND2X1 NAND2X1_36 ( .A(reset_n_bF_buf19), .B(core__abc_21302_new_n1180_), .Y(core__abc_21302_new_n1196_));
NAND2X1 NAND2X1_360 ( .A(core__abc_21302_new_n1705_), .B(core__abc_21302_new_n3097_), .Y(core__abc_21302_new_n3098_));
NAND2X1 NAND2X1_361 ( .A(core__abc_21302_new_n3100_), .B(core__abc_21302_new_n3098_), .Y(core__abc_21302_new_n3101_));
NAND2X1 NAND2X1_362 ( .A(core__abc_21302_new_n1341_), .B(core__abc_21302_new_n3103_), .Y(core__abc_21302_new_n3104_));
NAND2X1 NAND2X1_363 ( .A(core__abc_21302_new_n3113_), .B(core__abc_21302_new_n3115_), .Y(core__abc_21302_new_n3116_));
NAND2X1 NAND2X1_364 ( .A(core__abc_21302_new_n3111_), .B(core__abc_21302_new_n3116_), .Y(core__abc_21302_new_n3118_));
NAND2X1 NAND2X1_365 ( .A(core__abc_21302_new_n1716_), .B(core__abc_21302_new_n3132_), .Y(core__abc_21302_new_n3133_));
NAND2X1 NAND2X1_366 ( .A(core__abc_21302_new_n3135_), .B(core__abc_21302_new_n3133_), .Y(core__abc_21302_new_n3136_));
NAND2X1 NAND2X1_367 ( .A(core__abc_21302_new_n3137_), .B(core__abc_21302_new_n3138_), .Y(core__abc_21302_new_n3140_));
NAND2X1 NAND2X1_368 ( .A(core__abc_21302_new_n1917_), .B(core__abc_21302_new_n3141_), .Y(core__abc_21302_new_n3142_));
NAND2X1 NAND2X1_369 ( .A(core__abc_21302_new_n3140_), .B(core__abc_21302_new_n3139_), .Y(core__abc_21302_new_n3143_));
NAND2X1 NAND2X1_37 ( .A(core__abc_21302_new_n1186_), .B(core__abc_21302_new_n1179_), .Y(core__abc_21302_new_n1201_));
NAND2X1 NAND2X1_370 ( .A(core_v3_reg_61_), .B(core__abc_21302_new_n3143_), .Y(core__abc_21302_new_n3144_));
NAND2X1 NAND2X1_371 ( .A(core__abc_21302_new_n3144_), .B(core__abc_21302_new_n3142_), .Y(core__abc_21302_new_n3145_));
NAND2X1 NAND2X1_372 ( .A(core__abc_21302_new_n3145_), .B(core__abc_21302_new_n3136_), .Y(core__abc_21302_new_n3146_));
NAND2X1 NAND2X1_373 ( .A(core__abc_21302_new_n3109_), .B(core__abc_21302_new_n3090_), .Y(core__abc_21302_new_n3150_));
NAND2X1 NAND2X1_374 ( .A(core__abc_21302_new_n1853_), .B(core__abc_21302_new_n3161_), .Y(core__abc_21302_new_n3162_));
NAND2X1 NAND2X1_375 ( .A(core__abc_21302_new_n3162_), .B(core__abc_21302_new_n3163_), .Y(core__abc_21302_new_n3164_));
NAND2X1 NAND2X1_376 ( .A(core_v3_reg_40_), .B(core__abc_21302_new_n3164_), .Y(core__abc_21302_new_n3165_));
NAND2X1 NAND2X1_377 ( .A(core__abc_21302_new_n3165_), .B(core__abc_21302_new_n3166_), .Y(core__abc_21302_new_n3167_));
NAND2X1 NAND2X1_378 ( .A(core__abc_21302_new_n1705_), .B(core__abc_21302_new_n3134_), .Y(core__abc_21302_new_n3179_));
NAND2X1 NAND2X1_379 ( .A(core_v3_reg_62_), .B(core__abc_21302_new_n3195_), .Y(core__abc_21302_new_n3196_));
NAND2X1 NAND2X1_38 ( .A(core_finalize), .B(core__abc_21302_new_n1198_), .Y(core__abc_21302_new_n1204_));
NAND2X1 NAND2X1_380 ( .A(core__abc_21302_new_n3194_), .B(core__abc_21302_new_n3196_), .Y(core__abc_21302_new_n3197_));
NAND2X1 NAND2X1_381 ( .A(core__abc_21302_new_n1728_), .B(core__abc_21302_new_n3184_), .Y(core__abc_21302_new_n3199_));
NAND2X1 NAND2X1_382 ( .A(core__abc_21302_new_n3207_), .B(core__abc_21302_new_n3161_), .Y(core__abc_21302_new_n3208_));
NAND2X1 NAND2X1_383 ( .A(core_v3_reg_41_), .B(core__abc_21302_new_n3210_), .Y(core__abc_21302_new_n3211_));
NAND2X1 NAND2X1_384 ( .A(core__abc_21302_new_n3212_), .B(core__abc_21302_new_n3213_), .Y(core__abc_21302_new_n3214_));
NAND2X1 NAND2X1_385 ( .A(core__abc_21302_new_n3214_), .B(core__abc_21302_new_n3211_), .Y(core__abc_21302_new_n3215_));
NAND2X1 NAND2X1_386 ( .A(core_v3_reg_63_), .B(core__abc_21302_new_n3230_), .Y(core__abc_21302_new_n3231_));
NAND2X1 NAND2X1_387 ( .A(core__abc_21302_new_n3227_), .B(core__abc_21302_new_n3229_), .Y(core__abc_21302_new_n3233_));
NAND2X1 NAND2X1_388 ( .A(core__abc_21302_new_n3232_), .B(core__abc_21302_new_n3233_), .Y(core__abc_21302_new_n3234_));
NAND2X1 NAND2X1_389 ( .A(core__abc_21302_new_n3234_), .B(core__abc_21302_new_n3231_), .Y(core__abc_21302_new_n3240_));
NAND2X1 NAND2X1_39 ( .A(core_v1_reg_0_), .B(core_v0_reg_0_), .Y(core__abc_21302_new_n1209_));
NAND2X1 NAND2X1_390 ( .A(core__abc_21302_new_n3236_), .B(core__abc_21302_new_n3241_), .Y(core__abc_21302_new_n3242_));
NAND2X1 NAND2X1_391 ( .A(core__abc_21302_new_n3242_), .B(core__abc_21302_new_n3223_), .Y(core__abc_21302_new_n3244_));
NAND2X1 NAND2X1_392 ( .A(core__abc_21302_new_n3244_), .B(core__abc_21302_new_n3243_), .Y(core__abc_21302_new_n3245_));
NAND2X1 NAND2X1_393 ( .A(core__abc_21302_new_n3247_), .B(core__abc_21302_new_n3208_), .Y(core__abc_21302_new_n3248_));
NAND2X1 NAND2X1_394 ( .A(core__abc_21302_new_n1879_), .B(core__abc_21302_new_n3248_), .Y(core__abc_21302_new_n3253_));
NAND2X1 NAND2X1_395 ( .A(core__abc_21302_new_n3254_), .B(core__abc_21302_new_n3251_), .Y(core__abc_21302_new_n3255_));
NAND2X1 NAND2X1_396 ( .A(core__abc_21302_new_n3134_), .B(core__abc_21302_new_n3132_), .Y(core__abc_21302_new_n3267_));
NAND2X1 NAND2X1_397 ( .A(core__abc_21302_new_n3268_), .B(core__abc_21302_new_n3267_), .Y(core__abc_21302_new_n3269_));
NAND2X1 NAND2X1_398 ( .A(core__abc_21302_new_n3270_), .B(core__abc_21302_new_n3269_), .Y(core__abc_21302_new_n3271_));
NAND2X1 NAND2X1_399 ( .A(core__abc_21302_new_n3274_), .B(core__abc_21302_new_n3086_), .Y(core__abc_21302_new_n3276_));
NAND2X1 NAND2X1_4 ( .A(\addr[4] ), .B(_abc_19873_new_n887_), .Y(_abc_19873_new_n888_));
NAND2X1 NAND2X1_40 ( .A(core_v2_reg_0_), .B(core_v3_reg_0_), .Y(core__abc_21302_new_n1213_));
NAND2X1 NAND2X1_400 ( .A(core__abc_21302_new_n3224_), .B(core__abc_21302_new_n3226_), .Y(core__abc_21302_new_n3280_));
NAND2X1 NAND2X1_401 ( .A(core__abc_21302_new_n3202_), .B(core__abc_21302_new_n3241_), .Y(core__abc_21302_new_n3281_));
NAND2X1 NAND2X1_402 ( .A(core__abc_21302_new_n1739_), .B(core__abc_21302_new_n1728_), .Y(core__abc_21302_new_n3286_));
NAND2X1 NAND2X1_403 ( .A(core__abc_21302_new_n3095_), .B(core__abc_21302_new_n3287_), .Y(core__abc_21302_new_n3288_));
NAND2X1 NAND2X1_404 ( .A(core__abc_21302_new_n3289_), .B(core__abc_21302_new_n2927_), .Y(core__abc_21302_new_n3295_));
NAND2X1 NAND2X1_405 ( .A(core__abc_21302_new_n3300_), .B(core__abc_21302_new_n3303_), .Y(core__abc_21302_new_n3304_));
NAND2X1 NAND2X1_406 ( .A(core__abc_21302_new_n3304_), .B(core__abc_21302_new_n3302_), .Y(core__abc_21302_new_n3305_));
NAND2X1 NAND2X1_407 ( .A(core__abc_21302_new_n3306_), .B(core__abc_21302_new_n3285_), .Y(core__abc_21302_new_n3307_));
NAND2X1 NAND2X1_408 ( .A(core__abc_21302_new_n1750_), .B(core__abc_21302_new_n1761_), .Y(core__abc_21302_new_n3334_));
NAND2X1 NAND2X1_409 ( .A(core__abc_21302_new_n1761_), .B(core__abc_21302_new_n1751_), .Y(core__abc_21302_new_n3335_));
NAND2X1 NAND2X1_41 ( .A(core_v1_reg_1_), .B(core_v0_reg_1_), .Y(core__abc_21302_new_n1221_));
NAND2X1 NAND2X1_410 ( .A(core__abc_21302_new_n1388_), .B(core__abc_21302_new_n2548_), .Y(core__abc_21302_new_n3338_));
NAND2X1 NAND2X1_411 ( .A(core__abc_21302_new_n1385_), .B(core__abc_21302_new_n3338_), .Y(core__abc_21302_new_n3339_));
NAND2X1 NAND2X1_412 ( .A(core__abc_21302_new_n3341_), .B(core__abc_21302_new_n3337_), .Y(core__abc_21302_new_n3342_));
NAND2X1 NAND2X1_413 ( .A(core__abc_21302_new_n3342_), .B(core__abc_21302_new_n3344_), .Y(core__abc_21302_new_n3345_));
NAND2X1 NAND2X1_414 ( .A(core__abc_21302_new_n3304_), .B(core__abc_21302_new_n3346_), .Y(core__abc_21302_new_n3347_));
NAND2X1 NAND2X1_415 ( .A(core_v3_reg_44_), .B(core__abc_21302_new_n3358_), .Y(core__abc_21302_new_n3359_));
NAND2X1 NAND2X1_416 ( .A(core__abc_21302_new_n3356_), .B(core__abc_21302_new_n3359_), .Y(core__abc_21302_new_n3360_));
NAND2X1 NAND2X1_417 ( .A(core__abc_21302_new_n1905_), .B(core__abc_21302_new_n3353_), .Y(core__abc_21302_new_n3400_));
NAND2X1 NAND2X1_418 ( .A(core__abc_21302_new_n3402_), .B(core__abc_21302_new_n3406_), .Y(core__abc_21302_new_n3407_));
NAND2X1 NAND2X1_419 ( .A(core__abc_21302_new_n1424_), .B(core__abc_21302_new_n3420_), .Y(core__abc_21302_new_n3422_));
NAND2X1 NAND2X1_42 ( .A(core_v2_reg_1_), .B(core_v3_reg_1_), .Y(core__abc_21302_new_n1224_));
NAND2X1 NAND2X1_420 ( .A(core__abc_21302_new_n3423_), .B(core__abc_21302_new_n3427_), .Y(core__abc_21302_new_n3428_));
NAND2X1 NAND2X1_421 ( .A(core__abc_21302_new_n3435_), .B(core__abc_21302_new_n3416_), .Y(core__abc_21302_new_n3437_));
NAND2X1 NAND2X1_422 ( .A(core__abc_21302_new_n3437_), .B(core__abc_21302_new_n3436_), .Y(core__abc_21302_new_n3438_));
NAND2X1 NAND2X1_423 ( .A(core__abc_21302_new_n3448_), .B(core__abc_21302_new_n3447_), .Y(core__abc_21302_new_n3449_));
NAND2X1 NAND2X1_424 ( .A(core__abc_21302_new_n3419_), .B(core__abc_21302_new_n3417_), .Y(core__abc_21302_new_n3458_));
NAND2X1 NAND2X1_425 ( .A(core__abc_21302_new_n3381_), .B(core__abc_21302_new_n3469_), .Y(core__abc_21302_new_n3470_));
NAND2X1 NAND2X1_426 ( .A(core__abc_21302_new_n3471_), .B(core__abc_21302_new_n3470_), .Y(core__abc_21302_new_n3472_));
NAND2X1 NAND2X1_427 ( .A(core__abc_21302_new_n3378_), .B(core__abc_21302_new_n3469_), .Y(core__abc_21302_new_n3473_));
NAND2X1 NAND2X1_428 ( .A(core__abc_21302_new_n1436_), .B(core__abc_21302_new_n3478_), .Y(core__abc_21302_new_n3480_));
NAND2X1 NAND2X1_429 ( .A(core__abc_21302_new_n3480_), .B(core__abc_21302_new_n3479_), .Y(core__abc_21302_new_n3481_));
NAND2X1 NAND2X1_43 ( .A(core_v1_reg_3_), .B(core_v0_reg_3_), .Y(core__abc_21302_new_n1242_));
NAND2X1 NAND2X1_430 ( .A(core__abc_21302_new_n3476_), .B(core__abc_21302_new_n3482_), .Y(core__abc_21302_new_n3483_));
NAND2X1 NAND2X1_431 ( .A(core__abc_21302_new_n3483_), .B(core__abc_21302_new_n3484_), .Y(core__abc_21302_new_n3485_));
NAND2X1 NAND2X1_432 ( .A(core__abc_21302_new_n1811_), .B(core__abc_21302_new_n3505_), .Y(core__abc_21302_new_n3506_));
NAND2X1 NAND2X1_433 ( .A(core__abc_21302_new_n3507_), .B(core__abc_21302_new_n3509_), .Y(core__abc_21302_new_n3510_));
NAND2X1 NAND2X1_434 ( .A(core__abc_21302_new_n1448_), .B(core__abc_21302_new_n3508_), .Y(core__abc_21302_new_n3511_));
NAND2X1 NAND2X1_435 ( .A(core__abc_21302_new_n3511_), .B(core__abc_21302_new_n3510_), .Y(core__abc_21302_new_n3514_));
NAND2X1 NAND2X1_436 ( .A(core__abc_21302_new_n3513_), .B(core__abc_21302_new_n3514_), .Y(core__abc_21302_new_n3515_));
NAND2X1 NAND2X1_437 ( .A(core__abc_21302_new_n3512_), .B(core__abc_21302_new_n3515_), .Y(core__abc_21302_new_n3516_));
NAND2X1 NAND2X1_438 ( .A(core__abc_21302_new_n3506_), .B(core__abc_21302_new_n3503_), .Y(core__abc_21302_new_n3518_));
NAND2X1 NAND2X1_439 ( .A(core__abc_21302_new_n3486_), .B(core__abc_21302_new_n3520_), .Y(core__abc_21302_new_n3532_));
NAND2X1 NAND2X1_44 ( .A(core__abc_21302_new_n1242_), .B(core__abc_21302_new_n1241_), .Y(core__abc_21302_new_n1243_));
NAND2X1 NAND2X1_440 ( .A(core__abc_21302_new_n1797_), .B(core__abc_21302_new_n1811_), .Y(core__abc_21302_new_n3539_));
NAND2X1 NAND2X1_441 ( .A(core__abc_21302_new_n2575_), .B(core__abc_21302_new_n3549_), .Y(core__abc_21302_new_n3553_));
NAND2X1 NAND2X1_442 ( .A(core__abc_21302_new_n1821_), .B(core__abc_21302_new_n3546_), .Y(core__abc_21302_new_n3558_));
NAND2X1 NAND2X1_443 ( .A(core__abc_21302_new_n3555_), .B(core__abc_21302_new_n3552_), .Y(core__abc_21302_new_n3560_));
NAND2X1 NAND2X1_444 ( .A(core__abc_21302_new_n1834_), .B(core__abc_21302_new_n3578_), .Y(core__abc_21302_new_n3579_));
NAND2X1 NAND2X1_445 ( .A(core__abc_21302_new_n3582_), .B(core__abc_21302_new_n3586_), .Y(core__abc_21302_new_n3587_));
NAND2X1 NAND2X1_446 ( .A(core__abc_21302_new_n3576_), .B(core__abc_21302_new_n3578_), .Y(core__abc_21302_new_n3590_));
NAND2X1 NAND2X1_447 ( .A(core__abc_21302_new_n3592_), .B(core__abc_21302_new_n3575_), .Y(core__abc_21302_new_n3593_));
NAND2X1 NAND2X1_448 ( .A(core__abc_21302_new_n3593_), .B(core__abc_21302_new_n3594_), .Y(core__abc_21302_new_n3595_));
NAND2X1 NAND2X1_449 ( .A(core__abc_21302_new_n3561_), .B(core__abc_21302_new_n3557_), .Y(core__abc_21302_new_n3605_));
NAND2X1 NAND2X1_45 ( .A(core_v1_reg_4_), .B(core_v0_reg_4_), .Y(core__abc_21302_new_n1252_));
NAND2X1 NAND2X1_450 ( .A(core__abc_21302_new_n3534_), .B(core__abc_21302_new_n3606_), .Y(core__abc_21302_new_n3608_));
NAND2X1 NAND2X1_451 ( .A(core__abc_21302_new_n1821_), .B(core__abc_21302_new_n1834_), .Y(core__abc_21302_new_n3618_));
NAND2X1 NAND2X1_452 ( .A(core__abc_21302_new_n3637_), .B(core__abc_21302_new_n3635_), .Y(core__abc_21302_new_n3638_));
NAND2X1 NAND2X1_453 ( .A(core__abc_21302_new_n3639_), .B(core__abc_21302_new_n3642_), .Y(core__abc_21302_new_n3643_));
NAND2X1 NAND2X1_454 ( .A(core__abc_21302_new_n3643_), .B(core__abc_21302_new_n3641_), .Y(core__abc_21302_new_n3644_));
NAND2X1 NAND2X1_455 ( .A(core__abc_21302_new_n3659_), .B(core__abc_21302_new_n3658_), .Y(core__abc_21302_new_n3660_));
NAND2X1 NAND2X1_456 ( .A(core__abc_21302_new_n3661_), .B(core__abc_21302_new_n3664_), .Y(core__abc_21302_new_n3665_));
NAND2X1 NAND2X1_457 ( .A(core__abc_21302_new_n1490_), .B(core__abc_21302_new_n3663_), .Y(core__abc_21302_new_n3666_));
NAND2X1 NAND2X1_458 ( .A(core__abc_21302_new_n3666_), .B(core__abc_21302_new_n3665_), .Y(core__abc_21302_new_n3667_));
NAND2X1 NAND2X1_459 ( .A(core_v3_reg_9_), .B(core__abc_21302_new_n3667_), .Y(core__abc_21302_new_n3668_));
NAND2X1 NAND2X1_46 ( .A(core__abc_21302_new_n1252_), .B(core__abc_21302_new_n1251_), .Y(core__abc_21302_new_n1253_));
NAND2X1 NAND2X1_460 ( .A(core__abc_21302_new_n3670_), .B(core__abc_21302_new_n3668_), .Y(core__abc_21302_new_n3671_));
NAND2X1 NAND2X1_461 ( .A(core__abc_21302_new_n3660_), .B(core__abc_21302_new_n3672_), .Y(core__abc_21302_new_n3673_));
NAND2X1 NAND2X1_462 ( .A(core__abc_21302_new_n3671_), .B(core__abc_21302_new_n3674_), .Y(core__abc_21302_new_n3675_));
NAND2X1 NAND2X1_463 ( .A(core__abc_21302_new_n3673_), .B(core__abc_21302_new_n3675_), .Y(core__abc_21302_new_n3676_));
NAND2X1 NAND2X1_464 ( .A(core__abc_21302_new_n1874_), .B(core__abc_21302_new_n3699_), .Y(core__abc_21302_new_n3700_));
NAND2X1 NAND2X1_465 ( .A(core_v3_reg_10_), .B(core__abc_21302_new_n3708_), .Y(core__abc_21302_new_n3709_));
NAND2X1 NAND2X1_466 ( .A(core__abc_21302_new_n3707_), .B(core__abc_21302_new_n3709_), .Y(core__abc_21302_new_n3714_));
NAND2X1 NAND2X1_467 ( .A(core__abc_21302_new_n3715_), .B(core__abc_21302_new_n3711_), .Y(core__abc_21302_new_n3716_));
NAND2X1 NAND2X1_468 ( .A(core__abc_21302_new_n2551_), .B(core__abc_21302_new_n3704_), .Y(core__abc_21302_new_n3734_));
NAND2X1 NAND2X1_469 ( .A(core__abc_21302_new_n3738_), .B(core__abc_21302_new_n3741_), .Y(core__abc_21302_new_n3746_));
NAND2X1 NAND2X1_47 ( .A(core__abc_21302_new_n1261_), .B(core__abc_21302_new_n1262_), .Y(core__abc_21302_new_n1263_));
NAND2X1 NAND2X1_470 ( .A(core__abc_21302_new_n3748_), .B(core__abc_21302_new_n3729_), .Y(core__abc_21302_new_n3749_));
NAND2X1 NAND2X1_471 ( .A(core__abc_21302_new_n3749_), .B(core__abc_21302_new_n3750_), .Y(core__abc_21302_new_n3751_));
NAND2X1 NAND2X1_472 ( .A(core__abc_21302_new_n3769_), .B(core__abc_21302_new_n3695_), .Y(core__abc_21302_new_n3770_));
NAND2X1 NAND2X1_473 ( .A(core__abc_21302_new_n2887_), .B(core__abc_21302_new_n3782_), .Y(core__abc_21302_new_n3783_));
NAND2X1 NAND2X1_474 ( .A(core__abc_21302_new_n1899_), .B(core__abc_21302_new_n1914_), .Y(core__abc_21302_new_n3791_));
NAND2X1 NAND2X1_475 ( .A(core__abc_21302_new_n1900_), .B(core__abc_21302_new_n3773_), .Y(core__abc_21302_new_n3792_));
NAND2X1 NAND2X1_476 ( .A(core__abc_21302_new_n3807_), .B(core__abc_21302_new_n3776_), .Y(core__abc_21302_new_n3808_));
NAND2X1 NAND2X1_477 ( .A(core__abc_21302_new_n1539_), .B(core__abc_21302_new_n3810_), .Y(core__abc_21302_new_n3811_));
NAND2X1 NAND2X1_478 ( .A(core__abc_21302_new_n3812_), .B(core__abc_21302_new_n3815_), .Y(core__abc_21302_new_n3816_));
NAND2X1 NAND2X1_479 ( .A(core__abc_21302_new_n1551_), .B(core__abc_21302_new_n3837_), .Y(core__abc_21302_new_n3846_));
NAND2X1 NAND2X1_48 ( .A(core_v1_reg_5_), .B(core_v0_reg_5_), .Y(core__abc_21302_new_n1264_));
NAND2X1 NAND2X1_480 ( .A(core__abc_21302_new_n3847_), .B(core__abc_21302_new_n3840_), .Y(core__abc_21302_new_n3852_));
NAND2X1 NAND2X1_481 ( .A(core__abc_21302_new_n3853_), .B(core__abc_21302_new_n3849_), .Y(core__abc_21302_new_n3854_));
NAND2X1 NAND2X1_482 ( .A(core__abc_21302_new_n3778_), .B(core__abc_21302_new_n3774_), .Y(core__abc_21302_new_n3855_));
NAND2X1 NAND2X1_483 ( .A(core__abc_21302_new_n3859_), .B(core__abc_21302_new_n3860_), .Y(core__abc_21302_new_n3861_));
NAND2X1 NAND2X1_484 ( .A(core__abc_21302_new_n3863_), .B(core__abc_21302_new_n3767_), .Y(core__abc_21302_new_n3864_));
NAND2X1 NAND2X1_485 ( .A(core__abc_21302_new_n3857_), .B(core__abc_21302_new_n3864_), .Y(core__abc_21302_new_n3867_));
NAND2X1 NAND2X1_486 ( .A(core__abc_21302_new_n1937_), .B(core__abc_21302_new_n3881_), .Y(core__abc_21302_new_n3882_));
NAND2X1 NAND2X1_487 ( .A(core__abc_21302_new_n3879_), .B(core__abc_21302_new_n3881_), .Y(core__abc_21302_new_n3893_));
NAND2X1 NAND2X1_488 ( .A(core__abc_21302_new_n3886_), .B(core__abc_21302_new_n3889_), .Y(core__abc_21302_new_n3894_));
NAND2X1 NAND2X1_489 ( .A(core__abc_21302_new_n3895_), .B(core__abc_21302_new_n3891_), .Y(core__abc_21302_new_n3897_));
NAND2X1 NAND2X1_49 ( .A(core__abc_21302_new_n1264_), .B(core__abc_21302_new_n1263_), .Y(core__abc_21302_new_n1265_));
NAND2X1 NAND2X1_490 ( .A(core__abc_21302_new_n3898_), .B(core__abc_21302_new_n3896_), .Y(core__abc_21302_new_n3899_));
NAND2X1 NAND2X1_491 ( .A(core__abc_21302_new_n3853_), .B(core__abc_21302_new_n3895_), .Y(core__abc_21302_new_n3916_));
NAND2X1 NAND2X1_492 ( .A(core__abc_21302_new_n3891_), .B(core__abc_21302_new_n3916_), .Y(core__abc_21302_new_n3917_));
NAND2X1 NAND2X1_493 ( .A(core__abc_21302_new_n3914_), .B(core__abc_21302_new_n3919_), .Y(core__abc_21302_new_n3920_));
NAND2X1 NAND2X1_494 ( .A(core__abc_21302_new_n3924_), .B(core__abc_21302_new_n3922_), .Y(core__abc_21302_new_n3925_));
NAND2X1 NAND2X1_495 ( .A(core__abc_21302_new_n3930_), .B(core__abc_21302_new_n3932_), .Y(core__abc_21302_new_n3933_));
NAND2X1 NAND2X1_496 ( .A(core__abc_21302_new_n3059_), .B(core__abc_21302_new_n3933_), .Y(core__abc_21302_new_n3934_));
NAND2X1 NAND2X1_497 ( .A(core__abc_21302_new_n1210_), .B(core__abc_21302_new_n1223_), .Y(core__abc_21302_new_n3945_));
NAND2X1 NAND2X1_498 ( .A(core__abc_21302_new_n3946_), .B(core__abc_21302_new_n3945_), .Y(core__abc_21302_new_n3947_));
NAND2X1 NAND2X1_499 ( .A(core__abc_21302_new_n3949_), .B(core__abc_21302_new_n3950_), .Y(core__abc_21302_new_n3951_));
NAND2X1 NAND2X1_5 ( .A(\addr[1] ), .B(_abc_19873_new_n891_), .Y(_abc_19873_new_n892_));
NAND2X1 NAND2X1_50 ( .A(core_v1_reg_6_), .B(core_v0_reg_6_), .Y(core__abc_21302_new_n1274_));
NAND2X1 NAND2X1_500 ( .A(core__abc_21302_new_n1583_), .B(core__abc_21302_new_n3952_), .Y(core__abc_21302_new_n3953_));
NAND2X1 NAND2X1_501 ( .A(core__abc_21302_new_n3953_), .B(core__abc_21302_new_n3951_), .Y(core__abc_21302_new_n3954_));
NAND2X1 NAND2X1_502 ( .A(core__abc_21302_new_n3947_), .B(core__abc_21302_new_n3959_), .Y(core__abc_21302_new_n3960_));
NAND2X1 NAND2X1_503 ( .A(core__abc_21302_new_n3958_), .B(core__abc_21302_new_n3960_), .Y(core__abc_21302_new_n3961_));
NAND2X1 NAND2X1_504 ( .A(core__abc_21302_new_n1234_), .B(core__abc_21302_new_n2375_), .Y(core__abc_21302_new_n3976_));
NAND2X1 NAND2X1_505 ( .A(core__abc_21302_new_n3976_), .B(core__abc_21302_new_n3977_), .Y(core__abc_21302_new_n3978_));
NAND2X1 NAND2X1_506 ( .A(core__abc_21302_new_n3980_), .B(core__abc_21302_new_n3983_), .Y(core__abc_21302_new_n3984_));
NAND2X1 NAND2X1_507 ( .A(core__abc_21302_new_n3987_), .B(core__abc_21302_new_n3989_), .Y(core__abc_21302_new_n4001_));
NAND2X1 NAND2X1_508 ( .A(core__abc_21302_new_n3994_), .B(core__abc_21302_new_n3975_), .Y(core__abc_21302_new_n4002_));
NAND2X1 NAND2X1_509 ( .A(core__abc_21302_new_n1609_), .B(core__abc_21302_new_n4008_), .Y(core__abc_21302_new_n4009_));
NAND2X1 NAND2X1_51 ( .A(core__abc_21302_new_n1274_), .B(core__abc_21302_new_n1273_), .Y(core__abc_21302_new_n1275_));
NAND2X1 NAND2X1_510 ( .A(core__abc_21302_new_n4006_), .B(core__abc_21302_new_n4008_), .Y(core__abc_21302_new_n4012_));
NAND2X1 NAND2X1_511 ( .A(core__abc_21302_new_n4010_), .B(core__abc_21302_new_n4013_), .Y(core__abc_21302_new_n4014_));
NAND2X1 NAND2X1_512 ( .A(core__abc_21302_new_n4005_), .B(core__abc_21302_new_n4014_), .Y(core__abc_21302_new_n4015_));
NAND2X1 NAND2X1_513 ( .A(core__abc_21302_new_n4017_), .B(core__abc_21302_new_n4015_), .Y(core__abc_21302_new_n4018_));
NAND2X1 NAND2X1_514 ( .A(core__abc_21302_new_n4018_), .B(core__abc_21302_new_n4003_), .Y(core__abc_21302_new_n4020_));
NAND2X1 NAND2X1_515 ( .A(core__abc_21302_new_n4020_), .B(core__abc_21302_new_n4019_), .Y(core__abc_21302_new_n4021_));
NAND2X1 NAND2X1_516 ( .A(core__abc_21302_new_n2386_), .B(core__abc_21302_new_n2378_), .Y(core__abc_21302_new_n4041_));
NAND2X1 NAND2X1_517 ( .A(core__abc_21302_new_n1253_), .B(core__abc_21302_new_n2475_), .Y(core__abc_21302_new_n4042_));
NAND2X1 NAND2X1_518 ( .A(core__abc_21302_new_n4041_), .B(core__abc_21302_new_n4042_), .Y(core__abc_21302_new_n4043_));
NAND2X1 NAND2X1_519 ( .A(core_v3_reg_20_), .B(core__abc_21302_new_n4046_), .Y(core__abc_21302_new_n4047_));
NAND2X1 NAND2X1_52 ( .A(core_v1_reg_7_), .B(core_v0_reg_7_), .Y(core__abc_21302_new_n1284_));
NAND2X1 NAND2X1_520 ( .A(core__abc_21302_new_n1434_), .B(core__abc_21302_new_n4049_), .Y(core__abc_21302_new_n4050_));
NAND2X1 NAND2X1_521 ( .A(core__abc_21302_new_n4047_), .B(core__abc_21302_new_n4050_), .Y(core__abc_21302_new_n4052_));
NAND2X1 NAND2X1_522 ( .A(core__abc_21302_new_n4043_), .B(core__abc_21302_new_n4052_), .Y(core__abc_21302_new_n4053_));
NAND2X1 NAND2X1_523 ( .A(core__abc_21302_new_n4051_), .B(core__abc_21302_new_n4053_), .Y(core__abc_21302_new_n4054_));
NAND2X1 NAND2X1_524 ( .A(core__abc_21302_new_n4066_), .B(core__abc_21302_new_n4067_), .Y(core__abc_21302_new_n4068_));
NAND2X1 NAND2X1_525 ( .A(core__abc_21302_new_n4066_), .B(core__abc_21302_new_n4069_), .Y(core__abc_21302_new_n4073_));
NAND2X1 NAND2X1_526 ( .A(core__abc_21302_new_n4078_), .B(core__abc_21302_new_n4079_), .Y(core__abc_21302_new_n4081_));
NAND2X1 NAND2X1_527 ( .A(core__abc_21302_new_n4081_), .B(core__abc_21302_new_n4080_), .Y(core__abc_21302_new_n4083_));
NAND2X1 NAND2X1_528 ( .A(core__abc_21302_new_n3300_), .B(core__abc_21302_new_n4083_), .Y(core__abc_21302_new_n4084_));
NAND2X1 NAND2X1_529 ( .A(core__abc_21302_new_n4098_), .B(core__abc_21302_new_n4097_), .Y(core__abc_21302_new_n4099_));
NAND2X1 NAND2X1_53 ( .A(core__abc_21302_new_n1284_), .B(core__abc_21302_new_n1283_), .Y(core__abc_21302_new_n1285_));
NAND2X1 NAND2X1_530 ( .A(core__abc_21302_new_n4101_), .B(core__abc_21302_new_n4102_), .Y(core__abc_21302_new_n4103_));
NAND2X1 NAND2X1_531 ( .A(core_v3_reg_22_), .B(core__abc_21302_new_n4103_), .Y(core__abc_21302_new_n4104_));
NAND2X1 NAND2X1_532 ( .A(core__abc_21302_new_n1458_), .B(core__abc_21302_new_n4105_), .Y(core__abc_21302_new_n4106_));
NAND2X1 NAND2X1_533 ( .A(core__abc_21302_new_n1458_), .B(core__abc_21302_new_n4103_), .Y(core__abc_21302_new_n4109_));
NAND2X1 NAND2X1_534 ( .A(core_v3_reg_22_), .B(core__abc_21302_new_n4105_), .Y(core__abc_21302_new_n4110_));
NAND2X1 NAND2X1_535 ( .A(core__abc_21302_new_n4107_), .B(core__abc_21302_new_n4111_), .Y(core__abc_21302_new_n4112_));
NAND2X1 NAND2X1_536 ( .A(core__abc_21302_new_n4116_), .B(core__abc_21302_new_n4114_), .Y(core__abc_21302_new_n4117_));
NAND2X1 NAND2X1_537 ( .A(core__abc_21302_new_n3343_), .B(core__abc_21302_new_n4117_), .Y(core__abc_21302_new_n4118_));
NAND2X1 NAND2X1_538 ( .A(core__abc_21302_new_n2615_), .B(core__abc_21302_new_n4127_), .Y(core__abc_21302_new_n4132_));
NAND2X1 NAND2X1_539 ( .A(core__abc_21302_new_n4134_), .B(core__abc_21302_new_n4138_), .Y(core__abc_21302_new_n4139_));
NAND2X1 NAND2X1_54 ( .A(core_v2_reg_8_), .B(core_v3_reg_8_), .Y(core__abc_21302_new_n1294_));
NAND2X1 NAND2X1_540 ( .A(core_key_103_), .B(core__abc_21302_new_n2639__bF_buf1), .Y(core__abc_21302_new_n4147_));
NAND2X1 NAND2X1_541 ( .A(core__abc_21302_new_n4135_), .B(core__abc_21302_new_n4157_), .Y(core__abc_21302_new_n4158_));
NAND2X1 NAND2X1_542 ( .A(core__abc_21302_new_n4156_), .B(core__abc_21302_new_n4160_), .Y(core__abc_21302_new_n4161_));
NAND2X1 NAND2X1_543 ( .A(core__abc_21302_new_n4167_), .B(core__abc_21302_new_n4168_), .Y(core__abc_21302_new_n4169_));
NAND2X1 NAND2X1_544 ( .A(core__abc_21302_new_n2620_), .B(core__abc_21302_new_n2610_), .Y(core__abc_21302_new_n4174_));
NAND2X1 NAND2X1_545 ( .A(core__abc_21302_new_n4173_), .B(core__abc_21302_new_n4176_), .Y(core__abc_21302_new_n4178_));
NAND2X1 NAND2X1_546 ( .A(core__abc_21302_new_n4182_), .B(core__abc_21302_new_n4181_), .Y(core__abc_21302_new_n4183_));
NAND2X1 NAND2X1_547 ( .A(core__abc_21302_new_n4180_), .B(core__abc_21302_new_n4183_), .Y(core__abc_21302_new_n4184_));
NAND2X1 NAND2X1_548 ( .A(core__abc_21302_new_n1488_), .B(core__abc_21302_new_n4198_), .Y(core__abc_21302_new_n4199_));
NAND2X1 NAND2X1_549 ( .A(core_v3_reg_25_), .B(core__abc_21302_new_n4201_), .Y(core__abc_21302_new_n4202_));
NAND2X1 NAND2X1_55 ( .A(core__abc_21302_new_n1294_), .B(core__abc_21302_new_n1295_), .Y(core__abc_21302_new_n1296_));
NAND2X1 NAND2X1_550 ( .A(core__abc_21302_new_n4203_), .B(core__abc_21302_new_n4206_), .Y(core__abc_21302_new_n4207_));
NAND2X1 NAND2X1_551 ( .A(core__abc_21302_new_n3482_), .B(core__abc_21302_new_n4208_), .Y(core__abc_21302_new_n4209_));
NAND2X1 NAND2X1_552 ( .A(core__abc_21302_new_n4231_), .B(core__abc_21302_new_n4236_), .Y(core__abc_21302_new_n4237_));
NAND2X1 NAND2X1_553 ( .A(core__abc_21302_new_n1314_), .B(core__abc_21302_new_n4218_), .Y(core__abc_21302_new_n4250_));
NAND2X1 NAND2X1_554 ( .A(core__abc_21302_new_n2629_), .B(core__abc_21302_new_n2630_), .Y(core__abc_21302_new_n4255_));
NAND2X1 NAND2X1_555 ( .A(core__abc_21302_new_n1512_), .B(core__abc_21302_new_n4255_), .Y(core__abc_21302_new_n4256_));
NAND2X1 NAND2X1_556 ( .A(core__abc_21302_new_n4253_), .B(core__abc_21302_new_n4258_), .Y(core__abc_21302_new_n4259_));
NAND2X1 NAND2X1_557 ( .A(core__abc_21302_new_n4261_), .B(core__abc_21302_new_n4263_), .Y(core__abc_21302_new_n4264_));
NAND2X1 NAND2X1_558 ( .A(core__abc_21302_new_n4286_), .B(core__abc_21302_new_n2672_), .Y(core__abc_21302_new_n4287_));
NAND2X1 NAND2X1_559 ( .A(core__abc_21302_new_n4288_), .B(core__abc_21302_new_n4287_), .Y(core__abc_21302_new_n4289_));
NAND2X1 NAND2X1_56 ( .A(core_v2_reg_9_), .B(core_v3_reg_9_), .Y(core__abc_21302_new_n1304_));
NAND2X1 NAND2X1_560 ( .A(core_v3_reg_29_), .B(core__abc_21302_new_n2707_), .Y(core__abc_21302_new_n4301_));
NAND2X1 NAND2X1_561 ( .A(core__abc_21302_new_n1537_), .B(core__abc_21302_new_n2705_), .Y(core__abc_21302_new_n4302_));
NAND2X1 NAND2X1_562 ( .A(core__abc_21302_new_n1336_), .B(core__abc_21302_new_n4284_), .Y(core__abc_21302_new_n4303_));
NAND2X1 NAND2X1_563 ( .A(core__abc_21302_new_n2413_), .B(core__abc_21302_new_n4303_), .Y(core__abc_21302_new_n4304_));
NAND2X1 NAND2X1_564 ( .A(core__abc_21302_new_n4306_), .B(core__abc_21302_new_n4308_), .Y(core__abc_21302_new_n4309_));
NAND2X1 NAND2X1_565 ( .A(core__abc_21302_new_n4309_), .B(core__abc_21302_new_n4300_), .Y(core__abc_21302_new_n4311_));
NAND2X1 NAND2X1_566 ( .A(core__abc_21302_new_n4313_), .B(core__abc_21302_new_n4300_), .Y(core__abc_21302_new_n4315_));
NAND2X1 NAND2X1_567 ( .A(core__abc_21302_new_n4336_), .B(core__abc_21302_new_n4334_), .Y(core__abc_21302_new_n4337_));
NAND2X1 NAND2X1_568 ( .A(core__abc_21302_new_n4338_), .B(core__abc_21302_new_n4340_), .Y(core__abc_21302_new_n4341_));
NAND2X1 NAND2X1_569 ( .A(core__abc_21302_new_n3671_), .B(core__abc_21302_new_n4343_), .Y(core__abc_21302_new_n4344_));
NAND2X1 NAND2X1_57 ( .A(core__abc_21302_new_n1304_), .B(core__abc_21302_new_n1306_), .Y(core__abc_21302_new_n1307_));
NAND2X1 NAND2X1_570 ( .A(core__abc_21302_new_n4364_), .B(core__abc_21302_new_n4366_), .Y(core__abc_21302_new_n4367_));
NAND2X1 NAND2X1_571 ( .A(core_key_111_), .B(core__abc_21302_new_n2639__bF_buf6), .Y(core__abc_21302_new_n4379_));
NAND2X1 NAND2X1_572 ( .A(core__abc_21302_new_n4323_), .B(core__abc_21302_new_n4386_), .Y(core__abc_21302_new_n4389_));
NAND2X1 NAND2X1_573 ( .A(core__abc_21302_new_n4365_), .B(core__abc_21302_new_n2789_), .Y(core__abc_21302_new_n4391_));
NAND2X1 NAND2X1_574 ( .A(core__abc_21302_new_n4398_), .B(core__abc_21302_new_n2830_), .Y(core__abc_21302_new_n4401_));
NAND2X1 NAND2X1_575 ( .A(core__abc_21302_new_n4401_), .B(core__abc_21302_new_n4400_), .Y(core__abc_21302_new_n4402_));
NAND2X1 NAND2X1_576 ( .A(core__abc_21302_new_n4413_), .B(core__abc_21302_new_n2871_), .Y(core__abc_21302_new_n4414_));
NAND2X1 NAND2X1_577 ( .A(core__abc_21302_new_n4277_), .B(core__abc_21302_new_n4387_), .Y(core__abc_21302_new_n4428_));
NAND2X1 NAND2X1_578 ( .A(core__abc_21302_new_n4448_), .B(core__abc_21302_new_n4446_), .Y(core__abc_21302_new_n4449_));
NAND2X1 NAND2X1_579 ( .A(core__abc_21302_new_n4449_), .B(core__abc_21302_new_n2906_), .Y(core__abc_21302_new_n4452_));
NAND2X1 NAND2X1_58 ( .A(core_v2_reg_10_), .B(core_v3_reg_10_), .Y(core__abc_21302_new_n1315_));
NAND2X1 NAND2X1_580 ( .A(core__abc_21302_new_n4454_), .B(core__abc_21302_new_n4459_), .Y(core__abc_21302_new_n4460_));
NAND2X1 NAND2X1_581 ( .A(core__abc_21302_new_n4456_), .B(core__abc_21302_new_n4460_), .Y(core__abc_21302_new_n4461_));
NAND2X1 NAND2X1_582 ( .A(core__abc_21302_new_n3816_), .B(core__abc_21302_new_n4461_), .Y(core__abc_21302_new_n4462_));
NAND2X1 NAND2X1_583 ( .A(core__abc_21302_new_n1419_), .B(core__abc_21302_new_n4470_), .Y(core__abc_21302_new_n4473_));
NAND2X1 NAND2X1_584 ( .A(core__abc_21302_new_n4473_), .B(core__abc_21302_new_n4472_), .Y(core__abc_21302_new_n4474_));
NAND2X1 NAND2X1_585 ( .A(core__abc_21302_new_n4481_), .B(core__abc_21302_new_n4479_), .Y(core__abc_21302_new_n4482_));
NAND2X1 NAND2X1_586 ( .A(core__abc_21302_new_n3848_), .B(core__abc_21302_new_n4482_), .Y(core__abc_21302_new_n4483_));
NAND2X1 NAND2X1_587 ( .A(core__abc_21302_new_n4501_), .B(core__abc_21302_new_n4503_), .Y(core__abc_21302_new_n4504_));
NAND2X1 NAND2X1_588 ( .A(core__abc_21302_new_n4504_), .B(core__abc_21302_new_n2991_), .Y(core__abc_21302_new_n4506_));
NAND2X1 NAND2X1_589 ( .A(core__abc_21302_new_n4506_), .B(core__abc_21302_new_n4505_), .Y(core__abc_21302_new_n4507_));
NAND2X1 NAND2X1_59 ( .A(core__abc_21302_new_n1316_), .B(core__abc_21302_new_n1317_), .Y(core__abc_21302_new_n1318_));
NAND2X1 NAND2X1_590 ( .A(core__abc_21302_new_n4518_), .B(core__abc_21302_new_n4520_), .Y(core__abc_21302_new_n4521_));
NAND2X1 NAND2X1_591 ( .A(core__abc_21302_new_n4526_), .B(core__abc_21302_new_n4528_), .Y(core__abc_21302_new_n4531_));
NAND2X1 NAND2X1_592 ( .A(core__abc_21302_new_n4530_), .B(core__abc_21302_new_n4531_), .Y(core__abc_21302_new_n4532_));
NAND2X1 NAND2X1_593 ( .A(core__abc_21302_new_n4521_), .B(core__abc_21302_new_n3034_), .Y(core__abc_21302_new_n4541_));
NAND2X1 NAND2X1_594 ( .A(core__abc_21302_new_n1455_), .B(core__abc_21302_new_n4544_), .Y(core__abc_21302_new_n4545_));
NAND2X1 NAND2X1_595 ( .A(core__abc_21302_new_n4549_), .B(core__abc_21302_new_n4550_), .Y(core__abc_21302_new_n4551_));
NAND2X1 NAND2X1_596 ( .A(core__abc_21302_new_n3959_), .B(core__abc_21302_new_n4556_), .Y(core__abc_21302_new_n4557_));
NAND2X1 NAND2X1_597 ( .A(core__abc_21302_new_n4543_), .B(core__abc_21302_new_n4540_), .Y(core__abc_21302_new_n4565_));
NAND2X1 NAND2X1_598 ( .A(core__abc_21302_new_n4566_), .B(core__abc_21302_new_n4565_), .Y(core__abc_21302_new_n4567_));
NAND2X1 NAND2X1_599 ( .A(core__abc_21302_new_n4570_), .B(core__abc_21302_new_n4572_), .Y(core__abc_21302_new_n4573_));
NAND2X1 NAND2X1_6 ( .A(_abc_19873_new_n889__bF_buf4), .B(_abc_19873_new_n893__bF_buf4), .Y(_abc_19873_new_n894_));
NAND2X1 NAND2X1_60 ( .A(core__abc_21302_new_n1315_), .B(core__abc_21302_new_n1318_), .Y(core__abc_21302_new_n1319_));
NAND2X1 NAND2X1_600 ( .A(core__abc_21302_new_n4576_), .B(core__abc_21302_new_n4574_), .Y(core__abc_21302_new_n4577_));
NAND2X1 NAND2X1_601 ( .A(core_key_119_), .B(core__abc_21302_new_n2639__bF_buf4), .Y(core__abc_21302_new_n4587_));
NAND2X1 NAND2X1_602 ( .A(core__abc_21302_new_n4601_), .B(core__abc_21302_new_n4598_), .Y(core__abc_21302_new_n4602_));
NAND2X1 NAND2X1_603 ( .A(core__abc_21302_new_n1475_), .B(core__abc_21302_new_n4604_), .Y(core__abc_21302_new_n4605_));
NAND2X1 NAND2X1_604 ( .A(core__abc_21302_new_n4607_), .B(core__abc_21302_new_n4605_), .Y(core__abc_21302_new_n4608_));
NAND2X1 NAND2X1_605 ( .A(core__abc_21302_new_n3212_), .B(core__abc_21302_new_n3210_), .Y(core__abc_21302_new_n4621_));
NAND2X1 NAND2X1_606 ( .A(core_v3_reg_41_), .B(core__abc_21302_new_n3213_), .Y(core__abc_21302_new_n4622_));
NAND2X1 NAND2X1_607 ( .A(core__abc_21302_new_n4628_), .B(core__abc_21302_new_n4620_), .Y(core__abc_21302_new_n4630_));
NAND2X1 NAND2X1_608 ( .A(core_key_121_), .B(core__abc_21302_new_n2639__bF_buf2), .Y(core__abc_21302_new_n4636_));
NAND2X1 NAND2X1_609 ( .A(core__abc_21302_new_n4074_), .B(core__abc_21302_new_n4071_), .Y(core__abc_21302_new_n4642_));
NAND2X1 NAND2X1_61 ( .A(core_v2_reg_11_), .B(core_v3_reg_11_), .Y(core__abc_21302_new_n1327_));
NAND2X1 NAND2X1_610 ( .A(core__abc_21302_new_n4624_), .B(core__abc_21302_new_n3215_), .Y(core__abc_21302_new_n4643_));
NAND2X1 NAND2X1_611 ( .A(core__abc_21302_new_n4643_), .B(core__abc_21302_new_n4645_), .Y(core__abc_21302_new_n4646_));
NAND2X1 NAND2X1_612 ( .A(core__abc_21302_new_n4661_), .B(core__abc_21302_new_n4660_), .Y(core__abc_21302_new_n4662_));
NAND2X1 NAND2X1_613 ( .A(core__abc_21302_new_n4642_), .B(core__abc_21302_new_n4662_), .Y(core__abc_21302_new_n4663_));
NAND2X1 NAND2X1_614 ( .A(core__abc_21302_new_n4110_), .B(core__abc_21302_new_n4109_), .Y(core__abc_21302_new_n4671_));
NAND2X1 NAND2X1_615 ( .A(core__abc_21302_new_n4675_), .B(core__abc_21302_new_n4677_), .Y(core__abc_21302_new_n4678_));
NAND2X1 NAND2X1_616 ( .A(core__abc_21302_new_n4680_), .B(core__abc_21302_new_n4681_), .Y(core__abc_21302_new_n4682_));
NAND2X1 NAND2X1_617 ( .A(core__abc_21302_new_n4687_), .B(core__abc_21302_new_n4689_), .Y(core__abc_21302_new_n4690_));
NAND2X1 NAND2X1_618 ( .A(core__abc_21302_new_n2426_), .B(core__abc_21302_new_n4604_), .Y(core__abc_21302_new_n4707_));
NAND2X1 NAND2X1_619 ( .A(core__abc_21302_new_n4706_), .B(core__abc_21302_new_n4707_), .Y(core__abc_21302_new_n4708_));
NAND2X1 NAND2X1_62 ( .A(core__abc_21302_new_n1328_), .B(core__abc_21302_new_n1329_), .Y(core__abc_21302_new_n1330_));
NAND2X1 NAND2X1_620 ( .A(core__abc_21302_new_n1521_), .B(core__abc_21302_new_n4708_), .Y(core__abc_21302_new_n4709_));
NAND2X1 NAND2X1_621 ( .A(core__abc_21302_new_n2703_), .B(core__abc_21302_new_n3358_), .Y(core__abc_21302_new_n4715_));
NAND2X1 NAND2X1_622 ( .A(core__abc_21302_new_n4717_), .B(core__abc_21302_new_n4713_), .Y(core__abc_21302_new_n4718_));
NAND2X1 NAND2X1_623 ( .A(core__abc_21302_new_n4157_), .B(core__abc_21302_new_n4723_), .Y(core__abc_21302_new_n4724_));
NAND2X1 NAND2X1_624 ( .A(core__abc_21302_new_n4741_), .B(core__abc_21302_new_n4743_), .Y(core__abc_21302_new_n4744_));
NAND2X1 NAND2X1_625 ( .A(core__abc_21302_new_n4778_), .B(core__abc_21302_new_n4776_), .Y(core__abc_21302_new_n4779_));
NAND2X1 NAND2X1_626 ( .A(core__abc_21302_new_n4226_), .B(core__abc_21302_new_n4224_), .Y(core__abc_21302_new_n4795_));
NAND2X1 NAND2X1_627 ( .A(core__abc_21302_new_n4799_), .B(core__abc_21302_new_n4801_), .Y(core__abc_21302_new_n4802_));
NAND2X1 NAND2X1_628 ( .A(core__abc_21302_new_n4802_), .B(core__abc_21302_new_n3491_), .Y(core__abc_21302_new_n4803_));
NAND2X1 NAND2X1_629 ( .A(core__abc_21302_new_n4803_), .B(core__abc_21302_new_n4805_), .Y(core__abc_21302_new_n4806_));
NAND2X1 NAND2X1_63 ( .A(core__abc_21302_new_n1327_), .B(core__abc_21302_new_n1330_), .Y(core__abc_21302_new_n1331_));
NAND2X1 NAND2X1_630 ( .A(core__abc_21302_new_n3884_), .B(core__abc_21302_new_n3885_), .Y(core__abc_21302_new_n4823_));
NAND2X1 NAND2X1_631 ( .A(core__abc_21302_new_n4823_), .B(core__abc_21302_new_n4828_), .Y(core__abc_21302_new_n4829_));
NAND2X1 NAND2X1_632 ( .A(core__abc_21302_new_n4835_), .B(core__abc_21302_new_n4834_), .Y(core__abc_21302_new_n4836_));
NAND2X1 NAND2X1_633 ( .A(core__abc_21302_new_n3809_), .B(core__abc_21302_new_n3811_), .Y(core__abc_21302_new_n4839_));
NAND2X1 NAND2X1_634 ( .A(core_v1_reg_16_), .B(core__abc_21302_new_n4744_), .Y(core__abc_21302_new_n4842_));
NAND2X1 NAND2X1_635 ( .A(core_v1_reg_15_), .B(core__abc_21302_new_n4712_), .Y(core__abc_21302_new_n4849_));
NAND2X1 NAND2X1_636 ( .A(core__abc_21302_new_n4848_), .B(core__abc_21302_new_n4849_), .Y(core__abc_21302_new_n4850_));
NAND2X1 NAND2X1_637 ( .A(core__abc_21302_new_n3735_), .B(core__abc_21302_new_n3737_), .Y(core__abc_21302_new_n4854_));
NAND2X1 NAND2X1_638 ( .A(core__abc_21302_new_n4854_), .B(core__abc_21302_new_n4857_), .Y(core__abc_21302_new_n4858_));
NAND2X1 NAND2X1_639 ( .A(core__abc_21302_new_n3708_), .B(core__abc_21302_new_n4862_), .Y(core__abc_21302_new_n4863_));
NAND2X1 NAND2X1_64 ( .A(core_v2_reg_12_), .B(core_v3_reg_12_), .Y(core__abc_21302_new_n1337_));
NAND2X1 NAND2X1_640 ( .A(core__abc_21302_new_n4866_), .B(core__abc_21302_new_n4861_), .Y(core__abc_21302_new_n4867_));
NAND2X1 NAND2X1_641 ( .A(core__abc_21302_new_n3667_), .B(core__abc_21302_new_n4869_), .Y(core__abc_21302_new_n4870_));
NAND2X1 NAND2X1_642 ( .A(core__abc_21302_new_n4870_), .B(core__abc_21302_new_n4874_), .Y(core__abc_21302_new_n4875_));
NAND2X1 NAND2X1_643 ( .A(core__abc_21302_new_n4863_), .B(core__abc_21302_new_n4858_), .Y(core__abc_21302_new_n4876_));
NAND2X1 NAND2X1_644 ( .A(core__abc_21302_new_n3638_), .B(core__abc_21302_new_n4872_), .Y(core__abc_21302_new_n4891_));
NAND2X1 NAND2X1_645 ( .A(core__abc_21302_new_n4891_), .B(core__abc_21302_new_n4873_), .Y(core__abc_21302_new_n4892_));
NAND2X1 NAND2X1_646 ( .A(core__abc_21302_new_n3580_), .B(core__abc_21302_new_n3581_), .Y(core__abc_21302_new_n4895_));
NAND2X1 NAND2X1_647 ( .A(core_v1_reg_8_), .B(core__abc_21302_new_n4521_), .Y(core__abc_21302_new_n4919_));
NAND2X1 NAND2X1_648 ( .A(core__abc_21302_new_n3422_), .B(core__abc_21302_new_n3421_), .Y(core__abc_21302_new_n4932_));
NAND2X1 NAND2X1_649 ( .A(core__abc_21302_new_n4933_), .B(core__abc_21302_new_n4474_), .Y(core__abc_21302_new_n4934_));
NAND2X1 NAND2X1_65 ( .A(core__abc_21302_new_n1338_), .B(core__abc_21302_new_n1339_), .Y(core__abc_21302_new_n1340_));
NAND2X1 NAND2X1_650 ( .A(core__abc_21302_new_n4937_), .B(core__abc_21302_new_n4940_), .Y(core__abc_21302_new_n4941_));
NAND2X1 NAND2X1_651 ( .A(core__abc_21302_new_n4931_), .B(core__abc_21302_new_n4941_), .Y(core__abc_21302_new_n4942_));
NAND2X1 NAND2X1_652 ( .A(core__abc_21302_new_n2471_), .B(core__abc_21302_new_n4365_), .Y(core__abc_21302_new_n4964_));
NAND2X1 NAND2X1_653 ( .A(core_v1_reg_2_), .B(core__abc_21302_new_n4363_), .Y(core__abc_21302_new_n4965_));
NAND2X1 NAND2X1_654 ( .A(core__abc_21302_new_n4964_), .B(core__abc_21302_new_n4965_), .Y(core__abc_21302_new_n4967_));
NAND2X1 NAND2X1_655 ( .A(core__abc_21302_new_n3230_), .B(core__abc_21302_new_n4967_), .Y(core__abc_21302_new_n4968_));
NAND2X1 NAND2X1_656 ( .A(core__abc_21302_new_n3107_), .B(core__abc_21302_new_n4980_), .Y(core__abc_21302_new_n4981_));
NAND2X1 NAND2X1_657 ( .A(core__abc_21302_new_n3141_), .B(core__abc_21302_new_n4977_), .Y(core__abc_21302_new_n4988_));
NAND2X1 NAND2X1_658 ( .A(core__abc_21302_new_n3143_), .B(core__abc_21302_new_n4976_), .Y(core__abc_21302_new_n4989_));
NAND2X1 NAND2X1_659 ( .A(core__abc_21302_new_n4988_), .B(core__abc_21302_new_n4989_), .Y(core__abc_21302_new_n4990_));
NAND2X1 NAND2X1_66 ( .A(core_v2_reg_13_), .B(core_v3_reg_13_), .Y(core__abc_21302_new_n1349_));
NAND2X1 NAND2X1_660 ( .A(core__abc_21302_new_n4991_), .B(core__abc_21302_new_n4981_), .Y(core__abc_21302_new_n4992_));
NAND2X1 NAND2X1_661 ( .A(core__abc_21302_new_n4996_), .B(core__abc_21302_new_n4257_), .Y(core__abc_21302_new_n4997_));
NAND2X1 NAND2X1_662 ( .A(core_v1_reg_62_), .B(core__abc_21302_new_n4252_), .Y(core__abc_21302_new_n4998_));
NAND2X1 NAND2X1_663 ( .A(core__abc_21302_new_n4999_), .B(core__abc_21302_new_n4995_), .Y(core__abc_21302_new_n5000_));
NAND2X1 NAND2X1_664 ( .A(core__abc_21302_new_n4997_), .B(core__abc_21302_new_n4998_), .Y(core__abc_21302_new_n5003_));
NAND2X1 NAND2X1_665 ( .A(core__abc_21302_new_n3053_), .B(core__abc_21302_new_n5003_), .Y(core__abc_21302_new_n5004_));
NAND2X1 NAND2X1_666 ( .A(core__abc_21302_new_n5004_), .B(core__abc_21302_new_n5000_), .Y(core__abc_21302_new_n5005_));
NAND2X1 NAND2X1_667 ( .A(core__abc_21302_new_n3018_), .B(core__abc_21302_new_n5001_), .Y(core__abc_21302_new_n5007_));
NAND2X1 NAND2X1_668 ( .A(core__abc_21302_new_n5007_), .B(core__abc_21302_new_n5002_), .Y(core__abc_21302_new_n5008_));
NAND2X1 NAND2X1_669 ( .A(core__abc_21302_new_n2970_), .B(core__abc_21302_new_n5010_), .Y(core__abc_21302_new_n5011_));
NAND2X1 NAND2X1_67 ( .A(core__abc_21302_new_n1350_), .B(core__abc_21302_new_n1351_), .Y(core__abc_21302_new_n1352_));
NAND2X1 NAND2X1_670 ( .A(core__abc_21302_new_n2939_), .B(core__abc_21302_new_n5012_), .Y(core__abc_21302_new_n5013_));
NAND2X1 NAND2X1_671 ( .A(core__abc_21302_new_n2885_), .B(core__abc_21302_new_n5019_), .Y(core__abc_21302_new_n5020_));
NAND2X1 NAND2X1_672 ( .A(core__abc_21302_new_n2806_), .B(core__abc_21302_new_n5030_), .Y(core__abc_21302_new_n5032_));
NAND2X1 NAND2X1_673 ( .A(core__abc_21302_new_n2744_), .B(core__abc_21302_new_n5037_), .Y(core__abc_21302_new_n5038_));
NAND2X1 NAND2X1_674 ( .A(core_v1_reg_52_), .B(core__abc_21302_new_n3947_), .Y(core__abc_21302_new_n5043_));
NAND2X1 NAND2X1_675 ( .A(core__abc_21302_new_n1794_), .B(core__abc_21302_new_n3948_), .Y(core__abc_21302_new_n5044_));
NAND2X1 NAND2X1_676 ( .A(core__abc_21302_new_n2692_), .B(core__abc_21302_new_n5041_), .Y(core__abc_21302_new_n5051_));
NAND2X1 NAND2X1_677 ( .A(core__abc_21302_new_n5051_), .B(core__abc_21302_new_n5042_), .Y(core__abc_21302_new_n5052_));
NAND2X1 NAND2X1_678 ( .A(core__abc_21302_new_n2773_), .B(core__abc_21302_new_n5035_), .Y(core__abc_21302_new_n5055_));
NAND2X1 NAND2X1_679 ( .A(core__abc_21302_new_n5055_), .B(core__abc_21302_new_n5036_), .Y(core__abc_21302_new_n5056_));
NAND2X1 NAND2X1_68 ( .A(core_v2_reg_14_), .B(core_v3_reg_14_), .Y(core__abc_21302_new_n1361_));
NAND2X1 NAND2X1_680 ( .A(core__abc_21302_new_n5013_), .B(core__abc_21302_new_n5060_), .Y(core__abc_21302_new_n5061_));
NAND2X1 NAND2X1_681 ( .A(core__abc_21302_new_n3299_), .B(core__abc_21302_new_n4946_), .Y(core__abc_21302_new_n5066_));
NAND2X1 NAND2X1_682 ( .A(core__abc_21302_new_n5066_), .B(core__abc_21302_new_n4947_), .Y(core__abc_21302_new_n5067_));
NAND2X1 NAND2X1_683 ( .A(core__abc_21302_new_n3925_), .B(core__abc_21302_new_n5074_), .Y(core__abc_21302_new_n5076_));
NAND2X1 NAND2X1_684 ( .A(core__abc_21302_new_n2634__bF_buf5), .B(core__abc_21302_new_n5079_), .Y(core__abc_21302_new_n5080_));
NAND2X1 NAND2X1_685 ( .A(core_v2_reg_0_), .B(core__abc_21302_new_n5085__bF_buf5), .Y(core__abc_21302_new_n5086_));
NAND2X1 NAND2X1_686 ( .A(core__abc_21302_new_n2649_), .B(core__abc_21302_new_n2650_), .Y(core__abc_21302_new_n5088_));
NAND2X1 NAND2X1_687 ( .A(core__abc_21302_new_n5071_), .B(core__abc_21302_new_n4963_), .Y(core__abc_21302_new_n5093_));
NAND2X1 NAND2X1_688 ( .A(core__abc_21302_new_n5092_), .B(core__abc_21302_new_n5093_), .Y(core__abc_21302_new_n5094_));
NAND2X1 NAND2X1_689 ( .A(core_key_1_), .B(core__abc_21302_new_n2639__bF_buf1), .Y(core__abc_21302_new_n5099_));
NAND2X1 NAND2X1_69 ( .A(core__abc_21302_new_n1362_), .B(core__abc_21302_new_n1363_), .Y(core__abc_21302_new_n1364_));
NAND2X1 NAND2X1_690 ( .A(core_v2_reg_1_), .B(core__abc_21302_new_n5085__bF_buf4), .Y(core__abc_21302_new_n5102_));
NAND2X1 NAND2X1_691 ( .A(core__abc_21302_new_n5077_), .B(core__abc_21302_new_n5090_), .Y(core__abc_21302_new_n5105_));
NAND2X1 NAND2X1_692 ( .A(core__abc_21302_new_n5121_), .B(core__abc_21302_new_n5123_), .Y(core__abc_21302_new_n5124_));
NAND2X1 NAND2X1_693 ( .A(core_key_2_), .B(core__abc_21302_new_n2639__bF_buf0), .Y(core__abc_21302_new_n5126_));
NAND2X1 NAND2X1_694 ( .A(core__abc_21302_new_n5114_), .B(core__abc_21302_new_n5118_), .Y(core__abc_21302_new_n5133_));
NAND2X1 NAND2X1_695 ( .A(core__abc_21302_new_n4007_), .B(core__abc_21302_new_n4009_), .Y(core__abc_21302_new_n5135_));
NAND2X1 NAND2X1_696 ( .A(core__abc_21302_new_n5136_), .B(core__abc_21302_new_n2739_), .Y(core__abc_21302_new_n5137_));
NAND2X1 NAND2X1_697 ( .A(core__abc_21302_new_n5139_), .B(core__abc_21302_new_n5143_), .Y(core__abc_21302_new_n5144_));
NAND2X1 NAND2X1_698 ( .A(core__abc_21302_new_n2634__bF_buf4), .B(core__abc_21302_new_n5145_), .Y(core__abc_21302_new_n5146_));
NAND2X1 NAND2X1_699 ( .A(core_v2_reg_3_), .B(core__abc_21302_new_n5085__bF_buf2), .Y(core__abc_21302_new_n5149_));
NAND2X1 NAND2X1_7 ( .A(_abc_19873_new_n889__bF_buf3), .B(_abc_19873_new_n895__bF_buf4), .Y(_abc_19873_new_n896_));
NAND2X1 NAND2X1_70 ( .A(core_v2_reg_16_), .B(core_v3_reg_16_), .Y(core__abc_21302_new_n1385_));
NAND2X1 NAND2X1_700 ( .A(core__abc_21302_new_n4049_), .B(core__abc_21302_new_n5151_), .Y(core__abc_21302_new_n5152_));
NAND2X1 NAND2X1_701 ( .A(core__abc_21302_new_n5152_), .B(core__abc_21302_new_n5153_), .Y(core__abc_21302_new_n5154_));
NAND2X1 NAND2X1_702 ( .A(core__abc_21302_new_n5161_), .B(core__abc_21302_new_n5073_), .Y(core__abc_21302_new_n5162_));
NAND2X1 NAND2X1_703 ( .A(core__abc_21302_new_n5177_), .B(core__abc_21302_new_n5179_), .Y(core__abc_21302_new_n5180_));
NAND2X1 NAND2X1_704 ( .A(core_v2_reg_5_), .B(core__abc_21302_new_n5085__bF_buf0), .Y(core__abc_21302_new_n5185_));
NAND2X1 NAND2X1_705 ( .A(core__abc_21302_new_n4103_), .B(core__abc_21302_new_n5188_), .Y(core__abc_21302_new_n5189_));
NAND2X1 NAND2X1_706 ( .A(core__abc_21302_new_n4105_), .B(core__abc_21302_new_n5190_), .Y(core__abc_21302_new_n5191_));
NAND2X1 NAND2X1_707 ( .A(core__abc_21302_new_n5189_), .B(core__abc_21302_new_n5191_), .Y(core__abc_21302_new_n5192_));
NAND2X1 NAND2X1_708 ( .A(core__abc_21302_new_n5192_), .B(core__abc_21302_new_n5195_), .Y(core__abc_21302_new_n5198_));
NAND2X1 NAND2X1_709 ( .A(core__abc_21302_new_n2634__bF_buf3), .B(core__abc_21302_new_n5199_), .Y(core__abc_21302_new_n5200_));
NAND2X1 NAND2X1_71 ( .A(core_v2_reg_17_), .B(core_v3_reg_17_), .Y(core__abc_21302_new_n1396_));
NAND2X1 NAND2X1_710 ( .A(core_v2_reg_6_), .B(core__abc_21302_new_n5085__bF_buf5), .Y(core__abc_21302_new_n5203_));
NAND2X1 NAND2X1_711 ( .A(core__abc_21302_new_n4132_), .B(core__abc_21302_new_n4131_), .Y(core__abc_21302_new_n5207_));
NAND2X1 NAND2X1_712 ( .A(core__abc_21302_new_n5210_), .B(core__abc_21302_new_n2881_), .Y(core__abc_21302_new_n5213_));
NAND2X1 NAND2X1_713 ( .A(core_v1_reg_26_), .B(core__abc_21302_new_n2890_), .Y(core__abc_21302_new_n5214_));
NAND2X1 NAND2X1_714 ( .A(core__abc_21302_new_n5215_), .B(core__abc_21302_new_n5212_), .Y(core__abc_21302_new_n5216_));
NAND2X1 NAND2X1_715 ( .A(core__abc_21302_new_n5216_), .B(core__abc_21302_new_n5206_), .Y(core__abc_21302_new_n5217_));
NAND2X1 NAND2X1_716 ( .A(core_v2_reg_7_), .B(core__abc_21302_new_n5085__bF_buf4), .Y(core__abc_21302_new_n5224_));
NAND2X1 NAND2X1_717 ( .A(core__abc_21302_new_n5214_), .B(core__abc_21302_new_n5213_), .Y(core__abc_21302_new_n5231_));
NAND2X1 NAND2X1_718 ( .A(core__abc_21302_new_n5229_), .B(core__abc_21302_new_n5233_), .Y(core__abc_21302_new_n5234_));
NAND2X1 NAND2X1_719 ( .A(core__abc_21302_new_n5236_), .B(core__abc_21302_new_n5237_), .Y(core__abc_21302_new_n5238_));
NAND2X1 NAND2X1_72 ( .A(core__abc_21302_new_n1397_), .B(core__abc_21302_new_n1398_), .Y(core__abc_21302_new_n1399_));
NAND2X1 NAND2X1_720 ( .A(core__abc_21302_new_n5238_), .B(core__abc_21302_new_n5240_), .Y(core__abc_21302_new_n5241_));
NAND2X1 NAND2X1_721 ( .A(core__abc_21302_new_n5243_), .B(core__abc_21302_new_n5104__bF_buf6), .Y(core__abc_21302_new_n5244_));
NAND2X1 NAND2X1_722 ( .A(core__abc_21302_new_n5248_), .B(core__abc_21302_new_n2973_), .Y(core__abc_21302_new_n5249_));
NAND2X1 NAND2X1_723 ( .A(core_v1_reg_28_), .B(core__abc_21302_new_n2968_), .Y(core__abc_21302_new_n5250_));
NAND2X1 NAND2X1_724 ( .A(core__abc_21302_new_n5250_), .B(core__abc_21302_new_n5249_), .Y(core__abc_21302_new_n5252_));
NAND2X1 NAND2X1_725 ( .A(core__abc_21302_new_n4198_), .B(core__abc_21302_new_n5252_), .Y(core__abc_21302_new_n5253_));
NAND2X1 NAND2X1_726 ( .A(core__abc_21302_new_n5251_), .B(core__abc_21302_new_n5253_), .Y(core__abc_21302_new_n5254_));
NAND2X1 NAND2X1_727 ( .A(core__abc_21302_new_n2362__bF_buf9), .B(core__abc_21302_new_n5258_), .Y(core__abc_21302_new_n5259_));
NAND2X1 NAND2X1_728 ( .A(core__abc_21302_new_n2624_), .B(core__abc_21302_new_n4225_), .Y(core__abc_21302_new_n5267_));
NAND2X1 NAND2X1_729 ( .A(core_v1_reg_29_), .B(core__abc_21302_new_n3021_), .Y(core__abc_21302_new_n5270_));
NAND2X1 NAND2X1_73 ( .A(core__abc_21302_new_n1396_), .B(core__abc_21302_new_n1399_), .Y(core__abc_21302_new_n1400_));
NAND2X1 NAND2X1_730 ( .A(core__abc_21302_new_n5269_), .B(core__abc_21302_new_n5270_), .Y(core__abc_21302_new_n5271_));
NAND2X1 NAND2X1_731 ( .A(core__abc_21302_new_n5275_), .B(core__abc_21302_new_n5277_), .Y(core__abc_21302_new_n5278_));
NAND2X1 NAND2X1_732 ( .A(core__abc_21302_new_n5280_), .B(core__abc_21302_new_n5104__bF_buf2), .Y(core__abc_21302_new_n5281_));
NAND2X1 NAND2X1_733 ( .A(core_v1_reg_30_), .B(core__abc_21302_new_n3058_), .Y(core__abc_21302_new_n5288_));
NAND2X1 NAND2X1_734 ( .A(core__abc_21302_new_n5293_), .B(core__abc_21302_new_n5285_), .Y(core__abc_21302_new_n5295_));
NAND2X1 NAND2X1_735 ( .A(core__abc_21302_new_n5295_), .B(core__abc_21302_new_n5294_), .Y(core__abc_21302_new_n5296_));
NAND2X1 NAND2X1_736 ( .A(core__abc_21302_new_n2668_), .B(core__abc_21302_new_n5312_), .Y(core__abc_21302_new_n5314_));
NAND2X1 NAND2X1_737 ( .A(core__abc_21302_new_n5314_), .B(core__abc_21302_new_n5313_), .Y(core__abc_21302_new_n5315_));
NAND2X1 NAND2X1_738 ( .A(core__abc_21302_new_n2362__bF_buf8), .B(core__abc_21302_new_n5318_), .Y(core__abc_21302_new_n5319_));
NAND2X1 NAND2X1_739 ( .A(core__abc_21302_new_n5322_), .B(core__abc_21302_new_n5310_), .Y(core__abc_21302_new_n5323_));
NAND2X1 NAND2X1_74 ( .A(core_v2_reg_18_), .B(core_v3_reg_18_), .Y(core__abc_21302_new_n1408_));
NAND2X1 NAND2X1_740 ( .A(core__abc_21302_new_n5325_), .B(core__abc_21302_new_n3136_), .Y(core__abc_21302_new_n5326_));
NAND2X1 NAND2X1_741 ( .A(core_v1_reg_32_), .B(core__abc_21302_new_n3269_), .Y(core__abc_21302_new_n5327_));
NAND2X1 NAND2X1_742 ( .A(core__abc_21302_new_n5327_), .B(core__abc_21302_new_n5326_), .Y(core__abc_21302_new_n5328_));
NAND2X1 NAND2X1_743 ( .A(core__abc_21302_new_n2705_), .B(core__abc_21302_new_n5328_), .Y(core__abc_21302_new_n5329_));
NAND2X1 NAND2X1_744 ( .A(core__abc_21302_new_n2707_), .B(core__abc_21302_new_n5330_), .Y(core__abc_21302_new_n5331_));
NAND2X1 NAND2X1_745 ( .A(core__abc_21302_new_n5329_), .B(core__abc_21302_new_n5331_), .Y(core__abc_21302_new_n5332_));
NAND2X1 NAND2X1_746 ( .A(core__abc_21302_new_n5333_), .B(core__abc_21302_new_n5324_), .Y(core__abc_21302_new_n5334_));
NAND2X1 NAND2X1_747 ( .A(core__abc_21302_new_n5334_), .B(core__abc_21302_new_n5335_), .Y(core__abc_21302_new_n5336_));
NAND2X1 NAND2X1_748 ( .A(core__abc_21302_new_n2634__bF_buf7), .B(core__abc_21302_new_n5336_), .Y(core__abc_21302_new_n5337_));
NAND2X1 NAND2X1_749 ( .A(core__abc_21302_new_n2705_), .B(core__abc_21302_new_n5330_), .Y(core__abc_21302_new_n5342_));
NAND2X1 NAND2X1_75 ( .A(core__abc_21302_new_n1409_), .B(core__abc_21302_new_n1410_), .Y(core__abc_21302_new_n1411_));
NAND2X1 NAND2X1_750 ( .A(core__abc_21302_new_n2707_), .B(core__abc_21302_new_n5328_), .Y(core__abc_21302_new_n5343_));
NAND2X1 NAND2X1_751 ( .A(core__abc_21302_new_n5350_), .B(core__abc_21302_new_n5349_), .Y(core__abc_21302_new_n5351_));
NAND2X1 NAND2X1_752 ( .A(core__abc_21302_new_n5353_), .B(core__abc_21302_new_n5354_), .Y(core__abc_21302_new_n5355_));
NAND2X1 NAND2X1_753 ( .A(core__abc_21302_new_n5347_), .B(core__abc_21302_new_n5310_), .Y(core__abc_21302_new_n5359_));
NAND2X1 NAND2X1_754 ( .A(core__abc_21302_new_n5352_), .B(core__abc_21302_new_n5355_), .Y(core__abc_21302_new_n5360_));
NAND2X1 NAND2X1_755 ( .A(core__abc_21302_new_n5361_), .B(core__abc_21302_new_n5357_), .Y(core__abc_21302_new_n5362_));
NAND2X1 NAND2X1_756 ( .A(core__abc_21302_new_n2787_), .B(core__abc_21302_new_n2786_), .Y(core__abc_21302_new_n5368_));
NAND2X1 NAND2X1_757 ( .A(core__abc_21302_new_n5372_), .B(core__abc_21302_new_n5373_), .Y(core__abc_21302_new_n5374_));
NAND2X1 NAND2X1_758 ( .A(core__abc_21302_new_n5371_), .B(core__abc_21302_new_n5374_), .Y(core__abc_21302_new_n5375_));
NAND2X1 NAND2X1_759 ( .A(core__abc_21302_new_n5380_), .B(core__abc_21302_new_n5377_), .Y(core__abc_21302_new_n5381_));
NAND2X1 NAND2X1_76 ( .A(core__abc_21302_new_n1408_), .B(core__abc_21302_new_n1411_), .Y(core__abc_21302_new_n1412_));
NAND2X1 NAND2X1_760 ( .A(core__abc_21302_new_n5345_), .B(core__abc_21302_new_n5388_), .Y(core__abc_21302_new_n5390_));
NAND2X1 NAND2X1_761 ( .A(core__abc_21302_new_n5368_), .B(core__abc_21302_new_n5373_), .Y(core__abc_21302_new_n5391_));
NAND2X1 NAND2X1_762 ( .A(core__abc_21302_new_n5388_), .B(core__abc_21302_new_n5347_), .Y(core__abc_21302_new_n5396_));
NAND2X1 NAND2X1_763 ( .A(core__abc_21302_new_n2829_), .B(core__abc_21302_new_n5405_), .Y(core__abc_21302_new_n5406_));
NAND2X1 NAND2X1_764 ( .A(core__abc_21302_new_n5407_), .B(core__abc_21302_new_n5406_), .Y(core__abc_21302_new_n5408_));
NAND2X1 NAND2X1_765 ( .A(core__abc_21302_new_n2362__bF_buf7), .B(core__abc_21302_new_n5411_), .Y(core__abc_21302_new_n5412_));
NAND2X1 NAND2X1_766 ( .A(core__abc_21302_new_n5406_), .B(core__abc_21302_new_n5420_), .Y(core__abc_21302_new_n5421_));
NAND2X1 NAND2X1_767 ( .A(core__abc_21302_new_n2868_), .B(core__abc_21302_new_n5423_), .Y(core__abc_21302_new_n5424_));
NAND2X1 NAND2X1_768 ( .A(core__abc_21302_new_n5424_), .B(core__abc_21302_new_n5425_), .Y(core__abc_21302_new_n5426_));
NAND2X1 NAND2X1_769 ( .A(core__abc_21302_new_n2634__bF_buf5), .B(core__abc_21302_new_n5427_), .Y(core__abc_21302_new_n5428_));
NAND2X1 NAND2X1_77 ( .A(core_v2_reg_19_), .B(core_v3_reg_19_), .Y(core__abc_21302_new_n1420_));
NAND2X1 NAND2X1_770 ( .A(core_key_17_), .B(core__abc_21302_new_n2639__bF_buf3), .Y(core__abc_21302_new_n5429_));
NAND2X1 NAND2X1_771 ( .A(core__abc_21302_new_n3384_), .B(core__abc_21302_new_n3383_), .Y(core__abc_21302_new_n5434_));
NAND2X1 NAND2X1_772 ( .A(core__abc_21302_new_n2904_), .B(core__abc_21302_new_n5436_), .Y(core__abc_21302_new_n5437_));
NAND2X1 NAND2X1_773 ( .A(core__abc_21302_new_n5438_), .B(core__abc_21302_new_n5437_), .Y(core__abc_21302_new_n5439_));
NAND2X1 NAND2X1_774 ( .A(core__abc_21302_new_n5406_), .B(core__abc_21302_new_n5424_), .Y(core__abc_21302_new_n5441_));
NAND2X1 NAND2X1_775 ( .A(core__abc_21302_new_n5442_), .B(core__abc_21302_new_n5444_), .Y(core__abc_21302_new_n5445_));
NAND2X1 NAND2X1_776 ( .A(core__abc_21302_new_n5440_), .B(core__abc_21302_new_n5445_), .Y(core__abc_21302_new_n5446_));
NAND2X1 NAND2X1_777 ( .A(core__abc_21302_new_n5437_), .B(core__abc_21302_new_n5446_), .Y(core__abc_21302_new_n5454_));
NAND2X1 NAND2X1_778 ( .A(core__abc_21302_new_n5456_), .B(core__abc_21302_new_n5454_), .Y(core__abc_21302_new_n5458_));
NAND2X1 NAND2X1_779 ( .A(core__abc_21302_new_n5458_), .B(core__abc_21302_new_n5457_), .Y(core__abc_21302_new_n5459_));
NAND2X1 NAND2X1_78 ( .A(core__abc_21302_new_n1421_), .B(core__abc_21302_new_n1422_), .Y(core__abc_21302_new_n1423_));
NAND2X1 NAND2X1_780 ( .A(core__abc_21302_new_n5456_), .B(core__abc_21302_new_n5440_), .Y(core__abc_21302_new_n5469_));
NAND2X1 NAND2X1_781 ( .A(core__abc_21302_new_n5471_), .B(core__abc_21302_new_n5073_), .Y(core__abc_21302_new_n5472_));
NAND2X1 NAND2X1_782 ( .A(core__abc_21302_new_n2990_), .B(core__abc_21302_new_n5480_), .Y(core__abc_21302_new_n5483_));
NAND2X1 NAND2X1_783 ( .A(core__abc_21302_new_n2634__bF_buf3), .B(core__abc_21302_new_n5485_), .Y(core__abc_21302_new_n5486_));
NAND2X1 NAND2X1_784 ( .A(core_key_20_), .B(core__abc_21302_new_n2639__bF_buf2), .Y(core__abc_21302_new_n5487_));
NAND2X1 NAND2X1_785 ( .A(core__abc_21302_new_n5493_), .B(core__abc_21302_new_n3030_), .Y(core__abc_21302_new_n5494_));
NAND2X1 NAND2X1_786 ( .A(core__abc_21302_new_n5494_), .B(core__abc_21302_new_n5495_), .Y(core__abc_21302_new_n5496_));
NAND2X1 NAND2X1_787 ( .A(core__abc_21302_new_n5497_), .B(core__abc_21302_new_n5500_), .Y(core__abc_21302_new_n5501_));
NAND2X1 NAND2X1_788 ( .A(core__abc_21302_new_n3071_), .B(core__abc_21302_new_n5509_), .Y(core__abc_21302_new_n5510_));
NAND2X1 NAND2X1_789 ( .A(core__abc_21302_new_n5510_), .B(core__abc_21302_new_n5512_), .Y(core__abc_21302_new_n5513_));
NAND2X1 NAND2X1_79 ( .A(core__abc_21302_new_n1420_), .B(core__abc_21302_new_n1423_), .Y(core__abc_21302_new_n1424_));
NAND2X1 NAND2X1_790 ( .A(core__abc_21302_new_n5484_), .B(core__abc_21302_new_n5499_), .Y(core__abc_21302_new_n5514_));
NAND2X1 NAND2X1_791 ( .A(core__abc_21302_new_n5521_), .B(core__abc_21302_new_n5520_), .Y(core__abc_21302_new_n5522_));
NAND2X1 NAND2X1_792 ( .A(core__abc_21302_new_n3589_), .B(core__abc_21302_new_n3590_), .Y(core__abc_21302_new_n5529_));
NAND2X1 NAND2X1_793 ( .A(core__abc_21302_new_n3116_), .B(core__abc_21302_new_n5530_), .Y(core__abc_21302_new_n5531_));
NAND2X1 NAND2X1_794 ( .A(core__abc_21302_new_n5531_), .B(core__abc_21302_new_n5533_), .Y(core__abc_21302_new_n5534_));
NAND2X1 NAND2X1_795 ( .A(core__abc_21302_new_n5474_), .B(core__abc_21302_new_n5546_), .Y(core__abc_21302_new_n5552_));
NAND2X1 NAND2X1_796 ( .A(core__abc_21302_new_n5554_), .B(core__abc_21302_new_n3164_), .Y(core__abc_21302_new_n5557_));
NAND2X1 NAND2X1_797 ( .A(core__abc_21302_new_n5557_), .B(core__abc_21302_new_n5556_), .Y(core__abc_21302_new_n5558_));
NAND2X1 NAND2X1_798 ( .A(core__abc_21302_new_n5558_), .B(core__abc_21302_new_n5561_), .Y(core__abc_21302_new_n5562_));
NAND2X1 NAND2X1_799 ( .A(core__abc_21302_new_n5560_), .B(core__abc_21302_new_n5562_), .Y(core__abc_21302_new_n5563_));
NAND2X1 NAND2X1_8 ( .A(\addr[5] ), .B(_abc_19873_new_n899_), .Y(_abc_19873_new_n900_));
NAND2X1 NAND2X1_80 ( .A(core_v2_reg_20_), .B(core_v3_reg_20_), .Y(core__abc_21302_new_n1432_));
NAND2X1 NAND2X1_800 ( .A(core_key_24_), .B(core__abc_21302_new_n2639__bF_buf1), .Y(core__abc_21302_new_n5564_));
NAND2X1 NAND2X1_801 ( .A(core__abc_21302_new_n3253_), .B(core__abc_21302_new_n3252_), .Y(core__abc_21302_new_n5583_));
NAND2X1 NAND2X1_802 ( .A(core__abc_21302_new_n5586_), .B(core__abc_21302_new_n5585_), .Y(core__abc_21302_new_n5587_));
NAND2X1 NAND2X1_803 ( .A(core__abc_21302_new_n5559_), .B(core__abc_21302_new_n5576_), .Y(core__abc_21302_new_n5588_));
NAND2X1 NAND2X1_804 ( .A(core__abc_21302_new_n5594_), .B(core__abc_21302_new_n5593_), .Y(core__abc_21302_new_n5595_));
NAND2X1 NAND2X1_805 ( .A(core__abc_21302_new_n3731_), .B(core__abc_21302_new_n3733_), .Y(core__abc_21302_new_n5602_));
NAND2X1 NAND2X1_806 ( .A(core__abc_21302_new_n5604_), .B(core__abc_21302_new_n5606_), .Y(core__abc_21302_new_n5607_));
NAND2X1 NAND2X1_807 ( .A(core__abc_21302_new_n5617_), .B(core__abc_21302_new_n5589_), .Y(core__abc_21302_new_n5618_));
NAND2X1 NAND2X1_808 ( .A(core__abc_21302_new_n5626_), .B(core__abc_21302_new_n3358_), .Y(core__abc_21302_new_n5627_));
NAND2X1 NAND2X1_809 ( .A(core__abc_21302_new_n5628_), .B(core__abc_21302_new_n5627_), .Y(core__abc_21302_new_n5629_));
NAND2X1 NAND2X1_81 ( .A(core__abc_21302_new_n1433_), .B(core__abc_21302_new_n1434_), .Y(core__abc_21302_new_n1435_));
NAND2X1 NAND2X1_810 ( .A(core__abc_21302_new_n5637_), .B(core__abc_21302_new_n5630_), .Y(core__abc_21302_new_n5638_));
NAND2X1 NAND2X1_811 ( .A(core_key_28_), .B(core__abc_21302_new_n2639__bF_buf0), .Y(core__abc_21302_new_n5639_));
NAND2X1 NAND2X1_812 ( .A(core__abc_21302_new_n3401_), .B(core__abc_21302_new_n3397_), .Y(core__abc_21302_new_n5645_));
NAND2X1 NAND2X1_813 ( .A(core__abc_21302_new_n5647_), .B(core__abc_21302_new_n5645_), .Y(core__abc_21302_new_n5649_));
NAND2X1 NAND2X1_814 ( .A(core__abc_21302_new_n5649_), .B(core__abc_21302_new_n5648_), .Y(core__abc_21302_new_n5650_));
NAND2X1 NAND2X1_815 ( .A(core__abc_21302_new_n5636_), .B(core__abc_21302_new_n5652_), .Y(core__abc_21302_new_n5654_));
NAND2X1 NAND2X1_816 ( .A(core__abc_21302_new_n3445_), .B(core__abc_21302_new_n3444_), .Y(core__abc_21302_new_n5667_));
NAND2X1 NAND2X1_817 ( .A(core__abc_21302_new_n5670_), .B(core__abc_21302_new_n5667_), .Y(core__abc_21302_new_n5672_));
NAND2X1 NAND2X1_818 ( .A(core__abc_21302_new_n5672_), .B(core__abc_21302_new_n5671_), .Y(core__abc_21302_new_n5673_));
NAND2X1 NAND2X1_819 ( .A(core__abc_21302_new_n5675_), .B(core__abc_21302_new_n5676_), .Y(core__abc_21302_new_n5677_));
NAND2X1 NAND2X1_82 ( .A(core__abc_21302_new_n1432_), .B(core__abc_21302_new_n1435_), .Y(core__abc_21302_new_n1436_));
NAND2X1 NAND2X1_820 ( .A(core__abc_21302_new_n3880_), .B(core__abc_21302_new_n3882_), .Y(core__abc_21302_new_n5686_));
NAND2X1 NAND2X1_821 ( .A(core__abc_21302_new_n5049_), .B(core__abc_21302_new_n5708_), .Y(core__abc_21302_new_n5709_));
NAND2X1 NAND2X1_822 ( .A(core__abc_21302_new_n2634__bF_buf6), .B(core__abc_21302_new_n5714_), .Y(core__abc_21302_new_n5715_));
NAND2X1 NAND2X1_823 ( .A(core__abc_21302_new_n5038_), .B(core__abc_21302_new_n5040_), .Y(core__abc_21302_new_n5720_));
NAND2X1 NAND2X1_824 ( .A(core__abc_21302_new_n2634__bF_buf5), .B(core__abc_21302_new_n5721_), .Y(core__abc_21302_new_n5722_));
NAND2X1 NAND2X1_825 ( .A(core_key_36_), .B(core__abc_21302_new_n2639__bF_buf5), .Y(core__abc_21302_new_n5732_));
NAND2X1 NAND2X1_826 ( .A(core__abc_21302_new_n5032_), .B(core__abc_21302_new_n5031_), .Y(core__abc_21302_new_n5738_));
NAND2X1 NAND2X1_827 ( .A(core_v2_reg_37_), .B(core__abc_21302_new_n2365__bF_buf4), .Y(core__abc_21302_new_n5740_));
NAND2X1 NAND2X1_828 ( .A(core__abc_21302_new_n2634__bF_buf4), .B(core__abc_21302_new_n5745_), .Y(core__abc_21302_new_n5746_));
NAND2X1 NAND2X1_829 ( .A(core_v2_reg_38_), .B(core__abc_21302_new_n2365__bF_buf3), .Y(core__abc_21302_new_n5747_));
NAND2X1 NAND2X1_83 ( .A(core_v2_reg_21_), .B(core_v3_reg_21_), .Y(core__abc_21302_new_n1444_));
NAND2X1 NAND2X1_830 ( .A(core__abc_21302_new_n5020_), .B(core__abc_21302_new_n5023_), .Y(core__abc_21302_new_n5752_));
NAND2X1 NAND2X1_831 ( .A(core__abc_21302_new_n2634__bF_buf3), .B(core__abc_21302_new_n5756_), .Y(core__abc_21302_new_n5757_));
NAND2X1 NAND2X1_832 ( .A(core_v2_reg_39_), .B(core__abc_21302_new_n2365__bF_buf2), .Y(core__abc_21302_new_n5759_));
NAND2X1 NAND2X1_833 ( .A(core__abc_21302_new_n2634__bF_buf2), .B(core__abc_21302_new_n5764_), .Y(core__abc_21302_new_n5765_));
NAND2X1 NAND2X1_834 ( .A(core__abc_21302_new_n5013_), .B(core__abc_21302_new_n5773_), .Y(core__abc_21302_new_n5774_));
NAND2X1 NAND2X1_835 ( .A(core_v2_reg_41_), .B(core__abc_21302_new_n2365__bF_buf1), .Y(core__abc_21302_new_n5777_));
NAND2X1 NAND2X1_836 ( .A(core__abc_21302_new_n2634__bF_buf1), .B(core__abc_21302_new_n5783_), .Y(core__abc_21302_new_n5784_));
NAND2X1 NAND2X1_837 ( .A(core_v2_reg_42_), .B(core__abc_21302_new_n2365__bF_buf0), .Y(core__abc_21302_new_n5785_));
NAND2X1 NAND2X1_838 ( .A(core__abc_21302_new_n2634__bF_buf0), .B(core__abc_21302_new_n5791_), .Y(core__abc_21302_new_n5792_));
NAND2X1 NAND2X1_839 ( .A(core__abc_21302_new_n5797_), .B(core__abc_21302_new_n5800_), .Y(core__abc_21302_new_n5801_));
NAND2X1 NAND2X1_84 ( .A(core__abc_21302_new_n1445_), .B(core__abc_21302_new_n1446_), .Y(core__abc_21302_new_n1447_));
NAND2X1 NAND2X1_840 ( .A(core__abc_21302_new_n2634__bF_buf8), .B(core__abc_21302_new_n5804_), .Y(core__abc_21302_new_n5805_));
NAND2X1 NAND2X1_841 ( .A(core_key_44_), .B(core__abc_21302_new_n2639__bF_buf3), .Y(core__abc_21302_new_n5806_));
NAND2X1 NAND2X1_842 ( .A(core__abc_21302_new_n4981_), .B(core__abc_21302_new_n5801_), .Y(core__abc_21302_new_n5812_));
NAND2X1 NAND2X1_843 ( .A(core_v2_reg_45_), .B(core__abc_21302_new_n2365__bF_buf3), .Y(core__abc_21302_new_n5814_));
NAND2X1 NAND2X1_844 ( .A(core__abc_21302_new_n2634__bF_buf7), .B(core__abc_21302_new_n5820_), .Y(core__abc_21302_new_n5821_));
NAND2X1 NAND2X1_845 ( .A(core_v2_reg_46_), .B(core__abc_21302_new_n2365__bF_buf2), .Y(core__abc_21302_new_n5822_));
NAND2X1 NAND2X1_846 ( .A(core__abc_21302_new_n4966_), .B(core__abc_21302_new_n4968_), .Y(core__abc_21302_new_n5829_));
NAND2X1 NAND2X1_847 ( .A(core__abc_21302_new_n2634__bF_buf6), .B(core__abc_21302_new_n5832_), .Y(core__abc_21302_new_n5833_));
NAND2X1 NAND2X1_848 ( .A(core__abc_21302_new_n5839_), .B(core__abc_21302_new_n5800_), .Y(core__abc_21302_new_n5840_));
NAND2X1 NAND2X1_849 ( .A(core__abc_21302_new_n5838_), .B(core__abc_21302_new_n5840_), .Y(core__abc_21302_new_n5841_));
NAND2X1 NAND2X1_85 ( .A(core__abc_21302_new_n1444_), .B(core__abc_21302_new_n1447_), .Y(core__abc_21302_new_n1448_));
NAND2X1 NAND2X1_850 ( .A(core__abc_21302_new_n2634__bF_buf5), .B(core__abc_21302_new_n5842_), .Y(core__abc_21302_new_n5843_));
NAND2X1 NAND2X1_851 ( .A(core_key_49_), .B(core__abc_21302_new_n2639__bF_buf1), .Y(core__abc_21302_new_n5852_));
NAND2X1 NAND2X1_852 ( .A(core__abc_21302_new_n4931_), .B(core__abc_21302_new_n5859_), .Y(core__abc_21302_new_n5860_));
NAND2X1 NAND2X1_853 ( .A(core__abc_21302_new_n2634__bF_buf4), .B(core__abc_21302_new_n5863_), .Y(core__abc_21302_new_n5864_));
NAND2X1 NAND2X1_854 ( .A(core_v2_reg_50_), .B(core__abc_21302_new_n2365__bF_buf1), .Y(core__abc_21302_new_n5866_));
NAND2X1 NAND2X1_855 ( .A(core__abc_21302_new_n2362__bF_buf2), .B(core__abc_21302_new_n5874_), .Y(core__abc_21302_new_n5875_));
NAND2X1 NAND2X1_856 ( .A(core__abc_21302_new_n2362__bF_buf1), .B(core__abc_21302_new_n5885_), .Y(core__abc_21302_new_n5886_));
NAND2X1 NAND2X1_857 ( .A(core__abc_21302_new_n4923_), .B(core__abc_21302_new_n4920_), .Y(core__abc_21302_new_n5889_));
NAND2X1 NAND2X1_858 ( .A(core__abc_21302_new_n2362__bF_buf0), .B(core__abc_21302_new_n5895_), .Y(core__abc_21302_new_n5896_));
NAND2X1 NAND2X1_859 ( .A(core__abc_21302_new_n5899_), .B(core__abc_21302_new_n5900_), .Y(core__abc_21302_new_n5902_));
NAND2X1 NAND2X1_86 ( .A(core_v2_reg_22_), .B(core_v3_reg_22_), .Y(core__abc_21302_new_n1456_));
NAND2X1 NAND2X1_860 ( .A(core__abc_21302_new_n5902_), .B(core__abc_21302_new_n5901_), .Y(core__abc_21302_new_n5903_));
NAND2X1 NAND2X1_861 ( .A(core__abc_21302_new_n4900_), .B(core__abc_21302_new_n4904_), .Y(core__abc_21302_new_n5909_));
NAND2X1 NAND2X1_862 ( .A(core__abc_21302_new_n5910_), .B(core__abc_21302_new_n5911_), .Y(core__abc_21302_new_n5913_));
NAND2X1 NAND2X1_863 ( .A(core__abc_21302_new_n5913_), .B(core__abc_21302_new_n5912_), .Y(core__abc_21302_new_n5914_));
NAND2X1 NAND2X1_864 ( .A(core__abc_21302_new_n4892_), .B(core__abc_21302_new_n5072_), .Y(core__abc_21302_new_n5921_));
NAND2X1 NAND2X1_865 ( .A(core__abc_21302_new_n5921_), .B(core__abc_21302_new_n5922_), .Y(core__abc_21302_new_n5923_));
NAND2X1 NAND2X1_866 ( .A(core__abc_21302_new_n5925_), .B(core__abc_21302_new_n5104__bF_buf2), .Y(core__abc_21302_new_n5926_));
NAND2X1 NAND2X1_867 ( .A(core__abc_21302_new_n2634__bF_buf8), .B(core__abc_21302_new_n5931_), .Y(core__abc_21302_new_n5932_));
NAND2X1 NAND2X1_868 ( .A(core__abc_21302_new_n2362__bF_buf11), .B(core__abc_21302_new_n5940_), .Y(core__abc_21302_new_n5941_));
NAND2X1 NAND2X1_869 ( .A(core__abc_21302_new_n4866_), .B(core__abc_21302_new_n5937_), .Y(core__abc_21302_new_n5945_));
NAND2X1 NAND2X1_87 ( .A(core__abc_21302_new_n1457_), .B(core__abc_21302_new_n1458_), .Y(core__abc_21302_new_n1459_));
NAND2X1 NAND2X1_870 ( .A(core__abc_21302_new_n4863_), .B(core__abc_21302_new_n5945_), .Y(core__abc_21302_new_n5946_));
NAND2X1 NAND2X1_871 ( .A(core_v2_reg_59_), .B(core__abc_21302_new_n2365__bF_buf4), .Y(core__abc_21302_new_n5948_));
NAND2X1 NAND2X1_872 ( .A(core_key_60_), .B(core__abc_21302_new_n2639__bF_buf5), .Y(core__abc_21302_new_n5960_));
NAND2X1 NAND2X1_873 ( .A(core__abc_21302_new_n4846_), .B(core__abc_21302_new_n4843_), .Y(core__abc_21302_new_n5965_));
NAND2X1 NAND2X1_874 ( .A(core__abc_21302_new_n5966_), .B(core__abc_21302_new_n5969_), .Y(core__abc_21302_new_n5970_));
NAND2X1 NAND2X1_875 ( .A(core__abc_21302_new_n4837_), .B(core__abc_21302_new_n5976_), .Y(core__abc_21302_new_n5977_));
NAND2X1 NAND2X1_876 ( .A(core__abc_21302_new_n5977_), .B(core__abc_21302_new_n5978_), .Y(core__abc_21302_new_n5979_));
NAND2X1 NAND2X1_877 ( .A(core__abc_21302_new_n4831_), .B(core__abc_21302_new_n4829_), .Y(core__abc_21302_new_n5987_));
NAND2X1 NAND2X1_878 ( .A(core__abc_21302_new_n4883_), .B(core__abc_21302_new_n5977_), .Y(core__abc_21302_new_n5988_));
NAND2X1 NAND2X1_879 ( .A(core_v2_reg_63_), .B(core__abc_21302_new_n2365__bF_buf3), .Y(core__abc_21302_new_n5990_));
NAND2X1 NAND2X1_88 ( .A(core__abc_21302_new_n1456_), .B(core__abc_21302_new_n1459_), .Y(core__abc_21302_new_n1460_));
NAND2X1 NAND2X1_880 ( .A(core__abc_21302_new_n2634__bF_buf3), .B(core__abc_21302_new_n5730_), .Y(core__abc_21302_new_n6031_));
NAND2X1 NAND2X1_881 ( .A(core_key_68_), .B(core__abc_21302_new_n2639__bF_buf2), .Y(core__abc_21302_new_n6032_));
NAND2X1 NAND2X1_882 ( .A(core__abc_21302_new_n2362__bF_buf5), .B(core__abc_21302_new_n6035_), .Y(core__abc_21302_new_n6036_));
NAND2X1 NAND2X1_883 ( .A(core__abc_21302_new_n5511_), .B(core__abc_21302_new_n5757_), .Y(core__abc_21302_new_n6054_));
NAND2X1 NAND2X1_884 ( .A(core__abc_21302_new_n5532_), .B(core__abc_21302_new_n5765_), .Y(core__abc_21302_new_n6062_));
NAND2X1 NAND2X1_885 ( .A(core__abc_21302_new_n6061_), .B(core__abc_21302_new_n6062_), .Y(core__abc_21302_new_n6063_));
NAND2X1 NAND2X1_886 ( .A(core__abc_21302_new_n5043_), .B(core__abc_21302_new_n5044_), .Y(core__abc_21302_new_n6125_));
NAND2X1 NAND2X1_887 ( .A(core__abc_21302_new_n5037_), .B(core__abc_21302_new_n5883_), .Y(core__abc_21302_new_n6139_));
NAND2X1 NAND2X1_888 ( .A(core__abc_21302_new_n5019_), .B(core__abc_21302_new_n5924_), .Y(core__abc_21302_new_n6167_));
NAND2X1 NAND2X1_889 ( .A(core__abc_21302_new_n4984_), .B(core__abc_21302_new_n5079_), .Y(core__abc_21302_new_n6220_));
NAND2X1 NAND2X1_89 ( .A(core_v2_reg_25_), .B(core_v3_reg_25_), .Y(core__abc_21302_new_n1486_));
NAND2X1 NAND2X1_890 ( .A(core__abc_21302_new_n4956_), .B(core__abc_21302_new_n5199_), .Y(core__abc_21302_new_n6258_));
NAND2X1 NAND2X1_891 ( .A(core__abc_21302_new_n4907_), .B(core__abc_21302_new_n4909_), .Y(core__abc_21302_new_n6265_));
NAND2X1 NAND2X1_892 ( .A(core__abc_21302_new_n5219_), .B(core__abc_21302_new_n5217_), .Y(core__abc_21302_new_n6267_));
NAND2X1 NAND2X1_893 ( .A(core_v1_reg_40_), .B(core__abc_21302_new_n5998__bF_buf0), .Y(core__abc_21302_new_n6277_));
NAND2X1 NAND2X1_894 ( .A(core__abc_21302_new_n4857_), .B(core__abc_21302_new_n5316_), .Y(core__abc_21302_new_n6301_));
NAND2X1 NAND2X1_895 ( .A(core__abc_21302_new_n6009__bF_buf1), .B(core__abc_21302_new_n4379_), .Y(core__abc_21302_new_n6326_));
NAND2X1 NAND2X1_896 ( .A(core__abc_21302_new_n4828_), .B(core__abc_21302_new_n5409_), .Y(core__abc_21302_new_n6330_));
NAND2X1 NAND2X1_897 ( .A(core__abc_21302_new_n5577_), .B(core__abc_21302_new_n5575_), .Y(core__abc_21302_new_n6395_));
NAND2X1 NAND2X1_898 ( .A(core__abc_21302_new_n6394_), .B(core__abc_21302_new_n6396_), .Y(core__abc_21302_new_n6397_));
NAND2X1 NAND2X1_899 ( .A(core_v0_reg_0_), .B(core__abc_21302_new_n6450__bF_buf7), .Y(core__abc_21302_new_n6451_));
NAND2X1 NAND2X1_9 ( .A(\addr[0] ), .B(\addr[1] ), .Y(_abc_19873_new_n911_));
NAND2X1 NAND2X1_90 ( .A(core__abc_21302_new_n1487_), .B(core__abc_21302_new_n1488_), .Y(core__abc_21302_new_n1489_));
NAND2X1 NAND2X1_900 ( .A(core__abc_21302_new_n6452_), .B(core__abc_21302_new_n6449__bF_buf6), .Y(core__abc_21302_new_n6453_));
NAND2X1 NAND2X1_901 ( .A(core__abc_21302_new_n6458_), .B(core__abc_21302_new_n6449__bF_buf5), .Y(core__abc_21302_new_n6459_));
NAND2X1 NAND2X1_902 ( .A(core__abc_21302_new_n6459_), .B(core__abc_21302_new_n5099_), .Y(core__abc_21302_new_n6460_));
NAND2X1 NAND2X1_903 ( .A(core_v0_reg_1_), .B(core__abc_21302_new_n6450__bF_buf6), .Y(core__abc_21302_new_n6462_));
NAND2X1 NAND2X1_904 ( .A(core__abc_21302_new_n2634__bF_buf5), .B(core__abc_21302_new_n2700_), .Y(core__abc_21302_new_n6464_));
NAND2X1 NAND2X1_905 ( .A(core__abc_21302_new_n6466_), .B(core__abc_21302_new_n6449__bF_buf4), .Y(core__abc_21302_new_n6467_));
NAND2X1 NAND2X1_906 ( .A(core_v0_reg_2_), .B(core__abc_21302_new_n6450__bF_buf5), .Y(core__abc_21302_new_n6470_));
NAND2X1 NAND2X1_907 ( .A(core_v0_reg_3_), .B(core__abc_21302_new_n6450__bF_buf4), .Y(core__abc_21302_new_n6472_));
NAND2X1 NAND2X1_908 ( .A(core__abc_21302_new_n6473_), .B(core__abc_21302_new_n6449__bF_buf3), .Y(core__abc_21302_new_n6474_));
NAND2X1 NAND2X1_909 ( .A(core__abc_21302_new_n6479_), .B(core__abc_21302_new_n6449__bF_buf2), .Y(core__abc_21302_new_n6480_));
NAND2X1 NAND2X1_91 ( .A(core_v2_reg_26_), .B(core_v3_reg_26_), .Y(core__abc_21302_new_n1498_));
NAND2X1 NAND2X1_910 ( .A(core_v0_reg_4_), .B(core__abc_21302_new_n6450__bF_buf3), .Y(core__abc_21302_new_n6483_));
NAND2X1 NAND2X1_911 ( .A(core__abc_21302_new_n6486_), .B(core__abc_21302_new_n6449__bF_buf1), .Y(core__abc_21302_new_n6487_));
NAND2X1 NAND2X1_912 ( .A(core_v0_reg_5_), .B(core__abc_21302_new_n6450__bF_buf2), .Y(core__abc_21302_new_n6490_));
NAND2X1 NAND2X1_913 ( .A(core__abc_21302_new_n6493_), .B(core__abc_21302_new_n6449__bF_buf0), .Y(core__abc_21302_new_n6494_));
NAND2X1 NAND2X1_914 ( .A(core_v0_reg_6_), .B(core__abc_21302_new_n6450__bF_buf1), .Y(core__abc_21302_new_n6497_));
NAND2X1 NAND2X1_915 ( .A(core__abc_21302_new_n6500_), .B(core__abc_21302_new_n6449__bF_buf7), .Y(core__abc_21302_new_n6501_));
NAND2X1 NAND2X1_916 ( .A(core_v0_reg_7_), .B(core__abc_21302_new_n6450__bF_buf0), .Y(core__abc_21302_new_n6504_));
NAND2X1 NAND2X1_917 ( .A(core__abc_21302_new_n6507_), .B(core__abc_21302_new_n6449__bF_buf6), .Y(core__abc_21302_new_n6508_));
NAND2X1 NAND2X1_918 ( .A(core_v0_reg_8_), .B(core__abc_21302_new_n6450__bF_buf7), .Y(core__abc_21302_new_n6511_));
NAND2X1 NAND2X1_919 ( .A(core__abc_21302_new_n6515_), .B(core__abc_21302_new_n6449__bF_buf5), .Y(core__abc_21302_new_n6516_));
NAND2X1 NAND2X1_92 ( .A(core__abc_21302_new_n1499_), .B(core__abc_21302_new_n1500_), .Y(core__abc_21302_new_n1501_));
NAND2X1 NAND2X1_920 ( .A(core_v0_reg_9_), .B(core__abc_21302_new_n6450__bF_buf6), .Y(core__abc_21302_new_n6519_));
NAND2X1 NAND2X1_921 ( .A(core__abc_21302_new_n6522_), .B(core__abc_21302_new_n6449__bF_buf4), .Y(core__abc_21302_new_n6523_));
NAND2X1 NAND2X1_922 ( .A(core_v0_reg_10_), .B(core__abc_21302_new_n6450__bF_buf5), .Y(core__abc_21302_new_n6526_));
NAND2X1 NAND2X1_923 ( .A(core__abc_21302_new_n6529_), .B(core__abc_21302_new_n6449__bF_buf3), .Y(core__abc_21302_new_n6530_));
NAND2X1 NAND2X1_924 ( .A(core_v0_reg_11_), .B(core__abc_21302_new_n6450__bF_buf4), .Y(core__abc_21302_new_n6533_));
NAND2X1 NAND2X1_925 ( .A(core__abc_21302_new_n6537_), .B(core__abc_21302_new_n6449__bF_buf2), .Y(core__abc_21302_new_n6538_));
NAND2X1 NAND2X1_926 ( .A(core_v0_reg_12_), .B(core__abc_21302_new_n6450__bF_buf3), .Y(core__abc_21302_new_n6541_));
NAND2X1 NAND2X1_927 ( .A(core__abc_21302_new_n6544_), .B(core__abc_21302_new_n6449__bF_buf1), .Y(core__abc_21302_new_n6545_));
NAND2X1 NAND2X1_928 ( .A(core_v0_reg_13_), .B(core__abc_21302_new_n6450__bF_buf2), .Y(core__abc_21302_new_n6548_));
NAND2X1 NAND2X1_929 ( .A(core__abc_21302_new_n6551_), .B(core__abc_21302_new_n6449__bF_buf0), .Y(core__abc_21302_new_n6552_));
NAND2X1 NAND2X1_93 ( .A(core__abc_21302_new_n1498_), .B(core__abc_21302_new_n1501_), .Y(core__abc_21302_new_n1502_));
NAND2X1 NAND2X1_930 ( .A(core_v0_reg_14_), .B(core__abc_21302_new_n6450__bF_buf1), .Y(core__abc_21302_new_n6555_));
NAND2X1 NAND2X1_931 ( .A(core__abc_21302_new_n6558_), .B(core__abc_21302_new_n6449__bF_buf7), .Y(core__abc_21302_new_n6559_));
NAND2X1 NAND2X1_932 ( .A(core_v0_reg_15_), .B(core__abc_21302_new_n6450__bF_buf0), .Y(core__abc_21302_new_n6562_));
NAND2X1 NAND2X1_933 ( .A(core__abc_21302_new_n6565_), .B(core__abc_21302_new_n6449__bF_buf6), .Y(core__abc_21302_new_n6566_));
NAND2X1 NAND2X1_934 ( .A(core_v0_reg_16_), .B(core__abc_21302_new_n6450__bF_buf7), .Y(core__abc_21302_new_n6569_));
NAND2X1 NAND2X1_935 ( .A(core__abc_21302_new_n6572_), .B(core__abc_21302_new_n6449__bF_buf5), .Y(core__abc_21302_new_n6573_));
NAND2X1 NAND2X1_936 ( .A(core_v0_reg_17_), .B(core__abc_21302_new_n6450__bF_buf6), .Y(core__abc_21302_new_n6576_));
NAND2X1 NAND2X1_937 ( .A(core__abc_21302_new_n6580_), .B(core__abc_21302_new_n6449__bF_buf4), .Y(core__abc_21302_new_n6581_));
NAND2X1 NAND2X1_938 ( .A(core_v0_reg_18_), .B(core__abc_21302_new_n6450__bF_buf5), .Y(core__abc_21302_new_n6584_));
NAND2X1 NAND2X1_939 ( .A(core__abc_21302_new_n6587_), .B(core__abc_21302_new_n6449__bF_buf3), .Y(core__abc_21302_new_n6588_));
NAND2X1 NAND2X1_94 ( .A(core_v2_reg_27_), .B(core_v3_reg_27_), .Y(core__abc_21302_new_n1510_));
NAND2X1 NAND2X1_940 ( .A(core_v0_reg_19_), .B(core__abc_21302_new_n6450__bF_buf4), .Y(core__abc_21302_new_n6591_));
NAND2X1 NAND2X1_941 ( .A(core__abc_21302_new_n6594_), .B(core__abc_21302_new_n6449__bF_buf2), .Y(core__abc_21302_new_n6595_));
NAND2X1 NAND2X1_942 ( .A(core_v0_reg_20_), .B(core__abc_21302_new_n6450__bF_buf3), .Y(core__abc_21302_new_n6598_));
NAND2X1 NAND2X1_943 ( .A(core__abc_21302_new_n6601_), .B(core__abc_21302_new_n6449__bF_buf1), .Y(core__abc_21302_new_n6602_));
NAND2X1 NAND2X1_944 ( .A(core_v0_reg_21_), .B(core__abc_21302_new_n6450__bF_buf2), .Y(core__abc_21302_new_n6605_));
NAND2X1 NAND2X1_945 ( .A(core__abc_21302_new_n6608_), .B(core__abc_21302_new_n6449__bF_buf0), .Y(core__abc_21302_new_n6609_));
NAND2X1 NAND2X1_946 ( .A(core_v0_reg_22_), .B(core__abc_21302_new_n6450__bF_buf1), .Y(core__abc_21302_new_n6612_));
NAND2X1 NAND2X1_947 ( .A(core__abc_21302_new_n6615_), .B(core__abc_21302_new_n6449__bF_buf7), .Y(core__abc_21302_new_n6616_));
NAND2X1 NAND2X1_948 ( .A(core_v0_reg_23_), .B(core__abc_21302_new_n6450__bF_buf0), .Y(core__abc_21302_new_n6619_));
NAND2X1 NAND2X1_949 ( .A(core_v0_reg_24_), .B(core__abc_21302_new_n6450__bF_buf7), .Y(core__abc_21302_new_n6626_));
NAND2X1 NAND2X1_95 ( .A(core__abc_21302_new_n1511_), .B(core__abc_21302_new_n1512_), .Y(core__abc_21302_new_n1513_));
NAND2X1 NAND2X1_950 ( .A(core__abc_21302_new_n6630_), .B(core__abc_21302_new_n6449__bF_buf5), .Y(core__abc_21302_new_n6631_));
NAND2X1 NAND2X1_951 ( .A(core_v0_reg_25_), .B(core__abc_21302_new_n6450__bF_buf6), .Y(core__abc_21302_new_n6634_));
NAND2X1 NAND2X1_952 ( .A(core__abc_21302_new_n6638_), .B(core__abc_21302_new_n6449__bF_buf4), .Y(core__abc_21302_new_n6639_));
NAND2X1 NAND2X1_953 ( .A(core_v0_reg_26_), .B(core__abc_21302_new_n6450__bF_buf5), .Y(core__abc_21302_new_n6642_));
NAND2X1 NAND2X1_954 ( .A(core__abc_21302_new_n6646_), .B(core__abc_21302_new_n6449__bF_buf3), .Y(core__abc_21302_new_n6647_));
NAND2X1 NAND2X1_955 ( .A(core_v0_reg_27_), .B(core__abc_21302_new_n6450__bF_buf4), .Y(core__abc_21302_new_n6650_));
NAND2X1 NAND2X1_956 ( .A(core__abc_21302_new_n6653_), .B(core__abc_21302_new_n6449__bF_buf2), .Y(core__abc_21302_new_n6654_));
NAND2X1 NAND2X1_957 ( .A(core_v0_reg_28_), .B(core__abc_21302_new_n6450__bF_buf3), .Y(core__abc_21302_new_n6657_));
NAND2X1 NAND2X1_958 ( .A(core__abc_21302_new_n6660_), .B(core__abc_21302_new_n6449__bF_buf1), .Y(core__abc_21302_new_n6661_));
NAND2X1 NAND2X1_959 ( .A(core_v0_reg_29_), .B(core__abc_21302_new_n6450__bF_buf2), .Y(core__abc_21302_new_n6664_));
NAND2X1 NAND2X1_96 ( .A(core__abc_21302_new_n1510_), .B(core__abc_21302_new_n1513_), .Y(core__abc_21302_new_n1514_));
NAND2X1 NAND2X1_960 ( .A(core__abc_21302_new_n6667_), .B(core__abc_21302_new_n6449__bF_buf0), .Y(core__abc_21302_new_n6668_));
NAND2X1 NAND2X1_961 ( .A(core_v0_reg_30_), .B(core__abc_21302_new_n6450__bF_buf1), .Y(core__abc_21302_new_n6671_));
NAND2X1 NAND2X1_962 ( .A(core__abc_21302_new_n6674_), .B(core__abc_21302_new_n6449__bF_buf7), .Y(core__abc_21302_new_n6675_));
NAND2X1 NAND2X1_963 ( .A(core_v0_reg_31_), .B(core__abc_21302_new_n6450__bF_buf0), .Y(core__abc_21302_new_n6678_));
NAND2X1 NAND2X1_964 ( .A(core__abc_21302_new_n6680_), .B(core__abc_21302_new_n6449__bF_buf6), .Y(core__abc_21302_new_n6681_));
NAND2X1 NAND2X1_965 ( .A(core_v0_reg_32_), .B(core__abc_21302_new_n6450__bF_buf7), .Y(core__abc_21302_new_n6684_));
NAND2X1 NAND2X1_966 ( .A(core__abc_21302_new_n6686_), .B(core__abc_21302_new_n6449__bF_buf5), .Y(core__abc_21302_new_n6687_));
NAND2X1 NAND2X1_967 ( .A(core_v0_reg_33_), .B(core__abc_21302_new_n6450__bF_buf6), .Y(core__abc_21302_new_n6690_));
NAND2X1 NAND2X1_968 ( .A(core__abc_21302_new_n6693_), .B(core__abc_21302_new_n6449__bF_buf4), .Y(core__abc_21302_new_n6694_));
NAND2X1 NAND2X1_969 ( .A(core_v0_reg_34_), .B(core__abc_21302_new_n6450__bF_buf5), .Y(core__abc_21302_new_n6697_));
NAND2X1 NAND2X1_97 ( .A(core_v2_reg_28_), .B(core_v3_reg_28_), .Y(core__abc_21302_new_n1522_));
NAND2X1 NAND2X1_970 ( .A(core__abc_21302_new_n6700_), .B(core__abc_21302_new_n6449__bF_buf3), .Y(core__abc_21302_new_n6701_));
NAND2X1 NAND2X1_971 ( .A(core_v0_reg_35_), .B(core__abc_21302_new_n6450__bF_buf4), .Y(core__abc_21302_new_n6704_));
NAND2X1 NAND2X1_972 ( .A(core__abc_21302_new_n6707_), .B(core__abc_21302_new_n6449__bF_buf2), .Y(core__abc_21302_new_n6708_));
NAND2X1 NAND2X1_973 ( .A(core__abc_21302_new_n6708_), .B(core__abc_21302_new_n5732_), .Y(core__abc_21302_new_n6709_));
NAND2X1 NAND2X1_974 ( .A(core_v0_reg_36_), .B(core__abc_21302_new_n6450__bF_buf3), .Y(core__abc_21302_new_n6711_));
NAND2X1 NAND2X1_975 ( .A(core__abc_21302_new_n6713_), .B(core__abc_21302_new_n6449__bF_buf1), .Y(core__abc_21302_new_n6714_));
NAND2X1 NAND2X1_976 ( .A(core_v0_reg_37_), .B(core__abc_21302_new_n6450__bF_buf2), .Y(core__abc_21302_new_n6717_));
NAND2X1 NAND2X1_977 ( .A(core__abc_21302_new_n6720_), .B(core__abc_21302_new_n6449__bF_buf0), .Y(core__abc_21302_new_n6721_));
NAND2X1 NAND2X1_978 ( .A(core_v0_reg_38_), .B(core__abc_21302_new_n6450__bF_buf1), .Y(core__abc_21302_new_n6724_));
NAND2X1 NAND2X1_979 ( .A(core__abc_21302_new_n6727_), .B(core__abc_21302_new_n6449__bF_buf7), .Y(core__abc_21302_new_n6728_));
NAND2X1 NAND2X1_98 ( .A(core__abc_21302_new_n1523_), .B(core__abc_21302_new_n1524_), .Y(core__abc_21302_new_n1525_));
NAND2X1 NAND2X1_980 ( .A(core_v0_reg_39_), .B(core__abc_21302_new_n6450__bF_buf0), .Y(core__abc_21302_new_n6731_));
NAND2X1 NAND2X1_981 ( .A(core_v0_reg_40_), .B(core__abc_21302_new_n6450__bF_buf7), .Y(core__abc_21302_new_n6737_));
NAND2X1 NAND2X1_982 ( .A(core__abc_21302_new_n6741_), .B(core__abc_21302_new_n6449__bF_buf5), .Y(core__abc_21302_new_n6742_));
NAND2X1 NAND2X1_983 ( .A(core_v0_reg_41_), .B(core__abc_21302_new_n6450__bF_buf6), .Y(core__abc_21302_new_n6745_));
NAND2X1 NAND2X1_984 ( .A(core__abc_21302_new_n6748_), .B(core__abc_21302_new_n6449__bF_buf4), .Y(core__abc_21302_new_n6749_));
NAND2X1 NAND2X1_985 ( .A(core_v0_reg_42_), .B(core__abc_21302_new_n6450__bF_buf5), .Y(core__abc_21302_new_n6752_));
NAND2X1 NAND2X1_986 ( .A(core__abc_21302_new_n6755_), .B(core__abc_21302_new_n6449__bF_buf3), .Y(core__abc_21302_new_n6756_));
NAND2X1 NAND2X1_987 ( .A(core_v0_reg_43_), .B(core__abc_21302_new_n6450__bF_buf4), .Y(core__abc_21302_new_n6759_));
NAND2X1 NAND2X1_988 ( .A(core__abc_21302_new_n6762_), .B(core__abc_21302_new_n6449__bF_buf2), .Y(core__abc_21302_new_n6763_));
NAND2X1 NAND2X1_989 ( .A(core__abc_21302_new_n6763_), .B(core__abc_21302_new_n5806_), .Y(core__abc_21302_new_n6764_));
NAND2X1 NAND2X1_99 ( .A(core__abc_21302_new_n1522_), .B(core__abc_21302_new_n1525_), .Y(core__abc_21302_new_n1526_));
NAND2X1 NAND2X1_990 ( .A(core_v0_reg_44_), .B(core__abc_21302_new_n6450__bF_buf3), .Y(core__abc_21302_new_n6766_));
NAND2X1 NAND2X1_991 ( .A(core__abc_21302_new_n4311_), .B(core__abc_21302_new_n4310_), .Y(core__abc_21302_new_n6768_));
NAND2X1 NAND2X1_992 ( .A(core__abc_21302_new_n6769_), .B(core__abc_21302_new_n6449__bF_buf1), .Y(core__abc_21302_new_n6770_));
NAND2X1 NAND2X1_993 ( .A(core_v0_reg_45_), .B(core__abc_21302_new_n6450__bF_buf2), .Y(core__abc_21302_new_n6773_));
NAND2X1 NAND2X1_994 ( .A(core__abc_21302_new_n6776_), .B(core__abc_21302_new_n6449__bF_buf0), .Y(core__abc_21302_new_n6777_));
NAND2X1 NAND2X1_995 ( .A(core_v0_reg_46_), .B(core__abc_21302_new_n6450__bF_buf1), .Y(core__abc_21302_new_n6780_));
NAND2X1 NAND2X1_996 ( .A(core__abc_21302_new_n4376_), .B(core__abc_21302_new_n4375_), .Y(core__abc_21302_new_n6782_));
NAND2X1 NAND2X1_997 ( .A(core__abc_21302_new_n6783_), .B(core__abc_21302_new_n6449__bF_buf7), .Y(core__abc_21302_new_n6784_));
NAND2X1 NAND2X1_998 ( .A(core_v0_reg_47_), .B(core__abc_21302_new_n6450__bF_buf0), .Y(core__abc_21302_new_n6787_));
NAND2X1 NAND2X1_999 ( .A(core_v0_reg_48_), .B(core__abc_21302_new_n6450__bF_buf7), .Y(core__abc_21302_new_n6793_));
NAND3X1 NAND3X1_1 ( .A(core_ready), .B(_abc_19873_new_n877_), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n882_));
NAND3X1 NAND3X1_10 ( .A(word0_reg_1_), .B(_abc_19873_new_n905__bF_buf1), .C(_abc_19873_new_n901__bF_buf2), .Y(_abc_19873_new_n938_));
NAND3X1 NAND3X1_100 ( .A(_abc_19873_new_n1386_), .B(_abc_19873_new_n1384_), .C(_abc_19873_new_n1385_), .Y(_abc_19873_new_n1387_));
NAND3X1 NAND3X1_101 ( .A(core_mi_57_), .B(_abc_19873_new_n889__bF_buf3), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1400_));
NAND3X1 NAND3X1_102 ( .A(word1_reg_25_), .B(_abc_19873_new_n895__bF_buf0), .C(_abc_19873_new_n901__bF_buf2), .Y(_abc_19873_new_n1402_));
NAND3X1 NAND3X1_103 ( .A(word2_reg_25_), .B(_abc_19873_new_n901__bF_buf1), .C(_abc_19873_new_n893__bF_buf0), .Y(_abc_19873_new_n1403_));
NAND3X1 NAND3X1_104 ( .A(word3_reg_25_), .B(_abc_19873_new_n912__bF_buf3), .C(_abc_19873_new_n901__bF_buf0), .Y(_abc_19873_new_n1404_));
NAND3X1 NAND3X1_105 ( .A(_abc_19873_new_n1404_), .B(_abc_19873_new_n1402_), .C(_abc_19873_new_n1403_), .Y(_abc_19873_new_n1405_));
NAND3X1 NAND3X1_106 ( .A(core_mi_60_), .B(_abc_19873_new_n889__bF_buf2), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1456_));
NAND3X1 NAND3X1_107 ( .A(word1_reg_28_), .B(_abc_19873_new_n895__bF_buf4), .C(_abc_19873_new_n901__bF_buf7), .Y(_abc_19873_new_n1458_));
NAND3X1 NAND3X1_108 ( .A(word2_reg_28_), .B(_abc_19873_new_n901__bF_buf6), .C(_abc_19873_new_n893__bF_buf4), .Y(_abc_19873_new_n1459_));
NAND3X1 NAND3X1_109 ( .A(word3_reg_28_), .B(_abc_19873_new_n912__bF_buf2), .C(_abc_19873_new_n901__bF_buf5), .Y(_abc_19873_new_n1460_));
NAND3X1 NAND3X1_11 ( .A(_abc_19873_new_n938_), .B(_abc_19873_new_n936_), .C(_abc_19873_new_n937_), .Y(_abc_19873_new_n939_));
NAND3X1 NAND3X1_110 ( .A(_abc_19873_new_n1460_), .B(_abc_19873_new_n1458_), .C(_abc_19873_new_n1459_), .Y(_abc_19873_new_n1461_));
NAND3X1 NAND3X1_111 ( .A(core_mi_29_), .B(_abc_19873_new_n889__bF_buf1), .C(_abc_19873_new_n874_), .Y(_abc_19873_new_n1474_));
NAND3X1 NAND3X1_112 ( .A(core_mi_61_), .B(_abc_19873_new_n889__bF_buf0), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1475_));
NAND3X1 NAND3X1_113 ( .A(core_key_29_), .B(_abc_19873_new_n905__bF_buf3), .C(_abc_19873_new_n889__bF_buf4), .Y(_abc_19873_new_n1482_));
NAND3X1 NAND3X1_114 ( .A(core_key_125_), .B(_abc_19873_new_n912__bF_buf1), .C(_abc_19873_new_n889__bF_buf3), .Y(_abc_19873_new_n1483_));
NAND3X1 NAND3X1_115 ( .A(_abc_19873_new_n1482_), .B(_abc_19873_new_n1483_), .C(_abc_19873_new_n1481_), .Y(_abc_19873_new_n1484_));
NAND3X1 NAND3X1_116 ( .A(core_mi_62_), .B(_abc_19873_new_n889__bF_buf2), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1494_));
NAND3X1 NAND3X1_117 ( .A(word1_reg_30_), .B(_abc_19873_new_n895__bF_buf3), .C(_abc_19873_new_n901__bF_buf4), .Y(_abc_19873_new_n1496_));
NAND3X1 NAND3X1_118 ( .A(word2_reg_30_), .B(_abc_19873_new_n901__bF_buf3), .C(_abc_19873_new_n893__bF_buf2), .Y(_abc_19873_new_n1497_));
NAND3X1 NAND3X1_119 ( .A(word3_reg_30_), .B(_abc_19873_new_n912__bF_buf0), .C(_abc_19873_new_n901__bF_buf2), .Y(_abc_19873_new_n1498_));
NAND3X1 NAND3X1_12 ( .A(core_key_1_), .B(_abc_19873_new_n905__bF_buf0), .C(_abc_19873_new_n889__bF_buf2), .Y(_abc_19873_new_n945_));
NAND3X1 NAND3X1_120 ( .A(_abc_19873_new_n1498_), .B(_abc_19873_new_n1496_), .C(_abc_19873_new_n1497_), .Y(_abc_19873_new_n1499_));
NAND3X1 NAND3X1_121 ( .A(_abc_19873_new_n877_), .B(_abc_19873_new_n2284_), .C(_abc_19873_new_n2294_), .Y(_abc_19873_new_n2295_));
NAND3X1 NAND3X1_122 ( .A(core__abc_21302_new_n1136_), .B(core__abc_21302_new_n1140_), .C(core__abc_21302_new_n1134_), .Y(core__abc_21302_new_n1141_));
NAND3X1 NAND3X1_123 ( .A(core__abc_21302_new_n1170_), .B(core__abc_21302_new_n1173_), .C(core__abc_21302_new_n1168_), .Y(core__abc_21302_new_n1174_));
NAND3X1 NAND3X1_124 ( .A(core__abc_21302_new_n1146_), .B(core__abc_21302_new_n1159_), .C(core__abc_21302_new_n1178_), .Y(core__abc_21302_new_n1179_));
NAND3X1 NAND3X1_125 ( .A(core__abc_21302_new_n1191_), .B(core__abc_21302_new_n1192_), .C(core__abc_21302_new_n1187_), .Y(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_0_));
NAND3X1 NAND3X1_126 ( .A(core__abc_21302_new_n1186_), .B(core__abc_21302_new_n1205_), .C(core__abc_21302_new_n1179_), .Y(core__abc_21302_new_n1206_));
NAND3X1 NAND3X1_127 ( .A(core__abc_21302_new_n1234_), .B(core__abc_21302_new_n2374_), .C(core__abc_21302_new_n2375_), .Y(core__abc_21302_new_n2376_));
NAND3X1 NAND3X1_128 ( .A(core__abc_21302_new_n1360_), .B(core__abc_21302_new_n1372_), .C(core__abc_21302_new_n2415_), .Y(core__abc_21302_new_n2416_));
NAND3X1 NAND3X1_129 ( .A(core__abc_21302_new_n2431_), .B(core__abc_21302_new_n2432_), .C(core__abc_21302_new_n2430_), .Y(core__abc_21302_new_n2433_));
NAND3X1 NAND3X1_13 ( .A(word0_reg_2_), .B(_abc_19873_new_n905__bF_buf2), .C(_abc_19873_new_n901__bF_buf0), .Y(_abc_19873_new_n963_));
NAND3X1 NAND3X1_130 ( .A(core__abc_21302_new_n1546_), .B(core__abc_21302_new_n1558_), .C(core__abc_21302_new_n2462_), .Y(core__abc_21302_new_n2463_));
NAND3X1 NAND3X1_131 ( .A(core__abc_21302_new_n1293_), .B(core__abc_21302_new_n1303_), .C(core__abc_21302_new_n2484_), .Y(core__abc_21302_new_n2485_));
NAND3X1 NAND3X1_132 ( .A(core__abc_21302_new_n1237_), .B(core__abc_21302_new_n1246_), .C(core__abc_21302_new_n2517_), .Y(core__abc_21302_new_n2518_));
NAND3X1 NAND3X1_133 ( .A(core__abc_21302_new_n2549_), .B(core__abc_21302_new_n2550_), .C(core__abc_21302_new_n2555_), .Y(core__abc_21302_new_n2556_));
NAND3X1 NAND3X1_134 ( .A(core__abc_21302_new_n1683_), .B(core__abc_21302_new_n2513_), .C(core__abc_21302_new_n2624_), .Y(core__abc_21302_new_n2625_));
NAND3X1 NAND3X1_135 ( .A(core__abc_21302_new_n1683_), .B(core__abc_21302_new_n1697_), .C(core__abc_21302_new_n2624_), .Y(core__abc_21302_new_n2629_));
NAND3X1 NAND3X1_136 ( .A(core__abc_21302_new_n2649_), .B(core__abc_21302_new_n2653_), .C(core__abc_21302_new_n2650_), .Y(core__abc_21302_new_n2655_));
NAND3X1 NAND3X1_137 ( .A(core_v3_reg_30_), .B(core__abc_21302_new_n2729_), .C(core__abc_21302_new_n2730_), .Y(core__abc_21302_new_n2731_));
NAND3X1 NAND3X1_138 ( .A(core__abc_21302_new_n1591_), .B(core__abc_21302_new_n1604_), .C(core__abc_21302_new_n2687_), .Y(core__abc_21302_new_n2735_));
NAND3X1 NAND3X1_139 ( .A(core__abc_21302_new_n2682_), .B(core__abc_21302_new_n2737_), .C(core__abc_21302_new_n2684_), .Y(core__abc_21302_new_n2762_));
NAND3X1 NAND3X1_14 ( .A(word1_reg_2_), .B(_abc_19873_new_n895__bF_buf2), .C(_abc_19873_new_n901__bF_buf7), .Y(_abc_19873_new_n964_));
NAND3X1 NAND3X1_140 ( .A(core__abc_21302_new_n1730_), .B(core__abc_21302_new_n1743_), .C(core__abc_21302_new_n2729_), .Y(core__abc_21302_new_n2782_));
NAND3X1 NAND3X1_141 ( .A(core__abc_21302_new_n1730_), .B(core__abc_21302_new_n2783_), .C(core__abc_21302_new_n2729_), .Y(core__abc_21302_new_n2786_));
NAND3X1 NAND3X1_142 ( .A(core__abc_21302_new_n2803_), .B(core__abc_21302_new_n2807_), .C(core__abc_21302_new_n2802_), .Y(core__abc_21302_new_n2808_));
NAND3X1 NAND3X1_143 ( .A(core__abc_21302_new_n2720_), .B(core__abc_21302_new_n2814_), .C(core__abc_21302_new_n2662_), .Y(core__abc_21302_new_n2819_));
NAND3X1 NAND3X1_144 ( .A(core__abc_21302_new_n2857_), .B(core__abc_21302_new_n2891_), .C(core__abc_21302_new_n2888_), .Y(core__abc_21302_new_n2916_));
NAND3X1 NAND3X1_145 ( .A(core__abc_21302_new_n2944_), .B(core__abc_21302_new_n2972_), .C(core__abc_21302_new_n2975_), .Y(core__abc_21302_new_n3002_));
NAND3X1 NAND3X1_146 ( .A(core__abc_21302_new_n3046_), .B(core__abc_21302_new_n3048_), .C(core__abc_21302_new_n3056_), .Y(core__abc_21302_new_n3057_));
NAND3X1 NAND3X1_147 ( .A(core__abc_21302_new_n3024_), .B(core__abc_21302_new_n3060_), .C(core__abc_21302_new_n3057_), .Y(core__abc_21302_new_n3083_));
NAND3X1 NAND3X1_148 ( .A(core__abc_21302_new_n3112_), .B(core__abc_21302_new_n1839_), .C(core__abc_21302_new_n3067_), .Y(core__abc_21302_new_n3113_));
NAND3X1 NAND3X1_149 ( .A(core__abc_21302_new_n3199_), .B(core__abc_21302_new_n3200_), .C(core__abc_21302_new_n3201_), .Y(core__abc_21302_new_n3202_));
NAND3X1 NAND3X1_15 ( .A(word3_reg_2_), .B(_abc_19873_new_n912__bF_buf1), .C(_abc_19873_new_n901__bF_buf6), .Y(_abc_19873_new_n965_));
NAND3X1 NAND3X1_150 ( .A(core__abc_21302_new_n1726_), .B(core__abc_21302_new_n1739_), .C(core__abc_21302_new_n3199_), .Y(core__abc_21302_new_n3224_));
NAND3X1 NAND3X1_151 ( .A(core__abc_21302_new_n1361_), .B(core__abc_21302_new_n1377_), .C(core__abc_21302_new_n3192_), .Y(core__abc_21302_new_n3227_));
NAND3X1 NAND3X1_152 ( .A(core__abc_21302_new_n3224_), .B(core__abc_21302_new_n3226_), .C(core__abc_21302_new_n3235_), .Y(core__abc_21302_new_n3236_));
NAND3X1 NAND3X1_153 ( .A(core_v3_reg_42_), .B(core__abc_21302_new_n3253_), .C(core__abc_21302_new_n3252_), .Y(core__abc_21302_new_n3254_));
NAND3X1 NAND3X1_154 ( .A(core__abc_21302_new_n3109_), .B(core__abc_21302_new_n3146_), .C(core__abc_21302_new_n3271_), .Y(core__abc_21302_new_n3272_));
NAND3X1 NAND3X1_155 ( .A(core__abc_21302_new_n3236_), .B(core__abc_21302_new_n3241_), .C(core__abc_21302_new_n3203_), .Y(core__abc_21302_new_n3273_));
NAND3X1 NAND3X1_156 ( .A(core__abc_21302_new_n3088_), .B(core__abc_21302_new_n3274_), .C(core__abc_21302_new_n2919_), .Y(core__abc_21302_new_n3275_));
NAND3X1 NAND3X1_157 ( .A(core__abc_21302_new_n3276_), .B(core__abc_21302_new_n3275_), .C(core__abc_21302_new_n3284_), .Y(core__abc_21302_new_n3285_));
NAND3X1 NAND3X1_158 ( .A(core__abc_21302_new_n3312_), .B(core__abc_21302_new_n3313_), .C(core__abc_21302_new_n3253_), .Y(core__abc_21302_new_n3314_));
NAND3X1 NAND3X1_159 ( .A(core__abc_21302_new_n3383_), .B(core__abc_21302_new_n3384_), .C(core__abc_21302_new_n3388_), .Y(core__abc_21302_new_n3389_));
NAND3X1 NAND3X1_16 ( .A(_abc_19873_new_n963_), .B(_abc_19873_new_n965_), .C(_abc_19873_new_n964_), .Y(_abc_19873_new_n966_));
NAND3X1 NAND3X1_160 ( .A(core__abc_21302_new_n3398_), .B(core__abc_21302_new_n3399_), .C(core__abc_21302_new_n3400_), .Y(core__abc_21302_new_n3401_));
NAND3X1 NAND3X1_161 ( .A(core_v3_reg_45_), .B(core__abc_21302_new_n3401_), .C(core__abc_21302_new_n3397_), .Y(core__abc_21302_new_n3402_));
NAND3X1 NAND3X1_162 ( .A(core__abc_21302_new_n3398_), .B(core__abc_21302_new_n1919_), .C(core__abc_21302_new_n3400_), .Y(core__abc_21302_new_n3405_));
NAND3X1 NAND3X1_163 ( .A(core__abc_21302_new_n3403_), .B(core__abc_21302_new_n3405_), .C(core__abc_21302_new_n3404_), .Y(core__abc_21302_new_n3406_));
NAND3X1 NAND3X1_164 ( .A(core__abc_21302_new_n1771_), .B(core__abc_21302_new_n1785_), .C(core__abc_21302_new_n3383_), .Y(core__abc_21302_new_n3417_));
NAND3X1 NAND3X1_165 ( .A(core_v3_reg_3_), .B(core__abc_21302_new_n3422_), .C(core__abc_21302_new_n3421_), .Y(core__abc_21302_new_n3423_));
NAND3X1 NAND3X1_166 ( .A(core__abc_21302_new_n1771_), .B(core__abc_21302_new_n3418_), .C(core__abc_21302_new_n3383_), .Y(core__abc_21302_new_n3430_));
NAND3X1 NAND3X1_167 ( .A(core_v3_reg_46_), .B(core__abc_21302_new_n3445_), .C(core__abc_21302_new_n3444_), .Y(core__abc_21302_new_n3448_));
NAND3X1 NAND3X1_168 ( .A(core__abc_21302_new_n3394_), .B(core__abc_21302_new_n3465_), .C(core__abc_21302_new_n3434_), .Y(core__abc_21302_new_n3466_));
NAND3X1 NAND3X1_169 ( .A(core_v3_reg_5_), .B(core__abc_21302_new_n3511_), .C(core__abc_21302_new_n3510_), .Y(core__abc_21302_new_n3512_));
NAND3X1 NAND3X1_17 ( .A(core_finalize), .B(_abc_19873_new_n877_), .C(_abc_19873_new_n874_), .Y(_abc_19873_new_n972_));
NAND3X1 NAND3X1_170 ( .A(core__abc_21302_new_n3503_), .B(core__abc_21302_new_n3506_), .C(core__abc_21302_new_n3516_), .Y(core__abc_21302_new_n3533_));
NAND3X1 NAND3X1_171 ( .A(core__abc_21302_new_n2883_), .B(core__abc_21302_new_n3553_), .C(core__abc_21302_new_n3554_), .Y(core__abc_21302_new_n3555_));
NAND3X1 NAND3X1_172 ( .A(core__abc_21302_new_n3558_), .B(core__abc_21302_new_n3560_), .C(core__abc_21302_new_n3559_), .Y(core__abc_21302_new_n3561_));
NAND3X1 NAND3X1_173 ( .A(core__abc_21302_new_n1819_), .B(core__abc_21302_new_n3576_), .C(core__abc_21302_new_n3558_), .Y(core__abc_21302_new_n3577_));
NAND3X1 NAND3X1_174 ( .A(core__abc_21302_new_n1456_), .B(core__abc_21302_new_n2576_), .C(core__abc_21302_new_n3553_), .Y(core__abc_21302_new_n3580_));
NAND3X1 NAND3X1_175 ( .A(core_v3_reg_7_), .B(core__abc_21302_new_n3580_), .C(core__abc_21302_new_n3581_), .Y(core__abc_21302_new_n3582_));
NAND3X1 NAND3X1_176 ( .A(core__abc_21302_new_n1456_), .B(core__abc_21302_new_n1468_), .C(core__abc_21302_new_n3553_), .Y(core__abc_21302_new_n3584_));
NAND3X1 NAND3X1_177 ( .A(core__abc_21302_new_n3583_), .B(core__abc_21302_new_n3584_), .C(core__abc_21302_new_n3585_), .Y(core__abc_21302_new_n3586_));
NAND3X1 NAND3X1_178 ( .A(core__abc_21302_new_n1819_), .B(core__abc_21302_new_n1834_), .C(core__abc_21302_new_n3558_), .Y(core__abc_21302_new_n3589_));
NAND3X1 NAND3X1_179 ( .A(core__abc_21302_new_n3604_), .B(core__abc_21302_new_n3464_), .C(core__abc_21302_new_n3606_), .Y(core__abc_21302_new_n3607_));
NAND3X1 NAND3X1_18 ( .A(word0_reg_3_), .B(_abc_19873_new_n905__bF_buf0), .C(_abc_19873_new_n901__bF_buf5), .Y(_abc_19873_new_n985_));
NAND3X1 NAND3X1_180 ( .A(core__abc_21302_new_n3589_), .B(core__abc_21302_new_n3590_), .C(core__abc_21302_new_n3609_), .Y(core__abc_21302_new_n3610_));
NAND3X1 NAND3X1_181 ( .A(core__abc_21302_new_n3611_), .B(core__abc_21302_new_n3608_), .C(core__abc_21302_new_n3607_), .Y(core__abc_21302_new_n3612_));
NAND3X1 NAND3X1_182 ( .A(core__abc_21302_new_n3577_), .B(core__abc_21302_new_n3587_), .C(core__abc_21302_new_n3579_), .Y(core__abc_21302_new_n3613_));
NAND3X1 NAND3X1_183 ( .A(core__abc_21302_new_n3562_), .B(core__abc_21302_new_n3613_), .C(core__abc_21302_new_n3610_), .Y(core__abc_21302_new_n3614_));
NAND3X1 NAND3X1_184 ( .A(core__abc_21302_new_n3669_), .B(core__abc_21302_new_n3666_), .C(core__abc_21302_new_n3665_), .Y(core__abc_21302_new_n3670_));
NAND3X1 NAND3X1_185 ( .A(core__abc_21302_new_n3673_), .B(core__abc_21302_new_n3675_), .C(core__abc_21302_new_n3645_), .Y(core__abc_21302_new_n3690_));
NAND3X1 NAND3X1_186 ( .A(core__abc_21302_new_n3700_), .B(core__abc_21302_new_n3713_), .C(core__abc_21302_new_n3714_), .Y(core__abc_21302_new_n3715_));
NAND3X1 NAND3X1_187 ( .A(core__abc_21302_new_n3730_), .B(core__abc_21302_new_n1887_), .C(core__abc_21302_new_n3700_), .Y(core__abc_21302_new_n3731_));
NAND3X1 NAND3X1_188 ( .A(core__abc_21302_new_n1498_), .B(core__abc_21302_new_n2552_), .C(core__abc_21302_new_n3734_), .Y(core__abc_21302_new_n3735_));
NAND3X1 NAND3X1_189 ( .A(core_v3_reg_11_), .B(core__abc_21302_new_n3735_), .C(core__abc_21302_new_n3737_), .Y(core__abc_21302_new_n3738_));
NAND3X1 NAND3X1_19 ( .A(word1_reg_3_), .B(_abc_19873_new_n895__bF_buf1), .C(_abc_19873_new_n901__bF_buf4), .Y(_abc_19873_new_n986_));
NAND3X1 NAND3X1_190 ( .A(core__abc_21302_new_n1498_), .B(core__abc_21302_new_n1514_), .C(core__abc_21302_new_n3734_), .Y(core__abc_21302_new_n3739_));
NAND3X1 NAND3X1_191 ( .A(core__abc_21302_new_n1329_), .B(core__abc_21302_new_n3739_), .C(core__abc_21302_new_n3740_), .Y(core__abc_21302_new_n3741_));
NAND3X1 NAND3X1_192 ( .A(core__abc_21302_new_n3731_), .B(core__abc_21302_new_n3733_), .C(core__abc_21302_new_n3742_), .Y(core__abc_21302_new_n3743_));
NAND3X1 NAND3X1_193 ( .A(core__abc_21302_new_n3743_), .B(core__abc_21302_new_n3716_), .C(core__abc_21302_new_n3747_), .Y(core__abc_21302_new_n3761_));
NAND3X1 NAND3X1_194 ( .A(core__abc_21302_new_n1522_), .B(core__abc_21302_new_n3806_), .C(core__abc_21302_new_n3808_), .Y(core__abc_21302_new_n3809_));
NAND3X1 NAND3X1_195 ( .A(core_v3_reg_13_), .B(core__abc_21302_new_n3809_), .C(core__abc_21302_new_n3811_), .Y(core__abc_21302_new_n3812_));
NAND3X1 NAND3X1_196 ( .A(core__abc_21302_new_n3791_), .B(core__abc_21302_new_n3805_), .C(core__abc_21302_new_n3816_), .Y(core__abc_21302_new_n3818_));
NAND3X1 NAND3X1_197 ( .A(core__abc_21302_new_n1363_), .B(core__abc_21302_new_n3846_), .C(core__abc_21302_new_n3845_), .Y(core__abc_21302_new_n3847_));
NAND3X1 NAND3X1_198 ( .A(core__abc_21302_new_n3851_), .B(core__abc_21302_new_n3850_), .C(core__abc_21302_new_n3852_), .Y(core__abc_21302_new_n3853_));
NAND3X1 NAND3X1_199 ( .A(core__abc_21302_new_n3818_), .B(core__abc_21302_new_n3861_), .C(core__abc_21302_new_n3779_), .Y(core__abc_21302_new_n3862_));
NAND3X1 NAND3X1_2 ( .A(core_mi_32_), .B(_abc_19873_new_n889__bF_buf2), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n898_));
NAND3X1 NAND3X1_20 ( .A(word2_reg_3_), .B(_abc_19873_new_n901__bF_buf3), .C(_abc_19873_new_n893__bF_buf0), .Y(_abc_19873_new_n987_));
NAND3X1 NAND3X1_200 ( .A(core__abc_21302_new_n1925_), .B(core__abc_21302_new_n3879_), .C(core__abc_21302_new_n3850_), .Y(core__abc_21302_new_n3880_));
NAND3X1 NAND3X1_201 ( .A(core__abc_21302_new_n1547_), .B(core__abc_21302_new_n3883_), .C(core__abc_21302_new_n3845_), .Y(core__abc_21302_new_n3884_));
NAND3X1 NAND3X1_202 ( .A(core_v3_reg_15_), .B(core__abc_21302_new_n3884_), .C(core__abc_21302_new_n3885_), .Y(core__abc_21302_new_n3886_));
NAND3X1 NAND3X1_203 ( .A(core__abc_21302_new_n1547_), .B(core__abc_21302_new_n1559_), .C(core__abc_21302_new_n3845_), .Y(core__abc_21302_new_n3887_));
NAND3X1 NAND3X1_204 ( .A(core__abc_21302_new_n1374_), .B(core__abc_21302_new_n3887_), .C(core__abc_21302_new_n3888_), .Y(core__abc_21302_new_n3889_));
NAND3X1 NAND3X1_205 ( .A(core__abc_21302_new_n3880_), .B(core__abc_21302_new_n3882_), .C(core__abc_21302_new_n3890_), .Y(core__abc_21302_new_n3891_));
NAND3X1 NAND3X1_206 ( .A(core__abc_21302_new_n1925_), .B(core__abc_21302_new_n1937_), .C(core__abc_21302_new_n3850_), .Y(core__abc_21302_new_n3892_));
NAND3X1 NAND3X1_207 ( .A(core__abc_21302_new_n3894_), .B(core__abc_21302_new_n3892_), .C(core__abc_21302_new_n3893_), .Y(core__abc_21302_new_n3895_));
NAND3X1 NAND3X1_208 ( .A(core__abc_21302_new_n3891_), .B(core__abc_21302_new_n3895_), .C(core__abc_21302_new_n3878_), .Y(core__abc_21302_new_n3896_));
NAND3X1 NAND3X1_209 ( .A(core__abc_21302_new_n3615_), .B(core__abc_21302_new_n3910_), .C(core__abc_21302_new_n3911_), .Y(core__abc_21302_new_n3912_));
NAND3X1 NAND3X1_21 ( .A(_abc_19873_new_n985_), .B(_abc_19873_new_n986_), .C(_abc_19873_new_n987_), .Y(_abc_19873_new_n988_));
NAND3X1 NAND3X1_210 ( .A(core__abc_21302_new_n3910_), .B(core__abc_21302_new_n3911_), .C(core__abc_21302_new_n3612_), .Y(core__abc_21302_new_n3914_));
NAND3X1 NAND3X1_211 ( .A(core__abc_21302_new_n3891_), .B(core__abc_21302_new_n3895_), .C(core__abc_21302_new_n3866_), .Y(core__abc_21302_new_n3915_));
NAND3X1 NAND3X1_212 ( .A(core__abc_21302_new_n3958_), .B(core__abc_21302_new_n3929_), .C(core__abc_21302_new_n3960_), .Y(core__abc_21302_new_n3974_));
NAND3X1 NAND3X1_213 ( .A(core_v3_reg_18_), .B(core__abc_21302_new_n3984_), .C(core__abc_21302_new_n3988_), .Y(core__abc_21302_new_n3989_));
NAND3X1 NAND3X1_214 ( .A(core__abc_21302_new_n3979_), .B(core__abc_21302_new_n3987_), .C(core__abc_21302_new_n3989_), .Y(core__abc_21302_new_n3990_));
NAND3X1 NAND3X1_215 ( .A(core__abc_21302_new_n1410_), .B(core__abc_21302_new_n3984_), .C(core__abc_21302_new_n3988_), .Y(core__abc_21302_new_n3992_));
NAND3X1 NAND3X1_216 ( .A(core__abc_21302_new_n3978_), .B(core__abc_21302_new_n3991_), .C(core__abc_21302_new_n3992_), .Y(core__abc_21302_new_n3993_));
NAND3X1 NAND3X1_217 ( .A(core__abc_21302_new_n1596_), .B(core__abc_21302_new_n4006_), .C(core__abc_21302_new_n3984_), .Y(core__abc_21302_new_n4007_));
NAND3X1 NAND3X1_218 ( .A(core_v3_reg_19_), .B(core__abc_21302_new_n4007_), .C(core__abc_21302_new_n4009_), .Y(core__abc_21302_new_n4010_));
NAND3X1 NAND3X1_219 ( .A(core__abc_21302_new_n1596_), .B(core__abc_21302_new_n1609_), .C(core__abc_21302_new_n3984_), .Y(core__abc_21302_new_n4011_));
NAND3X1 NAND3X1_22 ( .A(core_key_35_), .B(_abc_19873_new_n889__bF_buf4), .C(_abc_19873_new_n895__bF_buf0), .Y(_abc_19873_new_n990_));
NAND3X1 NAND3X1_220 ( .A(core__abc_21302_new_n1422_), .B(core__abc_21302_new_n4011_), .C(core__abc_21302_new_n4012_), .Y(core__abc_21302_new_n4013_));
NAND3X1 NAND3X1_221 ( .A(core__abc_21302_new_n4016_), .B(core__abc_21302_new_n4010_), .C(core__abc_21302_new_n4013_), .Y(core__abc_21302_new_n4017_));
NAND3X1 NAND3X1_222 ( .A(core__abc_21302_new_n3994_), .B(core__abc_21302_new_n4017_), .C(core__abc_21302_new_n4015_), .Y(core__abc_21302_new_n4032_));
NAND3X1 NAND3X1_223 ( .A(core__abc_21302_new_n4044_), .B(core__abc_21302_new_n4047_), .C(core__abc_21302_new_n4050_), .Y(core__abc_21302_new_n4051_));
NAND3X1 NAND3X1_224 ( .A(core_v3_reg_21_), .B(core__abc_21302_new_n4068_), .C(core__abc_21302_new_n4070_), .Y(core__abc_21302_new_n4071_));
NAND3X1 NAND3X1_225 ( .A(core__abc_21302_new_n1446_), .B(core__abc_21302_new_n4072_), .C(core__abc_21302_new_n4073_), .Y(core__abc_21302_new_n4074_));
NAND3X1 NAND3X1_226 ( .A(core__abc_21302_new_n4065_), .B(core__abc_21302_new_n4074_), .C(core__abc_21302_new_n4071_), .Y(core__abc_21302_new_n4075_));
NAND3X1 NAND3X1_227 ( .A(core__abc_21302_new_n3301_), .B(core__abc_21302_new_n4081_), .C(core__abc_21302_new_n4080_), .Y(core__abc_21302_new_n4082_));
NAND3X1 NAND3X1_228 ( .A(core__abc_21302_new_n4099_), .B(core__abc_21302_new_n4106_), .C(core__abc_21302_new_n4104_), .Y(core__abc_21302_new_n4107_));
NAND3X1 NAND3X1_229 ( .A(core__abc_21302_new_n4108_), .B(core__abc_21302_new_n4110_), .C(core__abc_21302_new_n4109_), .Y(core__abc_21302_new_n4111_));
NAND3X1 NAND3X1_23 ( .A(word0_reg_4_), .B(_abc_19873_new_n905__bF_buf3), .C(_abc_19873_new_n901__bF_buf2), .Y(_abc_19873_new_n1006_));
NAND3X1 NAND3X1_230 ( .A(core__abc_21302_new_n4115_), .B(core__abc_21302_new_n4112_), .C(core__abc_21302_new_n4092_), .Y(core__abc_21302_new_n4116_));
NAND3X1 NAND3X1_231 ( .A(core_v3_reg_23_), .B(core__abc_21302_new_n4129_), .C(core__abc_21302_new_n4128_), .Y(core__abc_21302_new_n4130_));
NAND3X1 NAND3X1_232 ( .A(core__abc_21302_new_n1640_), .B(core__abc_21302_new_n1653_), .C(core__abc_21302_new_n4102_), .Y(core__abc_21302_new_n4131_));
NAND3X1 NAND3X1_233 ( .A(core__abc_21302_new_n2582_), .B(core__abc_21302_new_n4132_), .C(core__abc_21302_new_n4131_), .Y(core__abc_21302_new_n4133_));
NAND3X1 NAND3X1_234 ( .A(core__abc_21302_new_n4126_), .B(core__abc_21302_new_n4133_), .C(core__abc_21302_new_n4130_), .Y(core__abc_21302_new_n4134_));
NAND3X1 NAND3X1_235 ( .A(core__abc_21302_new_n4111_), .B(core__abc_21302_new_n4139_), .C(core__abc_21302_new_n4114_), .Y(core__abc_21302_new_n4140_));
NAND3X1 NAND3X1_236 ( .A(core__abc_21302_new_n3392_), .B(core__abc_21302_new_n4140_), .C(core__abc_21302_new_n4142_), .Y(core__abc_21302_new_n4143_));
NAND3X1 NAND3X1_237 ( .A(core__abc_21302_new_n2634__bF_buf7), .B(core__abc_21302_new_n4145_), .C(core__abc_21302_new_n4143_), .Y(core__abc_21302_new_n4146_));
NAND3X1 NAND3X1_238 ( .A(core__abc_21302_new_n4091_), .B(core__abc_21302_new_n4155_), .C(core__abc_21302_new_n4036_), .Y(core__abc_21302_new_n4156_));
NAND3X1 NAND3X1_239 ( .A(core__abc_21302_new_n3615_), .B(core__abc_21302_new_n4162_), .C(core__abc_21302_new_n3285_), .Y(core__abc_21302_new_n4163_));
NAND3X1 NAND3X1_24 ( .A(word1_reg_4_), .B(_abc_19873_new_n895__bF_buf4), .C(_abc_19873_new_n901__bF_buf1), .Y(_abc_19873_new_n1007_));
NAND3X1 NAND3X1_240 ( .A(core__abc_21302_new_n3863_), .B(core__abc_21302_new_n3764_), .C(core__abc_21302_new_n4166_), .Y(core__abc_21302_new_n4167_));
NAND3X1 NAND3X1_241 ( .A(core__abc_21302_new_n4091_), .B(core__abc_21302_new_n4037_), .C(core__abc_21302_new_n4155_), .Y(core__abc_21302_new_n4171_));
NAND3X1 NAND3X1_242 ( .A(core__abc_21302_new_n4195_), .B(core__abc_21302_new_n4199_), .C(core__abc_21302_new_n4202_), .Y(core__abc_21302_new_n4203_));
NAND3X1 NAND3X1_243 ( .A(core_v3_reg_26_), .B(core__abc_21302_new_n2624_), .C(core__abc_21302_new_n4225_), .Y(core__abc_21302_new_n4226_));
NAND3X1 NAND3X1_244 ( .A(core__abc_21302_new_n4220_), .B(core__abc_21302_new_n4226_), .C(core__abc_21302_new_n4224_), .Y(core__abc_21302_new_n4227_));
NAND3X1 NAND3X1_245 ( .A(core__abc_21302_new_n1500_), .B(core__abc_21302_new_n2624_), .C(core__abc_21302_new_n4225_), .Y(core__abc_21302_new_n4229_));
NAND3X1 NAND3X1_246 ( .A(core__abc_21302_new_n4219_), .B(core__abc_21302_new_n4229_), .C(core__abc_21302_new_n4228_), .Y(core__abc_21302_new_n4230_));
NAND3X1 NAND3X1_247 ( .A(core__abc_21302_new_n4203_), .B(core__abc_21302_new_n4206_), .C(core__abc_21302_new_n4179_), .Y(core__abc_21302_new_n4235_));
NAND3X1 NAND3X1_248 ( .A(core__abc_21302_new_n3512_), .B(core__abc_21302_new_n3515_), .C(core__abc_21302_new_n4241_), .Y(core__abc_21302_new_n4242_));
NAND3X1 NAND3X1_249 ( .A(core_v3_reg_27_), .B(core__abc_21302_new_n2629_), .C(core__abc_21302_new_n2630_), .Y(core__abc_21302_new_n4254_));
NAND3X1 NAND3X1_25 ( .A(word2_reg_4_), .B(_abc_19873_new_n901__bF_buf0), .C(_abc_19873_new_n893__bF_buf3), .Y(_abc_19873_new_n1008_));
NAND3X1 NAND3X1_250 ( .A(core__abc_21302_new_n4257_), .B(core__abc_21302_new_n4254_), .C(core__abc_21302_new_n4256_), .Y(core__abc_21302_new_n4258_));
NAND3X1 NAND3X1_251 ( .A(core__abc_21302_new_n4227_), .B(core__abc_21302_new_n4260_), .C(core__abc_21302_new_n4237_), .Y(core__abc_21302_new_n4261_));
NAND3X1 NAND3X1_252 ( .A(core__abc_21302_new_n4253_), .B(core__abc_21302_new_n4231_), .C(core__abc_21302_new_n4258_), .Y(core__abc_21302_new_n4274_));
NAND3X1 NAND3X1_253 ( .A(core__abc_21302_new_n2669_), .B(core__abc_21302_new_n4285_), .C(core__abc_21302_new_n2671_), .Y(core__abc_21302_new_n4288_));
NAND3X1 NAND3X1_254 ( .A(core__abc_21302_new_n4305_), .B(core__abc_21302_new_n4302_), .C(core__abc_21302_new_n4301_), .Y(core__abc_21302_new_n4306_));
NAND3X1 NAND3X1_255 ( .A(core__abc_21302_new_n3640_), .B(core__abc_21302_new_n4311_), .C(core__abc_21302_new_n4310_), .Y(core__abc_21302_new_n4312_));
NAND3X1 NAND3X1_256 ( .A(core__abc_21302_new_n3639_), .B(core__abc_21302_new_n4315_), .C(core__abc_21302_new_n4314_), .Y(core__abc_21302_new_n4316_));
NAND3X1 NAND3X1_257 ( .A(core__abc_21302_new_n4307_), .B(core__abc_21302_new_n4302_), .C(core__abc_21302_new_n4301_), .Y(core__abc_21302_new_n4326_));
NAND3X1 NAND3X1_258 ( .A(core__abc_21302_new_n1549_), .B(core__abc_21302_new_n2729_), .C(core__abc_21302_new_n2730_), .Y(core__abc_21302_new_n4332_));
NAND3X1 NAND3X1_259 ( .A(core__abc_21302_new_n4337_), .B(core__abc_21302_new_n4331_), .C(core__abc_21302_new_n4332_), .Y(core__abc_21302_new_n4338_));
NAND3X1 NAND3X1_26 ( .A(_abc_19873_new_n1006_), .B(_abc_19873_new_n1007_), .C(_abc_19873_new_n1008_), .Y(_abc_19873_new_n1009_));
NAND3X1 NAND3X1_260 ( .A(core__abc_21302_new_n4339_), .B(core__abc_21302_new_n2728_), .C(core__abc_21302_new_n2731_), .Y(core__abc_21302_new_n4340_));
NAND3X1 NAND3X1_261 ( .A(core__abc_21302_new_n3672_), .B(core__abc_21302_new_n4349_), .C(core__abc_21302_new_n4350_), .Y(core__abc_21302_new_n4351_));
NAND3X1 NAND3X1_262 ( .A(core_v3_reg_31_), .B(core__abc_21302_new_n2787_), .C(core__abc_21302_new_n2786_), .Y(core__abc_21302_new_n4358_));
NAND3X1 NAND3X1_263 ( .A(core__abc_21302_new_n2588_), .B(core__abc_21302_new_n2784_), .C(core__abc_21302_new_n2782_), .Y(core__abc_21302_new_n4359_));
NAND3X1 NAND3X1_264 ( .A(core__abc_21302_new_n4363_), .B(core__abc_21302_new_n4358_), .C(core__abc_21302_new_n4359_), .Y(core__abc_21302_new_n4364_));
NAND3X1 NAND3X1_265 ( .A(core__abc_21302_new_n4340_), .B(core__abc_21302_new_n4367_), .C(core__abc_21302_new_n4349_), .Y(core__abc_21302_new_n4368_));
NAND3X1 NAND3X1_266 ( .A(core__abc_21302_new_n3710_), .B(core__abc_21302_new_n4373_), .C(core__abc_21302_new_n4368_), .Y(core__abc_21302_new_n4374_));
NAND3X1 NAND3X1_267 ( .A(core__abc_21302_new_n4340_), .B(core__abc_21302_new_n4372_), .C(core__abc_21302_new_n4349_), .Y(core__abc_21302_new_n4375_));
NAND3X1 NAND3X1_268 ( .A(core__abc_21302_new_n3714_), .B(core__abc_21302_new_n4376_), .C(core__abc_21302_new_n4375_), .Y(core__abc_21302_new_n4377_));
NAND3X1 NAND3X1_269 ( .A(core__abc_21302_new_n4346_), .B(core__abc_21302_new_n4387_), .C(core__abc_21302_new_n4279_), .Y(core__abc_21302_new_n4388_));
NAND3X1 NAND3X1_27 ( .A(core_key_36_), .B(_abc_19873_new_n889__bF_buf3), .C(_abc_19873_new_n895__bF_buf3), .Y(_abc_19873_new_n1011_));
NAND3X1 NAND3X1_270 ( .A(core__abc_21302_new_n4346_), .B(core__abc_21302_new_n4387_), .C(core__abc_21302_new_n4161_), .Y(core__abc_21302_new_n4427_));
NAND3X1 NAND3X1_271 ( .A(core__abc_21302_new_n4428_), .B(core__abc_21302_new_n4393_), .C(core__abc_21302_new_n4427_), .Y(core__abc_21302_new_n4429_));
NAND3X1 NAND3X1_272 ( .A(core__abc_21302_new_n3860_), .B(core__abc_21302_new_n4456_), .C(core__abc_21302_new_n4460_), .Y(core__abc_21302_new_n4463_));
NAND3X1 NAND3X1_273 ( .A(core__abc_21302_new_n2955_), .B(core__abc_21302_new_n4474_), .C(core__abc_21302_new_n2954_), .Y(core__abc_21302_new_n4477_));
NAND3X1 NAND3X1_274 ( .A(core__abc_21302_new_n4451_), .B(core__abc_21302_new_n4478_), .C(core__abc_21302_new_n4456_), .Y(core__abc_21302_new_n4479_));
NAND3X1 NAND3X1_275 ( .A(core__abc_21302_new_n3852_), .B(core__abc_21302_new_n4481_), .C(core__abc_21302_new_n4479_), .Y(core__abc_21302_new_n4484_));
NAND3X1 NAND3X1_276 ( .A(core__abc_21302_new_n4477_), .B(core__abc_21302_new_n4453_), .C(core__abc_21302_new_n4476_), .Y(core__abc_21302_new_n4493_));
NAND3X1 NAND3X1_277 ( .A(core__abc_21302_new_n2446_), .B(core__abc_21302_new_n1443_), .C(core__abc_21302_new_n4501_), .Y(core__abc_21302_new_n4518_));
NAND3X1 NAND3X1_278 ( .A(core__abc_21302_new_n4505_), .B(core__abc_21302_new_n4525_), .C(core__abc_21302_new_n4517_), .Y(core__abc_21302_new_n4526_));
NAND3X1 NAND3X1_279 ( .A(core__abc_21302_new_n3926_), .B(core__abc_21302_new_n4526_), .C(core__abc_21302_new_n4528_), .Y(core__abc_21302_new_n4529_));
NAND3X1 NAND3X1_28 ( .A(core_mi_37_), .B(_abc_19873_new_n889__bF_buf2), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1023_));
NAND3X1 NAND3X1_280 ( .A(core__abc_21302_new_n3070_), .B(core__abc_21302_new_n4548_), .C(core__abc_21302_new_n3072_), .Y(core__abc_21302_new_n4549_));
NAND3X1 NAND3X1_281 ( .A(core__abc_21302_new_n4543_), .B(core__abc_21302_new_n4551_), .C(core__abc_21302_new_n4540_), .Y(core__abc_21302_new_n4553_));
NAND3X1 NAND3X1_282 ( .A(core__abc_21302_new_n4569_), .B(core__abc_21302_new_n1467_), .C(core__abc_21302_new_n4545_), .Y(core__abc_21302_new_n4570_));
NAND3X1 NAND3X1_283 ( .A(core__abc_21302_new_n3118_), .B(core__abc_21302_new_n4573_), .C(core__abc_21302_new_n4568_), .Y(core__abc_21302_new_n4574_));
NAND3X1 NAND3X1_284 ( .A(core__abc_21302_new_n4549_), .B(core__abc_21302_new_n4577_), .C(core__abc_21302_new_n4567_), .Y(core__abc_21302_new_n4578_));
NAND3X1 NAND3X1_285 ( .A(core__abc_21302_new_n4564_), .B(core__abc_21302_new_n4581_), .C(core__abc_21302_new_n4578_), .Y(core__abc_21302_new_n4582_));
NAND3X1 NAND3X1_286 ( .A(core__abc_21302_new_n4549_), .B(core__abc_21302_new_n4580_), .C(core__abc_21302_new_n4567_), .Y(core__abc_21302_new_n4583_));
NAND3X1 NAND3X1_287 ( .A(core__abc_21302_new_n4001_), .B(core__abc_21302_new_n4584_), .C(core__abc_21302_new_n4583_), .Y(core__abc_21302_new_n4585_));
NAND3X1 NAND3X1_288 ( .A(core__abc_21302_new_n4539_), .B(core__abc_21302_new_n4595_), .C(core__abc_21302_new_n4594_), .Y(core__abc_21302_new_n4596_));
NAND3X1 NAND3X1_289 ( .A(core__abc_21302_new_n4539_), .B(core__abc_21302_new_n4595_), .C(core__abc_21302_new_n4495_), .Y(core__abc_21302_new_n4598_));
NAND3X1 NAND3X1_29 ( .A(word2_reg_5_), .B(_abc_19873_new_n901__bF_buf7), .C(_abc_19873_new_n893__bF_buf2), .Y(_abc_19873_new_n1024_));
NAND3X1 NAND3X1_290 ( .A(core__abc_21302_new_n3118_), .B(core__abc_21302_new_n4575_), .C(core__abc_21302_new_n4568_), .Y(core__abc_21302_new_n4599_));
NAND3X1 NAND3X1_291 ( .A(core__abc_21302_new_n4052_), .B(core__abc_21302_new_n4630_), .C(core__abc_21302_new_n4633_), .Y(core__abc_21302_new_n4634_));
NAND3X1 NAND3X1_292 ( .A(core__abc_21302_new_n3214_), .B(core__abc_21302_new_n4626_), .C(core__abc_21302_new_n3211_), .Y(core__abc_21302_new_n4644_));
NAND3X1 NAND3X1_293 ( .A(core__abc_21302_new_n4609_), .B(core__abc_21302_new_n4644_), .C(core__abc_21302_new_n4643_), .Y(core__abc_21302_new_n4647_));
NAND3X1 NAND3X1_294 ( .A(core__abc_21302_new_n4652_), .B(core__abc_21302_new_n3254_), .C(core__abc_21302_new_n3251_), .Y(core__abc_21302_new_n4653_));
NAND3X1 NAND3X1_295 ( .A(core__abc_21302_new_n3246_), .B(core__abc_21302_new_n3253_), .C(core__abc_21302_new_n3252_), .Y(core__abc_21302_new_n4655_));
NAND3X1 NAND3X1_296 ( .A(core__abc_21302_new_n4651_), .B(core__abc_21302_new_n4655_), .C(core__abc_21302_new_n4654_), .Y(core__abc_21302_new_n4656_));
NAND3X1 NAND3X1_297 ( .A(core__abc_21302_new_n4646_), .B(core__abc_21302_new_n4658_), .C(core__abc_21302_new_n4649_), .Y(core__abc_21302_new_n4661_));
NAND3X1 NAND3X1_298 ( .A(core__abc_21302_new_n4664_), .B(core__abc_21302_new_n4661_), .C(core__abc_21302_new_n4660_), .Y(core__abc_21302_new_n4665_));
NAND3X1 NAND3X1_299 ( .A(core__abc_21302_new_n3311_), .B(core__abc_21302_new_n3314_), .C(core__abc_21302_new_n3315_), .Y(core__abc_21302_new_n4673_));
NAND3X1 NAND3X1_3 ( .A(word2_reg_0_), .B(_abc_19873_new_n901__bF_buf7), .C(_abc_19873_new_n893__bF_buf3), .Y(_abc_19873_new_n902_));
NAND3X1 NAND3X1_30 ( .A(word0_reg_5_), .B(_abc_19873_new_n905__bF_buf1), .C(_abc_19873_new_n901__bF_buf6), .Y(_abc_19873_new_n1025_));
NAND3X1 NAND3X1_300 ( .A(core__abc_21302_new_n4679_), .B(core__abc_21302_new_n4673_), .C(core__abc_21302_new_n4672_), .Y(core__abc_21302_new_n4680_));
NAND3X1 NAND3X1_301 ( .A(core__abc_21302_new_n4653_), .B(core__abc_21302_new_n4682_), .C(core__abc_21302_new_n4660_), .Y(core__abc_21302_new_n4683_));
NAND3X1 NAND3X1_302 ( .A(core__abc_21302_new_n4671_), .B(core__abc_21302_new_n4686_), .C(core__abc_21302_new_n4683_), .Y(core__abc_21302_new_n4687_));
NAND3X1 NAND3X1_303 ( .A(core__abc_21302_new_n4678_), .B(core__abc_21302_new_n4673_), .C(core__abc_21302_new_n4672_), .Y(core__abc_21302_new_n4699_));
NAND3X1 NAND3X1_304 ( .A(core__abc_21302_new_n4657_), .B(core__abc_21302_new_n4699_), .C(core__abc_21302_new_n4698_), .Y(core__abc_21302_new_n4700_));
NAND3X1 NAND3X1_305 ( .A(core__abc_21302_new_n3356_), .B(core__abc_21302_new_n4712_), .C(core__abc_21302_new_n3359_), .Y(core__abc_21302_new_n4713_));
NAND3X1 NAND3X1_306 ( .A(core__abc_21302_new_n4714_), .B(core__abc_21302_new_n4716_), .C(core__abc_21302_new_n4715_), .Y(core__abc_21302_new_n4717_));
NAND3X1 NAND3X1_307 ( .A(core__abc_21302_new_n4718_), .B(core__abc_21302_new_n4705_), .C(core__abc_21302_new_n4702_), .Y(core__abc_21302_new_n4720_));
NAND3X1 NAND3X1_308 ( .A(core__abc_21302_new_n2461_), .B(core__abc_21302_new_n1534_), .C(core__abc_21302_new_n4709_), .Y(core__abc_21302_new_n4741_));
NAND3X1 NAND3X1_309 ( .A(core__abc_21302_new_n4744_), .B(core__abc_21302_new_n3402_), .C(core__abc_21302_new_n3406_), .Y(core__abc_21302_new_n4745_));
NAND3X1 NAND3X1_31 ( .A(_abc_19873_new_n1025_), .B(_abc_19873_new_n1023_), .C(_abc_19873_new_n1024_), .Y(_abc_19873_new_n1026_));
NAND3X1 NAND3X1_310 ( .A(core__abc_21302_new_n4713_), .B(core__abc_21302_new_n4748_), .C(core__abc_21302_new_n4740_), .Y(core__abc_21302_new_n4749_));
NAND3X1 NAND3X1_311 ( .A(core__abc_21302_new_n4731_), .B(core__abc_21302_new_n4752_), .C(core__abc_21302_new_n4749_), .Y(core__abc_21302_new_n4753_));
NAND3X1 NAND3X1_312 ( .A(core__abc_21302_new_n4713_), .B(core__abc_21302_new_n4751_), .C(core__abc_21302_new_n4740_), .Y(core__abc_21302_new_n4754_));
NAND3X1 NAND3X1_313 ( .A(core__abc_21302_new_n4176_), .B(core__abc_21302_new_n4755_), .C(core__abc_21302_new_n4754_), .Y(core__abc_21302_new_n4756_));
NAND3X1 NAND3X1_314 ( .A(core__abc_21302_new_n3448_), .B(core__abc_21302_new_n4775_), .C(core__abc_21302_new_n3447_), .Y(core__abc_21302_new_n4776_));
NAND3X1 NAND3X1_315 ( .A(core__abc_21302_new_n4767_), .B(core__abc_21302_new_n4765_), .C(core__abc_21302_new_n4780_), .Y(core__abc_21302_new_n4781_));
NAND3X1 NAND3X1_316 ( .A(core__abc_21302_new_n4741_), .B(core__abc_21302_new_n4743_), .C(core__abc_21302_new_n3407_), .Y(core__abc_21302_new_n4782_));
NAND3X1 NAND3X1_317 ( .A(core__abc_21302_new_n4745_), .B(core__abc_21302_new_n4739_), .C(core__abc_21302_new_n4782_), .Y(core__abc_21302_new_n4783_));
NAND3X1 NAND3X1_318 ( .A(core__abc_21302_new_n4763_), .B(core__abc_21302_new_n4785_), .C(core__abc_21302_new_n4781_), .Y(core__abc_21302_new_n4786_));
NAND3X1 NAND3X1_319 ( .A(core__abc_21302_new_n4798_), .B(core__abc_21302_new_n1558_), .C(core__abc_21302_new_n4769_), .Y(core__abc_21302_new_n4799_));
NAND3X1 NAND3X1_32 ( .A(core_key_37_), .B(_abc_19873_new_n889__bF_buf1), .C(_abc_19873_new_n895__bF_buf1), .Y(_abc_19873_new_n1029_));
NAND3X1 NAND3X1_320 ( .A(core__abc_21302_new_n4799_), .B(core__abc_21302_new_n4801_), .C(core__abc_21302_new_n4804_), .Y(core__abc_21302_new_n4805_));
NAND3X1 NAND3X1_321 ( .A(core__abc_21302_new_n4797_), .B(core__abc_21302_new_n4785_), .C(core__abc_21302_new_n4806_), .Y(core__abc_21302_new_n4807_));
NAND3X1 NAND3X1_322 ( .A(core__abc_21302_new_n4795_), .B(core__abc_21302_new_n4807_), .C(core__abc_21302_new_n4809_), .Y(core__abc_21302_new_n4810_));
NAND3X1 NAND3X1_323 ( .A(core__abc_21302_new_n4797_), .B(core__abc_21302_new_n4785_), .C(core__abc_21302_new_n4808_), .Y(core__abc_21302_new_n4812_));
NAND3X1 NAND3X1_324 ( .A(core__abc_21302_new_n4811_), .B(core__abc_21302_new_n4813_), .C(core__abc_21302_new_n4812_), .Y(core__abc_21302_new_n4814_));
NAND3X1 NAND3X1_325 ( .A(core__abc_21302_new_n2634__bF_buf6), .B(core__abc_21302_new_n4810_), .C(core__abc_21302_new_n4814_), .Y(core__abc_21302_new_n4815_));
NAND3X1 NAND3X1_326 ( .A(core__abc_21302_new_n4824_), .B(core__abc_21302_new_n4799_), .C(core__abc_21302_new_n4801_), .Y(core__abc_21302_new_n4825_));
NAND3X1 NAND3X1_327 ( .A(core_v1_reg_17_), .B(core__abc_21302_new_n4769_), .C(core__abc_21302_new_n4772_), .Y(core__abc_21302_new_n4835_));
NAND3X1 NAND3X1_328 ( .A(core__abc_21302_new_n4831_), .B(core__abc_21302_new_n4837_), .C(core__abc_21302_new_n4829_), .Y(core__abc_21302_new_n4838_));
NAND3X1 NAND3X1_329 ( .A(core__abc_21302_new_n4839_), .B(core__abc_21302_new_n4842_), .C(core__abc_21302_new_n4841_), .Y(core__abc_21302_new_n4843_));
NAND3X1 NAND3X1_33 ( .A(word1_reg_6_), .B(_abc_19873_new_n895__bF_buf0), .C(_abc_19873_new_n901__bF_buf5), .Y(_abc_19873_new_n1048_));
NAND3X1 NAND3X1_330 ( .A(core__abc_21302_new_n4851_), .B(core__abc_21302_new_n4846_), .C(core__abc_21302_new_n4843_), .Y(core__abc_21302_new_n4852_));
NAND3X1 NAND3X1_331 ( .A(core__abc_21302_new_n3777_), .B(core__abc_21302_new_n4848_), .C(core__abc_21302_new_n4849_), .Y(core__abc_21302_new_n4880_));
NAND3X1 NAND3X1_332 ( .A(core__abc_21302_new_n4832_), .B(core__abc_21302_new_n4835_), .C(core__abc_21302_new_n4834_), .Y(core__abc_21302_new_n4883_));
NAND3X1 NAND3X1_333 ( .A(core__abc_21302_new_n4889_), .B(core__abc_21302_new_n4893_), .C(core__abc_21302_new_n4853_), .Y(core__abc_21302_new_n4894_));
NAND3X1 NAND3X1_334 ( .A(core__abc_21302_new_n4248_), .B(core__abc_21302_new_n4570_), .C(core__abc_21302_new_n4572_), .Y(core__abc_21302_new_n4896_));
NAND3X1 NAND3X1_335 ( .A(core__abc_21302_new_n4569_), .B(core__abc_21302_new_n4571_), .C(core__abc_21302_new_n4545_), .Y(core__abc_21302_new_n4897_));
NAND3X1 NAND3X1_336 ( .A(core_v1_reg_10_), .B(core__abc_21302_new_n4897_), .C(core__abc_21302_new_n4898_), .Y(core__abc_21302_new_n4899_));
NAND3X1 NAND3X1_337 ( .A(core__abc_21302_new_n4895_), .B(core__abc_21302_new_n4896_), .C(core__abc_21302_new_n4899_), .Y(core__abc_21302_new_n4900_));
NAND3X1 NAND3X1_338 ( .A(core_v1_reg_9_), .B(core__abc_21302_new_n4545_), .C(core__abc_21302_new_n4908_), .Y(core__abc_21302_new_n4909_));
NAND3X1 NAND3X1_339 ( .A(core__abc_21302_new_n4905_), .B(core__abc_21302_new_n4907_), .C(core__abc_21302_new_n4909_), .Y(core__abc_21302_new_n4910_));
NAND3X1 NAND3X1_34 ( .A(word2_reg_6_), .B(_abc_19873_new_n901__bF_buf4), .C(_abc_19873_new_n893__bF_buf1), .Y(_abc_19873_new_n1049_));
NAND3X1 NAND3X1_340 ( .A(core__abc_21302_new_n4906_), .B(core__abc_21302_new_n4545_), .C(core__abc_21302_new_n4908_), .Y(core__abc_21302_new_n4913_));
NAND3X1 NAND3X1_341 ( .A(core__abc_21302_new_n4911_), .B(core__abc_21302_new_n4912_), .C(core__abc_21302_new_n4913_), .Y(core__abc_21302_new_n4914_));
NAND3X1 NAND3X1_342 ( .A(core__abc_21302_new_n4900_), .B(core__abc_21302_new_n4915_), .C(core__abc_21302_new_n4904_), .Y(core__abc_21302_new_n4916_));
NAND3X1 NAND3X1_343 ( .A(core__abc_21302_new_n3514_), .B(core__abc_21302_new_n4919_), .C(core__abc_21302_new_n4918_), .Y(core__abc_21302_new_n4920_));
NAND3X1 NAND3X1_344 ( .A(core__abc_21302_new_n4926_), .B(core__abc_21302_new_n4923_), .C(core__abc_21302_new_n4920_), .Y(core__abc_21302_new_n4927_));
NAND3X1 NAND3X1_345 ( .A(core__abc_21302_new_n4938_), .B(core__abc_21302_new_n4934_), .C(core__abc_21302_new_n4939_), .Y(core__abc_21302_new_n4940_));
NAND3X1 NAND3X1_346 ( .A(core__abc_21302_new_n3233_), .B(core__abc_21302_new_n4964_), .C(core__abc_21302_new_n4965_), .Y(core__abc_21302_new_n4966_));
NAND3X1 NAND3X1_347 ( .A(core__abc_21302_new_n4966_), .B(core__abc_21302_new_n4974_), .C(core__abc_21302_new_n4968_), .Y(core__abc_21302_new_n4975_));
NAND3X1 NAND3X1_348 ( .A(core__abc_21302_new_n5028_), .B(core__abc_21302_new_n5020_), .C(core__abc_21302_new_n5023_), .Y(core__abc_21302_new_n5029_));
NAND3X1 NAND3X1_349 ( .A(core__abc_21302_new_n2651_), .B(core__abc_21302_new_n5043_), .C(core__abc_21302_new_n5044_), .Y(core__abc_21302_new_n5049_));
NAND3X1 NAND3X1_35 ( .A(word0_reg_6_), .B(_abc_19873_new_n905__bF_buf0), .C(_abc_19873_new_n901__bF_buf3), .Y(_abc_19873_new_n1050_));
NAND3X1 NAND3X1_350 ( .A(core__abc_21302_new_n5059_), .B(core__abc_21302_new_n5062_), .C(core__abc_21302_new_n5009_), .Y(core__abc_21302_new_n5063_));
NAND3X1 NAND3X1_351 ( .A(core__abc_21302_new_n4931_), .B(core__abc_21302_new_n5068_), .C(core__abc_21302_new_n4941_), .Y(core__abc_21302_new_n5069_));
NAND3X1 NAND3X1_352 ( .A(core__abc_21302_new_n4866_), .B(core__abc_21302_new_n4893_), .C(core__abc_21302_new_n4861_), .Y(core__abc_21302_new_n5091_));
NAND3X1 NAND3X1_353 ( .A(core__abc_21302_new_n5111_), .B(core__abc_21302_new_n5114_), .C(core__abc_21302_new_n5118_), .Y(core__abc_21302_new_n5119_));
NAND3X1 NAND3X1_354 ( .A(core__abc_21302_new_n5135_), .B(core__abc_21302_new_n5137_), .C(core__abc_21302_new_n5138_), .Y(core__abc_21302_new_n5139_));
NAND3X1 NAND3X1_355 ( .A(core__abc_21302_new_n5139_), .B(core__abc_21302_new_n5120_), .C(core__abc_21302_new_n5143_), .Y(core__abc_21302_new_n5158_));
NAND3X1 NAND3X1_356 ( .A(core__abc_21302_new_n4068_), .B(core__abc_21302_new_n4070_), .C(core__abc_21302_new_n5176_), .Y(core__abc_21302_new_n5177_));
NAND3X1 NAND3X1_357 ( .A(core__abc_21302_new_n4072_), .B(core__abc_21302_new_n4073_), .C(core__abc_21302_new_n5178_), .Y(core__abc_21302_new_n5179_));
NAND3X1 NAND3X1_358 ( .A(core__abc_21302_new_n5207_), .B(core__abc_21302_new_n5214_), .C(core__abc_21302_new_n5213_), .Y(core__abc_21302_new_n5215_));
NAND3X1 NAND3X1_359 ( .A(core__abc_21302_new_n5194_), .B(core__abc_21302_new_n5226_), .C(core__abc_21302_new_n5161_), .Y(core__abc_21302_new_n5227_));
NAND3X1 NAND3X1_36 ( .A(_abc_19873_new_n1050_), .B(_abc_19873_new_n1048_), .C(_abc_19873_new_n1049_), .Y(_abc_19873_new_n1051_));
NAND3X1 NAND3X1_360 ( .A(core__abc_21302_new_n5226_), .B(core__abc_21302_new_n5194_), .C(core__abc_21302_new_n5159_), .Y(core__abc_21302_new_n5229_));
NAND3X1 NAND3X1_361 ( .A(core__abc_21302_new_n4201_), .B(core__abc_21302_new_n5250_), .C(core__abc_21302_new_n5249_), .Y(core__abc_21302_new_n5251_));
NAND3X1 NAND3X1_362 ( .A(core__abc_21302_new_n4255_), .B(core__abc_21302_new_n5288_), .C(core__abc_21302_new_n5287_), .Y(core__abc_21302_new_n5289_));
NAND3X1 NAND3X1_363 ( .A(core__abc_21302_new_n5274_), .B(core__abc_21302_new_n5292_), .C(core__abc_21302_new_n5289_), .Y(core__abc_21302_new_n5303_));
NAND3X1 NAND3X1_364 ( .A(core__abc_21302_new_n5322_), .B(core__abc_21302_new_n5343_), .C(core__abc_21302_new_n5342_), .Y(core__abc_21302_new_n5346_));
NAND3X1 NAND3X1_365 ( .A(core_v1_reg_33_), .B(core__abc_21302_new_n3199_), .C(core__abc_21302_new_n3200_), .Y(core__abc_21302_new_n5350_));
NAND3X1 NAND3X1_366 ( .A(core__abc_21302_new_n5358_), .B(core__abc_21302_new_n5360_), .C(core__abc_21302_new_n5359_), .Y(core__abc_21302_new_n5361_));
NAND3X1 NAND3X1_367 ( .A(core__abc_21302_new_n5355_), .B(core__abc_21302_new_n5376_), .C(core__abc_21302_new_n5357_), .Y(core__abc_21302_new_n5377_));
NAND3X1 NAND3X1_368 ( .A(core__abc_21302_new_n5388_), .B(core__abc_21302_new_n5347_), .C(core__abc_21302_new_n5307_), .Y(core__abc_21302_new_n5389_));
NAND3X1 NAND3X1_369 ( .A(core__abc_21302_new_n5390_), .B(core__abc_21302_new_n5394_), .C(core__abc_21302_new_n5389_), .Y(core__abc_21302_new_n5395_));
NAND3X1 NAND3X1_37 ( .A(core_key_70_), .B(_abc_19873_new_n889__bF_buf0), .C(_abc_19873_new_n893__bF_buf0), .Y(_abc_19873_new_n1053_));
NAND3X1 NAND3X1_370 ( .A(core__abc_21302_new_n5393_), .B(core__abc_21302_new_n5356_), .C(core__abc_21302_new_n5391_), .Y(core__abc_21302_new_n5400_));
NAND3X1 NAND3X1_371 ( .A(core__abc_21302_new_n5399_), .B(core__abc_21302_new_n5228_), .C(core__abc_21302_new_n5401_), .Y(core__abc_21302_new_n5402_));
NAND3X1 NAND3X1_372 ( .A(core__abc_21302_new_n5399_), .B(core__abc_21302_new_n5401_), .C(core__abc_21302_new_n5234_), .Y(core__abc_21302_new_n5416_));
NAND3X1 NAND3X1_373 ( .A(core__abc_21302_new_n5389_), .B(core__abc_21302_new_n5415_), .C(core__abc_21302_new_n5416_), .Y(core__abc_21302_new_n5417_));
NAND3X1 NAND3X1_374 ( .A(core__abc_21302_new_n2634__bF_buf4), .B(core__abc_21302_new_n5446_), .C(core__abc_21302_new_n5448_), .Y(core__abc_21302_new_n5449_));
NAND3X1 NAND3X1_375 ( .A(core__abc_21302_new_n5482_), .B(core__abc_21302_new_n5496_), .C(core__abc_21302_new_n5492_), .Y(core__abc_21302_new_n5497_));
NAND3X1 NAND3X1_376 ( .A(core__abc_21302_new_n5513_), .B(core__abc_21302_new_n5518_), .C(core__abc_21302_new_n5516_), .Y(core__abc_21302_new_n5521_));
NAND3X1 NAND3X1_377 ( .A(core__abc_21302_new_n3113_), .B(core__abc_21302_new_n3115_), .C(core__abc_21302_new_n5532_), .Y(core__abc_21302_new_n5533_));
NAND3X1 NAND3X1_378 ( .A(core__abc_21302_new_n5510_), .B(core__abc_21302_new_n5534_), .C(core__abc_21302_new_n5520_), .Y(core__abc_21302_new_n5535_));
NAND3X1 NAND3X1_379 ( .A(core__abc_21302_new_n2634__bF_buf2), .B(core__abc_21302_new_n5538_), .C(core__abc_21302_new_n5535_), .Y(core__abc_21302_new_n5539_));
NAND3X1 NAND3X1_38 ( .A(word1_reg_7_), .B(_abc_19873_new_n895__bF_buf4), .C(_abc_19873_new_n901__bF_buf1), .Y(_abc_19873_new_n1067_));
NAND3X1 NAND3X1_380 ( .A(core__abc_21302_new_n2634__bF_buf1), .B(core__abc_21302_new_n5577_), .C(core__abc_21302_new_n5575_), .Y(core__abc_21302_new_n5578_));
NAND3X1 NAND3X1_381 ( .A(core__abc_21302_new_n5587_), .B(core__abc_21302_new_n5591_), .C(core__abc_21302_new_n5590_), .Y(core__abc_21302_new_n5594_));
NAND3X1 NAND3X1_382 ( .A(core__abc_21302_new_n3314_), .B(core__abc_21302_new_n5603_), .C(core__abc_21302_new_n3315_), .Y(core__abc_21302_new_n5604_));
NAND3X1 NAND3X1_383 ( .A(core__abc_21302_new_n5585_), .B(core__abc_21302_new_n5607_), .C(core__abc_21302_new_n5593_), .Y(core__abc_21302_new_n5608_));
NAND3X1 NAND3X1_384 ( .A(core__abc_21302_new_n2634__bF_buf0), .B(core__abc_21302_new_n5611_), .C(core__abc_21302_new_n5608_), .Y(core__abc_21302_new_n5612_));
NAND3X1 NAND3X1_385 ( .A(core__abc_21302_new_n5624_), .B(core__abc_21302_new_n5629_), .C(core__abc_21302_new_n5620_), .Y(core__abc_21302_new_n5630_));
NAND3X1 NAND3X1_386 ( .A(core__abc_21302_new_n5674_), .B(core__abc_21302_new_n5666_), .C(core__abc_21302_new_n5664_), .Y(core__abc_21302_new_n5675_));
NAND3X1 NAND3X1_387 ( .A(core__abc_21302_new_n5684_), .B(core__abc_21302_new_n5689_), .C(core__abc_21302_new_n5676_), .Y(core__abc_21302_new_n5690_));
NAND3X1 NAND3X1_388 ( .A(core__abc_21302_new_n2634__bF_buf8), .B(core__abc_21302_new_n5692_), .C(core__abc_21302_new_n5690_), .Y(core__abc_21302_new_n5693_));
NAND3X1 NAND3X1_389 ( .A(core__abc_21302_new_n5013_), .B(core__abc_21302_new_n5060_), .C(core__abc_21302_new_n5059_), .Y(core__abc_21302_new_n5773_));
NAND3X1 NAND3X1_39 ( .A(word2_reg_7_), .B(_abc_19873_new_n901__bF_buf0), .C(_abc_19873_new_n893__bF_buf4), .Y(_abc_19873_new_n1068_));
NAND3X1 NAND3X1_390 ( .A(core__abc_21302_new_n2634__bF_buf6), .B(core__abc_21302_new_n5954_), .C(core__abc_21302_new_n5958_), .Y(core__abc_21302_new_n5959_));
NAND3X1 NAND3X1_391 ( .A(core__abc_21302_new_n5965_), .B(core__abc_21302_new_n4880_), .C(core__abc_21302_new_n5954_), .Y(core__abc_21302_new_n5966_));
NAND3X1 NAND3X1_392 ( .A(core__abc_21302_new_n2634__bF_buf5), .B(core__abc_21302_new_n5701_), .C(core__abc_21302_new_n5373_), .Y(core__abc_21302_new_n6002_));
NAND3X1 NAND3X1_393 ( .A(core__abc_21302_new_n2634__bF_buf5), .B(core__abc_21302_new_n6139_), .C(core__abc_21302_new_n6140_), .Y(core__abc_21302_new_n6141_));
NAND3X1 NAND3X1_394 ( .A(core__abc_21302_new_n2634__bF_buf3), .B(core__abc_21302_new_n6168_), .C(core__abc_21302_new_n6167_), .Y(core__abc_21302_new_n6169_));
NAND3X1 NAND3X1_395 ( .A(core__abc_21302_new_n4999_), .B(core__abc_21302_new_n5954_), .C(core__abc_21302_new_n5958_), .Y(core__abc_21302_new_n6194_));
NAND3X1 NAND3X1_396 ( .A(core__abc_21302_new_n2634__bF_buf1), .B(core__abc_21302_new_n6195_), .C(core__abc_21302_new_n6194_), .Y(core__abc_21302_new_n6196_));
NAND3X1 NAND3X1_397 ( .A(core__abc_21302_new_n2634__bF_buf0), .B(core__abc_21302_new_n6220_), .C(core__abc_21302_new_n6221_), .Y(core__abc_21302_new_n6222_));
NAND3X1 NAND3X1_398 ( .A(core__abc_21302_new_n2634__bF_buf8), .B(core__abc_21302_new_n6258_), .C(core__abc_21302_new_n6259_), .Y(core__abc_21302_new_n6260_));
NAND3X1 NAND3X1_399 ( .A(core__abc_21302_new_n6265_), .B(core__abc_21302_new_n5219_), .C(core__abc_21302_new_n5217_), .Y(core__abc_21302_new_n6266_));
NAND3X1 NAND3X1_4 ( .A(word0_reg_0_), .B(_abc_19873_new_n905__bF_buf3), .C(_abc_19873_new_n901__bF_buf6), .Y(_abc_19873_new_n906_));
NAND3X1 NAND3X1_40 ( .A(word3_reg_7_), .B(_abc_19873_new_n912__bF_buf0), .C(_abc_19873_new_n901__bF_buf7), .Y(_abc_19873_new_n1069_));
NAND3X1 NAND3X1_400 ( .A(core__abc_21302_new_n4907_), .B(core__abc_21302_new_n4909_), .C(core__abc_21302_new_n6267_), .Y(core__abc_21302_new_n6268_));
NAND3X1 NAND3X1_401 ( .A(core__abc_21302_new_n2634__bF_buf7), .B(core__abc_21302_new_n6266_), .C(core__abc_21302_new_n6268_), .Y(core__abc_21302_new_n6269_));
NAND3X1 NAND3X1_402 ( .A(core__abc_21302_new_n2634__bF_buf5), .B(core__abc_21302_new_n6301_), .C(core__abc_21302_new_n6302_), .Y(core__abc_21302_new_n6303_));
NAND3X1 NAND3X1_403 ( .A(core__abc_21302_new_n4850_), .B(core__abc_21302_new_n5334_), .C(core__abc_21302_new_n5335_), .Y(core__abc_21302_new_n6309_));
NAND3X1 NAND3X1_404 ( .A(core__abc_21302_new_n4848_), .B(core__abc_21302_new_n4849_), .C(core__abc_21302_new_n5336_), .Y(core__abc_21302_new_n6310_));
NAND3X1 NAND3X1_405 ( .A(core__abc_21302_new_n2634__bF_buf4), .B(core__abc_21302_new_n6309_), .C(core__abc_21302_new_n6310_), .Y(core__abc_21302_new_n6311_));
NAND3X1 NAND3X1_406 ( .A(core__abc_21302_new_n5089_), .B(core__abc_21302_new_n5446_), .C(core__abc_21302_new_n5448_), .Y(core__abc_21302_new_n6344_));
NAND3X1 NAND3X1_407 ( .A(core__abc_21302_new_n2634__bF_buf2), .B(core__abc_21302_new_n6346_), .C(core__abc_21302_new_n6344_), .Y(core__abc_21302_new_n6347_));
NAND3X1 NAND3X1_408 ( .A(core__abc_21302_new_n5510_), .B(core__abc_21302_new_n5537_), .C(core__abc_21302_new_n5520_), .Y(core__abc_21302_new_n6378_));
NAND3X1 NAND3X1_409 ( .A(core__abc_21302_new_n5188_), .B(core__abc_21302_new_n6379_), .C(core__abc_21302_new_n6378_), .Y(core__abc_21302_new_n6380_));
NAND3X1 NAND3X1_41 ( .A(_abc_19873_new_n1069_), .B(_abc_19873_new_n1067_), .C(_abc_19873_new_n1068_), .Y(_abc_19873_new_n1070_));
NAND3X1 NAND3X1_410 ( .A(core__abc_21302_new_n5190_), .B(core__abc_21302_new_n5538_), .C(core__abc_21302_new_n5535_), .Y(core__abc_21302_new_n6381_));
NAND3X1 NAND3X1_411 ( .A(core__abc_21302_new_n2634__bF_buf0), .B(core__abc_21302_new_n6380_), .C(core__abc_21302_new_n6381_), .Y(core__abc_21302_new_n6382_));
NAND3X1 NAND3X1_412 ( .A(core__abc_21302_new_n6393_), .B(core__abc_21302_new_n5577_), .C(core__abc_21302_new_n5575_), .Y(core__abc_21302_new_n6394_));
NAND3X1 NAND3X1_413 ( .A(core__abc_21302_new_n5585_), .B(core__abc_21302_new_n5610_), .C(core__abc_21302_new_n5593_), .Y(core__abc_21302_new_n6408_));
NAND3X1 NAND3X1_414 ( .A(core__abc_21302_new_n5271_), .B(core__abc_21302_new_n6409_), .C(core__abc_21302_new_n6408_), .Y(core__abc_21302_new_n6410_));
NAND3X1 NAND3X1_415 ( .A(core__abc_21302_new_n6411_), .B(core__abc_21302_new_n5611_), .C(core__abc_21302_new_n5608_), .Y(core__abc_21302_new_n6412_));
NAND3X1 NAND3X1_416 ( .A(core__abc_21302_new_n2634__bF_buf8), .B(core__abc_21302_new_n6410_), .C(core__abc_21302_new_n6412_), .Y(core__abc_21302_new_n6413_));
NAND3X1 NAND3X1_417 ( .A(core__abc_21302_new_n5354_), .B(core__abc_21302_new_n5692_), .C(core__abc_21302_new_n5690_), .Y(core__abc_21302_new_n6439_));
NAND3X1 NAND3X1_418 ( .A(core__abc_21302_new_n5684_), .B(core__abc_21302_new_n5688_), .C(core__abc_21302_new_n5676_), .Y(core__abc_21302_new_n6441_));
NAND3X1 NAND3X1_419 ( .A(core__abc_21302_new_n5351_), .B(core__abc_21302_new_n6440_), .C(core__abc_21302_new_n6441_), .Y(core__abc_21302_new_n6442_));
NAND3X1 NAND3X1_42 ( .A(core_key_71_), .B(_abc_19873_new_n889__bF_buf4), .C(_abc_19873_new_n893__bF_buf3), .Y(_abc_19873_new_n1072_));
NAND3X1 NAND3X1_420 ( .A(core__abc_21302_new_n2634__bF_buf7), .B(core__abc_21302_new_n6439_), .C(core__abc_21302_new_n6442_), .Y(core__abc_21302_new_n6443_));
NAND3X1 NAND3X1_421 ( .A(reset_n_bF_buf44), .B(core__abc_21302_new_n1175_), .C(core__abc_21302_new_n1179_), .Y(core__abc_21302_new_n6906_));
NAND3X1 NAND3X1_43 ( .A(word3_reg_11_), .B(_abc_19873_new_n912__bF_buf3), .C(_abc_19873_new_n901__bF_buf6), .Y(_abc_19873_new_n1143_));
NAND3X1 NAND3X1_44 ( .A(word2_reg_11_), .B(_abc_19873_new_n901__bF_buf5), .C(_abc_19873_new_n893__bF_buf2), .Y(_abc_19873_new_n1144_));
NAND3X1 NAND3X1_45 ( .A(word1_reg_11_), .B(_abc_19873_new_n895__bF_buf2), .C(_abc_19873_new_n901__bF_buf4), .Y(_abc_19873_new_n1145_));
NAND3X1 NAND3X1_46 ( .A(_abc_19873_new_n1143_), .B(_abc_19873_new_n1144_), .C(_abc_19873_new_n1145_), .Y(_abc_19873_new_n1146_));
NAND3X1 NAND3X1_47 ( .A(core_key_43_), .B(_abc_19873_new_n889__bF_buf3), .C(_abc_19873_new_n895__bF_buf1), .Y(_abc_19873_new_n1148_));
NAND3X1 NAND3X1_48 ( .A(word1_reg_12_), .B(_abc_19873_new_n895__bF_buf0), .C(_abc_19873_new_n901__bF_buf3), .Y(_abc_19873_new_n1162_));
NAND3X1 NAND3X1_49 ( .A(word2_reg_12_), .B(_abc_19873_new_n901__bF_buf2), .C(_abc_19873_new_n893__bF_buf0), .Y(_abc_19873_new_n1163_));
NAND3X1 NAND3X1_5 ( .A(_abc_19873_new_n906_), .B(_abc_19873_new_n898_), .C(_abc_19873_new_n902_), .Y(_abc_19873_new_n907_));
NAND3X1 NAND3X1_50 ( .A(word3_reg_12_), .B(_abc_19873_new_n912__bF_buf2), .C(_abc_19873_new_n901__bF_buf1), .Y(_abc_19873_new_n1164_));
NAND3X1 NAND3X1_51 ( .A(_abc_19873_new_n1164_), .B(_abc_19873_new_n1162_), .C(_abc_19873_new_n1163_), .Y(_abc_19873_new_n1165_));
NAND3X1 NAND3X1_52 ( .A(core_key_44_), .B(_abc_19873_new_n889__bF_buf2), .C(_abc_19873_new_n895__bF_buf4), .Y(_abc_19873_new_n1167_));
NAND3X1 NAND3X1_53 ( .A(word0_reg_13_), .B(_abc_19873_new_n905__bF_buf1), .C(_abc_19873_new_n901__bF_buf0), .Y(_abc_19873_new_n1186_));
NAND3X1 NAND3X1_54 ( .A(word1_reg_13_), .B(_abc_19873_new_n895__bF_buf3), .C(_abc_19873_new_n901__bF_buf7), .Y(_abc_19873_new_n1187_));
NAND3X1 NAND3X1_55 ( .A(word3_reg_13_), .B(_abc_19873_new_n912__bF_buf1), .C(_abc_19873_new_n901__bF_buf6), .Y(_abc_19873_new_n1188_));
NAND3X1 NAND3X1_56 ( .A(_abc_19873_new_n1186_), .B(_abc_19873_new_n1188_), .C(_abc_19873_new_n1187_), .Y(_abc_19873_new_n1189_));
NAND3X1 NAND3X1_57 ( .A(core_mi_46_), .B(_abc_19873_new_n889__bF_buf1), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1199_));
NAND3X1 NAND3X1_58 ( .A(word1_reg_14_), .B(_abc_19873_new_n895__bF_buf2), .C(_abc_19873_new_n901__bF_buf5), .Y(_abc_19873_new_n1201_));
NAND3X1 NAND3X1_59 ( .A(word2_reg_14_), .B(_abc_19873_new_n901__bF_buf4), .C(_abc_19873_new_n893__bF_buf4), .Y(_abc_19873_new_n1202_));
NAND3X1 NAND3X1_6 ( .A(core_key_0_), .B(_abc_19873_new_n905__bF_buf2), .C(_abc_19873_new_n889__bF_buf4), .Y(_abc_19873_new_n919_));
NAND3X1 NAND3X1_60 ( .A(word3_reg_14_), .B(_abc_19873_new_n912__bF_buf0), .C(_abc_19873_new_n901__bF_buf3), .Y(_abc_19873_new_n1203_));
NAND3X1 NAND3X1_61 ( .A(_abc_19873_new_n1203_), .B(_abc_19873_new_n1201_), .C(_abc_19873_new_n1202_), .Y(_abc_19873_new_n1204_));
NAND3X1 NAND3X1_62 ( .A(core_mi_48_), .B(_abc_19873_new_n889__bF_buf0), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1236_));
NAND3X1 NAND3X1_63 ( .A(word1_reg_16_), .B(_abc_19873_new_n895__bF_buf1), .C(_abc_19873_new_n901__bF_buf2), .Y(_abc_19873_new_n1238_));
NAND3X1 NAND3X1_64 ( .A(word2_reg_16_), .B(_abc_19873_new_n901__bF_buf1), .C(_abc_19873_new_n893__bF_buf3), .Y(_abc_19873_new_n1239_));
NAND3X1 NAND3X1_65 ( .A(word3_reg_16_), .B(_abc_19873_new_n912__bF_buf3), .C(_abc_19873_new_n901__bF_buf0), .Y(_abc_19873_new_n1240_));
NAND3X1 NAND3X1_66 ( .A(_abc_19873_new_n1240_), .B(_abc_19873_new_n1238_), .C(_abc_19873_new_n1239_), .Y(_abc_19873_new_n1241_));
NAND3X1 NAND3X1_67 ( .A(word1_reg_17_), .B(_abc_19873_new_n895__bF_buf4), .C(_abc_19873_new_n901__bF_buf7), .Y(_abc_19873_new_n1257_));
NAND3X1 NAND3X1_68 ( .A(word2_reg_17_), .B(_abc_19873_new_n901__bF_buf6), .C(_abc_19873_new_n893__bF_buf1), .Y(_abc_19873_new_n1258_));
NAND3X1 NAND3X1_69 ( .A(word3_reg_17_), .B(_abc_19873_new_n912__bF_buf2), .C(_abc_19873_new_n901__bF_buf5), .Y(_abc_19873_new_n1259_));
NAND3X1 NAND3X1_7 ( .A(core_siphash_valid_reg), .B(_abc_19873_new_n877_), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n931_));
NAND3X1 NAND3X1_70 ( .A(_abc_19873_new_n1259_), .B(_abc_19873_new_n1257_), .C(_abc_19873_new_n1258_), .Y(_abc_19873_new_n1260_));
NAND3X1 NAND3X1_71 ( .A(core_mi_17_), .B(_abc_19873_new_n889__bF_buf4), .C(_abc_19873_new_n874_), .Y(_abc_19873_new_n1262_));
NAND3X1 NAND3X1_72 ( .A(word3_reg_18_), .B(_abc_19873_new_n912__bF_buf1), .C(_abc_19873_new_n901__bF_buf4), .Y(_abc_19873_new_n1272_));
NAND3X1 NAND3X1_73 ( .A(word2_reg_18_), .B(_abc_19873_new_n901__bF_buf3), .C(_abc_19873_new_n893__bF_buf0), .Y(_abc_19873_new_n1273_));
NAND3X1 NAND3X1_74 ( .A(word1_reg_18_), .B(_abc_19873_new_n895__bF_buf3), .C(_abc_19873_new_n901__bF_buf2), .Y(_abc_19873_new_n1274_));
NAND3X1 NAND3X1_75 ( .A(_abc_19873_new_n1272_), .B(_abc_19873_new_n1273_), .C(_abc_19873_new_n1274_), .Y(_abc_19873_new_n1275_));
NAND3X1 NAND3X1_76 ( .A(core_key_50_), .B(_abc_19873_new_n889__bF_buf3), .C(_abc_19873_new_n895__bF_buf2), .Y(_abc_19873_new_n1277_));
NAND3X1 NAND3X1_77 ( .A(core_mi_51_), .B(_abc_19873_new_n889__bF_buf2), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1291_));
NAND3X1 NAND3X1_78 ( .A(word1_reg_19_), .B(_abc_19873_new_n895__bF_buf1), .C(_abc_19873_new_n901__bF_buf1), .Y(_abc_19873_new_n1293_));
NAND3X1 NAND3X1_79 ( .A(word2_reg_19_), .B(_abc_19873_new_n901__bF_buf0), .C(_abc_19873_new_n893__bF_buf4), .Y(_abc_19873_new_n1294_));
NAND3X1 NAND3X1_8 ( .A(core_mi_33_), .B(_abc_19873_new_n889__bF_buf3), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n936_));
NAND3X1 NAND3X1_80 ( .A(word3_reg_19_), .B(_abc_19873_new_n912__bF_buf0), .C(_abc_19873_new_n901__bF_buf7), .Y(_abc_19873_new_n1295_));
NAND3X1 NAND3X1_81 ( .A(_abc_19873_new_n1295_), .B(_abc_19873_new_n1293_), .C(_abc_19873_new_n1294_), .Y(_abc_19873_new_n1296_));
NAND3X1 NAND3X1_82 ( .A(word3_reg_20_), .B(_abc_19873_new_n912__bF_buf3), .C(_abc_19873_new_n901__bF_buf6), .Y(_abc_19873_new_n1308_));
NAND3X1 NAND3X1_83 ( .A(word2_reg_20_), .B(_abc_19873_new_n901__bF_buf5), .C(_abc_19873_new_n893__bF_buf3), .Y(_abc_19873_new_n1309_));
NAND3X1 NAND3X1_84 ( .A(word1_reg_20_), .B(_abc_19873_new_n895__bF_buf0), .C(_abc_19873_new_n901__bF_buf4), .Y(_abc_19873_new_n1310_));
NAND3X1 NAND3X1_85 ( .A(_abc_19873_new_n1308_), .B(_abc_19873_new_n1309_), .C(_abc_19873_new_n1310_), .Y(_abc_19873_new_n1311_));
NAND3X1 NAND3X1_86 ( .A(core_key_52_), .B(_abc_19873_new_n889__bF_buf1), .C(_abc_19873_new_n895__bF_buf4), .Y(_abc_19873_new_n1313_));
NAND3X1 NAND3X1_87 ( .A(word3_reg_21_), .B(_abc_19873_new_n912__bF_buf2), .C(_abc_19873_new_n901__bF_buf3), .Y(_abc_19873_new_n1332_));
NAND3X1 NAND3X1_88 ( .A(word1_reg_21_), .B(_abc_19873_new_n895__bF_buf3), .C(_abc_19873_new_n901__bF_buf2), .Y(_abc_19873_new_n1333_));
NAND3X1 NAND3X1_89 ( .A(word0_reg_21_), .B(_abc_19873_new_n905__bF_buf0), .C(_abc_19873_new_n901__bF_buf1), .Y(_abc_19873_new_n1334_));
NAND3X1 NAND3X1_9 ( .A(word2_reg_1_), .B(_abc_19873_new_n901__bF_buf3), .C(_abc_19873_new_n893__bF_buf2), .Y(_abc_19873_new_n937_));
NAND3X1 NAND3X1_90 ( .A(_abc_19873_new_n1332_), .B(_abc_19873_new_n1334_), .C(_abc_19873_new_n1333_), .Y(_abc_19873_new_n1335_));
NAND3X1 NAND3X1_91 ( .A(core_mi_54_), .B(_abc_19873_new_n889__bF_buf0), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1345_));
NAND3X1 NAND3X1_92 ( .A(word1_reg_22_), .B(_abc_19873_new_n895__bF_buf2), .C(_abc_19873_new_n901__bF_buf0), .Y(_abc_19873_new_n1347_));
NAND3X1 NAND3X1_93 ( .A(word2_reg_22_), .B(_abc_19873_new_n901__bF_buf7), .C(_abc_19873_new_n893__bF_buf2), .Y(_abc_19873_new_n1348_));
NAND3X1 NAND3X1_94 ( .A(word3_reg_22_), .B(_abc_19873_new_n912__bF_buf1), .C(_abc_19873_new_n901__bF_buf6), .Y(_abc_19873_new_n1349_));
NAND3X1 NAND3X1_95 ( .A(_abc_19873_new_n1349_), .B(_abc_19873_new_n1347_), .C(_abc_19873_new_n1348_), .Y(_abc_19873_new_n1350_));
NAND3X1 NAND3X1_96 ( .A(core_mi_56_), .B(_abc_19873_new_n889__bF_buf4), .C(_abc_19873_new_n881_), .Y(_abc_19873_new_n1382_));
NAND3X1 NAND3X1_97 ( .A(word1_reg_24_), .B(_abc_19873_new_n895__bF_buf1), .C(_abc_19873_new_n901__bF_buf5), .Y(_abc_19873_new_n1384_));
NAND3X1 NAND3X1_98 ( .A(word2_reg_24_), .B(_abc_19873_new_n901__bF_buf4), .C(_abc_19873_new_n893__bF_buf1), .Y(_abc_19873_new_n1385_));
NAND3X1 NAND3X1_99 ( .A(word3_reg_24_), .B(_abc_19873_new_n912__bF_buf0), .C(_abc_19873_new_n901__bF_buf3), .Y(_abc_19873_new_n1386_));
NOR2X1 NOR2X1_1 ( .A(_abc_19873_new_n871_), .B(_abc_19873_new_n873_), .Y(_abc_19873_new_n874_));
NOR2X1 NOR2X1_10 ( .A(\addr[0] ), .B(\addr[1] ), .Y(_abc_19873_new_n904_));
NOR2X1 NOR2X1_100 ( .A(core_v1_reg_11_), .B(core_v0_reg_11_), .Y(core__abc_21302_new_n1324_));
NOR2X1 NOR2X1_101 ( .A(core__abc_21302_new_n1324_), .B(core__abc_21302_new_n1325_), .Y(core__abc_21302_new_n1326_));
NOR2X1 NOR2X1_102 ( .A(core_v1_reg_13_), .B(core_v0_reg_13_), .Y(core__abc_21302_new_n1346_));
NOR2X1 NOR2X1_103 ( .A(core__abc_21302_new_n1346_), .B(core__abc_21302_new_n1347_), .Y(core__abc_21302_new_n1348_));
NOR2X1 NOR2X1_104 ( .A(core_v1_reg_14_), .B(core_v0_reg_14_), .Y(core__abc_21302_new_n1358_));
NOR2X1 NOR2X1_105 ( .A(core__abc_21302_new_n1358_), .B(core__abc_21302_new_n1359_), .Y(core__abc_21302_new_n1360_));
NOR2X1 NOR2X1_106 ( .A(core_v1_reg_15_), .B(core_v0_reg_15_), .Y(core__abc_21302_new_n1370_));
NOR2X1 NOR2X1_107 ( .A(core__abc_21302_new_n1370_), .B(core__abc_21302_new_n1371_), .Y(core__abc_21302_new_n1372_));
NOR2X1 NOR2X1_108 ( .A(core__abc_21302_new_n1373_), .B(core__abc_21302_new_n1374_), .Y(core__abc_21302_new_n1375_));
NOR2X1 NOR2X1_109 ( .A(core_v2_reg_15_), .B(core_v3_reg_15_), .Y(core__abc_21302_new_n1376_));
NOR2X1 NOR2X1_11 ( .A(_abc_19873_new_n911_), .B(_abc_19873_new_n890_), .Y(_abc_19873_new_n912_));
NOR2X1 NOR2X1_110 ( .A(core__abc_21302_new_n1376_), .B(core__abc_21302_new_n1375_), .Y(core__abc_21302_new_n1377_));
NOR2X1 NOR2X1_111 ( .A(core_v1_reg_16_), .B(core_v0_reg_16_), .Y(core__abc_21302_new_n1382_));
NOR2X1 NOR2X1_112 ( .A(core_v2_reg_16_), .B(core_v3_reg_16_), .Y(core__abc_21302_new_n1387_));
NOR2X1 NOR2X1_113 ( .A(core__abc_21302_new_n1387_), .B(core__abc_21302_new_n1386_), .Y(core__abc_21302_new_n1388_));
NOR2X1 NOR2X1_114 ( .A(core_v1_reg_17_), .B(core_v0_reg_17_), .Y(core__abc_21302_new_n1393_));
NOR2X1 NOR2X1_115 ( .A(core_v1_reg_18_), .B(core_v0_reg_18_), .Y(core__abc_21302_new_n1405_));
NOR2X1 NOR2X1_116 ( .A(core__abc_21302_new_n1405_), .B(core__abc_21302_new_n1406_), .Y(core__abc_21302_new_n1407_));
NOR2X1 NOR2X1_117 ( .A(core_v1_reg_19_), .B(core_v0_reg_19_), .Y(core__abc_21302_new_n1417_));
NOR2X1 NOR2X1_118 ( .A(core__abc_21302_new_n1417_), .B(core__abc_21302_new_n1418_), .Y(core__abc_21302_new_n1419_));
NOR2X1 NOR2X1_119 ( .A(core_v1_reg_20_), .B(core_v0_reg_20_), .Y(core__abc_21302_new_n1429_));
NOR2X1 NOR2X1_12 ( .A(_abc_19873_new_n911_), .B(_abc_19873_new_n873_), .Y(_abc_19873_new_n917_));
NOR2X1 NOR2X1_120 ( .A(core__abc_21302_new_n1429_), .B(core__abc_21302_new_n1430_), .Y(core__abc_21302_new_n1431_));
NOR2X1 NOR2X1_121 ( .A(core_v1_reg_21_), .B(core_v0_reg_21_), .Y(core__abc_21302_new_n1441_));
NOR2X1 NOR2X1_122 ( .A(core__abc_21302_new_n1441_), .B(core__abc_21302_new_n1442_), .Y(core__abc_21302_new_n1443_));
NOR2X1 NOR2X1_123 ( .A(core_v1_reg_22_), .B(core_v0_reg_22_), .Y(core__abc_21302_new_n1453_));
NOR2X1 NOR2X1_124 ( .A(core__abc_21302_new_n1453_), .B(core__abc_21302_new_n1454_), .Y(core__abc_21302_new_n1455_));
NOR2X1 NOR2X1_125 ( .A(core_v1_reg_23_), .B(core_v0_reg_23_), .Y(core__abc_21302_new_n1465_));
NOR2X1 NOR2X1_126 ( .A(core__abc_21302_new_n1465_), .B(core__abc_21302_new_n1466_), .Y(core__abc_21302_new_n1467_));
NOR2X1 NOR2X1_127 ( .A(core_v1_reg_24_), .B(core_v0_reg_24_), .Y(core__abc_21302_new_n1473_));
NOR2X1 NOR2X1_128 ( .A(core__abc_21302_new_n1473_), .B(core__abc_21302_new_n1474_), .Y(core__abc_21302_new_n1475_));
NOR2X1 NOR2X1_129 ( .A(core__abc_21302_new_n1476_), .B(core__abc_21302_new_n1477_), .Y(core__abc_21302_new_n1478_));
NOR2X1 NOR2X1_13 ( .A(_abc_19873_new_n952_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n954_));
NOR2X1 NOR2X1_130 ( .A(core_v2_reg_24_), .B(core_v3_reg_24_), .Y(core__abc_21302_new_n1479_));
NOR2X1 NOR2X1_131 ( .A(core__abc_21302_new_n1479_), .B(core__abc_21302_new_n1478_), .Y(core__abc_21302_new_n1480_));
NOR2X1 NOR2X1_132 ( .A(core_v1_reg_26_), .B(core_v0_reg_26_), .Y(core__abc_21302_new_n1495_));
NOR2X1 NOR2X1_133 ( .A(core__abc_21302_new_n1495_), .B(core__abc_21302_new_n1496_), .Y(core__abc_21302_new_n1497_));
NOR2X1 NOR2X1_134 ( .A(core_v1_reg_27_), .B(core_v0_reg_27_), .Y(core__abc_21302_new_n1507_));
NOR2X1 NOR2X1_135 ( .A(core__abc_21302_new_n1507_), .B(core__abc_21302_new_n1508_), .Y(core__abc_21302_new_n1509_));
NOR2X1 NOR2X1_136 ( .A(core_v1_reg_28_), .B(core_v0_reg_28_), .Y(core__abc_21302_new_n1519_));
NOR2X1 NOR2X1_137 ( .A(core__abc_21302_new_n1519_), .B(core__abc_21302_new_n1520_), .Y(core__abc_21302_new_n1521_));
NOR2X1 NOR2X1_138 ( .A(core_v1_reg_29_), .B(core_v0_reg_29_), .Y(core__abc_21302_new_n1531_));
NOR2X1 NOR2X1_139 ( .A(core__abc_21302_new_n1531_), .B(core__abc_21302_new_n1533_), .Y(core__abc_21302_new_n1534_));
NOR2X1 NOR2X1_14 ( .A(_abc_19873_new_n976_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n977_));
NOR2X1 NOR2X1_140 ( .A(core_v1_reg_30_), .B(core_v0_reg_30_), .Y(core__abc_21302_new_n1544_));
NOR2X1 NOR2X1_141 ( .A(core__abc_21302_new_n1544_), .B(core__abc_21302_new_n1545_), .Y(core__abc_21302_new_n1546_));
NOR2X1 NOR2X1_142 ( .A(core_v1_reg_31_), .B(core_v0_reg_31_), .Y(core__abc_21302_new_n1556_));
NOR2X1 NOR2X1_143 ( .A(core__abc_21302_new_n1556_), .B(core__abc_21302_new_n1557_), .Y(core__abc_21302_new_n1558_));
NOR2X1 NOR2X1_144 ( .A(core_v1_reg_32_), .B(core_v0_reg_32_), .Y(core__abc_21302_new_n1564_));
NOR2X1 NOR2X1_145 ( .A(core__abc_21302_new_n1564_), .B(core__abc_21302_new_n1566_), .Y(core__abc_21302_new_n1567_));
NOR2X1 NOR2X1_146 ( .A(core_v2_reg_32_), .B(core_v3_reg_32_), .Y(core__abc_21302_new_n1570_));
NOR2X1 NOR2X1_147 ( .A(core_v1_reg_35_), .B(core_v0_reg_35_), .Y(core__abc_21302_new_n1602_));
NOR2X1 NOR2X1_148 ( .A(core_v1_reg_36_), .B(core_v0_reg_36_), .Y(core__abc_21302_new_n1614_));
NOR2X1 NOR2X1_149 ( .A(core__abc_21302_new_n1614_), .B(core__abc_21302_new_n1615_), .Y(core__abc_21302_new_n1616_));
NOR2X1 NOR2X1_15 ( .A(_abc_19873_new_n997_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n998_));
NOR2X1 NOR2X1_150 ( .A(core_v2_reg_36_), .B(core_v3_reg_36_), .Y(core__abc_21302_new_n1617_));
NOR2X1 NOR2X1_151 ( .A(core_v2_reg_37_), .B(core_v3_reg_37_), .Y(core__abc_21302_new_n1632_));
NOR2X1 NOR2X1_152 ( .A(core_v2_reg_38_), .B(core_v3_reg_38_), .Y(core__abc_21302_new_n1639_));
NOR2X1 NOR2X1_153 ( .A(core_v1_reg_39_), .B(core_v0_reg_39_), .Y(core__abc_21302_new_n1647_));
NOR2X1 NOR2X1_154 ( .A(core_v2_reg_39_), .B(core_v3_reg_39_), .Y(core__abc_21302_new_n1652_));
NOR2X1 NOR2X1_155 ( .A(core_v1_reg_40_), .B(core_v0_reg_40_), .Y(core__abc_21302_new_n1658_));
NOR2X1 NOR2X1_156 ( .A(core__abc_21302_new_n1658_), .B(core__abc_21302_new_n1659_), .Y(core__abc_21302_new_n1660_));
NOR2X1 NOR2X1_157 ( .A(core_v2_reg_40_), .B(core_v3_reg_40_), .Y(core__abc_21302_new_n1663_));
NOR2X1 NOR2X1_158 ( .A(core_v1_reg_41_), .B(core_v0_reg_41_), .Y(core__abc_21302_new_n1669_));
NOR2X1 NOR2X1_159 ( .A(core__abc_21302_new_n1669_), .B(core__abc_21302_new_n1670_), .Y(core__abc_21302_new_n1671_));
NOR2X1 NOR2X1_16 ( .A(_abc_19873_new_n1039_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1040_));
NOR2X1 NOR2X1_160 ( .A(core_v2_reg_41_), .B(core_v3_reg_41_), .Y(core__abc_21302_new_n1674_));
NOR2X1 NOR2X1_161 ( .A(core_v1_reg_42_), .B(core_v0_reg_42_), .Y(core__abc_21302_new_n1680_));
NOR2X1 NOR2X1_162 ( .A(core__abc_21302_new_n1680_), .B(core__abc_21302_new_n1681_), .Y(core__abc_21302_new_n1682_));
NOR2X1 NOR2X1_163 ( .A(core_v2_reg_42_), .B(core_v3_reg_42_), .Y(core__abc_21302_new_n1685_));
NOR2X1 NOR2X1_164 ( .A(core__abc_21302_new_n1685_), .B(core__abc_21302_new_n1684_), .Y(core__abc_21302_new_n1686_));
NOR2X1 NOR2X1_165 ( .A(core_v1_reg_43_), .B(core_v0_reg_43_), .Y(core__abc_21302_new_n1691_));
NOR2X1 NOR2X1_166 ( .A(core__abc_21302_new_n1691_), .B(core__abc_21302_new_n1692_), .Y(core__abc_21302_new_n1693_));
NOR2X1 NOR2X1_167 ( .A(core_v2_reg_43_), .B(core_v3_reg_43_), .Y(core__abc_21302_new_n1694_));
NOR2X1 NOR2X1_168 ( .A(core__abc_21302_new_n1694_), .B(core__abc_21302_new_n1696_), .Y(core__abc_21302_new_n1697_));
NOR2X1 NOR2X1_169 ( .A(core_v1_reg_44_), .B(core_v0_reg_44_), .Y(core__abc_21302_new_n1702_));
NOR2X1 NOR2X1_17 ( .A(_abc_19873_new_n1061_), .B(_abc_19873_new_n1065_), .Y(_abc_19873_new_n1066_));
NOR2X1 NOR2X1_170 ( .A(core__abc_21302_new_n1702_), .B(core__abc_21302_new_n1704_), .Y(core__abc_21302_new_n1705_));
NOR2X1 NOR2X1_171 ( .A(core_v2_reg_44_), .B(core_v3_reg_44_), .Y(core__abc_21302_new_n1706_));
NOR2X1 NOR2X1_172 ( .A(core__abc_21302_new_n1706_), .B(core__abc_21302_new_n1708_), .Y(core__abc_21302_new_n1709_));
NOR2X1 NOR2X1_173 ( .A(core_v2_reg_45_), .B(core_v3_reg_45_), .Y(core__abc_21302_new_n1717_));
NOR2X1 NOR2X1_174 ( .A(core__abc_21302_new_n1717_), .B(core__abc_21302_new_n1719_), .Y(core__abc_21302_new_n1720_));
NOR2X1 NOR2X1_175 ( .A(core_v1_reg_46_), .B(core_v0_reg_46_), .Y(core__abc_21302_new_n1725_));
NOR2X1 NOR2X1_176 ( .A(core__abc_21302_new_n1725_), .B(core__abc_21302_new_n1727_), .Y(core__abc_21302_new_n1728_));
NOR2X1 NOR2X1_177 ( .A(core_v2_reg_46_), .B(core_v3_reg_46_), .Y(core__abc_21302_new_n1729_));
NOR2X1 NOR2X1_178 ( .A(core_v1_reg_47_), .B(core_v0_reg_47_), .Y(core__abc_21302_new_n1737_));
NOR2X1 NOR2X1_179 ( .A(core__abc_21302_new_n1737_), .B(core__abc_21302_new_n1738_), .Y(core__abc_21302_new_n1739_));
NOR2X1 NOR2X1_18 ( .A(_abc_19873_new_n1079_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1080_));
NOR2X1 NOR2X1_180 ( .A(core_v2_reg_47_), .B(core_v3_reg_47_), .Y(core__abc_21302_new_n1740_));
NOR2X1 NOR2X1_181 ( .A(core_v1_reg_48_), .B(core_v0_reg_48_), .Y(core__abc_21302_new_n1748_));
NOR2X1 NOR2X1_182 ( .A(core__abc_21302_new_n1748_), .B(core__abc_21302_new_n1750_), .Y(core__abc_21302_new_n1751_));
NOR2X1 NOR2X1_183 ( .A(core_v2_reg_48_), .B(core_v3_reg_48_), .Y(core__abc_21302_new_n1752_));
NOR2X1 NOR2X1_184 ( .A(core__abc_21302_new_n1753_), .B(core__abc_21302_new_n1754_), .Y(core__abc_21302_new_n1755_));
NOR2X1 NOR2X1_185 ( .A(core__abc_21302_new_n1752_), .B(core__abc_21302_new_n1755_), .Y(core__abc_21302_new_n1756_));
NOR2X1 NOR2X1_186 ( .A(core_v2_reg_49_), .B(core_v3_reg_49_), .Y(core__abc_21302_new_n1762_));
NOR2X1 NOR2X1_187 ( .A(core__abc_21302_new_n1763_), .B(core__abc_21302_new_n1764_), .Y(core__abc_21302_new_n1765_));
NOR2X1 NOR2X1_188 ( .A(core__abc_21302_new_n1762_), .B(core__abc_21302_new_n1765_), .Y(core__abc_21302_new_n1766_));
NOR2X1 NOR2X1_189 ( .A(core_v1_reg_50_), .B(core_v0_reg_50_), .Y(core__abc_21302_new_n1770_));
NOR2X1 NOR2X1_19 ( .A(_abc_19873_new_n1088_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1089_));
NOR2X1 NOR2X1_190 ( .A(core__abc_21302_new_n1770_), .B(core__abc_21302_new_n1772_), .Y(core__abc_21302_new_n1773_));
NOR2X1 NOR2X1_191 ( .A(core_v2_reg_50_), .B(core_v3_reg_50_), .Y(core__abc_21302_new_n1774_));
NOR2X1 NOR2X1_192 ( .A(core__abc_21302_new_n1774_), .B(core__abc_21302_new_n1776_), .Y(core__abc_21302_new_n1777_));
NOR2X1 NOR2X1_193 ( .A(core_v1_reg_51_), .B(core_v0_reg_51_), .Y(core__abc_21302_new_n1782_));
NOR2X1 NOR2X1_194 ( .A(core__abc_21302_new_n1782_), .B(core__abc_21302_new_n1784_), .Y(core__abc_21302_new_n1785_));
NOR2X1 NOR2X1_195 ( .A(core_v2_reg_51_), .B(core_v3_reg_51_), .Y(core__abc_21302_new_n1786_));
NOR2X1 NOR2X1_196 ( .A(core__abc_21302_new_n1786_), .B(core__abc_21302_new_n1787_), .Y(core__abc_21302_new_n1788_));
NOR2X1 NOR2X1_197 ( .A(core_v1_reg_52_), .B(core_v0_reg_52_), .Y(core__abc_21302_new_n1793_));
NOR2X1 NOR2X1_198 ( .A(core__abc_21302_new_n1794_), .B(core__abc_21302_new_n1795_), .Y(core__abc_21302_new_n1796_));
NOR2X1 NOR2X1_199 ( .A(core__abc_21302_new_n1793_), .B(core__abc_21302_new_n1796_), .Y(core__abc_21302_new_n1797_));
NOR2X1 NOR2X1_2 ( .A(\addr[7] ), .B(\addr[6] ), .Y(_abc_19873_new_n875_));
NOR2X1 NOR2X1_20 ( .A(_abc_19873_new_n1098_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1099_));
NOR2X1 NOR2X1_200 ( .A(core_v2_reg_52_), .B(core_v3_reg_52_), .Y(core__abc_21302_new_n1798_));
NOR2X1 NOR2X1_201 ( .A(core__abc_21302_new_n1799_), .B(core__abc_21302_new_n1800_), .Y(core__abc_21302_new_n1801_));
NOR2X1 NOR2X1_202 ( .A(core__abc_21302_new_n1798_), .B(core__abc_21302_new_n1801_), .Y(core__abc_21302_new_n1802_));
NOR2X1 NOR2X1_203 ( .A(core__abc_21302_new_n1807_), .B(core__abc_21302_new_n1808_), .Y(core__abc_21302_new_n1809_));
NOR2X1 NOR2X1_204 ( .A(core_v1_reg_53_), .B(core_v0_reg_53_), .Y(core__abc_21302_new_n1810_));
NOR2X1 NOR2X1_205 ( .A(core__abc_21302_new_n1810_), .B(core__abc_21302_new_n1809_), .Y(core__abc_21302_new_n1811_));
NOR2X1 NOR2X1_206 ( .A(core_v2_reg_53_), .B(core_v3_reg_53_), .Y(core__abc_21302_new_n1812_));
NOR2X1 NOR2X1_207 ( .A(core__abc_21302_new_n1812_), .B(core__abc_21302_new_n1813_), .Y(core__abc_21302_new_n1814_));
NOR2X1 NOR2X1_208 ( .A(core_v1_reg_54_), .B(core_v0_reg_54_), .Y(core__abc_21302_new_n1818_));
NOR2X1 NOR2X1_209 ( .A(core__abc_21302_new_n1818_), .B(core__abc_21302_new_n1820_), .Y(core__abc_21302_new_n1821_));
NOR2X1 NOR2X1_21 ( .A(_abc_19873_new_n1107_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1108_));
NOR2X1 NOR2X1_210 ( .A(core_v2_reg_54_), .B(core_v3_reg_54_), .Y(core__abc_21302_new_n1822_));
NOR2X1 NOR2X1_211 ( .A(core__abc_21302_new_n1823_), .B(core__abc_21302_new_n1824_), .Y(core__abc_21302_new_n1825_));
NOR2X1 NOR2X1_212 ( .A(core__abc_21302_new_n1822_), .B(core__abc_21302_new_n1825_), .Y(core__abc_21302_new_n1826_));
NOR2X1 NOR2X1_213 ( .A(core_v1_reg_55_), .B(core_v0_reg_55_), .Y(core__abc_21302_new_n1831_));
NOR2X1 NOR2X1_214 ( .A(core__abc_21302_new_n1831_), .B(core__abc_21302_new_n1833_), .Y(core__abc_21302_new_n1834_));
NOR2X1 NOR2X1_215 ( .A(core_v2_reg_55_), .B(core_v3_reg_55_), .Y(core__abc_21302_new_n1835_));
NOR2X1 NOR2X1_216 ( .A(core__abc_21302_new_n1836_), .B(core__abc_21302_new_n1837_), .Y(core__abc_21302_new_n1838_));
NOR2X1 NOR2X1_217 ( .A(core__abc_21302_new_n1835_), .B(core__abc_21302_new_n1838_), .Y(core__abc_21302_new_n1839_));
NOR2X1 NOR2X1_218 ( .A(core_v1_reg_56_), .B(core_v0_reg_56_), .Y(core__abc_21302_new_n1844_));
NOR2X1 NOR2X1_219 ( .A(core__abc_21302_new_n1845_), .B(core__abc_21302_new_n1846_), .Y(core__abc_21302_new_n1847_));
NOR2X1 NOR2X1_22 ( .A(_abc_19873_new_n1117_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1118_));
NOR2X1 NOR2X1_220 ( .A(core__abc_21302_new_n1844_), .B(core__abc_21302_new_n1847_), .Y(core__abc_21302_new_n1848_));
NOR2X1 NOR2X1_221 ( .A(core_v2_reg_56_), .B(core_v3_reg_56_), .Y(core__abc_21302_new_n1849_));
NOR2X1 NOR2X1_222 ( .A(core__abc_21302_new_n1850_), .B(core__abc_21302_new_n1851_), .Y(core__abc_21302_new_n1852_));
NOR2X1 NOR2X1_223 ( .A(core__abc_21302_new_n1849_), .B(core__abc_21302_new_n1852_), .Y(core__abc_21302_new_n1853_));
NOR2X1 NOR2X1_224 ( .A(core_v1_reg_57_), .B(core_v0_reg_57_), .Y(core__abc_21302_new_n1858_));
NOR2X1 NOR2X1_225 ( .A(core__abc_21302_new_n1858_), .B(core__abc_21302_new_n1860_), .Y(core__abc_21302_new_n1861_));
NOR2X1 NOR2X1_226 ( .A(core_v2_reg_57_), .B(core_v3_reg_57_), .Y(core__abc_21302_new_n1862_));
NOR2X1 NOR2X1_227 ( .A(core__abc_21302_new_n1862_), .B(core__abc_21302_new_n1864_), .Y(core__abc_21302_new_n1865_));
NOR2X1 NOR2X1_228 ( .A(core_v1_reg_58_), .B(core_v0_reg_58_), .Y(core__abc_21302_new_n1870_));
NOR2X1 NOR2X1_229 ( .A(core__abc_21302_new_n1871_), .B(core__abc_21302_new_n1872_), .Y(core__abc_21302_new_n1873_));
NOR2X1 NOR2X1_23 ( .A(_abc_19873_new_n1126_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1127_));
NOR2X1 NOR2X1_230 ( .A(core__abc_21302_new_n1870_), .B(core__abc_21302_new_n1873_), .Y(core__abc_21302_new_n1874_));
NOR2X1 NOR2X1_231 ( .A(core_v2_reg_58_), .B(core_v3_reg_58_), .Y(core__abc_21302_new_n1875_));
NOR2X1 NOR2X1_232 ( .A(core__abc_21302_new_n1876_), .B(core__abc_21302_new_n1877_), .Y(core__abc_21302_new_n1878_));
NOR2X1 NOR2X1_233 ( .A(core__abc_21302_new_n1875_), .B(core__abc_21302_new_n1878_), .Y(core__abc_21302_new_n1879_));
NOR2X1 NOR2X1_234 ( .A(core_v1_reg_59_), .B(core_v0_reg_59_), .Y(core__abc_21302_new_n1884_));
NOR2X1 NOR2X1_235 ( .A(core__abc_21302_new_n1884_), .B(core__abc_21302_new_n1886_), .Y(core__abc_21302_new_n1887_));
NOR2X1 NOR2X1_236 ( .A(core_v2_reg_59_), .B(core_v3_reg_59_), .Y(core__abc_21302_new_n1888_));
NOR2X1 NOR2X1_237 ( .A(core__abc_21302_new_n1888_), .B(core__abc_21302_new_n1890_), .Y(core__abc_21302_new_n1891_));
NOR2X1 NOR2X1_238 ( .A(core_v1_reg_60_), .B(core_v0_reg_60_), .Y(core__abc_21302_new_n1896_));
NOR2X1 NOR2X1_239 ( .A(core__abc_21302_new_n1897_), .B(core__abc_21302_new_n1898_), .Y(core__abc_21302_new_n1899_));
NOR2X1 NOR2X1_24 ( .A(_abc_19873_new_n1141_), .B(_abc_19873_new_n1138_), .Y(_abc_19873_new_n1142_));
NOR2X1 NOR2X1_240 ( .A(core__abc_21302_new_n1896_), .B(core__abc_21302_new_n1899_), .Y(core__abc_21302_new_n1900_));
NOR2X1 NOR2X1_241 ( .A(core_v2_reg_60_), .B(core_v3_reg_60_), .Y(core__abc_21302_new_n1901_));
NOR2X1 NOR2X1_242 ( .A(core__abc_21302_new_n1902_), .B(core__abc_21302_new_n1903_), .Y(core__abc_21302_new_n1904_));
NOR2X1 NOR2X1_243 ( .A(core__abc_21302_new_n1901_), .B(core__abc_21302_new_n1904_), .Y(core__abc_21302_new_n1905_));
NOR2X1 NOR2X1_244 ( .A(core_v1_reg_61_), .B(core_v0_reg_61_), .Y(core__abc_21302_new_n1910_));
NOR2X1 NOR2X1_245 ( .A(core__abc_21302_new_n1911_), .B(core__abc_21302_new_n1912_), .Y(core__abc_21302_new_n1913_));
NOR2X1 NOR2X1_246 ( .A(core__abc_21302_new_n1910_), .B(core__abc_21302_new_n1913_), .Y(core__abc_21302_new_n1914_));
NOR2X1 NOR2X1_247 ( .A(core_v2_reg_61_), .B(core_v3_reg_61_), .Y(core__abc_21302_new_n1915_));
NOR2X1 NOR2X1_248 ( .A(core__abc_21302_new_n1916_), .B(core__abc_21302_new_n1917_), .Y(core__abc_21302_new_n1918_));
NOR2X1 NOR2X1_249 ( .A(core__abc_21302_new_n1915_), .B(core__abc_21302_new_n1918_), .Y(core__abc_21302_new_n1919_));
NOR2X1 NOR2X1_25 ( .A(_abc_19873_new_n1160_), .B(_abc_19873_new_n1157_), .Y(_abc_19873_new_n1161_));
NOR2X1 NOR2X1_250 ( .A(core_v1_reg_62_), .B(core_v0_reg_62_), .Y(core__abc_21302_new_n1924_));
NOR2X1 NOR2X1_251 ( .A(core__abc_21302_new_n1924_), .B(core__abc_21302_new_n1926_), .Y(core__abc_21302_new_n1927_));
NOR2X1 NOR2X1_252 ( .A(core_v2_reg_62_), .B(core_v3_reg_62_), .Y(core__abc_21302_new_n1928_));
NOR2X1 NOR2X1_253 ( .A(core__abc_21302_new_n1929_), .B(core__abc_21302_new_n1930_), .Y(core__abc_21302_new_n1931_));
NOR2X1 NOR2X1_254 ( .A(core__abc_21302_new_n1928_), .B(core__abc_21302_new_n1931_), .Y(core__abc_21302_new_n1932_));
NOR2X1 NOR2X1_255 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_ctrl_reg_2_), .Y(core__abc_21302_new_n1943_));
NOR2X1 NOR2X1_256 ( .A(core__abc_21302_new_n1944_), .B(core__abc_21302_new_n1155_), .Y(core__abc_21302_new_n1945_));
NOR2X1 NOR2X1_257 ( .A(core__abc_21302_new_n1185__bF_buf10), .B(core__abc_21302_new_n1947_), .Y(core__0siphash_word0_reg_63_0__0_));
NOR2X1 NOR2X1_258 ( .A(core__abc_21302_new_n1185__bF_buf9), .B(core__abc_21302_new_n1950_), .Y(core__0siphash_word0_reg_63_0__1_));
NOR2X1 NOR2X1_259 ( .A(core__abc_21302_new_n1185__bF_buf8), .B(core__abc_21302_new_n1953_), .Y(core__0siphash_word0_reg_63_0__2_));
NOR2X1 NOR2X1_26 ( .A(_abc_19873_new_n1177_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1178_));
NOR2X1 NOR2X1_260 ( .A(core__abc_21302_new_n1185__bF_buf7), .B(core__abc_21302_new_n1956_), .Y(core__0siphash_word0_reg_63_0__3_));
NOR2X1 NOR2X1_261 ( .A(core__abc_21302_new_n1185__bF_buf6), .B(core__abc_21302_new_n1959_), .Y(core__0siphash_word0_reg_63_0__4_));
NOR2X1 NOR2X1_262 ( .A(core__abc_21302_new_n1185__bF_buf5), .B(core__abc_21302_new_n1962_), .Y(core__0siphash_word0_reg_63_0__5_));
NOR2X1 NOR2X1_263 ( .A(core__abc_21302_new_n1185__bF_buf4), .B(core__abc_21302_new_n1965_), .Y(core__0siphash_word0_reg_63_0__6_));
NOR2X1 NOR2X1_264 ( .A(core__abc_21302_new_n1185__bF_buf3), .B(core__abc_21302_new_n1968_), .Y(core__0siphash_word0_reg_63_0__7_));
NOR2X1 NOR2X1_265 ( .A(core__abc_21302_new_n1185__bF_buf2), .B(core__abc_21302_new_n1971_), .Y(core__0siphash_word0_reg_63_0__8_));
NOR2X1 NOR2X1_266 ( .A(core__abc_21302_new_n1185__bF_buf1), .B(core__abc_21302_new_n1974_), .Y(core__0siphash_word0_reg_63_0__9_));
NOR2X1 NOR2X1_267 ( .A(core__abc_21302_new_n1185__bF_buf0), .B(core__abc_21302_new_n1977_), .Y(core__0siphash_word0_reg_63_0__10_));
NOR2X1 NOR2X1_268 ( .A(core__abc_21302_new_n1185__bF_buf13), .B(core__abc_21302_new_n1980_), .Y(core__0siphash_word0_reg_63_0__11_));
NOR2X1 NOR2X1_269 ( .A(core__abc_21302_new_n1185__bF_buf12), .B(core__abc_21302_new_n1983_), .Y(core__0siphash_word0_reg_63_0__12_));
NOR2X1 NOR2X1_27 ( .A(_abc_19873_new_n1196_), .B(_abc_19873_new_n1194_), .Y(_abc_19873_new_n1197_));
NOR2X1 NOR2X1_270 ( .A(core__abc_21302_new_n1185__bF_buf11), .B(core__abc_21302_new_n1986_), .Y(core__0siphash_word0_reg_63_0__13_));
NOR2X1 NOR2X1_271 ( .A(core__abc_21302_new_n1185__bF_buf10), .B(core__abc_21302_new_n1989_), .Y(core__0siphash_word0_reg_63_0__14_));
NOR2X1 NOR2X1_272 ( .A(core__abc_21302_new_n1185__bF_buf9), .B(core__abc_21302_new_n1992_), .Y(core__0siphash_word0_reg_63_0__15_));
NOR2X1 NOR2X1_273 ( .A(core__abc_21302_new_n1185__bF_buf8), .B(core__abc_21302_new_n1995_), .Y(core__0siphash_word0_reg_63_0__16_));
NOR2X1 NOR2X1_274 ( .A(core__abc_21302_new_n1185__bF_buf7), .B(core__abc_21302_new_n1998_), .Y(core__0siphash_word0_reg_63_0__17_));
NOR2X1 NOR2X1_275 ( .A(core__abc_21302_new_n1185__bF_buf6), .B(core__abc_21302_new_n2001_), .Y(core__0siphash_word0_reg_63_0__18_));
NOR2X1 NOR2X1_276 ( .A(core__abc_21302_new_n1185__bF_buf5), .B(core__abc_21302_new_n2004_), .Y(core__0siphash_word0_reg_63_0__19_));
NOR2X1 NOR2X1_277 ( .A(core__abc_21302_new_n1185__bF_buf4), .B(core__abc_21302_new_n2007_), .Y(core__0siphash_word0_reg_63_0__20_));
NOR2X1 NOR2X1_278 ( .A(core__abc_21302_new_n1185__bF_buf3), .B(core__abc_21302_new_n2010_), .Y(core__0siphash_word0_reg_63_0__21_));
NOR2X1 NOR2X1_279 ( .A(core__abc_21302_new_n1185__bF_buf2), .B(core__abc_21302_new_n2013_), .Y(core__0siphash_word0_reg_63_0__22_));
NOR2X1 NOR2X1_28 ( .A(_abc_19873_new_n1210_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1211_));
NOR2X1 NOR2X1_280 ( .A(core__abc_21302_new_n1185__bF_buf1), .B(core__abc_21302_new_n2016_), .Y(core__0siphash_word0_reg_63_0__23_));
NOR2X1 NOR2X1_281 ( .A(core__abc_21302_new_n1185__bF_buf0), .B(core__abc_21302_new_n2019_), .Y(core__0siphash_word0_reg_63_0__24_));
NOR2X1 NOR2X1_282 ( .A(core__abc_21302_new_n1185__bF_buf13), .B(core__abc_21302_new_n2022_), .Y(core__0siphash_word0_reg_63_0__25_));
NOR2X1 NOR2X1_283 ( .A(core__abc_21302_new_n1185__bF_buf12), .B(core__abc_21302_new_n2025_), .Y(core__0siphash_word0_reg_63_0__26_));
NOR2X1 NOR2X1_284 ( .A(core__abc_21302_new_n1185__bF_buf11), .B(core__abc_21302_new_n2028_), .Y(core__0siphash_word0_reg_63_0__27_));
NOR2X1 NOR2X1_285 ( .A(core__abc_21302_new_n1185__bF_buf10), .B(core__abc_21302_new_n2031_), .Y(core__0siphash_word0_reg_63_0__28_));
NOR2X1 NOR2X1_286 ( .A(core__abc_21302_new_n1185__bF_buf9), .B(core__abc_21302_new_n2034_), .Y(core__0siphash_word0_reg_63_0__29_));
NOR2X1 NOR2X1_287 ( .A(core__abc_21302_new_n1185__bF_buf8), .B(core__abc_21302_new_n2037_), .Y(core__0siphash_word0_reg_63_0__30_));
NOR2X1 NOR2X1_288 ( .A(core__abc_21302_new_n1185__bF_buf7), .B(core__abc_21302_new_n2040_), .Y(core__0siphash_word0_reg_63_0__31_));
NOR2X1 NOR2X1_289 ( .A(core__abc_21302_new_n1185__bF_buf6), .B(core__abc_21302_new_n2043_), .Y(core__0siphash_word0_reg_63_0__32_));
NOR2X1 NOR2X1_29 ( .A(_abc_19873_new_n1219_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1220_));
NOR2X1 NOR2X1_290 ( .A(core__abc_21302_new_n1185__bF_buf5), .B(core__abc_21302_new_n2046_), .Y(core__0siphash_word0_reg_63_0__33_));
NOR2X1 NOR2X1_291 ( .A(core__abc_21302_new_n1185__bF_buf4), .B(core__abc_21302_new_n2049_), .Y(core__0siphash_word0_reg_63_0__34_));
NOR2X1 NOR2X1_292 ( .A(core__abc_21302_new_n1185__bF_buf3), .B(core__abc_21302_new_n2052_), .Y(core__0siphash_word0_reg_63_0__35_));
NOR2X1 NOR2X1_293 ( .A(core__abc_21302_new_n1185__bF_buf2), .B(core__abc_21302_new_n2055_), .Y(core__0siphash_word0_reg_63_0__36_));
NOR2X1 NOR2X1_294 ( .A(core__abc_21302_new_n1185__bF_buf1), .B(core__abc_21302_new_n2058_), .Y(core__0siphash_word0_reg_63_0__37_));
NOR2X1 NOR2X1_295 ( .A(core__abc_21302_new_n1185__bF_buf0), .B(core__abc_21302_new_n2061_), .Y(core__0siphash_word0_reg_63_0__38_));
NOR2X1 NOR2X1_296 ( .A(core__abc_21302_new_n1185__bF_buf13), .B(core__abc_21302_new_n2064_), .Y(core__0siphash_word0_reg_63_0__39_));
NOR2X1 NOR2X1_297 ( .A(core__abc_21302_new_n1185__bF_buf12), .B(core__abc_21302_new_n2067_), .Y(core__0siphash_word0_reg_63_0__40_));
NOR2X1 NOR2X1_298 ( .A(core__abc_21302_new_n1185__bF_buf11), .B(core__abc_21302_new_n2070_), .Y(core__0siphash_word0_reg_63_0__41_));
NOR2X1 NOR2X1_299 ( .A(core__abc_21302_new_n1185__bF_buf10), .B(core__abc_21302_new_n2073_), .Y(core__0siphash_word0_reg_63_0__42_));
NOR2X1 NOR2X1_3 ( .A(\addr[4] ), .B(\addr[5] ), .Y(_abc_19873_new_n876_));
NOR2X1 NOR2X1_30 ( .A(_abc_19873_new_n1233_), .B(_abc_19873_new_n1231_), .Y(_abc_19873_new_n1234_));
NOR2X1 NOR2X1_300 ( .A(core__abc_21302_new_n1185__bF_buf9), .B(core__abc_21302_new_n2076_), .Y(core__0siphash_word0_reg_63_0__43_));
NOR2X1 NOR2X1_301 ( .A(core__abc_21302_new_n1185__bF_buf8), .B(core__abc_21302_new_n2079_), .Y(core__0siphash_word0_reg_63_0__44_));
NOR2X1 NOR2X1_302 ( .A(core__abc_21302_new_n1185__bF_buf7), .B(core__abc_21302_new_n2082_), .Y(core__0siphash_word0_reg_63_0__45_));
NOR2X1 NOR2X1_303 ( .A(core__abc_21302_new_n1185__bF_buf6), .B(core__abc_21302_new_n2085_), .Y(core__0siphash_word0_reg_63_0__46_));
NOR2X1 NOR2X1_304 ( .A(core__abc_21302_new_n1185__bF_buf5), .B(core__abc_21302_new_n2088_), .Y(core__0siphash_word0_reg_63_0__47_));
NOR2X1 NOR2X1_305 ( .A(core__abc_21302_new_n1185__bF_buf4), .B(core__abc_21302_new_n2091_), .Y(core__0siphash_word0_reg_63_0__48_));
NOR2X1 NOR2X1_306 ( .A(core__abc_21302_new_n1185__bF_buf3), .B(core__abc_21302_new_n2094_), .Y(core__0siphash_word0_reg_63_0__49_));
NOR2X1 NOR2X1_307 ( .A(core__abc_21302_new_n1185__bF_buf2), .B(core__abc_21302_new_n2097_), .Y(core__0siphash_word0_reg_63_0__50_));
NOR2X1 NOR2X1_308 ( .A(core__abc_21302_new_n1185__bF_buf1), .B(core__abc_21302_new_n2100_), .Y(core__0siphash_word0_reg_63_0__51_));
NOR2X1 NOR2X1_309 ( .A(core__abc_21302_new_n1185__bF_buf0), .B(core__abc_21302_new_n2103_), .Y(core__0siphash_word0_reg_63_0__52_));
NOR2X1 NOR2X1_31 ( .A(_abc_19873_new_n1252_), .B(_abc_19873_new_n1249_), .Y(_abc_19873_new_n1253_));
NOR2X1 NOR2X1_310 ( .A(core__abc_21302_new_n1185__bF_buf13), .B(core__abc_21302_new_n2106_), .Y(core__0siphash_word0_reg_63_0__53_));
NOR2X1 NOR2X1_311 ( .A(core__abc_21302_new_n1185__bF_buf12), .B(core__abc_21302_new_n2109_), .Y(core__0siphash_word0_reg_63_0__54_));
NOR2X1 NOR2X1_312 ( .A(core__abc_21302_new_n1185__bF_buf11), .B(core__abc_21302_new_n2112_), .Y(core__0siphash_word0_reg_63_0__55_));
NOR2X1 NOR2X1_313 ( .A(core__abc_21302_new_n1185__bF_buf10), .B(core__abc_21302_new_n2115_), .Y(core__0siphash_word0_reg_63_0__56_));
NOR2X1 NOR2X1_314 ( .A(core__abc_21302_new_n1185__bF_buf9), .B(core__abc_21302_new_n2118_), .Y(core__0siphash_word0_reg_63_0__57_));
NOR2X1 NOR2X1_315 ( .A(core__abc_21302_new_n1185__bF_buf8), .B(core__abc_21302_new_n2121_), .Y(core__0siphash_word0_reg_63_0__58_));
NOR2X1 NOR2X1_316 ( .A(core__abc_21302_new_n1185__bF_buf7), .B(core__abc_21302_new_n2124_), .Y(core__0siphash_word0_reg_63_0__59_));
NOR2X1 NOR2X1_317 ( .A(core__abc_21302_new_n1185__bF_buf6), .B(core__abc_21302_new_n2127_), .Y(core__0siphash_word0_reg_63_0__60_));
NOR2X1 NOR2X1_318 ( .A(core__abc_21302_new_n1185__bF_buf5), .B(core__abc_21302_new_n2130_), .Y(core__0siphash_word0_reg_63_0__61_));
NOR2X1 NOR2X1_319 ( .A(core__abc_21302_new_n1185__bF_buf4), .B(core__abc_21302_new_n2133_), .Y(core__0siphash_word0_reg_63_0__62_));
NOR2X1 NOR2X1_32 ( .A(_abc_19873_new_n1270_), .B(_abc_19873_new_n1268_), .Y(_abc_19873_new_n1271_));
NOR2X1 NOR2X1_320 ( .A(core__abc_21302_new_n1185__bF_buf3), .B(core__abc_21302_new_n2136_), .Y(core__0siphash_word0_reg_63_0__63_));
NOR2X1 NOR2X1_321 ( .A(core_siphash_ctrl_reg_5_), .B(core__abc_21302_new_n1155_), .Y(core__abc_21302_new_n2138_));
NOR2X1 NOR2X1_322 ( .A(core__abc_21302_new_n2143_), .B(core__abc_21302_new_n2144_), .Y(core__abc_21302_new_n2145_));
NOR2X1 NOR2X1_323 ( .A(core__abc_21302_new_n1137_), .B(core__abc_21302_new_n2145_), .Y(core__abc_21302_new_n2146_));
NOR2X1 NOR2X1_324 ( .A(core__abc_21302_new_n2147_), .B(core__abc_21302_new_n2146_), .Y(core__0loop_ctr_reg_3_0__0_));
NOR2X1 NOR2X1_325 ( .A(core__abc_21302_new_n2156_), .B(core__abc_21302_new_n2142_), .Y(core__abc_21302_new_n2157_));
NOR2X1 NOR2X1_326 ( .A(core__abc_21302_new_n2159_), .B(core__abc_21302_new_n2155_), .Y(core__0loop_ctr_reg_3_0__2_));
NOR2X1 NOR2X1_327 ( .A(core__abc_21302_new_n1155_), .B(core__abc_21302_new_n1177_), .Y(core__abc_21302_new_n2165_));
NOR2X1 NOR2X1_328 ( .A(core__abc_21302_new_n1200_), .B(core__abc_21302_new_n2166_), .Y(core__abc_21302_new_n2167_));
NOR2X1 NOR2X1_329 ( .A(core_siphash_ctrl_reg_2_), .B(core__abc_21302_new_n1150_), .Y(core__abc_21302_new_n2361_));
NOR2X1 NOR2X1_33 ( .A(_abc_19873_new_n1288_), .B(_abc_19873_new_n1286_), .Y(_abc_19873_new_n1289_));
NOR2X1 NOR2X1_330 ( .A(core_siphash_ctrl_reg_2_), .B(core__abc_21302_new_n2365__bF_buf4), .Y(core__abc_21302_new_n2366_));
NOR2X1 NOR2X1_331 ( .A(core__abc_21302_new_n2363__bF_buf5), .B(core__abc_21302_new_n2368__bF_buf4), .Y(core__abc_21302_new_n2369_));
NOR2X1 NOR2X1_332 ( .A(core_v1_reg_3_), .B(core_v0_reg_3_), .Y(core__abc_21302_new_n2372_));
NOR2X1 NOR2X1_333 ( .A(core__abc_21302_new_n2372_), .B(core__abc_21302_new_n2373_), .Y(core__abc_21302_new_n2374_));
NOR2X1 NOR2X1_334 ( .A(core_v1_reg_6_), .B(core_v0_reg_6_), .Y(core__abc_21302_new_n2379_));
NOR2X1 NOR2X1_335 ( .A(core__abc_21302_new_n2379_), .B(core__abc_21302_new_n2380_), .Y(core__abc_21302_new_n2381_));
NOR2X1 NOR2X1_336 ( .A(core_v1_reg_7_), .B(core_v0_reg_7_), .Y(core__abc_21302_new_n2382_));
NOR2X1 NOR2X1_337 ( .A(core__abc_21302_new_n2382_), .B(core__abc_21302_new_n2383_), .Y(core__abc_21302_new_n2384_));
NOR2X1 NOR2X1_338 ( .A(core_v1_reg_5_), .B(core_v0_reg_5_), .Y(core__abc_21302_new_n2387_));
NOR2X1 NOR2X1_339 ( .A(core__abc_21302_new_n2387_), .B(core__abc_21302_new_n2388_), .Y(core__abc_21302_new_n2389_));
NOR2X1 NOR2X1_34 ( .A(_abc_19873_new_n1306_), .B(_abc_19873_new_n1304_), .Y(_abc_19873_new_n1307_));
NOR2X1 NOR2X1_340 ( .A(core__abc_21302_new_n2385_), .B(core__abc_21302_new_n2390_), .Y(core__abc_21302_new_n2391_));
NOR2X1 NOR2X1_341 ( .A(core__abc_21302_new_n2398_), .B(core__abc_21302_new_n2399_), .Y(core__abc_21302_new_n2400_));
NOR2X1 NOR2X1_342 ( .A(core__abc_21302_new_n2401_), .B(core__abc_21302_new_n2402_), .Y(core__abc_21302_new_n2403_));
NOR2X1 NOR2X1_343 ( .A(core__abc_21302_new_n2421_), .B(core__abc_21302_new_n2422_), .Y(core__abc_21302_new_n2423_));
NOR2X1 NOR2X1_344 ( .A(core__abc_21302_new_n2424_), .B(core__abc_21302_new_n2425_), .Y(core__abc_21302_new_n2426_));
NOR2X1 NOR2X1_345 ( .A(core__abc_21302_new_n2428_), .B(core__abc_21302_new_n2429_), .Y(core__abc_21302_new_n2430_));
NOR2X1 NOR2X1_346 ( .A(core__abc_21302_new_n1384_), .B(core__abc_21302_new_n1395_), .Y(core__abc_21302_new_n2431_));
NOR2X1 NOR2X1_347 ( .A(core__abc_21302_new_n2433_), .B(core__abc_21302_new_n2427_), .Y(core__abc_21302_new_n2434_));
NOR2X1 NOR2X1_348 ( .A(core__abc_21302_new_n2371_), .B(core__abc_21302_new_n2467_), .Y(core__abc_21302_new_n2468_));
NOR2X1 NOR2X1_349 ( .A(core__abc_21302_new_n1275_), .B(core__abc_21302_new_n1285_), .Y(core__abc_21302_new_n2476_));
NOR2X1 NOR2X1_35 ( .A(_abc_19873_new_n1320_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1321_));
NOR2X1 NOR2X1_350 ( .A(core__abc_21302_new_n1253_), .B(core__abc_21302_new_n1265_), .Y(core__abc_21302_new_n2477_));
NOR2X1 NOR2X1_351 ( .A(core__abc_21302_new_n2483_), .B(core__abc_21302_new_n2485_), .Y(core__abc_21302_new_n2486_));
NOR2X1 NOR2X1_352 ( .A(core__abc_21302_new_n2495_), .B(core__abc_21302_new_n2494_), .Y(core__abc_21302_new_n2496_));
NOR2X1 NOR2X1_353 ( .A(core__abc_21302_new_n1567_), .B(core__abc_21302_new_n2505_), .Y(core__abc_21302_new_n2506_));
NOR2X1 NOR2X1_354 ( .A(core__abc_21302_new_n2468_), .B(core__abc_21302_new_n2506_), .Y(core__abc_21302_new_n2509_));
NOR2X1 NOR2X1_355 ( .A(core__abc_21302_new_n2520_), .B(core__abc_21302_new_n2521_), .Y(core__abc_21302_new_n2522_));
NOR2X1 NOR2X1_356 ( .A(core__abc_21302_new_n2528_), .B(core__abc_21302_new_n2527_), .Y(core__abc_21302_new_n2529_));
NOR2X1 NOR2X1_357 ( .A(core__abc_21302_new_n1296_), .B(core__abc_21302_new_n1307_), .Y(core__abc_21302_new_n2530_));
NOR2X1 NOR2X1_358 ( .A(core__abc_21302_new_n1319_), .B(core__abc_21302_new_n1331_), .Y(core__abc_21302_new_n2531_));
NOR2X1 NOR2X1_359 ( .A(core__abc_21302_new_n1361_), .B(core__abc_21302_new_n1376_), .Y(core__abc_21302_new_n2544_));
NOR2X1 NOR2X1_36 ( .A(_abc_19873_new_n1342_), .B(_abc_19873_new_n1340_), .Y(_abc_19873_new_n1343_));
NOR2X1 NOR2X1_360 ( .A(core__abc_21302_new_n1375_), .B(core__abc_21302_new_n2544_), .Y(core__abc_21302_new_n2545_));
NOR2X1 NOR2X1_361 ( .A(core__abc_21302_new_n1559_), .B(core__abc_21302_new_n1551_), .Y(core__abc_21302_new_n2549_));
NOR2X1 NOR2X1_362 ( .A(core__abc_21302_new_n1526_), .B(core__abc_21302_new_n1539_), .Y(core__abc_21302_new_n2550_));
NOR2X1 NOR2X1_363 ( .A(core__abc_21302_new_n2553_), .B(core__abc_21302_new_n2554_), .Y(core__abc_21302_new_n2555_));
NOR2X1 NOR2X1_364 ( .A(core__abc_21302_new_n1468_), .B(core__abc_21302_new_n1460_), .Y(core__abc_21302_new_n2557_));
NOR2X1 NOR2X1_365 ( .A(core__abc_21302_new_n1436_), .B(core__abc_21302_new_n1448_), .Y(core__abc_21302_new_n2558_));
NOR2X1 NOR2X1_366 ( .A(core__abc_21302_new_n2564_), .B(core__abc_21302_new_n2562_), .Y(core__abc_21302_new_n2565_));
NOR2X1 NOR2X1_367 ( .A(core__abc_21302_new_n2566_), .B(core__abc_21302_new_n2556_), .Y(core__abc_21302_new_n2567_));
NOR2X1 NOR2X1_368 ( .A(core__abc_21302_new_n1412_), .B(core__abc_21302_new_n1424_), .Y(core__abc_21302_new_n2570_));
NOR2X1 NOR2X1_369 ( .A(core__abc_21302_new_n2569_), .B(core__abc_21302_new_n2573_), .Y(core__abc_21302_new_n2574_));
NOR2X1 NOR2X1_37 ( .A(_abc_19873_new_n1356_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1357_));
NOR2X1 NOR2X1_370 ( .A(core__abc_21302_new_n2581_), .B(core__abc_21302_new_n2582_), .Y(core__abc_21302_new_n2583_));
NOR2X1 NOR2X1_371 ( .A(core__abc_21302_new_n2585_), .B(core__abc_21302_new_n2574_), .Y(core__abc_21302_new_n2586_));
NOR2X1 NOR2X1_372 ( .A(core__abc_21302_new_n1502_), .B(core__abc_21302_new_n1514_), .Y(core__abc_21302_new_n2593_));
NOR2X1 NOR2X1_373 ( .A(core__abc_21302_new_n2591_), .B(core__abc_21302_new_n2600_), .Y(core__abc_21302_new_n2601_));
NOR2X1 NOR2X1_374 ( .A(core__abc_21302_new_n1642_), .B(core__abc_21302_new_n1653_), .Y(core__abc_21302_new_n2603_));
NOR2X1 NOR2X1_375 ( .A(core__abc_21302_new_n1620_), .B(core__abc_21302_new_n1633_), .Y(core__abc_21302_new_n2604_));
NOR2X1 NOR2X1_376 ( .A(core__abc_21302_new_n1583_), .B(core__abc_21302_new_n1571_), .Y(core__abc_21302_new_n2606_));
NOR2X1 NOR2X1_377 ( .A(core__abc_21302_new_n1597_), .B(core__abc_21302_new_n1609_), .Y(core__abc_21302_new_n2607_));
NOR2X1 NOR2X1_378 ( .A(core__abc_21302_new_n2608_), .B(core__abc_21302_new_n2605_), .Y(core__abc_21302_new_n2609_));
NOR2X1 NOR2X1_379 ( .A(core__abc_21302_new_n2613_), .B(core__abc_21302_new_n2605_), .Y(core__abc_21302_new_n2614_));
NOR2X1 NOR2X1_38 ( .A(_abc_19873_new_n1365_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1366_));
NOR2X1 NOR2X1_380 ( .A(core__abc_21302_new_n2619_), .B(core__abc_21302_new_n2614_), .Y(core__abc_21302_new_n2620_));
NOR2X1 NOR2X1_381 ( .A(core__abc_21302_new_n1664_), .B(core__abc_21302_new_n1675_), .Y(core__abc_21302_new_n2621_));
NOR2X1 NOR2X1_382 ( .A(core__abc_21302_new_n2631_), .B(core__abc_21302_new_n2628_), .Y(core__abc_21302_new_n2632_));
NOR2X1 NOR2X1_383 ( .A(core__abc_21302_new_n2138_), .B(core__abc_21302_new_n2633_), .Y(core__abc_21302_new_n2634_));
NOR2X1 NOR2X1_384 ( .A(core__abc_21302_new_n2139_), .B(core__abc_21302_new_n2638_), .Y(core__abc_21302_new_n2639_));
NOR2X1 NOR2X1_385 ( .A(core_key_64_), .B(core__abc_21302_new_n2640__bF_buf11), .Y(core__abc_21302_new_n2641_));
NOR2X1 NOR2X1_386 ( .A(core__abc_21302_new_n1566_), .B(core__abc_21302_new_n2647_), .Y(core__abc_21302_new_n2648_));
NOR2X1 NOR2X1_387 ( .A(core__abc_21302_new_n2654_), .B(core__abc_21302_new_n2656_), .Y(core__abc_21302_new_n2657_));
NOR2X1 NOR2X1_388 ( .A(core__abc_21302_new_n2662_), .B(core__abc_21302_new_n2664_), .Y(core__abc_21302_new_n2665_));
NOR2X1 NOR2X1_389 ( .A(core__abc_21302_new_n2370_), .B(core__abc_21302_new_n2677_), .Y(core__abc_21302_new_n2678_));
NOR2X1 NOR2X1_39 ( .A(_abc_19873_new_n1379_), .B(_abc_19873_new_n1377_), .Y(_abc_19873_new_n1380_));
NOR2X1 NOR2X1_390 ( .A(core__abc_21302_new_n2682_), .B(core__abc_21302_new_n2686_), .Y(core__abc_21302_new_n2689_));
NOR2X1 NOR2X1_391 ( .A(core__abc_21302_new_n2693_), .B(core__abc_21302_new_n2696_), .Y(core__abc_21302_new_n2697_));
NOR2X1 NOR2X1_392 ( .A(core__abc_21302_new_n1537_), .B(core__abc_21302_new_n2705_), .Y(core__abc_21302_new_n2706_));
NOR2X1 NOR2X1_393 ( .A(core_v3_reg_29_), .B(core__abc_21302_new_n2707_), .Y(core__abc_21302_new_n2708_));
NOR2X1 NOR2X1_394 ( .A(core__abc_21302_new_n2706_), .B(core__abc_21302_new_n2708_), .Y(core__abc_21302_new_n2709_));
NOR2X1 NOR2X1_395 ( .A(core__abc_21302_new_n2725_), .B(core__abc_21302_new_n2726_), .Y(core__abc_21302_new_n2727_));
NOR2X1 NOR2X1_396 ( .A(core__abc_21302_new_n2673__bF_buf8), .B(core__abc_21302_new_n2751_), .Y(core__abc_21302_new_n2754_));
NOR2X1 NOR2X1_397 ( .A(core__abc_21302_new_n1616_), .B(core__abc_21302_new_n2767_), .Y(core__abc_21302_new_n2769_));
NOR2X1 NOR2X1_398 ( .A(core__abc_21302_new_n2769_), .B(core__abc_21302_new_n2768_), .Y(core__abc_21302_new_n2777_));
NOR2X1 NOR2X1_399 ( .A(core__abc_21302_new_n2785_), .B(core__abc_21302_new_n2788_), .Y(core__abc_21302_new_n2789_));
NOR2X1 NOR2X1_4 ( .A(_abc_19873_new_n873_), .B(_abc_19873_new_n880_), .Y(_abc_19873_new_n881_));
NOR2X1 NOR2X1_40 ( .A(_abc_19873_new_n1397_), .B(_abc_19873_new_n1395_), .Y(_abc_19873_new_n1398_));
NOR2X1 NOR2X1_400 ( .A(core__abc_21302_new_n1185__bF_buf2), .B(core__abc_21302_new_n2796_), .Y(core__0v3_reg_63_0__4_));
NOR2X1 NOR2X1_401 ( .A(core__abc_21302_new_n1615_), .B(core__abc_21302_new_n2768_), .Y(core__abc_21302_new_n2801_));
NOR2X1 NOR2X1_402 ( .A(core__abc_21302_new_n1732_), .B(core__abc_21302_new_n1743_), .Y(core__abc_21302_new_n2814_));
NOR2X1 NOR2X1_403 ( .A(core__abc_21302_new_n2815_), .B(core__abc_21302_new_n2663_), .Y(core__abc_21302_new_n2816_));
NOR2X1 NOR2X1_404 ( .A(core__abc_21302_new_n1756_), .B(core__abc_21302_new_n2825_), .Y(core__abc_21302_new_n2826_));
NOR2X1 NOR2X1_405 ( .A(core__abc_21302_new_n2828_), .B(core__abc_21302_new_n2826_), .Y(core__abc_21302_new_n2829_));
NOR2X1 NOR2X1_406 ( .A(core__abc_21302_new_n1185__bF_buf1), .B(core__abc_21302_new_n2837_), .Y(core__0v3_reg_63_0__5_));
NOR2X1 NOR2X1_407 ( .A(core__abc_21302_new_n1638_), .B(core__abc_21302_new_n2842_), .Y(core__abc_21302_new_n2843_));
NOR2X1 NOR2X1_408 ( .A(core__abc_21302_new_n2521_), .B(core__abc_21302_new_n2770_), .Y(core__abc_21302_new_n2845_));
NOR2X1 NOR2X1_409 ( .A(core__abc_21302_new_n2846_), .B(core__abc_21302_new_n2845_), .Y(core__abc_21302_new_n2848_));
NOR2X1 NOR2X1_41 ( .A(_abc_19873_new_n1411_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1412_));
NOR2X1 NOR2X1_410 ( .A(core__abc_21302_new_n2843_), .B(core__abc_21302_new_n2844_), .Y(core__abc_21302_new_n2853_));
NOR2X1 NOR2X1_411 ( .A(core__abc_21302_new_n2807_), .B(core__abc_21302_new_n2809_), .Y(core__abc_21302_new_n2859_));
NOR2X1 NOR2X1_412 ( .A(core_v3_reg_33_), .B(core__abc_21302_new_n2868_), .Y(core__abc_21302_new_n2869_));
NOR2X1 NOR2X1_413 ( .A(core__abc_21302_new_n2869_), .B(core__abc_21302_new_n2870_), .Y(core__abc_21302_new_n2871_));
NOR2X1 NOR2X1_414 ( .A(core__abc_21302_new_n2879_), .B(core__abc_21302_new_n2843_), .Y(core__abc_21302_new_n2880_));
NOR2X1 NOR2X1_415 ( .A(core__abc_21302_new_n2827_), .B(core__abc_21302_new_n2896_), .Y(core__abc_21302_new_n2897_));
NOR2X1 NOR2X1_416 ( .A(core__abc_21302_new_n2864_), .B(core__abc_21302_new_n2896_), .Y(core__abc_21302_new_n2898_));
NOR2X1 NOR2X1_417 ( .A(core__abc_21302_new_n2895_), .B(core__abc_21302_new_n2900_), .Y(core__abc_21302_new_n2902_));
NOR2X1 NOR2X1_418 ( .A(core__abc_21302_new_n2902_), .B(core__abc_21302_new_n2901_), .Y(core__abc_21302_new_n2904_));
NOR2X1 NOR2X1_419 ( .A(core__abc_21302_new_n1185__bF_buf0), .B(core__abc_21302_new_n2913_), .Y(core__0v3_reg_63_0__7_));
NOR2X1 NOR2X1_42 ( .A(_abc_19873_new_n1420_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1421_));
NOR2X1 NOR2X1_420 ( .A(core_key_72_), .B(core__abc_21302_new_n2640__bF_buf4), .Y(core__abc_21302_new_n2915_));
NOR2X1 NOR2X1_421 ( .A(core__abc_21302_new_n1638_), .B(core__abc_21302_new_n1649_), .Y(core__abc_21302_new_n2921_));
NOR2X1 NOR2X1_422 ( .A(core__abc_21302_new_n2922_), .B(core__abc_21302_new_n2766_), .Y(core__abc_21302_new_n2927_));
NOR2X1 NOR2X1_423 ( .A(core__abc_21302_new_n2920_), .B(core__abc_21302_new_n2928_), .Y(core__abc_21302_new_n2929_));
NOR2X1 NOR2X1_424 ( .A(core__abc_21302_new_n1660_), .B(core__abc_21302_new_n2935_), .Y(core__abc_21302_new_n2936_));
NOR2X1 NOR2X1_425 ( .A(core__abc_21302_new_n2936_), .B(core__abc_21302_new_n2929_), .Y(core__abc_21302_new_n2937_));
NOR2X1 NOR2X1_426 ( .A(core__abc_21302_new_n2944_), .B(core__abc_21302_new_n2919_), .Y(core__abc_21302_new_n2945_));
NOR2X1 NOR2X1_427 ( .A(core__abc_21302_new_n2945_), .B(core__abc_21302_new_n2946_), .Y(core__abc_21302_new_n2947_));
NOR2X1 NOR2X1_428 ( .A(core__abc_21302_new_n1659_), .B(core__abc_21302_new_n2929_), .Y(core__abc_21302_new_n2964_));
NOR2X1 NOR2X1_429 ( .A(core__abc_21302_new_n2977_), .B(core__abc_21302_new_n2946_), .Y(core__abc_21302_new_n2978_));
NOR2X1 NOR2X1_43 ( .A(_abc_19873_new_n1430_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1431_));
NOR2X1 NOR2X1_430 ( .A(core__abc_21302_new_n2948_), .B(core__abc_21302_new_n2895_), .Y(core__abc_21302_new_n2981_));
NOR2X1 NOR2X1_431 ( .A(core__abc_21302_new_n2986_), .B(core__abc_21302_new_n2983_), .Y(core__abc_21302_new_n2987_));
NOR2X1 NOR2X1_432 ( .A(core__abc_21302_new_n1185__bF_buf13), .B(core__abc_21302_new_n2998_), .Y(core__0v3_reg_63_0__9_));
NOR2X1 NOR2X1_433 ( .A(core_key_74_), .B(core__abc_21302_new_n2640__bF_buf3), .Y(core__abc_21302_new_n3000_));
NOR2X1 NOR2X1_434 ( .A(core__abc_21302_new_n3006_), .B(core__abc_21302_new_n3012_), .Y(core__abc_21302_new_n3013_));
NOR2X1 NOR2X1_435 ( .A(core__abc_21302_new_n3013_), .B(core__abc_21302_new_n3014_), .Y(core__abc_21302_new_n3021_));
NOR2X1 NOR2X1_436 ( .A(core__abc_21302_new_n1681_), .B(core__abc_21302_new_n3013_), .Y(core__abc_21302_new_n3045_));
NOR2X1 NOR2X1_437 ( .A(core__abc_21302_new_n1826_), .B(core__abc_21302_new_n3066_), .Y(core__abc_21302_new_n3069_));
NOR2X1 NOR2X1_438 ( .A(core__abc_21302_new_n3069_), .B(core__abc_21302_new_n3068_), .Y(core__abc_21302_new_n3071_));
NOR2X1 NOR2X1_439 ( .A(core__abc_21302_new_n3002_), .B(core__abc_21302_new_n3083_), .Y(core__abc_21302_new_n3088_));
NOR2X1 NOR2X1_44 ( .A(_abc_19873_new_n1439_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1440_));
NOR2X1 NOR2X1_440 ( .A(core__abc_21302_new_n3007_), .B(core__abc_21302_new_n3091_), .Y(core__abc_21302_new_n3095_));
NOR2X1 NOR2X1_441 ( .A(core__abc_21302_new_n1341_), .B(core__abc_21302_new_n3103_), .Y(core__abc_21302_new_n3106_));
NOR2X1 NOR2X1_442 ( .A(core__abc_21302_new_n3106_), .B(core__abc_21302_new_n3105_), .Y(core__abc_21302_new_n3107_));
NOR2X1 NOR2X1_443 ( .A(core__abc_21302_new_n3111_), .B(core__abc_21302_new_n3116_), .Y(core__abc_21302_new_n3117_));
NOR2X1 NOR2X1_444 ( .A(core__abc_21302_new_n3117_), .B(core__abc_21302_new_n3119_), .Y(core__abc_21302_new_n3120_));
NOR2X1 NOR2X1_445 ( .A(core_key_77_), .B(core__abc_21302_new_n2640__bF_buf2), .Y(core__abc_21302_new_n3129_));
NOR2X1 NOR2X1_446 ( .A(core__abc_21302_new_n3130_), .B(core__abc_21302_new_n3099_), .Y(core__abc_21302_new_n3131_));
NOR2X1 NOR2X1_447 ( .A(core__abc_21302_new_n1704_), .B(core__abc_21302_new_n3131_), .Y(core__abc_21302_new_n3132_));
NOR2X1 NOR2X1_448 ( .A(core__abc_21302_new_n3145_), .B(core__abc_21302_new_n3136_), .Y(core__abc_21302_new_n3148_));
NOR2X1 NOR2X1_449 ( .A(core__abc_21302_new_n3148_), .B(core__abc_21302_new_n3147_), .Y(core__abc_21302_new_n3149_));
NOR2X1 NOR2X1_45 ( .A(_abc_19873_new_n1453_), .B(_abc_19873_new_n1451_), .Y(_abc_19873_new_n1454_));
NOR2X1 NOR2X1_450 ( .A(core__abc_21302_new_n3149_), .B(core__abc_21302_new_n3151_), .Y(core__abc_21302_new_n3152_));
NOR2X1 NOR2X1_451 ( .A(core__abc_21302_new_n3152_), .B(core__abc_21302_new_n3153_), .Y(core__abc_21302_new_n3154_));
NOR2X1 NOR2X1_452 ( .A(core__abc_21302_new_n3157_), .B(core__abc_21302_new_n3159_), .Y(core__abc_21302_new_n3160_));
NOR2X1 NOR2X1_453 ( .A(core_key_78_), .B(core__abc_21302_new_n2640__bF_buf1), .Y(core__abc_21302_new_n3175_));
NOR2X1 NOR2X1_454 ( .A(core__abc_21302_new_n3148_), .B(core__abc_21302_new_n3153_), .Y(core__abc_21302_new_n3176_));
NOR2X1 NOR2X1_455 ( .A(core__abc_21302_new_n3177_), .B(core__abc_21302_new_n3181_), .Y(core__abc_21302_new_n3182_));
NOR2X1 NOR2X1_456 ( .A(core__abc_21302_new_n1728_), .B(core__abc_21302_new_n3184_), .Y(core__abc_21302_new_n3185_));
NOR2X1 NOR2X1_457 ( .A(core__abc_21302_new_n3187_), .B(core__abc_21302_new_n3189_), .Y(core__abc_21302_new_n3190_));
NOR2X1 NOR2X1_458 ( .A(core__abc_21302_new_n3193_), .B(core__abc_21302_new_n3191_), .Y(core__abc_21302_new_n3195_));
NOR2X1 NOR2X1_459 ( .A(core__abc_21302_new_n3237_), .B(core__abc_21302_new_n3225_), .Y(core__abc_21302_new_n3238_));
NOR2X1 NOR2X1_46 ( .A(_abc_19873_new_n1469_), .B(_abc_19873_new_n1472_), .Y(_abc_19873_new_n1473_));
NOR2X1 NOR2X1_460 ( .A(core__abc_21302_new_n1879_), .B(core__abc_21302_new_n3248_), .Y(core__abc_21302_new_n3249_));
NOR2X1 NOR2X1_461 ( .A(core__abc_21302_new_n3261_), .B(core__abc_21302_new_n3259_), .Y(core__abc_21302_new_n3262_));
NOR2X1 NOR2X1_462 ( .A(core__abc_21302_new_n3272_), .B(core__abc_21302_new_n3273_), .Y(core__abc_21302_new_n3274_));
NOR2X1 NOR2X1_463 ( .A(core__abc_21302_new_n3286_), .B(core__abc_21302_new_n3179_), .Y(core__abc_21302_new_n3287_));
NOR2X1 NOR2X1_464 ( .A(core__abc_21302_new_n1751_), .B(core__abc_21302_new_n3296_), .Y(core__abc_21302_new_n3298_));
NOR2X1 NOR2X1_465 ( .A(core__abc_21302_new_n3298_), .B(core__abc_21302_new_n3297_), .Y(core__abc_21302_new_n3303_));
NOR2X1 NOR2X1_466 ( .A(core__abc_21302_new_n3306_), .B(core__abc_21302_new_n3285_), .Y(core__abc_21302_new_n3309_));
NOR2X1 NOR2X1_467 ( .A(core__abc_21302_new_n3309_), .B(core__abc_21302_new_n3308_), .Y(core__abc_21302_new_n3310_));
NOR2X1 NOR2X1_468 ( .A(core__abc_21302_new_n3317_), .B(core__abc_21302_new_n3250_), .Y(core__abc_21302_new_n3318_));
NOR2X1 NOR2X1_469 ( .A(core__abc_21302_new_n3316_), .B(core__abc_21302_new_n3320_), .Y(core__abc_21302_new_n3321_));
NOR2X1 NOR2X1_47 ( .A(_abc_19873_new_n1491_), .B(_abc_19873_new_n1489_), .Y(_abc_19873_new_n1492_));
NOR2X1 NOR2X1_470 ( .A(core__abc_21302_new_n3288_), .B(core__abc_21302_new_n2934_), .Y(core__abc_21302_new_n3330_));
NOR2X1 NOR2X1_471 ( .A(core__abc_21302_new_n1761_), .B(core__abc_21302_new_n3332_), .Y(core__abc_21302_new_n3333_));
NOR2X1 NOR2X1_472 ( .A(core__abc_21302_new_n3336_), .B(core__abc_21302_new_n3333_), .Y(core__abc_21302_new_n3337_));
NOR2X1 NOR2X1_473 ( .A(core__abc_21302_new_n3347_), .B(core__abc_21302_new_n3308_), .Y(core__abc_21302_new_n3348_));
NOR2X1 NOR2X1_474 ( .A(core__abc_21302_new_n3349_), .B(core__abc_21302_new_n3348_), .Y(core__abc_21302_new_n3350_));
NOR2X1 NOR2X1_475 ( .A(core__abc_21302_new_n1905_), .B(core__abc_21302_new_n3353_), .Y(core__abc_21302_new_n3355_));
NOR2X1 NOR2X1_476 ( .A(core_key_82_), .B(core__abc_21302_new_n2640__bF_buf0), .Y(core__abc_21302_new_n3368_));
NOR2X1 NOR2X1_477 ( .A(core__abc_21302_new_n3346_), .B(core__abc_21302_new_n3307_), .Y(core__abc_21302_new_n3369_));
NOR2X1 NOR2X1_478 ( .A(core__abc_21302_new_n3341_), .B(core__abc_21302_new_n3371_), .Y(core__abc_21302_new_n3372_));
NOR2X1 NOR2X1_479 ( .A(core__abc_21302_new_n3375_), .B(core__abc_21302_new_n3369_), .Y(core__abc_21302_new_n3376_));
NOR2X1 NOR2X1_48 ( .A(_abc_19873_new_n1505_), .B(_abc_19873_new_n924_), .Y(_abc_19873_new_n1506_));
NOR2X1 NOR2X1_480 ( .A(core__abc_21302_new_n3377_), .B(core__abc_21302_new_n3382_), .Y(core__abc_21302_new_n3390_));
NOR2X1 NOR2X1_481 ( .A(core__abc_21302_new_n1424_), .B(core__abc_21302_new_n3420_), .Y(core__abc_21302_new_n3425_));
NOR2X1 NOR2X1_482 ( .A(core__abc_21302_new_n3357_), .B(core__abc_21302_new_n3399_), .Y(core__abc_21302_new_n3441_));
NOR2X1 NOR2X1_483 ( .A(core__abc_21302_new_n3440_), .B(core__abc_21302_new_n3442_), .Y(core__abc_21302_new_n3443_));
NOR2X1 NOR2X1_484 ( .A(core__abc_21302_new_n1185__bF_buf11), .B(core__abc_21302_new_n3456_), .Y(core__0v3_reg_63_0__19_));
NOR2X1 NOR2X1_485 ( .A(core__abc_21302_new_n3428_), .B(core__abc_21302_new_n3458_), .Y(core__abc_21302_new_n3459_));
NOR2X1 NOR2X1_486 ( .A(core__abc_21302_new_n3461_), .B(core__abc_21302_new_n3462_), .Y(core__abc_21302_new_n3463_));
NOR2X1 NOR2X1_487 ( .A(core__abc_21302_new_n3377_), .B(core__abc_21302_new_n3418_), .Y(core__abc_21302_new_n3469_));
NOR2X1 NOR2X1_488 ( .A(core__abc_21302_new_n2370_), .B(core__abc_21302_new_n3495_), .Y(core__abc_21302_new_n3496_));
NOR2X1 NOR2X1_489 ( .A(core_key_85_), .B(core__abc_21302_new_n2640__bF_buf9), .Y(core__abc_21302_new_n3499_));
NOR2X1 NOR2X1_49 ( .A(_abc_19873_new_n1514_), .B(_abc_19873_new_n953_), .Y(_abc_19873_new_n1515_));
NOR2X1 NOR2X1_490 ( .A(core__abc_21302_new_n3517_), .B(core__abc_21302_new_n3519_), .Y(core__abc_21302_new_n3520_));
NOR2X1 NOR2X1_491 ( .A(core_key_86_), .B(core__abc_21302_new_n2640__bF_buf8), .Y(core__abc_21302_new_n3531_));
NOR2X1 NOR2X1_492 ( .A(core__abc_21302_new_n3537_), .B(core__abc_21302_new_n3542_), .Y(core__abc_21302_new_n3543_));
NOR2X1 NOR2X1_493 ( .A(core__abc_21302_new_n1821_), .B(core__abc_21302_new_n3546_), .Y(core__abc_21302_new_n3547_));
NOR2X1 NOR2X1_494 ( .A(core__abc_21302_new_n2575_), .B(core__abc_21302_new_n3549_), .Y(core__abc_21302_new_n3551_));
NOR2X1 NOR2X1_495 ( .A(core__abc_21302_new_n3562_), .B(core__abc_21302_new_n3536_), .Y(core__abc_21302_new_n3564_));
NOR2X1 NOR2X1_496 ( .A(core__abc_21302_new_n3564_), .B(core__abc_21302_new_n3563_), .Y(core__abc_21302_new_n3565_));
NOR2X1 NOR2X1_497 ( .A(core__abc_21302_new_n3574_), .B(core__abc_21302_new_n3563_), .Y(core__abc_21302_new_n3575_));
NOR2X1 NOR2X1_498 ( .A(core__abc_21302_new_n3591_), .B(core__abc_21302_new_n3588_), .Y(core__abc_21302_new_n3592_));
NOR2X1 NOR2X1_499 ( .A(core__abc_21302_new_n3600_), .B(core__abc_21302_new_n3598_), .Y(core__abc_21302_new_n3601_));
NOR2X1 NOR2X1_5 ( .A(_abc_19873_new_n886_), .B(_abc_19873_new_n888_), .Y(_abc_19873_new_n889_));
NOR2X1 NOR2X1_50 ( .A(_abc_19873_new_n1848_), .B(_abc_19873_new_n918_), .Y(_abc_19873_new_n2265_));
NOR2X1 NOR2X1_500 ( .A(core__abc_21302_new_n3618_), .B(core__abc_21302_new_n3539_), .Y(core__abc_21302_new_n3619_));
NOR2X1 NOR2X1_501 ( .A(core__abc_21302_new_n3473_), .B(core__abc_21302_new_n3620_), .Y(core__abc_21302_new_n3621_));
NOR2X1 NOR2X1_502 ( .A(core__abc_21302_new_n3620_), .B(core__abc_21302_new_n3500_), .Y(core__abc_21302_new_n3622_));
NOR2X1 NOR2X1_503 ( .A(core__abc_21302_new_n3617_), .B(core__abc_21302_new_n3626_), .Y(core__abc_21302_new_n3627_));
NOR2X1 NOR2X1_504 ( .A(core__abc_21302_new_n3624_), .B(core__abc_21302_new_n3622_), .Y(core__abc_21302_new_n3629_));
NOR2X1 NOR2X1_505 ( .A(core__abc_21302_new_n1848_), .B(core__abc_21302_new_n3630_), .Y(core__abc_21302_new_n3631_));
NOR2X1 NOR2X1_506 ( .A(core__abc_21302_new_n3627_), .B(core__abc_21302_new_n3631_), .Y(core__abc_21302_new_n3642_));
NOR2X1 NOR2X1_507 ( .A(core__abc_21302_new_n1185__bF_buf10), .B(core__abc_21302_new_n3653_), .Y(core__0v3_reg_63_0__24_));
NOR2X1 NOR2X1_508 ( .A(core__abc_21302_new_n3687_), .B(core__abc_21302_new_n2640__bF_buf5), .Y(core__abc_21302_new_n3688_));
NOR2X1 NOR2X1_509 ( .A(core__abc_21302_new_n3694_), .B(core__abc_21302_new_n3617_), .Y(core__abc_21302_new_n3695_));
NOR2X1 NOR2X1_51 ( .A(_abc_19873_new_n878_), .B(_abc_19873_new_n2287_), .Y(_0ctrl_reg_2_0__0_));
NOR2X1 NOR2X1_510 ( .A(core__abc_21302_new_n1874_), .B(core__abc_21302_new_n3699_), .Y(core__abc_21302_new_n3702_));
NOR2X1 NOR2X1_511 ( .A(core__abc_21302_new_n2551_), .B(core__abc_21302_new_n3704_), .Y(core__abc_21302_new_n3705_));
NOR2X1 NOR2X1_512 ( .A(core__abc_21302_new_n3702_), .B(core__abc_21302_new_n3701_), .Y(core__abc_21302_new_n3725_));
NOR2X1 NOR2X1_513 ( .A(core__abc_21302_new_n3727_), .B(core__abc_21302_new_n3693_), .Y(core__abc_21302_new_n3728_));
NOR2X1 NOR2X1_514 ( .A(core__abc_21302_new_n3726_), .B(core__abc_21302_new_n3728_), .Y(core__abc_21302_new_n3729_));
NOR2X1 NOR2X1_515 ( .A(core__abc_21302_new_n3779_), .B(core__abc_21302_new_n3767_), .Y(core__abc_21302_new_n3781_));
NOR2X1 NOR2X1_516 ( .A(core__abc_21302_new_n3781_), .B(core__abc_21302_new_n3780_), .Y(core__abc_21302_new_n3782_));
NOR2X1 NOR2X1_517 ( .A(core__abc_21302_new_n1899_), .B(core__abc_21302_new_n1914_), .Y(core__abc_21302_new_n3793_));
NOR2X1 NOR2X1_518 ( .A(core__abc_21302_new_n3768_), .B(core__abc_21302_new_n3801_), .Y(core__abc_21302_new_n3802_));
NOR2X1 NOR2X1_519 ( .A(core__abc_21302_new_n1539_), .B(core__abc_21302_new_n3810_), .Y(core__abc_21302_new_n3813_));
NOR2X1 NOR2X1_52 ( .A(_abc_19873_new_n878_), .B(_abc_19873_new_n2289_), .Y(_0ctrl_reg_2_0__1_));
NOR2X1 NOR2X1_520 ( .A(core__abc_21302_new_n3817_), .B(core__abc_21302_new_n3819_), .Y(core__abc_21302_new_n3820_));
NOR2X1 NOR2X1_521 ( .A(core__abc_21302_new_n1185__bF_buf8), .B(core__abc_21302_new_n3828_), .Y(core__0v3_reg_63_0__29_));
NOR2X1 NOR2X1_522 ( .A(core_key_94_), .B(core__abc_21302_new_n2640__bF_buf1), .Y(core__abc_21302_new_n3830_));
NOR2X1 NOR2X1_523 ( .A(core__abc_21302_new_n3831_), .B(core__abc_21302_new_n3833_), .Y(core__abc_21302_new_n3834_));
NOR2X1 NOR2X1_524 ( .A(core__abc_21302_new_n1551_), .B(core__abc_21302_new_n3837_), .Y(core__abc_21302_new_n3838_));
NOR2X1 NOR2X1_525 ( .A(core__abc_21302_new_n3866_), .B(core__abc_21302_new_n3867_), .Y(core__abc_21302_new_n3868_));
NOR2X1 NOR2X1_526 ( .A(core__abc_21302_new_n3865_), .B(core__abc_21302_new_n3868_), .Y(core__abc_21302_new_n3869_));
NOR2X1 NOR2X1_527 ( .A(core__abc_21302_new_n3877_), .B(core__abc_21302_new_n3865_), .Y(core__abc_21302_new_n3878_));
NOR2X1 NOR2X1_528 ( .A(core__abc_21302_new_n3904_), .B(core__abc_21302_new_n3902_), .Y(core__abc_21302_new_n3905_));
NOR2X1 NOR2X1_529 ( .A(core__abc_21302_new_n3761_), .B(core__abc_21302_new_n3690_), .Y(core__abc_21302_new_n3910_));
NOR2X1 NOR2X1_53 ( .A(_abc_19873_new_n878_), .B(_abc_19873_new_n2291_), .Y(_0ctrl_reg_2_0__2_));
NOR2X1 NOR2X1_530 ( .A(core__abc_21302_new_n2602_), .B(core__abc_21302_new_n2568_), .Y(core__abc_21302_new_n3921_));
NOR2X1 NOR2X1_531 ( .A(core__abc_21302_new_n1211_), .B(core__abc_21302_new_n3926_), .Y(core__abc_21302_new_n3928_));
NOR2X1 NOR2X1_532 ( .A(core__abc_21302_new_n3928_), .B(core__abc_21302_new_n3927_), .Y(core__abc_21302_new_n3929_));
NOR2X1 NOR2X1_533 ( .A(core__abc_21302_new_n3913_), .B(core__abc_21302_new_n3920_), .Y(core__abc_21302_new_n3931_));
NOR2X1 NOR2X1_534 ( .A(core__abc_21302_new_n1398_), .B(core__abc_21302_new_n3954_), .Y(core__abc_21302_new_n3955_));
NOR2X1 NOR2X1_535 ( .A(core_v3_reg_17_), .B(core__abc_21302_new_n3956_), .Y(core__abc_21302_new_n3957_));
NOR2X1 NOR2X1_536 ( .A(core__abc_21302_new_n3955_), .B(core__abc_21302_new_n3957_), .Y(core__abc_21302_new_n3959_));
NOR2X1 NOR2X1_537 ( .A(core__abc_21302_new_n2673__bF_buf10), .B(core__abc_21302_new_n3963_), .Y(core__abc_21302_new_n3964_));
NOR2X1 NOR2X1_538 ( .A(core__abc_21302_new_n3980_), .B(core__abc_21302_new_n3983_), .Y(core__abc_21302_new_n3986_));
NOR2X1 NOR2X1_539 ( .A(core__abc_21302_new_n3974_), .B(core__abc_21302_new_n4032_), .Y(core__abc_21302_new_n4037_));
NOR2X1 NOR2X1_54 ( .A(_abc_19873_new_n873_), .B(_abc_19873_new_n892_), .Y(_abc_19873_new_n2294_));
NOR2X1 NOR2X1_540 ( .A(core__abc_21302_new_n4038_), .B(core__abc_21302_new_n3931_), .Y(core__abc_21302_new_n4039_));
NOR2X1 NOR2X1_541 ( .A(core__abc_21302_new_n4036_), .B(core__abc_21302_new_n4039_), .Y(core__abc_21302_new_n4040_));
NOR2X1 NOR2X1_542 ( .A(core__abc_21302_new_n4077_), .B(core__abc_21302_new_n4076_), .Y(core__abc_21302_new_n4078_));
NOR2X1 NOR2X1_543 ( .A(core__abc_21302_new_n2370_), .B(core__abc_21302_new_n4149_), .Y(core__abc_21302_new_n4150_));
NOR2X1 NOR2X1_544 ( .A(core__abc_21302_new_n4136_), .B(core__abc_21302_new_n4137_), .Y(core__abc_21302_new_n4157_));
NOR2X1 NOR2X1_545 ( .A(core__abc_21302_new_n4161_), .B(core__abc_21302_new_n4172_), .Y(core__abc_21302_new_n4181_));
NOR2X1 NOR2X1_546 ( .A(core__abc_21302_new_n2514_), .B(core__abc_21302_new_n2623_), .Y(core__abc_21302_new_n4222_));
NOR2X1 NOR2X1_547 ( .A(core__abc_21302_new_n4205_), .B(core__abc_21302_new_n4204_), .Y(core__abc_21302_new_n4232_));
NOR2X1 NOR2X1_548 ( .A(core__abc_21302_new_n4231_), .B(core__abc_21302_new_n4236_), .Y(core__abc_21302_new_n4239_));
NOR2X1 NOR2X1_549 ( .A(core__abc_21302_new_n4239_), .B(core__abc_21302_new_n4238_), .Y(core__abc_21302_new_n4241_));
NOR2X1 NOR2X1_55 ( .A(core_compression_rounds_1_), .B(core_compression_rounds_0_), .Y(core__abc_21302_new_n1130_));
NOR2X1 NOR2X1_550 ( .A(core__abc_21302_new_n4277_), .B(core__abc_21302_new_n4282_), .Y(core__abc_21302_new_n4283_));
NOR2X1 NOR2X1_551 ( .A(core__abc_21302_new_n2673__bF_buf0), .B(core__abc_21302_new_n4292_), .Y(core__abc_21302_new_n4293_));
NOR2X1 NOR2X1_552 ( .A(core_key_112_), .B(core__abc_21302_new_n2640__bF_buf1), .Y(core__abc_21302_new_n4385_));
NOR2X1 NOR2X1_553 ( .A(core__abc_21302_new_n4281_), .B(core__abc_21302_new_n4389_), .Y(core__abc_21302_new_n4390_));
NOR2X1 NOR2X1_554 ( .A(core__abc_21302_new_n4398_), .B(core__abc_21302_new_n2830_), .Y(core__abc_21302_new_n4399_));
NOR2X1 NOR2X1_555 ( .A(core__abc_21302_new_n4418_), .B(core__abc_21302_new_n4415_), .Y(core__abc_21302_new_n4419_));
NOR2X1 NOR2X1_556 ( .A(core__abc_21302_new_n4419_), .B(core__abc_21302_new_n4423_), .Y(core__abc_21302_new_n4424_));
NOR2X1 NOR2X1_557 ( .A(core__abc_21302_new_n4449_), .B(core__abc_21302_new_n2906_), .Y(core__abc_21302_new_n4450_));
NOR2X1 NOR2X1_558 ( .A(core__abc_21302_new_n4458_), .B(core__abc_21302_new_n4457_), .Y(core__abc_21302_new_n4459_));
NOR2X1 NOR2X1_559 ( .A(core__abc_21302_new_n2495_), .B(core__abc_21302_new_n2492_), .Y(core__abc_21302_new_n4500_));
NOR2X1 NOR2X1_56 ( .A(core_compression_rounds_2_), .B(core__abc_21302_new_n1131_), .Y(core__abc_21302_new_n1132_));
NOR2X1 NOR2X1_560 ( .A(core__abc_21302_new_n2445_), .B(core__abc_21302_new_n4500_), .Y(core__abc_21302_new_n4502_));
NOR2X1 NOR2X1_561 ( .A(core__abc_21302_new_n4522_), .B(core__abc_21302_new_n3033_), .Y(core__abc_21302_new_n4523_));
NOR2X1 NOR2X1_562 ( .A(core__abc_21302_new_n4524_), .B(core__abc_21302_new_n4523_), .Y(core__abc_21302_new_n4525_));
NOR2X1 NOR2X1_563 ( .A(core__abc_21302_new_n1455_), .B(core__abc_21302_new_n4544_), .Y(core__abc_21302_new_n4547_));
NOR2X1 NOR2X1_564 ( .A(core__abc_21302_new_n4547_), .B(core__abc_21302_new_n4546_), .Y(core__abc_21302_new_n4548_));
NOR2X1 NOR2X1_565 ( .A(core__abc_21302_new_n4552_), .B(core__abc_21302_new_n4554_), .Y(core__abc_21302_new_n4556_));
NOR2X1 NOR2X1_566 ( .A(core__abc_21302_new_n4497_), .B(core__abc_21302_new_n4493_), .Y(core__abc_21302_new_n4594_));
NOR2X1 NOR2X1_567 ( .A(core__abc_21302_new_n4602_), .B(core__abc_21302_new_n4597_), .Y(core__abc_21302_new_n4603_));
NOR2X1 NOR2X1_568 ( .A(core__abc_21302_new_n4625_), .B(core__abc_21302_new_n4627_), .Y(core__abc_21302_new_n4628_));
NOR2X1 NOR2X1_569 ( .A(core__abc_21302_new_n4628_), .B(core__abc_21302_new_n4620_), .Y(core__abc_21302_new_n4629_));
NOR2X1 NOR2X1_57 ( .A(core__abc_21302_new_n1144_), .B(core__abc_21302_new_n1141_), .Y(core__abc_21302_new_n1145_));
NOR2X1 NOR2X1_570 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n4688_), .Y(core__abc_21302_new_n4689_));
NOR2X1 NOR2X1_571 ( .A(core__abc_21302_new_n4647_), .B(core__abc_21302_new_n4700_), .Y(core__abc_21302_new_n4701_));
NOR2X1 NOR2X1_572 ( .A(core__abc_21302_new_n4700_), .B(core__abc_21302_new_n4646_), .Y(core__abc_21302_new_n4703_));
NOR2X1 NOR2X1_573 ( .A(core__abc_21302_new_n1521_), .B(core__abc_21302_new_n4708_), .Y(core__abc_21302_new_n4711_));
NOR2X1 NOR2X1_574 ( .A(core__abc_21302_new_n4711_), .B(core__abc_21302_new_n4710_), .Y(core__abc_21302_new_n4712_));
NOR2X1 NOR2X1_575 ( .A(core__abc_21302_new_n4719_), .B(core__abc_21302_new_n4721_), .Y(core__abc_21302_new_n4723_));
NOR2X1 NOR2X1_576 ( .A(core__abc_21302_new_n4747_), .B(core__abc_21302_new_n4746_), .Y(core__abc_21302_new_n4748_));
NOR2X1 NOR2X1_577 ( .A(core__abc_21302_new_n2462_), .B(core__abc_21302_new_n4768_), .Y(core__abc_21302_new_n4771_));
NOR2X1 NOR2X1_578 ( .A(core__abc_21302_new_n4770_), .B(core__abc_21302_new_n4773_), .Y(core__abc_21302_new_n4774_));
NOR2X1 NOR2X1_579 ( .A(core__abc_21302_new_n4775_), .B(core__abc_21302_new_n3449_), .Y(core__abc_21302_new_n4796_));
NOR2X1 NOR2X1_58 ( .A(core_siphash_word1_we_bF_buf10), .B(core_siphash_ctrl_reg_1_), .Y(core__abc_21302_new_n1150_));
NOR2X1 NOR2X1_580 ( .A(core_key_0_), .B(core__abc_21302_new_n2640__bF_buf1), .Y(core__abc_21302_new_n4822_));
NOR2X1 NOR2X1_581 ( .A(core__abc_21302_new_n4827_), .B(core__abc_21302_new_n4826_), .Y(core__abc_21302_new_n4828_));
NOR2X1 NOR2X1_582 ( .A(core__abc_21302_new_n3838_), .B(core__abc_21302_new_n3839_), .Y(core__abc_21302_new_n4832_));
NOR2X1 NOR2X1_583 ( .A(core_v1_reg_16_), .B(core__abc_21302_new_n4744_), .Y(core__abc_21302_new_n4840_));
NOR2X1 NOR2X1_584 ( .A(core__abc_21302_new_n4852_), .B(core__abc_21302_new_n4838_), .Y(core__abc_21302_new_n4853_));
NOR2X1 NOR2X1_585 ( .A(core_v1_reg_14_), .B(core__abc_21302_new_n4679_), .Y(core__abc_21302_new_n4855_));
NOR2X1 NOR2X1_586 ( .A(core__abc_21302_new_n4360_), .B(core__abc_21302_new_n4678_), .Y(core__abc_21302_new_n4856_));
NOR2X1 NOR2X1_587 ( .A(core__abc_21302_new_n4856_), .B(core__abc_21302_new_n4855_), .Y(core__abc_21302_new_n4857_));
NOR2X1 NOR2X1_588 ( .A(core__abc_21302_new_n4892_), .B(core__abc_21302_new_n4890_), .Y(core__abc_21302_new_n4893_));
NOR2X1 NOR2X1_589 ( .A(core__abc_21302_new_n3551_), .B(core__abc_21302_new_n3550_), .Y(core__abc_21302_new_n4905_));
NOR2X1 NOR2X1_59 ( .A(core_siphash_ctrl_reg_3_), .B(core_siphash_ctrl_reg_6_), .Y(core__abc_21302_new_n1152_));
NOR2X1 NOR2X1_590 ( .A(core_v1_reg_8_), .B(core__abc_21302_new_n4521_), .Y(core__abc_21302_new_n4917_));
NOR2X1 NOR2X1_591 ( .A(core__abc_21302_new_n4927_), .B(core__abc_21302_new_n4916_), .Y(core__abc_21302_new_n4928_));
NOR2X1 NOR2X1_592 ( .A(core__abc_21302_new_n4933_), .B(core__abc_21302_new_n4474_), .Y(core__abc_21302_new_n4936_));
NOR2X1 NOR2X1_593 ( .A(core__abc_21302_new_n4936_), .B(core__abc_21302_new_n4935_), .Y(core__abc_21302_new_n4950_));
NOR2X1 NOR2X1_594 ( .A(core__abc_21302_new_n4917_), .B(core__abc_21302_new_n4922_), .Y(core__abc_21302_new_n4956_));
NOR2X1 NOR2X1_595 ( .A(core__abc_21302_new_n5008_), .B(core__abc_21302_new_n5005_), .Y(core__abc_21302_new_n5009_));
NOR2X1 NOR2X1_596 ( .A(core_v1_reg_58_), .B(core__abc_21302_new_n4126_), .Y(core__abc_21302_new_n5017_));
NOR2X1 NOR2X1_597 ( .A(core__abc_21302_new_n1871_), .B(core__abc_21302_new_n4135_), .Y(core__abc_21302_new_n5018_));
NOR2X1 NOR2X1_598 ( .A(core__abc_21302_new_n5017_), .B(core__abc_21302_new_n5018_), .Y(core__abc_21302_new_n5019_));
NOR2X1 NOR2X1_599 ( .A(core__abc_21302_new_n2850_), .B(core__abc_21302_new_n5025_), .Y(core__abc_21302_new_n5026_));
NOR2X1 NOR2X1_6 ( .A(_abc_19873_new_n890_), .B(_abc_19873_new_n892_), .Y(_abc_19873_new_n893_));
NOR2X1 NOR2X1_60 ( .A(core_siphash_ctrl_reg_4_), .B(core__abc_21302_new_n1153_), .Y(core__abc_21302_new_n1154_));
NOR2X1 NOR2X1_600 ( .A(core__abc_21302_new_n5046_), .B(core__abc_21302_new_n5047_), .Y(core__abc_21302_new_n5048_));
NOR2X1 NOR2X1_601 ( .A(core__abc_21302_new_n5061_), .B(core__abc_21302_new_n5014_), .Y(core__abc_21302_new_n5062_));
NOR2X1 NOR2X1_602 ( .A(core__abc_21302_new_n5067_), .B(core__abc_21302_new_n5065_), .Y(core__abc_21302_new_n5068_));
NOR2X1 NOR2X1_603 ( .A(core__abc_21302_new_n2673__bF_buf5), .B(core__abc_21302_new_n5097_), .Y(core__abc_21302_new_n5098_));
NOR2X1 NOR2X1_604 ( .A(core__abc_21302_new_n5105_), .B(core__abc_21302_new_n5095_), .Y(core__abc_21302_new_n5106_));
NOR2X1 NOR2X1_605 ( .A(core__abc_21302_new_n3986_), .B(core__abc_21302_new_n3985_), .Y(core__abc_21302_new_n5111_));
NOR2X1 NOR2X1_606 ( .A(core__abc_21302_new_n5113_), .B(core__abc_21302_new_n2696_), .Y(core__abc_21302_new_n5116_));
NOR2X1 NOR2X1_607 ( .A(core__abc_21302_new_n2673__bF_buf4), .B(core__abc_21302_new_n5124_), .Y(core__abc_21302_new_n5125_));
NOR2X1 NOR2X1_608 ( .A(core__abc_21302_new_n5131_), .B(core__abc_21302_new_n2640__bF_buf11), .Y(core__abc_21302_new_n5132_));
NOR2X1 NOR2X1_609 ( .A(core__abc_21302_new_n5141_), .B(core__abc_21302_new_n5142_), .Y(core__abc_21302_new_n5155_));
NOR2X1 NOR2X1_61 ( .A(core__abc_21302_new_n1151_), .B(core__abc_21302_new_n1155_), .Y(core__abc_21302_new_n1156_));
NOR2X1 NOR2X1_610 ( .A(core__abc_21302_new_n5105_), .B(core__abc_21302_new_n5158_), .Y(core__abc_21302_new_n5161_));
NOR2X1 NOR2X1_611 ( .A(core__abc_21302_new_n5164_), .B(core__abc_21302_new_n5166_), .Y(core__abc_21302_new_n5167_));
NOR2X1 NOR2X1_612 ( .A(core__abc_21302_new_n1185__bF_buf5), .B(core__abc_21302_new_n5172_), .Y(core__0v2_reg_63_0__4_));
NOR2X1 NOR2X1_613 ( .A(core__abc_21302_new_n2673__bF_buf2), .B(core__abc_21302_new_n5181_), .Y(core__abc_21302_new_n5182_));
NOR2X1 NOR2X1_614 ( .A(core_key_6_), .B(core__abc_21302_new_n2640__bF_buf9), .Y(core__abc_21302_new_n5187_));
NOR2X1 NOR2X1_615 ( .A(core__abc_21302_new_n5154_), .B(core__abc_21302_new_n5180_), .Y(core__abc_21302_new_n5194_));
NOR2X1 NOR2X1_616 ( .A(core__abc_21302_new_n5192_), .B(core__abc_21302_new_n5195_), .Y(core__abc_21302_new_n5196_));
NOR2X1 NOR2X1_617 ( .A(core__abc_21302_new_n5205_), .B(core__abc_21302_new_n5196_), .Y(core__abc_21302_new_n5206_));
NOR2X1 NOR2X1_618 ( .A(core_v1_reg_26_), .B(core__abc_21302_new_n2890_), .Y(core__abc_21302_new_n5209_));
NOR2X1 NOR2X1_619 ( .A(core__abc_21302_new_n5210_), .B(core__abc_21302_new_n2881_), .Y(core__abc_21302_new_n5211_));
NOR2X1 NOR2X1_62 ( .A(core__abc_21302_new_n1148_), .B(core__abc_21302_new_n1157_), .Y(core__abc_21302_new_n1158_));
NOR2X1 NOR2X1_620 ( .A(core__abc_21302_new_n5236_), .B(core__abc_21302_new_n5237_), .Y(core__abc_21302_new_n5239_));
NOR2X1 NOR2X1_621 ( .A(core__abc_21302_new_n5246_), .B(core__abc_21302_new_n5245_), .Y(core__0v2_reg_63_0__8_));
NOR2X1 NOR2X1_622 ( .A(core__abc_21302_new_n5262_), .B(core__abc_21302_new_n5235_), .Y(core__abc_21302_new_n5263_));
NOR2X1 NOR2X1_623 ( .A(core__abc_21302_new_n5283_), .B(core__abc_21302_new_n5282_), .Y(core__0v2_reg_63_0__10_));
NOR2X1 NOR2X1_624 ( .A(core_v1_reg_30_), .B(core__abc_21302_new_n3058_), .Y(core__abc_21302_new_n5286_));
NOR2X1 NOR2X1_625 ( .A(core__abc_21302_new_n5298_), .B(core__abc_21302_new_n5085__bF_buf3), .Y(core__abc_21302_new_n5299_));
NOR2X1 NOR2X1_626 ( .A(core__abc_21302_new_n1185__bF_buf1), .B(core__abc_21302_new_n5301_), .Y(core__0v2_reg_63_0__11_));
NOR2X1 NOR2X1_627 ( .A(core__abc_21302_new_n5338_), .B(core__abc_21302_new_n5085__bF_buf2), .Y(core__abc_21302_new_n5339_));
NOR2X1 NOR2X1_628 ( .A(core__abc_21302_new_n2724_), .B(core__abc_21302_new_n2727_), .Y(core__abc_21302_new_n5353_));
NOR2X1 NOR2X1_629 ( .A(core__abc_21302_new_n5363_), .B(core__abc_21302_new_n5085__bF_buf1), .Y(core__abc_21302_new_n5364_));
NOR2X1 NOR2X1_63 ( .A(core_final_rounds_1_), .B(core_final_rounds_0_), .Y(core__abc_21302_new_n1161_));
NOR2X1 NOR2X1_630 ( .A(core__abc_21302_new_n1185__bF_buf0), .B(core__abc_21302_new_n5366_), .Y(core__0v2_reg_63_0__14_));
NOR2X1 NOR2X1_631 ( .A(core_v1_reg_34_), .B(core__abc_21302_new_n3280_), .Y(core__abc_21302_new_n5369_));
NOR2X1 NOR2X1_632 ( .A(core__abc_21302_new_n5370_), .B(core__abc_21302_new_n5369_), .Y(core__abc_21302_new_n5373_));
NOR2X1 NOR2X1_633 ( .A(core__abc_21302_new_n5383_), .B(core__abc_21302_new_n5085__bF_buf0), .Y(core__abc_21302_new_n5384_));
NOR2X1 NOR2X1_634 ( .A(core__abc_21302_new_n1185__bF_buf13), .B(core__abc_21302_new_n5386_), .Y(core__0v2_reg_63_0__15_));
NOR2X1 NOR2X1_635 ( .A(core__abc_21302_new_n5309_), .B(core__abc_21302_new_n5396_), .Y(core__abc_21302_new_n5397_));
NOR2X1 NOR2X1_636 ( .A(core__abc_21302_new_n5303_), .B(core__abc_21302_new_n5262_), .Y(core__abc_21302_new_n5399_));
NOR2X1 NOR2X1_637 ( .A(core__abc_21302_new_n5346_), .B(core__abc_21302_new_n5400_), .Y(core__abc_21302_new_n5401_));
NOR2X1 NOR2X1_638 ( .A(core__abc_21302_new_n5430_), .B(core__abc_21302_new_n5085__bF_buf5), .Y(core__abc_21302_new_n5431_));
NOR2X1 NOR2X1_639 ( .A(core__abc_21302_new_n5408_), .B(core__abc_21302_new_n5426_), .Y(core__abc_21302_new_n5443_));
NOR2X1 NOR2X1_64 ( .A(core_final_rounds_3_), .B(core__abc_21302_new_n1162_), .Y(core__abc_21302_new_n1169_));
NOR2X1 NOR2X1_640 ( .A(core__abc_21302_new_n5440_), .B(core__abc_21302_new_n5445_), .Y(core__abc_21302_new_n5447_));
NOR2X1 NOR2X1_641 ( .A(core__abc_21302_new_n5450_), .B(core__abc_21302_new_n5085__bF_buf4), .Y(core__abc_21302_new_n5451_));
NOR2X1 NOR2X1_642 ( .A(core__abc_21302_new_n5461_), .B(core__abc_21302_new_n5085__bF_buf3), .Y(core__abc_21302_new_n5462_));
NOR2X1 NOR2X1_643 ( .A(core__abc_21302_new_n1185__bF_buf12), .B(core__abc_21302_new_n5464_), .Y(core__0v2_reg_63_0__19_));
NOR2X1 NOR2X1_644 ( .A(core__abc_21302_new_n5469_), .B(core__abc_21302_new_n5473_), .Y(core__abc_21302_new_n5474_));
NOR2X1 NOR2X1_645 ( .A(core__abc_21302_new_n5470_), .B(core__abc_21302_new_n5476_), .Y(core__abc_21302_new_n5477_));
NOR2X1 NOR2X1_646 ( .A(core__abc_21302_new_n2990_), .B(core__abc_21302_new_n5480_), .Y(core__abc_21302_new_n5481_));
NOR2X1 NOR2X1_647 ( .A(core__abc_21302_new_n5488_), .B(core__abc_21302_new_n5085__bF_buf2), .Y(core__abc_21302_new_n5489_));
NOR2X1 NOR2X1_648 ( .A(core__abc_21302_new_n5502_), .B(core__abc_21302_new_n5085__bF_buf1), .Y(core__abc_21302_new_n5503_));
NOR2X1 NOR2X1_649 ( .A(core__abc_21302_new_n1185__bF_buf11), .B(core__abc_21302_new_n5505_), .Y(core__0v2_reg_63_0__21_));
NOR2X1 NOR2X1_65 ( .A(core__abc_21302_new_n1174_), .B(core__abc_21302_new_n1165_), .Y(core__abc_21302_new_n1175_));
NOR2X1 NOR2X1_650 ( .A(core__abc_21302_new_n3547_), .B(core__abc_21302_new_n3543_), .Y(core__abc_21302_new_n5508_));
NOR2X1 NOR2X1_651 ( .A(core__abc_21302_new_n5523_), .B(core__abc_21302_new_n5085__bF_buf0), .Y(core__abc_21302_new_n5524_));
NOR2X1 NOR2X1_652 ( .A(core__abc_21302_new_n1185__bF_buf10), .B(core__abc_21302_new_n5526_), .Y(core__0v2_reg_63_0__22_));
NOR2X1 NOR2X1_653 ( .A(core__abc_21302_new_n5541_), .B(core__abc_21302_new_n5085__bF_buf5), .Y(core__abc_21302_new_n5542_));
NOR2X1 NOR2X1_654 ( .A(core__abc_21302_new_n5514_), .B(core__abc_21302_new_n5545_), .Y(core__abc_21302_new_n5546_));
NOR2X1 NOR2X1_655 ( .A(core__abc_21302_new_n5554_), .B(core__abc_21302_new_n3164_), .Y(core__abc_21302_new_n5555_));
NOR2X1 NOR2X1_656 ( .A(core__abc_21302_new_n5551_), .B(core__abc_21302_new_n5553_), .Y(core__abc_21302_new_n5561_));
NOR2X1 NOR2X1_657 ( .A(core__abc_21302_new_n5565_), .B(core__abc_21302_new_n5085__bF_buf4), .Y(core__abc_21302_new_n5566_));
NOR2X1 NOR2X1_658 ( .A(core__abc_21302_new_n1185__bF_buf9), .B(core__abc_21302_new_n5568_), .Y(core__0v2_reg_63_0__24_));
NOR2X1 NOR2X1_659 ( .A(core__abc_21302_new_n5555_), .B(core__abc_21302_new_n5570_), .Y(core__abc_21302_new_n5571_));
NOR2X1 NOR2X1_66 ( .A(core_siphash_ctrl_reg_5_), .B(core__abc_21302_new_n1151_), .Y(core__abc_21302_new_n1176_));
NOR2X1 NOR2X1_660 ( .A(core__abc_21302_new_n5572_), .B(core__abc_21302_new_n3210_), .Y(core__abc_21302_new_n5574_));
NOR2X1 NOR2X1_661 ( .A(core__abc_21302_new_n5574_), .B(core__abc_21302_new_n5573_), .Y(core__abc_21302_new_n5576_));
NOR2X1 NOR2X1_662 ( .A(core__abc_21302_new_n5579_), .B(core__abc_21302_new_n5085__bF_buf3), .Y(core__abc_21302_new_n5580_));
NOR2X1 NOR2X1_663 ( .A(core__abc_21302_new_n5596_), .B(core__abc_21302_new_n5085__bF_buf2), .Y(core__abc_21302_new_n5597_));
NOR2X1 NOR2X1_664 ( .A(core__abc_21302_new_n1185__bF_buf8), .B(core__abc_21302_new_n5599_), .Y(core__0v2_reg_63_0__26_));
NOR2X1 NOR2X1_665 ( .A(core__abc_21302_new_n5613_), .B(core__abc_21302_new_n5085__bF_buf1), .Y(core__abc_21302_new_n5614_));
NOR2X1 NOR2X1_666 ( .A(core__abc_21302_new_n5607_), .B(core__abc_21302_new_n5587_), .Y(core__abc_21302_new_n5617_));
NOR2X1 NOR2X1_667 ( .A(core__abc_21302_new_n5591_), .B(core__abc_21302_new_n5621_), .Y(core__abc_21302_new_n5622_));
NOR2X1 NOR2X1_668 ( .A(core__abc_21302_new_n5623_), .B(core__abc_21302_new_n5622_), .Y(core__abc_21302_new_n5624_));
NOR2X1 NOR2X1_669 ( .A(core__abc_21302_new_n5550_), .B(core__abc_21302_new_n5547_), .Y(core__abc_21302_new_n5631_));
NOR2X1 NOR2X1_67 ( .A(core_finalize), .B(core_compress), .Y(core__abc_21302_new_n1181_));
NOR2X1 NOR2X1_670 ( .A(core__abc_21302_new_n5640_), .B(core__abc_21302_new_n5085__bF_buf0), .Y(core__abc_21302_new_n5641_));
NOR2X1 NOR2X1_671 ( .A(core__abc_21302_new_n1185__bF_buf7), .B(core__abc_21302_new_n5643_), .Y(core__0v2_reg_63_0__28_));
NOR2X1 NOR2X1_672 ( .A(core__abc_21302_new_n5651_), .B(core__abc_21302_new_n5652_), .Y(core__abc_21302_new_n5653_));
NOR2X1 NOR2X1_673 ( .A(core__abc_21302_new_n5658_), .B(core__abc_21302_new_n5085__bF_buf5), .Y(core__abc_21302_new_n5659_));
NOR2X1 NOR2X1_674 ( .A(core__abc_21302_new_n1185__bF_buf6), .B(core__abc_21302_new_n5661_), .Y(core__0v2_reg_63_0__29_));
NOR2X1 NOR2X1_675 ( .A(core__abc_21302_new_n5629_), .B(core__abc_21302_new_n5650_), .Y(core__abc_21302_new_n5663_));
NOR2X1 NOR2X1_676 ( .A(core__abc_21302_new_n3834_), .B(core__abc_21302_new_n3835_), .Y(core__abc_21302_new_n5668_));
NOR2X1 NOR2X1_677 ( .A(core__abc_21302_new_n5678_), .B(core__abc_21302_new_n5085__bF_buf4), .Y(core__abc_21302_new_n5679_));
NOR2X1 NOR2X1_678 ( .A(core__abc_21302_new_n1185__bF_buf5), .B(core__abc_21302_new_n5681_), .Y(core__0v2_reg_63_0__30_));
NOR2X1 NOR2X1_679 ( .A(core__abc_21302_new_n5669_), .B(core__abc_21302_new_n5667_), .Y(core__abc_21302_new_n5683_));
NOR2X1 NOR2X1_68 ( .A(core__abc_21302_new_n1184_), .B(core__abc_21302_new_n1185__bF_buf13), .Y(core__abc_21302_new_n1186_));
NOR2X1 NOR2X1_680 ( .A(core__abc_21302_new_n5695_), .B(core__abc_21302_new_n5085__bF_buf3), .Y(core__abc_21302_new_n5696_));
NOR2X1 NOR2X1_681 ( .A(core_key_32_), .B(core__abc_21302_new_n2640__bF_buf1), .Y(core__abc_21302_new_n5699_));
NOR2X1 NOR2X1_682 ( .A(core__abc_21302_new_n5701_), .B(core__abc_21302_new_n2673__bF_buf1), .Y(core__abc_21302_new_n5702_));
NOR2X1 NOR2X1_683 ( .A(core__abc_21302_new_n5716_), .B(core__abc_21302_new_n5085__bF_buf0), .Y(core__abc_21302_new_n5717_));
NOR2X1 NOR2X1_684 ( .A(core__abc_21302_new_n5724_), .B(core__abc_21302_new_n5085__bF_buf5), .Y(core__abc_21302_new_n5725_));
NOR2X1 NOR2X1_685 ( .A(core__abc_21302_new_n2673__bF_buf0), .B(core__abc_21302_new_n5730_), .Y(core__abc_21302_new_n5731_));
NOR2X1 NOR2X1_686 ( .A(core_key_37_), .B(core__abc_21302_new_n2640__bF_buf10), .Y(core__abc_21302_new_n5737_));
NOR2X1 NOR2X1_687 ( .A(core__abc_21302_new_n5748_), .B(core__abc_21302_new_n5085__bF_buf2), .Y(core__abc_21302_new_n5749_));
NOR2X1 NOR2X1_688 ( .A(core__abc_21302_new_n5760_), .B(core__abc_21302_new_n5085__bF_buf1), .Y(core__abc_21302_new_n5761_));
NOR2X1 NOR2X1_689 ( .A(core__abc_21302_new_n5085__bF_buf0), .B(core__abc_21302_new_n5768_), .Y(core__abc_21302_new_n5769_));
NOR2X1 NOR2X1_69 ( .A(core__abc_21302_new_n1188_), .B(core__abc_21302_new_n1145_), .Y(core__abc_21302_new_n1189_));
NOR2X1 NOR2X1_690 ( .A(core_key_41_), .B(core__abc_21302_new_n2640__bF_buf6), .Y(core__abc_21302_new_n5772_));
NOR2X1 NOR2X1_691 ( .A(core__abc_21302_new_n5786_), .B(core__abc_21302_new_n5085__bF_buf5), .Y(core__abc_21302_new_n5787_));
NOR2X1 NOR2X1_692 ( .A(core__abc_21302_new_n5797_), .B(core__abc_21302_new_n5800_), .Y(core__abc_21302_new_n5803_));
NOR2X1 NOR2X1_693 ( .A(core__abc_21302_new_n5803_), .B(core__abc_21302_new_n5802_), .Y(core__abc_21302_new_n5804_));
NOR2X1 NOR2X1_694 ( .A(core__abc_21302_new_n5807_), .B(core__abc_21302_new_n5085__bF_buf4), .Y(core__abc_21302_new_n5808_));
NOR2X1 NOR2X1_695 ( .A(core_key_45_), .B(core__abc_21302_new_n2640__bF_buf4), .Y(core__abc_21302_new_n5811_));
NOR2X1 NOR2X1_696 ( .A(core__abc_21302_new_n5823_), .B(core__abc_21302_new_n5085__bF_buf3), .Y(core__abc_21302_new_n5824_));
NOR2X1 NOR2X1_697 ( .A(core__abc_21302_new_n4993_), .B(core__abc_21302_new_n4975_), .Y(core__abc_21302_new_n5839_));
NOR2X1 NOR2X1_698 ( .A(core__abc_21302_new_n5085__bF_buf2), .B(core__abc_21302_new_n5845_), .Y(core__abc_21302_new_n5846_));
NOR2X1 NOR2X1_699 ( .A(core__abc_21302_new_n5853_), .B(core__abc_21302_new_n5085__bF_buf1), .Y(core__abc_21302_new_n5854_));
NOR2X1 NOR2X1_7 ( .A(_abc_19873_new_n890_), .B(_abc_19873_new_n880_), .Y(_abc_19873_new_n895_));
NOR2X1 NOR2X1_70 ( .A(core__abc_21302_new_n1185__bF_buf12), .B(core__abc_21302_new_n1151_), .Y(core__abc_21302_new_n1192_));
NOR2X1 NOR2X1_700 ( .A(core__abc_21302_new_n1185__bF_buf2), .B(core__abc_21302_new_n5856_), .Y(core__0v2_reg_63_0__49_));
NOR2X1 NOR2X1_701 ( .A(core__abc_21302_new_n4931_), .B(core__abc_21302_new_n5859_), .Y(core__abc_21302_new_n5862_));
NOR2X1 NOR2X1_702 ( .A(core__abc_21302_new_n5862_), .B(core__abc_21302_new_n5861_), .Y(core__abc_21302_new_n5863_));
NOR2X1 NOR2X1_703 ( .A(core__abc_21302_new_n5867_), .B(core__abc_21302_new_n5085__bF_buf0), .Y(core__abc_21302_new_n5868_));
NOR2X1 NOR2X1_704 ( .A(core__abc_21302_new_n5069_), .B(core__abc_21302_new_n5849_), .Y(core__abc_21302_new_n5878_));
NOR2X1 NOR2X1_705 ( .A(core__abc_21302_new_n4926_), .B(core__abc_21302_new_n5881_), .Y(core__abc_21302_new_n5882_));
NOR2X1 NOR2X1_706 ( .A(core__abc_21302_new_n5880_), .B(core__abc_21302_new_n5882_), .Y(core__abc_21302_new_n5883_));
NOR2X1 NOR2X1_707 ( .A(core__abc_21302_new_n5904_), .B(core__abc_21302_new_n5085__bF_buf5), .Y(core__abc_21302_new_n5905_));
NOR2X1 NOR2X1_708 ( .A(core__abc_21302_new_n1185__bF_buf1), .B(core__abc_21302_new_n5907_), .Y(core__0v2_reg_63_0__54_));
NOR2X1 NOR2X1_709 ( .A(core__abc_21302_new_n5916_), .B(core__abc_21302_new_n5085__bF_buf4), .Y(core__abc_21302_new_n5917_));
NOR2X1 NOR2X1_71 ( .A(core_initalize), .B(core__abc_21302_new_n1198_), .Y(core__abc_21302_new_n1199_));
NOR2X1 NOR2X1_710 ( .A(core__abc_21302_new_n1185__bF_buf0), .B(core__abc_21302_new_n5919_), .Y(core__0v2_reg_63_0__55_));
NOR2X1 NOR2X1_711 ( .A(core__abc_21302_new_n5928_), .B(core__abc_21302_new_n5927_), .Y(core__0v2_reg_63_0__56_));
NOR2X1 NOR2X1_712 ( .A(core_key_59_), .B(core__abc_21302_new_n2640__bF_buf6), .Y(core__abc_21302_new_n5944_));
NOR2X1 NOR2X1_713 ( .A(core__abc_21302_new_n5091_), .B(core__abc_21302_new_n5072_), .Y(core__abc_21302_new_n5953_));
NOR2X1 NOR2X1_714 ( .A(core__abc_21302_new_n4878_), .B(core__abc_21302_new_n5953_), .Y(core__abc_21302_new_n5955_));
NOR2X1 NOR2X1_715 ( .A(core__abc_21302_new_n4851_), .B(core__abc_21302_new_n5956_), .Y(core__abc_21302_new_n5957_));
NOR2X1 NOR2X1_716 ( .A(core__abc_21302_new_n5961_), .B(core__abc_21302_new_n5085__bF_buf3), .Y(core__abc_21302_new_n5962_));
NOR2X1 NOR2X1_717 ( .A(core__abc_21302_new_n5971_), .B(core__abc_21302_new_n5085__bF_buf2), .Y(core__abc_21302_new_n5972_));
NOR2X1 NOR2X1_718 ( .A(core__abc_21302_new_n1185__bF_buf13), .B(core__abc_21302_new_n5974_), .Y(core__0v2_reg_63_0__61_));
NOR2X1 NOR2X1_719 ( .A(core__abc_21302_new_n5980_), .B(core__abc_21302_new_n5085__bF_buf1), .Y(core__abc_21302_new_n5981_));
NOR2X1 NOR2X1_72 ( .A(core_initalize), .B(core__abc_21302_new_n1204_), .Y(core__abc_21302_new_n1205_));
NOR2X1 NOR2X1_720 ( .A(core__abc_21302_new_n1185__bF_buf12), .B(core__abc_21302_new_n5983_), .Y(core__0v2_reg_63_0__62_));
NOR2X1 NOR2X1_721 ( .A(core__abc_21302_new_n5985_), .B(core__abc_21302_new_n2640__bF_buf3), .Y(core__abc_21302_new_n5986_));
NOR2X1 NOR2X1_722 ( .A(core__abc_21302_new_n2138_), .B(core__abc_21302_new_n2638_), .Y(core__abc_21302_new_n5998_));
NOR2X1 NOR2X1_723 ( .A(core__abc_21302_new_n2363__bF_buf4), .B(core__abc_21302_new_n5995_), .Y(core__abc_21302_new_n6009_));
NOR2X1 NOR2X1_724 ( .A(core__abc_21302_new_n2673__bF_buf0), .B(core__abc_21302_new_n5714_), .Y(core__abc_21302_new_n6015_));
NOR2X1 NOR2X1_725 ( .A(core__abc_21302_new_n6047_), .B(core__abc_21302_new_n2640__bF_buf1), .Y(core__abc_21302_new_n6048_));
NOR2X1 NOR2X1_726 ( .A(core__abc_21302_new_n1185__bF_buf5), .B(core__abc_21302_new_n6098_), .Y(core__0v1_reg_63_0__13_));
NOR2X1 NOR2X1_727 ( .A(core__abc_21302_new_n5030_), .B(core__abc_21302_new_n5903_), .Y(core__abc_21302_new_n6154_));
NOR2X1 NOR2X1_728 ( .A(core__abc_21302_new_n3598_), .B(core__abc_21302_new_n6163_), .Y(core__abc_21302_new_n6164_));
NOR2X1 NOR2X1_729 ( .A(core__abc_21302_new_n1185__bF_buf4), .B(core__abc_21302_new_n6186_), .Y(core__0v1_reg_63_0__26_));
NOR2X1 NOR2X1_73 ( .A(core_v1_reg_0_), .B(core_v0_reg_0_), .Y(core__abc_21302_new_n1208_));
NOR2X1 NOR2X1_730 ( .A(core__abc_21302_new_n3902_), .B(core__abc_21302_new_n6216_), .Y(core__abc_21302_new_n6217_));
NOR2X1 NOR2X1_731 ( .A(core__abc_21302_new_n4902_), .B(core__abc_21302_new_n4903_), .Y(core__abc_21302_new_n6274_));
NOR2X1 NOR2X1_732 ( .A(core__abc_21302_new_n4840_), .B(core__abc_21302_new_n4845_), .Y(core__abc_21302_new_n6316_));
NOR2X1 NOR2X1_733 ( .A(core__abc_21302_new_n4492_), .B(core__abc_21302_new_n6361_), .Y(core__abc_21302_new_n6362_));
NOR2X1 NOR2X1_734 ( .A(core__abc_21302_new_n1185__bF_buf3), .B(core__abc_21302_new_n6364_), .Y(core__0v1_reg_63_0__52_));
NOR2X1 NOR2X1_735 ( .A(core__abc_21302_new_n4593_), .B(core__abc_21302_new_n6389_), .Y(core__abc_21302_new_n6390_));
NOR2X1 NOR2X1_736 ( .A(core__abc_21302_new_n5286_), .B(core__abc_21302_new_n5291_), .Y(core__abc_21302_new_n6418_));
NOR2X1 NOR2X1_737 ( .A(core__abc_21302_new_n6448_), .B(core__abc_21302_new_n2366_), .Y(core__abc_21302_new_n6449_));
NOR2X1 NOR2X1_738 ( .A(core__abc_21302_new_n2673__bF_buf10), .B(core__abc_21302_new_n2781_), .Y(core__abc_21302_new_n6478_));
NOR2X1 NOR2X1_739 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n2813_), .Y(core__abc_21302_new_n6485_));
NOR2X1 NOR2X1_74 ( .A(core__abc_21302_new_n1208_), .B(core__abc_21302_new_n1210_), .Y(core__abc_21302_new_n1211_));
NOR2X1 NOR2X1_740 ( .A(core__abc_21302_new_n2673__bF_buf7), .B(core__abc_21302_new_n2894_), .Y(core__abc_21302_new_n6499_));
NOR2X1 NOR2X1_741 ( .A(core__abc_21302_new_n2673__bF_buf6), .B(core__abc_21302_new_n2979_), .Y(core__abc_21302_new_n6513_));
NOR2X1 NOR2X1_742 ( .A(core__abc_21302_new_n2673__bF_buf5), .B(core__abc_21302_new_n3205_), .Y(core__abc_21302_new_n6550_));
NOR2X1 NOR2X1_743 ( .A(core__abc_21302_new_n2673__bF_buf3), .B(core__abc_21302_new_n3351_), .Y(core__abc_21302_new_n6571_));
NOR2X1 NOR2X1_744 ( .A(core__abc_21302_new_n2673__bF_buf2), .B(core__abc_21302_new_n3396_), .Y(core__abc_21302_new_n6578_));
NOR2X1 NOR2X1_745 ( .A(core__abc_21302_new_n2673__bF_buf0), .B(core__abc_21302_new_n3488_), .Y(core__abc_21302_new_n6593_));
NOR2X1 NOR2X1_746 ( .A(core__abc_21302_new_n2673__bF_buf11), .B(core__abc_21302_new_n3522_), .Y(core__abc_21302_new_n6600_));
NOR2X1 NOR2X1_747 ( .A(core__abc_21302_new_n2673__bF_buf8), .B(core__abc_21302_new_n3678_), .Y(core__abc_21302_new_n6628_));
NOR2X1 NOR2X1_748 ( .A(core__abc_21302_new_n2673__bF_buf6), .B(core__abc_21302_new_n3821_), .Y(core__abc_21302_new_n6659_));
NOR2X1 NOR2X1_749 ( .A(core__abc_21302_new_n2673__bF_buf0), .B(core__abc_21302_new_n4117_), .Y(core__abc_21302_new_n6719_));
NOR2X1 NOR2X1_75 ( .A(core_v2_reg_0_), .B(core_v3_reg_0_), .Y(core__abc_21302_new_n1212_));
NOR2X1 NOR2X1_750 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n4208_), .Y(core__abc_21302_new_n6739_));
NOR2X1 NOR2X1_751 ( .A(core__abc_21302_new_n2673__bF_buf6), .B(core__abc_21302_new_n4343_), .Y(core__abc_21302_new_n6775_));
NOR2X1 NOR2X1_752 ( .A(core__abc_21302_new_n2673__bF_buf3), .B(core__abc_21302_new_n4434_), .Y(core__abc_21302_new_n6795_));
NOR2X1 NOR2X1_753 ( .A(core__abc_21302_new_n2673__bF_buf2), .B(core__abc_21302_new_n4461_), .Y(core__abc_21302_new_n6802_));
NOR2X1 NOR2X1_754 ( .A(core__abc_21302_new_n2673__bF_buf10), .B(core__abc_21302_new_n6852_), .Y(core__abc_21302_new_n6853_));
NOR2X1 NOR2X1_755 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n4662_), .Y(core__abc_21302_new_n6860_));
NOR2X1 NOR2X1_756 ( .A(core__abc_21302_new_n2673__bF_buf6), .B(core__abc_21302_new_n6890_), .Y(core__abc_21302_new_n6891_));
NOR2X1 NOR2X1_757 ( .A(core__abc_21302_new_n1185__bF_buf8), .B(core__abc_21302_new_n1146_), .Y(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1474));
NOR2X1 NOR2X1_758 ( .A(core_long), .B(core__abc_21302_new_n6907_), .Y(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1470));
NOR2X1 NOR2X1_759 ( .A(core__abc_21302_new_n6909_), .B(core__abc_21302_new_n6907_), .Y(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1496));
NOR2X1 NOR2X1_76 ( .A(core__abc_21302_new_n1212_), .B(core__abc_21302_new_n1214_), .Y(core__abc_21302_new_n1215_));
NOR2X1 NOR2X1_760 ( .A(core__abc_21302_new_n1195_), .B(core__abc_21302_new_n6906_), .Y(core__abc_15204_auto_fsm_map_cc_118_implement_pattern_cache_1509));
NOR2X1 NOR2X1_77 ( .A(core_v1_reg_1_), .B(core_v0_reg_1_), .Y(core__abc_21302_new_n1220_));
NOR2X1 NOR2X1_78 ( .A(core__abc_21302_new_n1220_), .B(core__abc_21302_new_n1222_), .Y(core__abc_21302_new_n1223_));
NOR2X1 NOR2X1_79 ( .A(core_v2_reg_1_), .B(core_v3_reg_1_), .Y(core__abc_21302_new_n1226_));
NOR2X1 NOR2X1_8 ( .A(_abc_19873_new_n886_), .B(_abc_19873_new_n900_), .Y(_abc_19873_new_n901_));
NOR2X1 NOR2X1_80 ( .A(core__abc_21302_new_n1226_), .B(core__abc_21302_new_n1225_), .Y(core__abc_21302_new_n1227_));
NOR2X1 NOR2X1_81 ( .A(core_v1_reg_2_), .B(core_v0_reg_2_), .Y(core__abc_21302_new_n1233_));
NOR2X1 NOR2X1_82 ( .A(core__abc_21302_new_n1233_), .B(core__abc_21302_new_n1232_), .Y(core__abc_21302_new_n1234_));
NOR2X1 NOR2X1_83 ( .A(core_v2_reg_2_), .B(core_v3_reg_2_), .Y(core__abc_21302_new_n1236_));
NOR2X1 NOR2X1_84 ( .A(core__abc_21302_new_n1236_), .B(core__abc_21302_new_n1235_), .Y(core__abc_21302_new_n1237_));
NOR2X1 NOR2X1_85 ( .A(core_v2_reg_3_), .B(core_v3_reg_3_), .Y(core__abc_21302_new_n1245_));
NOR2X1 NOR2X1_86 ( .A(core__abc_21302_new_n1245_), .B(core__abc_21302_new_n1244_), .Y(core__abc_21302_new_n1246_));
NOR2X1 NOR2X1_87 ( .A(core_v2_reg_4_), .B(core_v3_reg_4_), .Y(core__abc_21302_new_n1255_));
NOR2X1 NOR2X1_88 ( .A(core__abc_21302_new_n1255_), .B(core__abc_21302_new_n1254_), .Y(core__abc_21302_new_n1256_));
NOR2X1 NOR2X1_89 ( .A(core_v2_reg_5_), .B(core_v3_reg_5_), .Y(core__abc_21302_new_n1267_));
NOR2X1 NOR2X1_9 ( .A(\addr[3] ), .B(\addr[2] ), .Y(_abc_19873_new_n903_));
NOR2X1 NOR2X1_90 ( .A(core__abc_21302_new_n1267_), .B(core__abc_21302_new_n1266_), .Y(core__abc_21302_new_n1268_));
NOR2X1 NOR2X1_91 ( .A(core_v2_reg_6_), .B(core_v3_reg_6_), .Y(core__abc_21302_new_n1277_));
NOR2X1 NOR2X1_92 ( .A(core__abc_21302_new_n1277_), .B(core__abc_21302_new_n1276_), .Y(core__abc_21302_new_n1278_));
NOR2X1 NOR2X1_93 ( .A(core_v2_reg_7_), .B(core_v3_reg_7_), .Y(core__abc_21302_new_n1287_));
NOR2X1 NOR2X1_94 ( .A(core__abc_21302_new_n1287_), .B(core__abc_21302_new_n1286_), .Y(core__abc_21302_new_n1288_));
NOR2X1 NOR2X1_95 ( .A(core_v1_reg_9_), .B(core_v0_reg_9_), .Y(core__abc_21302_new_n1301_));
NOR2X1 NOR2X1_96 ( .A(core__abc_21302_new_n1301_), .B(core__abc_21302_new_n1302_), .Y(core__abc_21302_new_n1303_));
NOR2X1 NOR2X1_97 ( .A(core_v2_reg_9_), .B(core_v3_reg_9_), .Y(core__abc_21302_new_n1305_));
NOR2X1 NOR2X1_98 ( .A(core_v1_reg_10_), .B(core_v0_reg_10_), .Y(core__abc_21302_new_n1312_));
NOR2X1 NOR2X1_99 ( .A(core__abc_21302_new_n1312_), .B(core__abc_21302_new_n1313_), .Y(core__abc_21302_new_n1314_));
NOR3X1 NOR3X1_1 ( .A(_abc_19873_new_n883_), .B(_abc_19873_new_n897_), .C(_abc_19873_new_n907_), .Y(_abc_19873_new_n908_));
NOR3X1 NOR3X1_10 ( .A(_abc_19873_new_n1012_), .B(_abc_19873_new_n1015_), .C(_abc_19873_new_n1009_), .Y(_abc_19873_new_n1016_));
NOR3X1 NOR3X1_11 ( .A(_abc_19873_new_n1019_), .B(_abc_19873_new_n1022_), .C(_abc_19873_new_n1026_), .Y(_abc_19873_new_n1027_));
NOR3X1 NOR3X1_12 ( .A(_abc_19873_new_n1030_), .B(_abc_19873_new_n1033_), .C(_abc_19873_new_n1036_), .Y(_abc_19873_new_n1037_));
NOR3X1 NOR3X1_13 ( .A(_abc_19873_new_n1040_), .B(_abc_19873_new_n1046_), .C(_abc_19873_new_n1043_), .Y(_abc_19873_new_n1047_));
NOR3X1 NOR3X1_14 ( .A(_abc_19873_new_n1054_), .B(_abc_19873_new_n1056_), .C(_abc_19873_new_n1051_), .Y(_abc_19873_new_n1057_));
NOR3X1 NOR3X1_15 ( .A(_abc_19873_new_n1073_), .B(_abc_19873_new_n1076_), .C(_abc_19873_new_n1070_), .Y(_abc_19873_new_n1077_));
NOR3X1 NOR3X1_16 ( .A(_abc_19873_new_n1080_), .B(_abc_19873_new_n1083_), .C(_abc_19873_new_n1086_), .Y(_abc_19873_new_n1087_));
NOR3X1 NOR3X1_17 ( .A(_abc_19873_new_n1089_), .B(_abc_19873_new_n1092_), .C(_abc_19873_new_n1095_), .Y(_abc_19873_new_n1096_));
NOR3X1 NOR3X1_18 ( .A(_abc_19873_new_n1099_), .B(_abc_19873_new_n1102_), .C(_abc_19873_new_n1105_), .Y(_abc_19873_new_n1106_));
NOR3X1 NOR3X1_19 ( .A(_abc_19873_new_n1108_), .B(_abc_19873_new_n1111_), .C(_abc_19873_new_n1114_), .Y(_abc_19873_new_n1115_));
NOR3X1 NOR3X1_2 ( .A(_abc_19873_new_n920_), .B(_abc_19873_new_n915_), .C(_abc_19873_new_n925_), .Y(_abc_19873_new_n926_));
NOR3X1 NOR3X1_20 ( .A(_abc_19873_new_n1118_), .B(_abc_19873_new_n1121_), .C(_abc_19873_new_n1124_), .Y(_abc_19873_new_n1125_));
NOR3X1 NOR3X1_21 ( .A(_abc_19873_new_n1127_), .B(_abc_19873_new_n1130_), .C(_abc_19873_new_n1133_), .Y(_abc_19873_new_n1134_));
NOR3X1 NOR3X1_22 ( .A(_abc_19873_new_n1149_), .B(_abc_19873_new_n1152_), .C(_abc_19873_new_n1146_), .Y(_abc_19873_new_n1153_));
NOR3X1 NOR3X1_23 ( .A(_abc_19873_new_n1168_), .B(_abc_19873_new_n1171_), .C(_abc_19873_new_n1165_), .Y(_abc_19873_new_n1172_));
NOR3X1 NOR3X1_24 ( .A(_abc_19873_new_n1178_), .B(_abc_19873_new_n1176_), .C(_abc_19873_new_n1181_), .Y(_abc_19873_new_n1182_));
NOR3X1 NOR3X1_25 ( .A(_abc_19873_new_n1019_), .B(_abc_19873_new_n1185_), .C(_abc_19873_new_n1189_), .Y(_abc_19873_new_n1190_));
NOR3X1 NOR3X1_26 ( .A(_abc_19873_new_n1200_), .B(_abc_19873_new_n1207_), .C(_abc_19873_new_n1204_), .Y(_abc_19873_new_n1208_));
NOR3X1 NOR3X1_27 ( .A(_abc_19873_new_n1211_), .B(_abc_19873_new_n1214_), .C(_abc_19873_new_n1217_), .Y(_abc_19873_new_n1218_));
NOR3X1 NOR3X1_28 ( .A(_abc_19873_new_n1220_), .B(_abc_19873_new_n1223_), .C(_abc_19873_new_n1226_), .Y(_abc_19873_new_n1227_));
NOR3X1 NOR3X1_29 ( .A(_abc_19873_new_n1237_), .B(_abc_19873_new_n1244_), .C(_abc_19873_new_n1241_), .Y(_abc_19873_new_n1245_));
NOR3X1 NOR3X1_3 ( .A(_abc_19873_new_n932_), .B(_abc_19873_new_n935_), .C(_abc_19873_new_n939_), .Y(_abc_19873_new_n940_));
NOR3X1 NOR3X1_30 ( .A(_abc_19873_new_n1263_), .B(_abc_19873_new_n1256_), .C(_abc_19873_new_n1260_), .Y(_abc_19873_new_n1264_));
NOR3X1 NOR3X1_31 ( .A(_abc_19873_new_n1278_), .B(_abc_19873_new_n1281_), .C(_abc_19873_new_n1275_), .Y(_abc_19873_new_n1282_));
NOR3X1 NOR3X1_32 ( .A(_abc_19873_new_n1292_), .B(_abc_19873_new_n1299_), .C(_abc_19873_new_n1296_), .Y(_abc_19873_new_n1300_));
NOR3X1 NOR3X1_33 ( .A(_abc_19873_new_n1314_), .B(_abc_19873_new_n1317_), .C(_abc_19873_new_n1311_), .Y(_abc_19873_new_n1318_));
NOR3X1 NOR3X1_34 ( .A(_abc_19873_new_n1321_), .B(_abc_19873_new_n1324_), .C(_abc_19873_new_n1327_), .Y(_abc_19873_new_n1328_));
NOR3X1 NOR3X1_35 ( .A(_abc_19873_new_n1019_), .B(_abc_19873_new_n1331_), .C(_abc_19873_new_n1335_), .Y(_abc_19873_new_n1336_));
NOR3X1 NOR3X1_36 ( .A(_abc_19873_new_n1346_), .B(_abc_19873_new_n1353_), .C(_abc_19873_new_n1350_), .Y(_abc_19873_new_n1354_));
NOR3X1 NOR3X1_37 ( .A(_abc_19873_new_n1357_), .B(_abc_19873_new_n1360_), .C(_abc_19873_new_n1363_), .Y(_abc_19873_new_n1364_));
NOR3X1 NOR3X1_38 ( .A(_abc_19873_new_n1366_), .B(_abc_19873_new_n1369_), .C(_abc_19873_new_n1372_), .Y(_abc_19873_new_n1373_));
NOR3X1 NOR3X1_39 ( .A(_abc_19873_new_n1383_), .B(_abc_19873_new_n1390_), .C(_abc_19873_new_n1387_), .Y(_abc_19873_new_n1391_));
NOR3X1 NOR3X1_4 ( .A(_abc_19873_new_n946_), .B(_abc_19873_new_n943_), .C(_abc_19873_new_n949_), .Y(_abc_19873_new_n950_));
NOR3X1 NOR3X1_40 ( .A(_abc_19873_new_n1401_), .B(_abc_19873_new_n1408_), .C(_abc_19873_new_n1405_), .Y(_abc_19873_new_n1409_));
NOR3X1 NOR3X1_41 ( .A(_abc_19873_new_n1412_), .B(_abc_19873_new_n1415_), .C(_abc_19873_new_n1418_), .Y(_abc_19873_new_n1419_));
NOR3X1 NOR3X1_42 ( .A(_abc_19873_new_n1421_), .B(_abc_19873_new_n1424_), .C(_abc_19873_new_n1427_), .Y(_abc_19873_new_n1428_));
NOR3X1 NOR3X1_43 ( .A(_abc_19873_new_n1431_), .B(_abc_19873_new_n1434_), .C(_abc_19873_new_n1437_), .Y(_abc_19873_new_n1438_));
NOR3X1 NOR3X1_44 ( .A(_abc_19873_new_n1440_), .B(_abc_19873_new_n1443_), .C(_abc_19873_new_n1446_), .Y(_abc_19873_new_n1447_));
NOR3X1 NOR3X1_45 ( .A(_abc_19873_new_n1457_), .B(_abc_19873_new_n1464_), .C(_abc_19873_new_n1461_), .Y(_abc_19873_new_n1465_));
NOR3X1 NOR3X1_46 ( .A(_abc_19873_new_n1476_), .B(_abc_19873_new_n1479_), .C(_abc_19873_new_n1484_), .Y(_abc_19873_new_n1485_));
NOR3X1 NOR3X1_47 ( .A(_abc_19873_new_n1495_), .B(_abc_19873_new_n1502_), .C(_abc_19873_new_n1499_), .Y(_abc_19873_new_n1503_));
NOR3X1 NOR3X1_48 ( .A(_abc_19873_new_n1506_), .B(_abc_19873_new_n1509_), .C(_abc_19873_new_n1512_), .Y(_abc_19873_new_n1513_));
NOR3X1 NOR3X1_49 ( .A(_abc_19873_new_n1515_), .B(_abc_19873_new_n1518_), .C(_abc_19873_new_n1521_), .Y(_abc_19873_new_n1522_));
NOR3X1 NOR3X1_5 ( .A(_abc_19873_new_n954_), .B(_abc_19873_new_n957_), .C(_abc_19873_new_n961_), .Y(_abc_19873_new_n962_));
NOR3X1 NOR3X1_50 ( .A(core_v3_reg_43_), .B(core__abc_21302_new_n3319_), .C(core__abc_21302_new_n3318_), .Y(core__abc_21302_new_n3320_));
NOR3X1 NOR3X1_51 ( .A(core__abc_21302_new_n3517_), .B(core__abc_21302_new_n3485_), .C(core__abc_21302_new_n3519_), .Y(core__abc_21302_new_n3604_));
NOR3X1 NOR3X1_52 ( .A(core__abc_21302_new_n3605_), .B(core__abc_21302_new_n3591_), .C(core__abc_21302_new_n3588_), .Y(core__abc_21302_new_n3606_));
NOR3X1 NOR3X1_53 ( .A(core__abc_21302_new_n3614_), .B(core__abc_21302_new_n3466_), .C(core__abc_21302_new_n3532_), .Y(core__abc_21302_new_n3615_));
NOR3X1 NOR3X1_54 ( .A(core__abc_21302_new_n3854_), .B(core__abc_21302_new_n3862_), .C(core__abc_21302_new_n3897_), .Y(core__abc_21302_new_n3911_));
NOR3X1 NOR3X1_55 ( .A(core__abc_21302_new_n4077_), .B(core__abc_21302_new_n4054_), .C(core__abc_21302_new_n4076_), .Y(core__abc_21302_new_n4091_));
NOR3X1 NOR3X1_56 ( .A(core__abc_21302_new_n3862_), .B(core__abc_21302_new_n3915_), .C(core__abc_21302_new_n3766_), .Y(core__abc_21302_new_n4162_));
NOR3X1 NOR3X1_57 ( .A(core__abc_21302_new_n4165_), .B(core__abc_21302_new_n3854_), .C(core__abc_21302_new_n4164_), .Y(core__abc_21302_new_n4166_));
NOR3X1 NOR3X1_58 ( .A(core__abc_21302_new_n4171_), .B(core__abc_21302_new_n4281_), .C(core__abc_21302_new_n4389_), .Y(core__abc_21302_new_n4420_));
NOR3X1 NOR3X1_59 ( .A(core__abc_21302_new_n4402_), .B(core__abc_21302_new_n4418_), .C(core__abc_21302_new_n4415_), .Y(core__abc_21302_new_n4430_));
NOR3X1 NOR3X1_6 ( .A(_abc_19873_new_n973_), .B(_abc_19873_new_n970_), .C(_abc_19873_new_n966_), .Y(_abc_19873_new_n974_));
NOR3X1 NOR3X1_60 ( .A(core__abc_21302_new_n4507_), .B(core__abc_21302_new_n4524_), .C(core__abc_21302_new_n4523_), .Y(core__abc_21302_new_n4539_));
NOR3X1 NOR3X1_61 ( .A(core__abc_21302_new_n4718_), .B(core__abc_21302_new_n4747_), .C(core__abc_21302_new_n4746_), .Y(core__abc_21302_new_n4764_));
NOR3X1 NOR3X1_62 ( .A(core__abc_21302_new_n4766_), .B(core__abc_21302_new_n4779_), .C(core__abc_21302_new_n4784_), .Y(core__abc_21302_new_n4787_));
NOR3X1 NOR3X1_63 ( .A(core__abc_21302_new_n4927_), .B(core__abc_21302_new_n5069_), .C(core__abc_21302_new_n4916_), .Y(core__abc_21302_new_n5070_));
NOR3X1 NOR3X1_64 ( .A(core__abc_21302_new_n4852_), .B(core__abc_21302_new_n4838_), .C(core__abc_21302_new_n5091_), .Y(core__abc_21302_new_n5092_));
NOR3X1 NOR3X1_65 ( .A(core__abc_21302_new_n5290_), .B(core__abc_21302_new_n5286_), .C(core__abc_21302_new_n5291_), .Y(core__abc_21302_new_n5305_));
NOR3X1 NOR3X1_66 ( .A(core__abc_21302_new_n5227_), .B(core__abc_21302_new_n5309_), .C(core__abc_21302_new_n5396_), .Y(core__abc_21302_new_n5471_));
NOR3X1 NOR3X1_7 ( .A(_abc_19873_new_n977_), .B(_abc_19873_new_n983_), .C(_abc_19873_new_n980_), .Y(_abc_19873_new_n984_));
NOR3X1 NOR3X1_8 ( .A(_abc_19873_new_n991_), .B(_abc_19873_new_n994_), .C(_abc_19873_new_n988_), .Y(_abc_19873_new_n995_));
NOR3X1 NOR3X1_9 ( .A(_abc_19873_new_n998_), .B(_abc_19873_new_n1004_), .C(_abc_19873_new_n1001_), .Y(_abc_19873_new_n1005_));
OAI21X1 OAI21X1_1 ( .A(_abc_19873_new_n870_), .B(_abc_19873_new_n878_), .C(_abc_19873_new_n882_), .Y(_abc_19873_new_n883_));
OAI21X1 OAI21X1_10 ( .A(_abc_19873_new_n905__bF_buf2), .B(_abc_19873_new_n895__bF_buf2), .C(_abc_19873_new_n877_), .Y(_abc_19873_new_n1018_));
OAI21X1 OAI21X1_100 ( .A(core_siphash_word_88_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf13), .Y(_abc_19873_new_n1671_));
OAI21X1 OAI21X1_1000 ( .A(core__abc_21302_new_n2485_), .B(core__abc_21302_new_n2397_), .C(core__abc_21302_new_n2489_), .Y(core__abc_21302_new_n4284_));
OAI21X1 OAI21X1_1001 ( .A(core__abc_21302_new_n4296_), .B(core__abc_21302_new_n4293_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n4297_));
OAI21X1 OAI21X1_1002 ( .A(core__abc_21302_new_n2363__bF_buf4), .B(core__abc_21302_new_n2368__bF_buf1), .C(core_v3_reg_45_), .Y(core__abc_21302_new_n4299_));
OAI21X1 OAI21X1_1003 ( .A(core__abc_21302_new_n4289_), .B(core__abc_21302_new_n4283_), .C(core__abc_21302_new_n4287_), .Y(core__abc_21302_new_n4300_));
OAI21X1 OAI21X1_1004 ( .A(core__abc_21302_new_n2706_), .B(core__abc_21302_new_n2708_), .C(core__abc_21302_new_n4307_), .Y(core__abc_21302_new_n4308_));
OAI21X1 OAI21X1_1005 ( .A(core__abc_21302_new_n4319_), .B(core__abc_21302_new_n4317_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n4320_));
OAI21X1 OAI21X1_1006 ( .A(core__abc_21302_new_n2363__bF_buf3), .B(core__abc_21302_new_n2368__bF_buf0), .C(core_v3_reg_46_), .Y(core__abc_21302_new_n4322_));
OAI21X1 OAI21X1_1007 ( .A(core__abc_21302_new_n2706_), .B(core__abc_21302_new_n2708_), .C(core__abc_21302_new_n4305_), .Y(core__abc_21302_new_n4325_));
OAI21X1 OAI21X1_1008 ( .A(core__abc_21302_new_n4324_), .B(core__abc_21302_new_n4283_), .C(core__abc_21302_new_n4329_), .Y(core__abc_21302_new_n4330_));
OAI21X1 OAI21X1_1009 ( .A(core__abc_21302_new_n2724_), .B(core__abc_21302_new_n2727_), .C(core_v3_reg_30_), .Y(core__abc_21302_new_n4331_));
OAI21X1 OAI21X1_101 ( .A(core_siphash_word_89_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf12), .Y(_abc_19873_new_n1674_));
OAI21X1 OAI21X1_1010 ( .A(core__abc_21302_new_n2415_), .B(core__abc_21302_new_n4333_), .C(core__abc_21302_new_n1360_), .Y(core__abc_21302_new_n4334_));
OAI21X1 OAI21X1_1011 ( .A(core__abc_21302_new_n1358_), .B(core__abc_21302_new_n1359_), .C(core__abc_21302_new_n4335_), .Y(core__abc_21302_new_n4336_));
OAI21X1 OAI21X1_1012 ( .A(core__abc_21302_new_n4161_), .B(core__abc_21302_new_n4172_), .C(core__abc_21302_new_n4346_), .Y(core__abc_21302_new_n4347_));
OAI21X1 OAI21X1_1013 ( .A(core__abc_21302_new_n4328_), .B(core__abc_21302_new_n4348_), .C(core__abc_21302_new_n4342_), .Y(core__abc_21302_new_n4349_));
OAI21X1 OAI21X1_1014 ( .A(core__abc_21302_new_n4354_), .B(core__abc_21302_new_n4352_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n4355_));
OAI21X1 OAI21X1_1015 ( .A(core__abc_21302_new_n2363__bF_buf2), .B(core__abc_21302_new_n2368__bF_buf4), .C(core_v3_reg_47_), .Y(core__abc_21302_new_n4357_));
OAI21X1 OAI21X1_1016 ( .A(core__abc_21302_new_n4360_), .B(core__abc_21302_new_n4361_), .C(core__abc_21302_new_n4334_), .Y(core__abc_21302_new_n4362_));
OAI21X1 OAI21X1_1017 ( .A(core__abc_21302_new_n2785_), .B(core__abc_21302_new_n2788_), .C(core__abc_21302_new_n4365_), .Y(core__abc_21302_new_n4366_));
OAI21X1 OAI21X1_1018 ( .A(core__abc_21302_new_n4277_), .B(core__abc_21302_new_n4282_), .C(core__abc_21302_new_n4323_), .Y(core__abc_21302_new_n4370_));
OAI21X1 OAI21X1_1019 ( .A(core__abc_21302_new_n4369_), .B(core__abc_21302_new_n4371_), .C(core__abc_21302_new_n4372_), .Y(core__abc_21302_new_n4373_));
OAI21X1 OAI21X1_102 ( .A(core_siphash_word_90_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf11), .Y(_abc_19873_new_n1676_));
OAI21X1 OAI21X1_1020 ( .A(core__abc_21302_new_n4369_), .B(core__abc_21302_new_n4371_), .C(core__abc_21302_new_n4367_), .Y(core__abc_21302_new_n4376_));
OAI21X1 OAI21X1_1021 ( .A(core__abc_21302_new_n2168__bF_buf5), .B(core__abc_21302_new_n4380_), .C(core__abc_21302_new_n4379_), .Y(core__abc_21302_new_n4381_));
OAI21X1 OAI21X1_1022 ( .A(core__abc_21302_new_n4381_), .B(core__abc_21302_new_n4378_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n4382_));
OAI21X1 OAI21X1_1023 ( .A(core__abc_21302_new_n2363__bF_buf1), .B(core__abc_21302_new_n2368__bF_buf3), .C(core_v3_reg_48_), .Y(core__abc_21302_new_n4384_));
OAI21X1 OAI21X1_1024 ( .A(core__abc_21302_new_n4365_), .B(core__abc_21302_new_n2789_), .C(core__abc_21302_new_n4340_), .Y(core__abc_21302_new_n4392_));
OAI21X1 OAI21X1_1025 ( .A(core__abc_21302_new_n4389_), .B(core__abc_21302_new_n4345_), .C(core__abc_21302_new_n4393_), .Y(core__abc_21302_new_n4394_));
OAI21X1 OAI21X1_1026 ( .A(core__abc_21302_new_n4388_), .B(core__abc_21302_new_n3931_), .C(core__abc_21302_new_n4395_), .Y(core__abc_21302_new_n4396_));
OAI21X1 OAI21X1_1027 ( .A(core__abc_21302_new_n4385_), .B(core__abc_21302_new_n4407_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n4408_));
OAI21X1 OAI21X1_1028 ( .A(core__abc_21302_new_n2363__bF_buf0), .B(core__abc_21302_new_n2368__bF_buf2), .C(core_v3_reg_49_), .Y(core__abc_21302_new_n4410_));
OAI21X1 OAI21X1_1029 ( .A(core__abc_21302_new_n1382_), .B(core__abc_21302_new_n2492_), .C(core__abc_21302_new_n4411_), .Y(core__abc_21302_new_n4412_));
OAI21X1 OAI21X1_103 ( .A(core_siphash_word_91_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf10), .Y(_abc_19873_new_n1678_));
OAI21X1 OAI21X1_1030 ( .A(core__abc_21302_new_n2869_), .B(core__abc_21302_new_n2870_), .C(core__abc_21302_new_n4416_), .Y(core__abc_21302_new_n4417_));
OAI21X1 OAI21X1_1031 ( .A(core__abc_21302_new_n3913_), .B(core__abc_21302_new_n3920_), .C(core__abc_21302_new_n4420_), .Y(core__abc_21302_new_n4421_));
OAI21X1 OAI21X1_1032 ( .A(core__abc_21302_new_n4402_), .B(core__abc_21302_new_n4422_), .C(core__abc_21302_new_n4400_), .Y(core__abc_21302_new_n4423_));
OAI21X1 OAI21X1_1033 ( .A(core__abc_21302_new_n4429_), .B(core__abc_21302_new_n4426_), .C(core__abc_21302_new_n4430_), .Y(core__abc_21302_new_n4431_));
OAI21X1 OAI21X1_1034 ( .A(core__abc_21302_new_n4400_), .B(core__abc_21302_new_n4425_), .C(core__abc_21302_new_n4431_), .Y(core__abc_21302_new_n4432_));
OAI21X1 OAI21X1_1035 ( .A(core__abc_21302_new_n4432_), .B(core__abc_21302_new_n4424_), .C(core__abc_21302_new_n3778_), .Y(core__abc_21302_new_n4433_));
OAI21X1 OAI21X1_1036 ( .A(core__abc_21302_new_n4439_), .B(core__abc_21302_new_n4436_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n4440_));
OAI21X1 OAI21X1_1037 ( .A(core__abc_21302_new_n2363__bF_buf5), .B(core__abc_21302_new_n2368__bF_buf1), .C(core_v3_reg_50_), .Y(core__abc_21302_new_n4442_));
OAI21X1 OAI21X1_1038 ( .A(core__abc_21302_new_n4444_), .B(core__abc_21302_new_n4445_), .C(core__abc_21302_new_n1407_), .Y(core__abc_21302_new_n4446_));
OAI21X1 OAI21X1_1039 ( .A(core__abc_21302_new_n1405_), .B(core__abc_21302_new_n1406_), .C(core__abc_21302_new_n4447_), .Y(core__abc_21302_new_n4448_));
OAI21X1 OAI21X1_104 ( .A(core_siphash_word_92_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf9), .Y(_abc_19873_new_n1681_));
OAI21X1 OAI21X1_1040 ( .A(core__abc_21302_new_n4466_), .B(core__abc_21302_new_n4464_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n4467_));
OAI21X1 OAI21X1_1041 ( .A(core__abc_21302_new_n2363__bF_buf4), .B(core__abc_21302_new_n2368__bF_buf0), .C(core_v3_reg_51_), .Y(core__abc_21302_new_n4469_));
OAI21X1 OAI21X1_1042 ( .A(core__abc_21302_new_n1405_), .B(core__abc_21302_new_n4447_), .C(core__abc_21302_new_n2441_), .Y(core__abc_21302_new_n4470_));
OAI21X1 OAI21X1_1043 ( .A(core__abc_21302_new_n1417_), .B(core__abc_21302_new_n1418_), .C(core__abc_21302_new_n4471_), .Y(core__abc_21302_new_n4472_));
OAI21X1 OAI21X1_1044 ( .A(core__abc_21302_new_n4450_), .B(core__abc_21302_new_n4455_), .C(core__abc_21302_new_n4480_), .Y(core__abc_21302_new_n4481_));
OAI21X1 OAI21X1_1045 ( .A(core__abc_21302_new_n4488_), .B(core__abc_21302_new_n4485_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n4489_));
OAI21X1 OAI21X1_1046 ( .A(core__abc_21302_new_n2363__bF_buf3), .B(core__abc_21302_new_n2368__bF_buf4), .C(core_v3_reg_52_), .Y(core__abc_21302_new_n4491_));
OAI21X1 OAI21X1_1047 ( .A(core__abc_21302_new_n4443_), .B(core__abc_21302_new_n4493_), .C(core__abc_21302_new_n4494_), .Y(core__abc_21302_new_n4495_));
OAI21X1 OAI21X1_1048 ( .A(core__abc_21302_new_n4498_), .B(core__abc_21302_new_n4422_), .C(core__abc_21302_new_n4496_), .Y(core__abc_21302_new_n4499_));
OAI21X1 OAI21X1_1049 ( .A(core__abc_21302_new_n2445_), .B(core__abc_21302_new_n4500_), .C(core__abc_21302_new_n1431_), .Y(core__abc_21302_new_n4501_));
OAI21X1 OAI21X1_105 ( .A(core_siphash_word_93_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf8), .Y(_abc_19873_new_n1683_));
OAI21X1 OAI21X1_1050 ( .A(core__abc_21302_new_n1429_), .B(core__abc_21302_new_n1430_), .C(core__abc_21302_new_n4502_), .Y(core__abc_21302_new_n4503_));
OAI21X1 OAI21X1_1051 ( .A(core__abc_21302_new_n4492_), .B(core__abc_21302_new_n4511_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n4512_));
OAI21X1 OAI21X1_1052 ( .A(core__abc_21302_new_n2363__bF_buf2), .B(core__abc_21302_new_n2368__bF_buf3), .C(core_v3_reg_53_), .Y(core__abc_21302_new_n4514_));
OAI21X1 OAI21X1_1053 ( .A(core__abc_21302_new_n4495_), .B(core__abc_21302_new_n4515_), .C(core__abc_21302_new_n4516_), .Y(core__abc_21302_new_n4517_));
OAI21X1 OAI21X1_1054 ( .A(core__abc_21302_new_n1429_), .B(core__abc_21302_new_n4502_), .C(core__abc_21302_new_n2446_), .Y(core__abc_21302_new_n4519_));
OAI21X1 OAI21X1_1055 ( .A(core__abc_21302_new_n1441_), .B(core__abc_21302_new_n1442_), .C(core__abc_21302_new_n4519_), .Y(core__abc_21302_new_n4520_));
OAI21X1 OAI21X1_1056 ( .A(core__abc_21302_new_n2991_), .B(core__abc_21302_new_n4504_), .C(core__abc_21302_new_n4517_), .Y(core__abc_21302_new_n4527_));
OAI21X1 OAI21X1_1057 ( .A(core__abc_21302_new_n4523_), .B(core__abc_21302_new_n4524_), .C(core__abc_21302_new_n4527_), .Y(core__abc_21302_new_n4528_));
OAI21X1 OAI21X1_1058 ( .A(core__abc_21302_new_n4535_), .B(core__abc_21302_new_n4533_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n4536_));
OAI21X1 OAI21X1_1059 ( .A(core__abc_21302_new_n2363__bF_buf1), .B(core__abc_21302_new_n2368__bF_buf2), .C(core_v3_reg_54_), .Y(core__abc_21302_new_n4538_));
OAI21X1 OAI21X1_106 ( .A(core_siphash_word_94_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf7), .Y(_abc_19873_new_n1686_));
OAI21X1 OAI21X1_1060 ( .A(core__abc_21302_new_n4495_), .B(core__abc_21302_new_n4515_), .C(core__abc_21302_new_n4539_), .Y(core__abc_21302_new_n4540_));
OAI21X1 OAI21X1_1061 ( .A(core__abc_21302_new_n4505_), .B(core__abc_21302_new_n4524_), .C(core__abc_21302_new_n4541_), .Y(core__abc_21302_new_n4542_));
OAI21X1 OAI21X1_1062 ( .A(core__abc_21302_new_n2429_), .B(core__abc_21302_new_n4502_), .C(core__abc_21302_new_n2449_), .Y(core__abc_21302_new_n4544_));
OAI21X1 OAI21X1_1063 ( .A(core__abc_21302_new_n4546_), .B(core__abc_21302_new_n4547_), .C(core__abc_21302_new_n3073_), .Y(core__abc_21302_new_n4550_));
OAI21X1 OAI21X1_1064 ( .A(core__abc_21302_new_n4552_), .B(core__abc_21302_new_n4554_), .C(core__abc_21302_new_n3971_), .Y(core__abc_21302_new_n4555_));
OAI21X1 OAI21X1_1065 ( .A(core__abc_21302_new_n4560_), .B(core__abc_21302_new_n4558_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n4561_));
OAI21X1 OAI21X1_1066 ( .A(core__abc_21302_new_n2363__bF_buf0), .B(core__abc_21302_new_n2368__bF_buf1), .C(core_v3_reg_55_), .Y(core__abc_21302_new_n4563_));
OAI21X1 OAI21X1_1067 ( .A(core__abc_21302_new_n1454_), .B(core__abc_21302_new_n4546_), .C(core__abc_21302_new_n4571_), .Y(core__abc_21302_new_n4572_));
OAI21X1 OAI21X1_1068 ( .A(core__abc_21302_new_n3117_), .B(core__abc_21302_new_n3119_), .C(core__abc_21302_new_n4575_), .Y(core__abc_21302_new_n4576_));
OAI21X1 OAI21X1_1069 ( .A(core__abc_21302_new_n4579_), .B(core__abc_21302_new_n4552_), .C(core__abc_21302_new_n4580_), .Y(core__abc_21302_new_n4581_));
OAI21X1 OAI21X1_107 ( .A(core_siphash_word_95_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf6), .Y(_abc_19873_new_n1688_));
OAI21X1 OAI21X1_1070 ( .A(core__abc_21302_new_n4579_), .B(core__abc_21302_new_n4552_), .C(core__abc_21302_new_n4577_), .Y(core__abc_21302_new_n4584_));
OAI21X1 OAI21X1_1071 ( .A(core__abc_21302_new_n2168__bF_buf10), .B(core__abc_21302_new_n4588_), .C(core__abc_21302_new_n4587_), .Y(core__abc_21302_new_n4589_));
OAI21X1 OAI21X1_1072 ( .A(core__abc_21302_new_n4589_), .B(core__abc_21302_new_n4586_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n4590_));
OAI21X1 OAI21X1_1073 ( .A(core__abc_21302_new_n2363__bF_buf5), .B(core__abc_21302_new_n2368__bF_buf0), .C(core_v3_reg_56_), .Y(core__abc_21302_new_n4592_));
OAI21X1 OAI21X1_1074 ( .A(core__abc_21302_new_n4575_), .B(core__abc_21302_new_n3120_), .C(core__abc_21302_new_n4549_), .Y(core__abc_21302_new_n4600_));
OAI21X1 OAI21X1_1075 ( .A(core__abc_21302_new_n2433_), .B(core__abc_21302_new_n2492_), .C(core__abc_21302_new_n2452_), .Y(core__abc_21302_new_n4604_));
OAI21X1 OAI21X1_1076 ( .A(core__abc_21302_new_n1473_), .B(core__abc_21302_new_n1474_), .C(core__abc_21302_new_n4606_), .Y(core__abc_21302_new_n4607_));
OAI21X1 OAI21X1_1077 ( .A(core__abc_21302_new_n4593_), .B(core__abc_21302_new_n4613_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n4614_));
OAI21X1 OAI21X1_1078 ( .A(core__abc_21302_new_n2363__bF_buf4), .B(core__abc_21302_new_n2368__bF_buf4), .C(core_v3_reg_57_), .Y(core__abc_21302_new_n4616_));
OAI21X1 OAI21X1_1079 ( .A(core__abc_21302_new_n4602_), .B(core__abc_21302_new_n4597_), .C(core__abc_21302_new_n4609_), .Y(core__abc_21302_new_n4619_));
OAI21X1 OAI21X1_108 ( .A(core_siphash_word_32_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf5), .Y(_abc_19873_new_n1690_));
OAI21X1 OAI21X1_1080 ( .A(core__abc_21302_new_n4618_), .B(core__abc_21302_new_n4608_), .C(core__abc_21302_new_n4619_), .Y(core__abc_21302_new_n4620_));
OAI21X1 OAI21X1_1081 ( .A(core__abc_21302_new_n2453_), .B(core__abc_21302_new_n2454_), .C(core__abc_21302_new_n4605_), .Y(core__abc_21302_new_n4623_));
OAI21X1 OAI21X1_1082 ( .A(core__abc_21302_new_n4629_), .B(core__abc_21302_new_n4631_), .C(core__abc_21302_new_n4617_), .Y(core__abc_21302_new_n4632_));
OAI21X1 OAI21X1_1083 ( .A(core__abc_21302_new_n2168__bF_buf8), .B(core__abc_21302_new_n4637_), .C(core__abc_21302_new_n4636_), .Y(core__abc_21302_new_n4638_));
OAI21X1 OAI21X1_1084 ( .A(core__abc_21302_new_n4638_), .B(core__abc_21302_new_n4635_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n4639_));
OAI21X1 OAI21X1_1085 ( .A(core__abc_21302_new_n2363__bF_buf3), .B(core__abc_21302_new_n2368__bF_buf3), .C(core_v3_reg_58_), .Y(core__abc_21302_new_n4641_));
OAI21X1 OAI21X1_1086 ( .A(core__abc_21302_new_n4618_), .B(core__abc_21302_new_n4608_), .C(core__abc_21302_new_n4644_), .Y(core__abc_21302_new_n4645_));
OAI21X1 OAI21X1_1087 ( .A(core__abc_21302_new_n4602_), .B(core__abc_21302_new_n4597_), .C(core__abc_21302_new_n4648_), .Y(core__abc_21302_new_n4649_));
OAI21X1 OAI21X1_1088 ( .A(core__abc_21302_new_n2424_), .B(core__abc_21302_new_n4606_), .C(core__abc_21302_new_n2457_), .Y(core__abc_21302_new_n4650_));
OAI21X1 OAI21X1_1089 ( .A(core__abc_21302_new_n3249_), .B(core__abc_21302_new_n3250_), .C(core_v3_reg_42_), .Y(core__abc_21302_new_n4654_));
OAI21X1 OAI21X1_109 ( .A(core_siphash_word_33_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf4), .Y(_abc_19873_new_n1692_));
OAI21X1 OAI21X1_1090 ( .A(core__abc_21302_new_n4668_), .B(core__abc_21302_new_n4666_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n4669_));
OAI21X1 OAI21X1_1091 ( .A(core__abc_21302_new_n3319_), .B(core__abc_21302_new_n3318_), .C(core_v3_reg_43_), .Y(core__abc_21302_new_n4672_));
OAI21X1 OAI21X1_1092 ( .A(core__abc_21302_new_n1507_), .B(core__abc_21302_new_n1508_), .C(core__abc_21302_new_n4674_), .Y(core__abc_21302_new_n4675_));
OAI21X1 OAI21X1_1093 ( .A(core__abc_21302_new_n1496_), .B(core__abc_21302_new_n4676_), .C(core__abc_21302_new_n1509_), .Y(core__abc_21302_new_n4677_));
OAI21X1 OAI21X1_1094 ( .A(core__abc_21302_new_n3316_), .B(core__abc_21302_new_n3320_), .C(core__abc_21302_new_n4678_), .Y(core__abc_21302_new_n4681_));
OAI21X1 OAI21X1_1095 ( .A(core__abc_21302_new_n4684_), .B(core__abc_21302_new_n4659_), .C(core__abc_21302_new_n4685_), .Y(core__abc_21302_new_n4686_));
OAI21X1 OAI21X1_1096 ( .A(core__abc_21302_new_n4692_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n2369__bF_buf0), .Y(core__abc_21302_new_n4693_));
OAI21X1 OAI21X1_1097 ( .A(core_v3_reg_59_), .B(core__abc_21302_new_n2369__bF_buf7), .C(reset_n_bF_buf0), .Y(core__abc_21302_new_n4695_));
OAI21X1 OAI21X1_1098 ( .A(core__abc_21302_new_n2363__bF_buf2), .B(core__abc_21302_new_n2368__bF_buf2), .C(core_v3_reg_60_), .Y(core__abc_21302_new_n4697_));
OAI21X1 OAI21X1_1099 ( .A(core__abc_21302_new_n3316_), .B(core__abc_21302_new_n3320_), .C(core__abc_21302_new_n4679_), .Y(core__abc_21302_new_n4698_));
OAI21X1 OAI21X1_11 ( .A(_abc_19873_new_n1028_), .B(_abc_19873_new_n960__bF_buf1), .C(_abc_19873_new_n1029_), .Y(_abc_19873_new_n1030_));
OAI21X1 OAI21X1_110 ( .A(core_siphash_word_34_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf3), .Y(_abc_19873_new_n1695_));
OAI21X1 OAI21X1_1100 ( .A(core__abc_21302_new_n4602_), .B(core__abc_21302_new_n4597_), .C(core__abc_21302_new_n4701_), .Y(core__abc_21302_new_n4702_));
OAI21X1 OAI21X1_1101 ( .A(core__abc_21302_new_n3255_), .B(core__abc_21302_new_n4651_), .C(core__abc_21302_new_n4698_), .Y(core__abc_21302_new_n4704_));
OAI21X1 OAI21X1_1102 ( .A(core__abc_21302_new_n3355_), .B(core__abc_21302_new_n3354_), .C(core_v3_reg_44_), .Y(core__abc_21302_new_n4714_));
OAI21X1 OAI21X1_1103 ( .A(core__abc_21302_new_n4727_), .B(core__abc_21302_new_n4725_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n4728_));
OAI21X1 OAI21X1_1104 ( .A(core__abc_21302_new_n2363__bF_buf1), .B(core__abc_21302_new_n2368__bF_buf1), .C(core_v3_reg_61_), .Y(core__abc_21302_new_n4730_));
OAI21X1 OAI21X1_1105 ( .A(core__abc_21302_new_n4429_), .B(core__abc_21302_new_n4426_), .C(core__abc_21302_new_n4732_), .Y(core__abc_21302_new_n4733_));
OAI21X1 OAI21X1_1106 ( .A(core__abc_21302_new_n4679_), .B(core__abc_21302_new_n3322_), .C(core__abc_21302_new_n4704_), .Y(core__abc_21302_new_n4737_));
OAI21X1 OAI21X1_1107 ( .A(core__abc_21302_new_n4646_), .B(core__abc_21302_new_n4700_), .C(core__abc_21302_new_n4737_), .Y(core__abc_21302_new_n4738_));
OAI21X1 OAI21X1_1108 ( .A(core__abc_21302_new_n4738_), .B(core__abc_21302_new_n4736_), .C(core__abc_21302_new_n4739_), .Y(core__abc_21302_new_n4740_));
OAI21X1 OAI21X1_1109 ( .A(core__abc_21302_new_n1520_), .B(core__abc_21302_new_n4710_), .C(core__abc_21302_new_n4742_), .Y(core__abc_21302_new_n4743_));
OAI21X1 OAI21X1_111 ( .A(core_siphash_word_35_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf2), .Y(_abc_19873_new_n1698_));
OAI21X1 OAI21X1_1110 ( .A(core__abc_21302_new_n4750_), .B(core__abc_21302_new_n4719_), .C(core__abc_21302_new_n4751_), .Y(core__abc_21302_new_n4752_));
OAI21X1 OAI21X1_1111 ( .A(core__abc_21302_new_n4750_), .B(core__abc_21302_new_n4719_), .C(core__abc_21302_new_n4748_), .Y(core__abc_21302_new_n4755_));
OAI21X1 OAI21X1_1112 ( .A(core__abc_21302_new_n4759_), .B(core__abc_21302_new_n4757_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n4760_));
OAI21X1 OAI21X1_1113 ( .A(core__abc_21302_new_n2363__bF_buf0), .B(core__abc_21302_new_n2368__bF_buf0), .C(core_v3_reg_62_), .Y(core__abc_21302_new_n4762_));
OAI21X1 OAI21X1_1114 ( .A(core__abc_21302_new_n4738_), .B(core__abc_21302_new_n4736_), .C(core__abc_21302_new_n4764_), .Y(core__abc_21302_new_n4765_));
OAI21X1 OAI21X1_1115 ( .A(core__abc_21302_new_n4713_), .B(core__abc_21302_new_n4747_), .C(core__abc_21302_new_n4745_), .Y(core__abc_21302_new_n4766_));
OAI21X1 OAI21X1_1116 ( .A(core__abc_21302_new_n2462_), .B(core__abc_21302_new_n4768_), .C(core__abc_21302_new_n1546_), .Y(core__abc_21302_new_n4769_));
OAI21X1 OAI21X1_1117 ( .A(core__abc_21302_new_n1544_), .B(core__abc_21302_new_n1545_), .C(core__abc_21302_new_n4771_), .Y(core__abc_21302_new_n4772_));
OAI21X1 OAI21X1_1118 ( .A(core__abc_21302_new_n3446_), .B(core__abc_21302_new_n4777_), .C(core__abc_21302_new_n4774_), .Y(core__abc_21302_new_n4778_));
OAI21X1 OAI21X1_1119 ( .A(core__abc_21302_new_n4766_), .B(core__abc_21302_new_n4784_), .C(core__abc_21302_new_n4779_), .Y(core__abc_21302_new_n4785_));
OAI21X1 OAI21X1_112 ( .A(core_siphash_word_36_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf1), .Y(_abc_19873_new_n1701_));
OAI21X1 OAI21X1_1120 ( .A(core__abc_21302_new_n4787_), .B(core__abc_21302_new_n4788_), .C(core__abc_21302_new_n4232_), .Y(core__abc_21302_new_n4789_));
OAI21X1 OAI21X1_1121 ( .A(core__abc_21302_new_n4792_), .B(core__abc_21302_new_n4790_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n4793_));
OAI21X1 OAI21X1_1122 ( .A(core__abc_21302_new_n1544_), .B(core__abc_21302_new_n4771_), .C(core__abc_21302_new_n4798_), .Y(core__abc_21302_new_n4800_));
OAI21X1 OAI21X1_1123 ( .A(core__abc_21302_new_n1556_), .B(core__abc_21302_new_n1557_), .C(core__abc_21302_new_n4800_), .Y(core__abc_21302_new_n4801_));
OAI21X1 OAI21X1_1124 ( .A(core__abc_21302_new_n4796_), .B(core__abc_21302_new_n4788_), .C(core__abc_21302_new_n4808_), .Y(core__abc_21302_new_n4809_));
OAI21X1 OAI21X1_1125 ( .A(core__abc_21302_new_n4796_), .B(core__abc_21302_new_n4788_), .C(core__abc_21302_new_n4806_), .Y(core__abc_21302_new_n4813_));
OAI21X1 OAI21X1_1126 ( .A(core__abc_21302_new_n4817_), .B(core__abc_21302_new_n2640__bF_buf2), .C(core__abc_21302_new_n2369__bF_buf6), .Y(core__abc_21302_new_n4818_));
OAI21X1 OAI21X1_1127 ( .A(core_v3_reg_63_), .B(core__abc_21302_new_n2369__bF_buf5), .C(reset_n_bF_buf69), .Y(core__abc_21302_new_n4820_));
OAI21X1 OAI21X1_1128 ( .A(core__abc_21302_new_n4827_), .B(core__abc_21302_new_n4826_), .C(core__abc_21302_new_n4830_), .Y(core__abc_21302_new_n4831_));
OAI21X1 OAI21X1_1129 ( .A(core__abc_21302_new_n4770_), .B(core__abc_21302_new_n4773_), .C(core__abc_21302_new_n4833_), .Y(core__abc_21302_new_n4834_));
OAI21X1 OAI21X1_113 ( .A(core_siphash_word_37_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf0), .Y(_abc_19873_new_n1703_));
OAI21X1 OAI21X1_1130 ( .A(core__abc_21302_new_n4840_), .B(core__abc_21302_new_n4845_), .C(core__abc_21302_new_n4844_), .Y(core__abc_21302_new_n4846_));
OAI21X1 OAI21X1_1131 ( .A(core__abc_21302_new_n4711_), .B(core__abc_21302_new_n4710_), .C(core__abc_21302_new_n4847_), .Y(core__abc_21302_new_n4848_));
OAI21X1 OAI21X1_1132 ( .A(core__abc_21302_new_n4856_), .B(core__abc_21302_new_n4855_), .C(core__abc_21302_new_n4859_), .Y(core__abc_21302_new_n4860_));
OAI21X1 OAI21X1_1133 ( .A(core__abc_21302_new_n3705_), .B(core__abc_21302_new_n3706_), .C(core__abc_21302_new_n4864_), .Y(core__abc_21302_new_n4865_));
OAI21X1 OAI21X1_1134 ( .A(core__abc_21302_new_n3667_), .B(core__abc_21302_new_n4869_), .C(core__abc_21302_new_n4873_), .Y(core__abc_21302_new_n4874_));
OAI21X1 OAI21X1_1135 ( .A(core__abc_21302_new_n4854_), .B(core__abc_21302_new_n4857_), .C(core__abc_21302_new_n4876_), .Y(core__abc_21302_new_n4877_));
OAI21X1 OAI21X1_1136 ( .A(core__abc_21302_new_n4875_), .B(core__abc_21302_new_n4867_), .C(core__abc_21302_new_n4877_), .Y(core__abc_21302_new_n4878_));
OAI21X1 OAI21X1_1137 ( .A(core__abc_21302_new_n4881_), .B(core__abc_21302_new_n4879_), .C(core__abc_21302_new_n4846_), .Y(core__abc_21302_new_n4882_));
OAI21X1 OAI21X1_1138 ( .A(core__abc_21302_new_n4823_), .B(core__abc_21302_new_n4828_), .C(core__abc_21302_new_n4884_), .Y(core__abc_21302_new_n4885_));
OAI21X1 OAI21X1_1139 ( .A(core__abc_21302_new_n4838_), .B(core__abc_21302_new_n4882_), .C(core__abc_21302_new_n4886_), .Y(core__abc_21302_new_n4887_));
OAI21X1 OAI21X1_114 ( .A(core_siphash_word_38_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf69), .Y(_abc_19873_new_n1706_));
OAI21X1 OAI21X1_1140 ( .A(core__abc_21302_new_n1454_), .B(core__abc_21302_new_n4546_), .C(core__abc_21302_new_n1467_), .Y(core__abc_21302_new_n4898_));
OAI21X1 OAI21X1_1141 ( .A(core__abc_21302_new_n4902_), .B(core__abc_21302_new_n4903_), .C(core__abc_21302_new_n4901_), .Y(core__abc_21302_new_n4904_));
OAI21X1 OAI21X1_1142 ( .A(core__abc_21302_new_n4547_), .B(core__abc_21302_new_n4546_), .C(core__abc_21302_new_n4906_), .Y(core__abc_21302_new_n4907_));
OAI21X1 OAI21X1_1143 ( .A(core__abc_21302_new_n4547_), .B(core__abc_21302_new_n4546_), .C(core_v1_reg_9_), .Y(core__abc_21302_new_n4912_));
OAI21X1 OAI21X1_1144 ( .A(core__abc_21302_new_n4917_), .B(core__abc_21302_new_n4922_), .C(core__abc_21302_new_n4921_), .Y(core__abc_21302_new_n4923_));
OAI21X1 OAI21X1_1145 ( .A(core__abc_21302_new_n4936_), .B(core__abc_21302_new_n4935_), .C(core__abc_21302_new_n4932_), .Y(core__abc_21302_new_n4937_));
OAI21X1 OAI21X1_1146 ( .A(core__abc_21302_new_n3340_), .B(core__abc_21302_new_n4945_), .C(core__abc_21302_new_n4947_), .Y(core__abc_21302_new_n4948_));
OAI21X1 OAI21X1_1147 ( .A(core__abc_21302_new_n4943_), .B(core__abc_21302_new_n4944_), .C(core__abc_21302_new_n4948_), .Y(core__abc_21302_new_n4949_));
OAI21X1 OAI21X1_1148 ( .A(core__abc_21302_new_n3425_), .B(core__abc_21302_new_n3426_), .C(core__abc_21302_new_n4950_), .Y(core__abc_21302_new_n4952_));
OAI21X1 OAI21X1_1149 ( .A(core__abc_21302_new_n4929_), .B(core__abc_21302_new_n4951_), .C(core__abc_21302_new_n4952_), .Y(core__abc_21302_new_n4953_));
OAI21X1 OAI21X1_115 ( .A(core_siphash_word_39_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf68), .Y(_abc_19873_new_n1709_));
OAI21X1 OAI21X1_1150 ( .A(core__abc_21302_new_n4932_), .B(core__abc_21302_new_n4950_), .C(core__abc_21302_new_n4953_), .Y(core__abc_21302_new_n4954_));
OAI21X1 OAI21X1_1151 ( .A(core__abc_21302_new_n4949_), .B(core__abc_21302_new_n4942_), .C(core__abc_21302_new_n4954_), .Y(core__abc_21302_new_n4955_));
OAI21X1 OAI21X1_1152 ( .A(core__abc_21302_new_n3481_), .B(core__abc_21302_new_n4925_), .C(core__abc_21302_new_n4920_), .Y(core__abc_21302_new_n4957_));
OAI21X1 OAI21X1_1153 ( .A(core__abc_21302_new_n3514_), .B(core__abc_21302_new_n4956_), .C(core__abc_21302_new_n4957_), .Y(core__abc_21302_new_n4958_));
OAI21X1 OAI21X1_1154 ( .A(core__abc_21302_new_n4916_), .B(core__abc_21302_new_n4958_), .C(core__abc_21302_new_n4961_), .Y(core__abc_21302_new_n4962_));
OAI21X1 OAI21X1_1155 ( .A(core__abc_21302_new_n3191_), .B(core__abc_21302_new_n3193_), .C(core__abc_21302_new_n4971_), .Y(core__abc_21302_new_n4973_));
OAI21X1 OAI21X1_1156 ( .A(core__abc_21302_new_n3141_), .B(core__abc_21302_new_n4977_), .C(core__abc_21302_new_n4981_), .Y(core__abc_21302_new_n4982_));
OAI21X1 OAI21X1_1157 ( .A(core__abc_21302_new_n3143_), .B(core__abc_21302_new_n4976_), .C(core__abc_21302_new_n4982_), .Y(core__abc_21302_new_n4983_));
OAI21X1 OAI21X1_1158 ( .A(core__abc_21302_new_n4983_), .B(core__abc_21302_new_n4975_), .C(core__abc_21302_new_n4986_), .Y(core__abc_21302_new_n4987_));
OAI21X1 OAI21X1_1159 ( .A(core__abc_21302_new_n3105_), .B(core__abc_21302_new_n3106_), .C(core__abc_21302_new_n4979_), .Y(core__abc_21302_new_n4991_));
OAI21X1 OAI21X1_116 ( .A(core_siphash_word_40_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf67), .Y(_abc_19873_new_n1711_));
OAI21X1 OAI21X1_1160 ( .A(core__abc_21302_new_n5002_), .B(core__abc_21302_new_n5005_), .C(core__abc_21302_new_n5000_), .Y(core__abc_21302_new_n5006_));
OAI21X1 OAI21X1_1161 ( .A(core__abc_21302_new_n5013_), .B(core__abc_21302_new_n5014_), .C(core__abc_21302_new_n5011_), .Y(core__abc_21302_new_n5015_));
OAI21X1 OAI21X1_1162 ( .A(core__abc_21302_new_n5018_), .B(core__abc_21302_new_n5017_), .C(core__abc_21302_new_n5022_), .Y(core__abc_21302_new_n5023_));
OAI21X1 OAI21X1_1163 ( .A(core__abc_21302_new_n5050_), .B(core__abc_21302_new_n5052_), .C(core__abc_21302_new_n5042_), .Y(core__abc_21302_new_n5053_));
OAI21X1 OAI21X1_1164 ( .A(core__abc_21302_new_n5056_), .B(core__abc_21302_new_n5054_), .C(core__abc_21302_new_n5036_), .Y(core__abc_21302_new_n5057_));
OAI21X1 OAI21X1_1165 ( .A(core__abc_21302_new_n5033_), .B(core__abc_21302_new_n5057_), .C(core__abc_21302_new_n5031_), .Y(core__abc_21302_new_n5058_));
OAI21X1 OAI21X1_1166 ( .A(core__abc_21302_new_n5029_), .B(core__abc_21302_new_n5058_), .C(core__abc_21302_new_n5027_), .Y(core__abc_21302_new_n5059_));
OAI21X1 OAI21X1_1167 ( .A(core__abc_21302_new_n4987_), .B(core__abc_21302_new_n5064_), .C(core__abc_21302_new_n5070_), .Y(core__abc_21302_new_n5071_));
OAI21X1 OAI21X1_1168 ( .A(core__abc_21302_new_n4894_), .B(core__abc_21302_new_n5072_), .C(core__abc_21302_new_n4888_), .Y(core__abc_21302_new_n5073_));
OAI21X1 OAI21X1_1169 ( .A(core__abc_21302_new_n2364__bF_buf4), .B(core__abc_21302_new_n5081_), .C(core__abc_21302_new_n5080_), .Y(core__abc_21302_new_n5082_));
OAI21X1 OAI21X1_117 ( .A(core_siphash_word_41_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf66), .Y(_abc_19873_new_n1713_));
OAI21X1 OAI21X1_1170 ( .A(core__abc_21302_new_n4822_), .B(core__abc_21302_new_n5082_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n5083_));
OAI21X1 OAI21X1_1171 ( .A(core__abc_21302_new_n2138_), .B(core__abc_21302_new_n2633_), .C(core__abc_21302_new_n2640__bF_buf0), .Y(core__abc_21302_new_n5084_));
OAI21X1 OAI21X1_1172 ( .A(core__abc_21302_new_n2365__bF_buf3), .B(core__abc_21302_new_n5084_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n5085_));
OAI21X1 OAI21X1_1173 ( .A(core__abc_21302_new_n5078_), .B(core__abc_21302_new_n5095_), .C(core__abc_21302_new_n5075_), .Y(core__abc_21302_new_n5096_));
OAI21X1 OAI21X1_1174 ( .A(core_v2_reg_1_), .B(core__abc_21302_new_n2364__bF_buf3), .C(core__abc_21302_new_n5099_), .Y(core__abc_21302_new_n5100_));
OAI21X1 OAI21X1_1175 ( .A(core__abc_21302_new_n5100_), .B(core__abc_21302_new_n5098_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n5101_));
OAI21X1 OAI21X1_1176 ( .A(core__abc_21302_new_n3956_), .B(core__abc_21302_new_n5107_), .C(core__abc_21302_new_n5075_), .Y(core__abc_21302_new_n5108_));
OAI21X1 OAI21X1_1177 ( .A(core__abc_21302_new_n3954_), .B(core__abc_21302_new_n5089_), .C(core__abc_21302_new_n5108_), .Y(core__abc_21302_new_n5109_));
OAI21X1 OAI21X1_1178 ( .A(core__abc_21302_new_n2689_), .B(core__abc_21302_new_n2688_), .C(core__abc_21302_new_n5113_), .Y(core__abc_21302_new_n5114_));
OAI21X1 OAI21X1_1179 ( .A(core__abc_21302_new_n5115_), .B(core__abc_21302_new_n5116_), .C(core__abc_21302_new_n5112_), .Y(core__abc_21302_new_n5117_));
OAI21X1 OAI21X1_118 ( .A(core_siphash_word_42_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf65), .Y(_abc_19873_new_n1715_));
OAI21X1 OAI21X1_1180 ( .A(core__abc_21302_new_n5110_), .B(core__abc_21302_new_n5106_), .C(core__abc_21302_new_n5120_), .Y(core__abc_21302_new_n5121_));
OAI21X1 OAI21X1_1181 ( .A(core__abc_21302_new_n5105_), .B(core__abc_21302_new_n5095_), .C(core__abc_21302_new_n5109_), .Y(core__abc_21302_new_n5122_));
OAI21X1 OAI21X1_1182 ( .A(core_v2_reg_2_), .B(core__abc_21302_new_n2364__bF_buf2), .C(core__abc_21302_new_n5126_), .Y(core__abc_21302_new_n5127_));
OAI21X1 OAI21X1_1183 ( .A(core__abc_21302_new_n5127_), .B(core__abc_21302_new_n5125_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n5128_));
OAI21X1 OAI21X1_1184 ( .A(core__abc_21302_new_n2741_), .B(core__abc_21302_new_n5104__bF_buf7), .C(core__abc_21302_new_n5128_), .Y(core__abc_21302_new_n5129_));
OAI21X1 OAI21X1_1185 ( .A(core__abc_21302_new_n5112_), .B(core__abc_21302_new_n5133_), .C(core__abc_21302_new_n5121_), .Y(core__abc_21302_new_n5134_));
OAI21X1 OAI21X1_1186 ( .A(core__abc_21302_new_n5141_), .B(core__abc_21302_new_n5142_), .C(core__abc_21302_new_n5140_), .Y(core__abc_21302_new_n5143_));
OAI21X1 OAI21X1_1187 ( .A(core_v2_reg_3_), .B(core__abc_21302_new_n2364__bF_buf1), .C(core__abc_21302_new_n5146_), .Y(core__abc_21302_new_n5147_));
OAI21X1 OAI21X1_1188 ( .A(core__abc_21302_new_n5132_), .B(core__abc_21302_new_n5147_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n5148_));
OAI21X1 OAI21X1_1189 ( .A(core__abc_21302_new_n5112_), .B(core__abc_21302_new_n5133_), .C(core__abc_21302_new_n5139_), .Y(core__abc_21302_new_n5156_));
OAI21X1 OAI21X1_119 ( .A(core_siphash_word_43_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf64), .Y(_abc_19873_new_n1718_));
OAI21X1 OAI21X1_1190 ( .A(core__abc_21302_new_n5135_), .B(core__abc_21302_new_n5155_), .C(core__abc_21302_new_n5156_), .Y(core__abc_21302_new_n5157_));
OAI21X1 OAI21X1_1191 ( .A(core__abc_21302_new_n5109_), .B(core__abc_21302_new_n5158_), .C(core__abc_21302_new_n5157_), .Y(core__abc_21302_new_n5159_));
OAI21X1 OAI21X1_1192 ( .A(core__abc_21302_new_n5165_), .B(core__abc_21302_new_n5095_), .C(core__abc_21302_new_n5160_), .Y(core__abc_21302_new_n5166_));
OAI21X1 OAI21X1_1193 ( .A(core__abc_21302_new_n2673__bF_buf3), .B(core__abc_21302_new_n5168_), .C(core__abc_21302_new_n5170_), .Y(core__abc_21302_new_n5171_));
OAI21X1 OAI21X1_1194 ( .A(core__abc_21302_new_n5154_), .B(core__abc_21302_new_n5174_), .C(core__abc_21302_new_n5153_), .Y(core__abc_21302_new_n5175_));
OAI21X1 OAI21X1_1195 ( .A(core__abc_21302_new_n5183_), .B(core__abc_21302_new_n5182_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n5184_));
OAI21X1 OAI21X1_1196 ( .A(core__abc_21302_new_n5153_), .B(core__abc_21302_new_n5180_), .C(core__abc_21302_new_n5179_), .Y(core__abc_21302_new_n5193_));
OAI21X1 OAI21X1_1197 ( .A(core_v2_reg_6_), .B(core__abc_21302_new_n2364__bF_buf5), .C(core__abc_21302_new_n5200_), .Y(core__abc_21302_new_n5201_));
OAI21X1 OAI21X1_1198 ( .A(core__abc_21302_new_n5187_), .B(core__abc_21302_new_n5201_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n5202_));
OAI21X1 OAI21X1_1199 ( .A(core__abc_21302_new_n5209_), .B(core__abc_21302_new_n5211_), .C(core__abc_21302_new_n5208_), .Y(core__abc_21302_new_n5212_));
OAI21X1 OAI21X1_12 ( .A(_abc_19873_new_n1052_), .B(_abc_19873_new_n913__bF_buf3), .C(_abc_19873_new_n1053_), .Y(_abc_19873_new_n1054_));
OAI21X1 OAI21X1_120 ( .A(core_siphash_word_44_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf63), .Y(_abc_19873_new_n1721_));
OAI21X1 OAI21X1_1200 ( .A(core__abc_21302_new_n5205_), .B(core__abc_21302_new_n5196_), .C(core__abc_21302_new_n5218_), .Y(core__abc_21302_new_n5219_));
OAI21X1 OAI21X1_1201 ( .A(core__abc_21302_new_n5222_), .B(core__abc_21302_new_n5220_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n5223_));
OAI21X1 OAI21X1_1202 ( .A(core__abc_21302_new_n5209_), .B(core__abc_21302_new_n5211_), .C(core__abc_21302_new_n5207_), .Y(core__abc_21302_new_n5230_));
OAI21X1 OAI21X1_1203 ( .A(core__abc_21302_new_n5207_), .B(core__abc_21302_new_n5231_), .C(core__abc_21302_new_n5191_), .Y(core__abc_21302_new_n5232_));
OAI21X1 OAI21X1_1204 ( .A(core_v2_reg_8_), .B(core__abc_21302_new_n5104__bF_buf5), .C(reset_n_bF_buf67), .Y(core__abc_21302_new_n5246_));
OAI21X1 OAI21X1_1205 ( .A(core__abc_21302_new_n5241_), .B(core__abc_21302_new_n5235_), .C(core__abc_21302_new_n5240_), .Y(core__abc_21302_new_n5255_));
OAI21X1 OAI21X1_1206 ( .A(core_key_9_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n5257_), .Y(core__abc_21302_new_n5258_));
OAI21X1 OAI21X1_1207 ( .A(core_v2_reg_9_), .B(core__abc_21302_new_n5104__bF_buf4), .C(reset_n_bF_buf66), .Y(core__abc_21302_new_n5260_));
OAI21X1 OAI21X1_1208 ( .A(core__abc_21302_new_n3013_), .B(core__abc_21302_new_n3014_), .C(core__abc_21302_new_n5268_), .Y(core__abc_21302_new_n5269_));
OAI21X1 OAI21X1_1209 ( .A(core__abc_21302_new_n2626_), .B(core__abc_21302_new_n4223_), .C(core__abc_21302_new_n5271_), .Y(core__abc_21302_new_n5273_));
OAI21X1 OAI21X1_121 ( .A(core_siphash_word_45_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf62), .Y(_abc_19873_new_n1724_));
OAI21X1 OAI21X1_1210 ( .A(core__abc_21302_new_n5266_), .B(core__abc_21302_new_n5263_), .C(core__abc_21302_new_n5274_), .Y(core__abc_21302_new_n5275_));
OAI21X1 OAI21X1_1211 ( .A(core__abc_21302_new_n5262_), .B(core__abc_21302_new_n5235_), .C(core__abc_21302_new_n5265_), .Y(core__abc_21302_new_n5276_));
OAI21X1 OAI21X1_1212 ( .A(core_v2_reg_10_), .B(core__abc_21302_new_n5104__bF_buf1), .C(reset_n_bF_buf65), .Y(core__abc_21302_new_n5283_));
OAI21X1 OAI21X1_1213 ( .A(core__abc_21302_new_n5267_), .B(core__abc_21302_new_n5271_), .C(core__abc_21302_new_n5275_), .Y(core__abc_21302_new_n5285_));
OAI21X1 OAI21X1_1214 ( .A(core__abc_21302_new_n5286_), .B(core__abc_21302_new_n5291_), .C(core__abc_21302_new_n5290_), .Y(core__abc_21302_new_n5292_));
OAI21X1 OAI21X1_1215 ( .A(core__abc_21302_new_n2673__bF_buf0), .B(core__abc_21302_new_n5296_), .C(core__abc_21302_new_n5299_), .Y(core__abc_21302_new_n5300_));
OAI21X1 OAI21X1_1216 ( .A(core_v2_reg_11_), .B(core__abc_21302_new_n5104__bF_buf0), .C(core__abc_21302_new_n5300_), .Y(core__abc_21302_new_n5301_));
OAI21X1 OAI21X1_1217 ( .A(core__abc_21302_new_n5265_), .B(core__abc_21302_new_n5303_), .C(core__abc_21302_new_n5306_), .Y(core__abc_21302_new_n5307_));
OAI21X1 OAI21X1_1218 ( .A(core__abc_21302_new_n5309_), .B(core__abc_21302_new_n5235_), .C(core__abc_21302_new_n5308_), .Y(core__abc_21302_new_n5310_));
OAI21X1 OAI21X1_1219 ( .A(core_key_12_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n5317_), .Y(core__abc_21302_new_n5318_));
OAI21X1 OAI21X1_122 ( .A(core_siphash_word_46_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf61), .Y(_abc_19873_new_n1727_));
OAI21X1 OAI21X1_1220 ( .A(core_v2_reg_12_), .B(core__abc_21302_new_n5104__bF_buf7), .C(reset_n_bF_buf64), .Y(core__abc_21302_new_n5320_));
OAI21X1 OAI21X1_1221 ( .A(core__abc_21302_new_n2668_), .B(core__abc_21302_new_n5312_), .C(core__abc_21302_new_n5323_), .Y(core__abc_21302_new_n5324_));
OAI21X1 OAI21X1_1222 ( .A(core_v2_reg_13_), .B(core__abc_21302_new_n5104__bF_buf5), .C(reset_n_bF_buf63), .Y(core__abc_21302_new_n5340_));
OAI21X1 OAI21X1_1223 ( .A(core__abc_21302_new_n3185_), .B(core__abc_21302_new_n3182_), .C(core__abc_21302_new_n1576_), .Y(core__abc_21302_new_n5349_));
OAI21X1 OAI21X1_1224 ( .A(core__abc_21302_new_n2724_), .B(core__abc_21302_new_n2727_), .C(core__abc_21302_new_n5351_), .Y(core__abc_21302_new_n5352_));
OAI21X1 OAI21X1_1225 ( .A(core__abc_21302_new_n5345_), .B(core__abc_21302_new_n5348_), .C(core__abc_21302_new_n5356_), .Y(core__abc_21302_new_n5357_));
OAI21X1 OAI21X1_1226 ( .A(core__abc_21302_new_n2673__bF_buf11), .B(core__abc_21302_new_n5362_), .C(core__abc_21302_new_n5364_), .Y(core__abc_21302_new_n5365_));
OAI21X1 OAI21X1_1227 ( .A(core_v2_reg_14_), .B(core__abc_21302_new_n5104__bF_buf4), .C(core__abc_21302_new_n5365_), .Y(core__abc_21302_new_n5366_));
OAI21X1 OAI21X1_1228 ( .A(core__abc_21302_new_n5370_), .B(core__abc_21302_new_n5369_), .C(core__abc_21302_new_n5368_), .Y(core__abc_21302_new_n5371_));
OAI21X1 OAI21X1_1229 ( .A(core__abc_21302_new_n5378_), .B(core__abc_21302_new_n5379_), .C(core__abc_21302_new_n5375_), .Y(core__abc_21302_new_n5380_));
OAI21X1 OAI21X1_123 ( .A(core_siphash_word_47_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf60), .Y(_abc_19873_new_n1729_));
OAI21X1 OAI21X1_1230 ( .A(core__abc_21302_new_n2673__bF_buf10), .B(core__abc_21302_new_n5381_), .C(core__abc_21302_new_n5384_), .Y(core__abc_21302_new_n5385_));
OAI21X1 OAI21X1_1231 ( .A(core_v2_reg_15_), .B(core__abc_21302_new_n5104__bF_buf3), .C(core__abc_21302_new_n5385_), .Y(core__abc_21302_new_n5386_));
OAI21X1 OAI21X1_1232 ( .A(core__abc_21302_new_n5370_), .B(core__abc_21302_new_n5369_), .C(core__abc_21302_new_n5372_), .Y(core__abc_21302_new_n5393_));
OAI21X1 OAI21X1_1233 ( .A(core__abc_21302_new_n5402_), .B(core__abc_21302_new_n5095_), .C(core__abc_21302_new_n5398_), .Y(core__abc_21302_new_n5403_));
OAI21X1 OAI21X1_1234 ( .A(core__abc_21302_new_n2826_), .B(core__abc_21302_new_n2828_), .C(core__abc_21302_new_n5404_), .Y(core__abc_21302_new_n5407_));
OAI21X1 OAI21X1_1235 ( .A(core_key_16_), .B(core__abc_21302_new_n2640__bF_buf1), .C(core__abc_21302_new_n5410_), .Y(core__abc_21302_new_n5411_));
OAI21X1 OAI21X1_1236 ( .A(core_v2_reg_16_), .B(core__abc_21302_new_n5104__bF_buf2), .C(reset_n_bF_buf62), .Y(core__abc_21302_new_n5413_));
OAI21X1 OAI21X1_1237 ( .A(core__abc_21302_new_n5418_), .B(core__abc_21302_new_n5417_), .C(core__abc_21302_new_n5419_), .Y(core__abc_21302_new_n5420_));
OAI21X1 OAI21X1_1238 ( .A(core__abc_21302_new_n1397_), .B(core__abc_21302_new_n2364__bF_buf5), .C(core__abc_21302_new_n5429_), .Y(core__abc_21302_new_n5430_));
OAI21X1 OAI21X1_1239 ( .A(core_v2_reg_17_), .B(core__abc_21302_new_n5104__bF_buf0), .C(reset_n_bF_buf61), .Y(core__abc_21302_new_n5432_));
OAI21X1 OAI21X1_124 ( .A(core_siphash_word_48_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf59), .Y(_abc_19873_new_n1732_));
OAI21X1 OAI21X1_1240 ( .A(core__abc_21302_new_n2901_), .B(core__abc_21302_new_n2902_), .C(core__abc_21302_new_n5435_), .Y(core__abc_21302_new_n5438_));
OAI21X1 OAI21X1_1241 ( .A(core__abc_21302_new_n2868_), .B(core__abc_21302_new_n5423_), .C(core__abc_21302_new_n5441_), .Y(core__abc_21302_new_n5442_));
OAI21X1 OAI21X1_1242 ( .A(core__abc_21302_new_n5418_), .B(core__abc_21302_new_n5417_), .C(core__abc_21302_new_n5443_), .Y(core__abc_21302_new_n5444_));
OAI21X1 OAI21X1_1243 ( .A(core_v2_reg_18_), .B(core__abc_21302_new_n5104__bF_buf7), .C(reset_n_bF_buf60), .Y(core__abc_21302_new_n5452_));
OAI21X1 OAI21X1_1244 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n5459_), .C(core__abc_21302_new_n5462_), .Y(core__abc_21302_new_n5463_));
OAI21X1 OAI21X1_1245 ( .A(core_v2_reg_19_), .B(core__abc_21302_new_n5104__bF_buf6), .C(core__abc_21302_new_n5463_), .Y(core__abc_21302_new_n5464_));
OAI21X1 OAI21X1_1246 ( .A(core__abc_21302_new_n2953_), .B(core__abc_21302_new_n5466_), .C(core__abc_21302_new_n5437_), .Y(core__abc_21302_new_n5467_));
OAI21X1 OAI21X1_1247 ( .A(core__abc_21302_new_n2952_), .B(core__abc_21302_new_n5455_), .C(core__abc_21302_new_n5467_), .Y(core__abc_21302_new_n5468_));
OAI21X1 OAI21X1_1248 ( .A(core__abc_21302_new_n5442_), .B(core__abc_21302_new_n5469_), .C(core__abc_21302_new_n5468_), .Y(core__abc_21302_new_n5470_));
OAI21X1 OAI21X1_1249 ( .A(core__abc_21302_new_n1433_), .B(core__abc_21302_new_n2364__bF_buf2), .C(core__abc_21302_new_n5487_), .Y(core__abc_21302_new_n5488_));
OAI21X1 OAI21X1_125 ( .A(core_siphash_word_49_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf58), .Y(_abc_19873_new_n1735_));
OAI21X1 OAI21X1_1250 ( .A(core_v2_reg_20_), .B(core__abc_21302_new_n5104__bF_buf5), .C(reset_n_bF_buf59), .Y(core__abc_21302_new_n5490_));
OAI21X1 OAI21X1_1251 ( .A(core__abc_21302_new_n5470_), .B(core__abc_21302_new_n5476_), .C(core__abc_21302_new_n5484_), .Y(core__abc_21302_new_n5492_));
OAI21X1 OAI21X1_1252 ( .A(core__abc_21302_new_n5481_), .B(core__abc_21302_new_n5498_), .C(core__abc_21302_new_n5499_), .Y(core__abc_21302_new_n5500_));
OAI21X1 OAI21X1_1253 ( .A(core__abc_21302_new_n2673__bF_buf8), .B(core__abc_21302_new_n5501_), .C(core__abc_21302_new_n5503_), .Y(core__abc_21302_new_n5504_));
OAI21X1 OAI21X1_1254 ( .A(core_v2_reg_21_), .B(core__abc_21302_new_n5104__bF_buf4), .C(core__abc_21302_new_n5504_), .Y(core__abc_21302_new_n5505_));
OAI21X1 OAI21X1_1255 ( .A(core__abc_21302_new_n3068_), .B(core__abc_21302_new_n3069_), .C(core__abc_21302_new_n5511_), .Y(core__abc_21302_new_n5512_));
OAI21X1 OAI21X1_1256 ( .A(core__abc_21302_new_n5470_), .B(core__abc_21302_new_n5476_), .C(core__abc_21302_new_n5515_), .Y(core__abc_21302_new_n5516_));
OAI21X1 OAI21X1_1257 ( .A(core__abc_21302_new_n5482_), .B(core__abc_21302_new_n5496_), .C(core__abc_21302_new_n5494_), .Y(core__abc_21302_new_n5517_));
OAI21X1 OAI21X1_1258 ( .A(core__abc_21302_new_n2673__bF_buf7), .B(core__abc_21302_new_n5522_), .C(core__abc_21302_new_n5524_), .Y(core__abc_21302_new_n5525_));
OAI21X1 OAI21X1_1259 ( .A(core_v2_reg_22_), .B(core__abc_21302_new_n5104__bF_buf3), .C(core__abc_21302_new_n5525_), .Y(core__abc_21302_new_n5526_));
OAI21X1 OAI21X1_126 ( .A(core_siphash_word_50_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf57), .Y(_abc_19873_new_n1738_));
OAI21X1 OAI21X1_1260 ( .A(core__abc_21302_new_n5536_), .B(core__abc_21302_new_n5519_), .C(core__abc_21302_new_n5537_), .Y(core__abc_21302_new_n5538_));
OAI21X1 OAI21X1_1261 ( .A(core_v2_reg_23_), .B(core__abc_21302_new_n5104__bF_buf2), .C(reset_n_bF_buf58), .Y(core__abc_21302_new_n5543_));
OAI21X1 OAI21X1_1262 ( .A(core__abc_21302_new_n5518_), .B(core__abc_21302_new_n5545_), .C(core__abc_21302_new_n5549_), .Y(core__abc_21302_new_n5550_));
OAI21X1 OAI21X1_1263 ( .A(core__abc_21302_new_n5551_), .B(core__abc_21302_new_n5553_), .C(core__abc_21302_new_n5559_), .Y(core__abc_21302_new_n5560_));
OAI21X1 OAI21X1_1264 ( .A(core__abc_21302_new_n1476_), .B(core__abc_21302_new_n2364__bF_buf4), .C(core__abc_21302_new_n5564_), .Y(core__abc_21302_new_n5565_));
OAI21X1 OAI21X1_1265 ( .A(core__abc_21302_new_n2673__bF_buf6), .B(core__abc_21302_new_n5563_), .C(core__abc_21302_new_n5566_), .Y(core__abc_21302_new_n5567_));
OAI21X1 OAI21X1_1266 ( .A(core_v2_reg_24_), .B(core__abc_21302_new_n5104__bF_buf1), .C(core__abc_21302_new_n5567_), .Y(core__abc_21302_new_n5568_));
OAI21X1 OAI21X1_1267 ( .A(core__abc_21302_new_n5573_), .B(core__abc_21302_new_n5574_), .C(core__abc_21302_new_n5571_), .Y(core__abc_21302_new_n5575_));
OAI21X1 OAI21X1_1268 ( .A(core__abc_21302_new_n5555_), .B(core__abc_21302_new_n5570_), .C(core__abc_21302_new_n5576_), .Y(core__abc_21302_new_n5577_));
OAI21X1 OAI21X1_1269 ( .A(core_v2_reg_25_), .B(core__abc_21302_new_n5104__bF_buf0), .C(reset_n_bF_buf57), .Y(core__abc_21302_new_n5581_));
OAI21X1 OAI21X1_127 ( .A(core_siphash_word_51_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf56), .Y(_abc_19873_new_n1741_));
OAI21X1 OAI21X1_1270 ( .A(core__abc_21302_new_n3249_), .B(core__abc_21302_new_n3250_), .C(core__abc_21302_new_n5584_), .Y(core__abc_21302_new_n5586_));
OAI21X1 OAI21X1_1271 ( .A(core__abc_21302_new_n5551_), .B(core__abc_21302_new_n5553_), .C(core__abc_21302_new_n5589_), .Y(core__abc_21302_new_n5590_));
OAI21X1 OAI21X1_1272 ( .A(core__abc_21302_new_n2673__bF_buf5), .B(core__abc_21302_new_n5595_), .C(core__abc_21302_new_n5597_), .Y(core__abc_21302_new_n5598_));
OAI21X1 OAI21X1_1273 ( .A(core_v2_reg_26_), .B(core__abc_21302_new_n5104__bF_buf7), .C(core__abc_21302_new_n5598_), .Y(core__abc_21302_new_n5599_));
OAI21X1 OAI21X1_1274 ( .A(core__abc_21302_new_n3319_), .B(core__abc_21302_new_n3318_), .C(core__abc_21302_new_n5605_), .Y(core__abc_21302_new_n5606_));
OAI21X1 OAI21X1_1275 ( .A(core__abc_21302_new_n5609_), .B(core__abc_21302_new_n5592_), .C(core__abc_21302_new_n5610_), .Y(core__abc_21302_new_n5611_));
OAI21X1 OAI21X1_1276 ( .A(core_v2_reg_27_), .B(core__abc_21302_new_n5104__bF_buf6), .C(reset_n_bF_buf56), .Y(core__abc_21302_new_n5615_));
OAI21X1 OAI21X1_1277 ( .A(core__abc_21302_new_n5551_), .B(core__abc_21302_new_n5553_), .C(core__abc_21302_new_n5619_), .Y(core__abc_21302_new_n5620_));
OAI21X1 OAI21X1_1278 ( .A(core__abc_21302_new_n5585_), .B(core__abc_21302_new_n5607_), .C(core__abc_21302_new_n5604_), .Y(core__abc_21302_new_n5623_));
OAI21X1 OAI21X1_1279 ( .A(core__abc_21302_new_n3355_), .B(core__abc_21302_new_n3354_), .C(core__abc_21302_new_n5625_), .Y(core__abc_21302_new_n5628_));
OAI21X1 OAI21X1_128 ( .A(core_siphash_word_52_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf55), .Y(_abc_19873_new_n1744_));
OAI21X1 OAI21X1_1280 ( .A(core__abc_21302_new_n5418_), .B(core__abc_21302_new_n5417_), .C(core__abc_21302_new_n5632_), .Y(core__abc_21302_new_n5633_));
OAI21X1 OAI21X1_1281 ( .A(core__abc_21302_new_n5635_), .B(core__abc_21302_new_n5634_), .C(core__abc_21302_new_n5636_), .Y(core__abc_21302_new_n5637_));
OAI21X1 OAI21X1_1282 ( .A(core__abc_21302_new_n1523_), .B(core__abc_21302_new_n2364__bF_buf0), .C(core__abc_21302_new_n5639_), .Y(core__abc_21302_new_n5640_));
OAI21X1 OAI21X1_1283 ( .A(core__abc_21302_new_n2673__bF_buf4), .B(core__abc_21302_new_n5638_), .C(core__abc_21302_new_n5641_), .Y(core__abc_21302_new_n5642_));
OAI21X1 OAI21X1_1284 ( .A(core_v2_reg_28_), .B(core__abc_21302_new_n5104__bF_buf5), .C(core__abc_21302_new_n5642_), .Y(core__abc_21302_new_n5643_));
OAI21X1 OAI21X1_1285 ( .A(core__abc_21302_new_n5627_), .B(core__abc_21302_new_n5650_), .C(core__abc_21302_new_n5656_), .Y(core__abc_21302_new_n5657_));
OAI21X1 OAI21X1_1286 ( .A(core__abc_21302_new_n2673__bF_buf3), .B(core__abc_21302_new_n5657_), .C(core__abc_21302_new_n5659_), .Y(core__abc_21302_new_n5660_));
OAI21X1 OAI21X1_1287 ( .A(core_v2_reg_29_), .B(core__abc_21302_new_n5104__bF_buf4), .C(core__abc_21302_new_n5660_), .Y(core__abc_21302_new_n5661_));
OAI21X1 OAI21X1_1288 ( .A(core__abc_21302_new_n5635_), .B(core__abc_21302_new_n5634_), .C(core__abc_21302_new_n5663_), .Y(core__abc_21302_new_n5664_));
OAI21X1 OAI21X1_1289 ( .A(core__abc_21302_new_n5627_), .B(core__abc_21302_new_n5650_), .C(core__abc_21302_new_n5648_), .Y(core__abc_21302_new_n5665_));
OAI21X1 OAI21X1_129 ( .A(core_siphash_word_53_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf54), .Y(_abc_19873_new_n1747_));
OAI21X1 OAI21X1_1290 ( .A(core__abc_21302_new_n5665_), .B(core__abc_21302_new_n5655_), .C(core__abc_21302_new_n5673_), .Y(core__abc_21302_new_n5676_));
OAI21X1 OAI21X1_1291 ( .A(core__abc_21302_new_n2673__bF_buf2), .B(core__abc_21302_new_n5677_), .C(core__abc_21302_new_n5679_), .Y(core__abc_21302_new_n5680_));
OAI21X1 OAI21X1_1292 ( .A(core_v2_reg_30_), .B(core__abc_21302_new_n5104__bF_buf3), .C(core__abc_21302_new_n5680_), .Y(core__abc_21302_new_n5681_));
OAI21X1 OAI21X1_1293 ( .A(core__abc_21302_new_n5683_), .B(core__abc_21302_new_n5691_), .C(core__abc_21302_new_n5688_), .Y(core__abc_21302_new_n5692_));
OAI21X1 OAI21X1_1294 ( .A(core_v2_reg_31_), .B(core__abc_21302_new_n5104__bF_buf2), .C(reset_n_bF_buf55), .Y(core__abc_21302_new_n5697_));
OAI21X1 OAI21X1_1295 ( .A(core__abc_21302_new_n5699_), .B(core__abc_21302_new_n5702_), .C(core__abc_21302_new_n5104__bF_buf1), .Y(core__abc_21302_new_n5703_));
OAI21X1 OAI21X1_1296 ( .A(core__abc_21302_new_n2365__bF_buf1), .B(core__abc_21302_new_n5085__bF_buf2), .C(core_v2_reg_32_), .Y(core__abc_21302_new_n5704_));
OAI21X1 OAI21X1_1297 ( .A(core__abc_21302_new_n2365__bF_buf0), .B(core__abc_21302_new_n5085__bF_buf1), .C(core_v2_reg_33_), .Y(core__abc_21302_new_n5706_));
OAI21X1 OAI21X1_1298 ( .A(core__abc_21302_new_n5707_), .B(core__abc_21302_new_n5711_), .C(core__abc_21302_new_n5104__bF_buf0), .Y(core__abc_21302_new_n5712_));
OAI21X1 OAI21X1_1299 ( .A(core_v2_reg_34_), .B(core__abc_21302_new_n5104__bF_buf7), .C(reset_n_bF_buf54), .Y(core__abc_21302_new_n5718_));
OAI21X1 OAI21X1_13 ( .A(_abc_19873_new_n1055_), .B(_abc_19873_new_n896__bF_buf1), .C(_abc_19873_new_n982_), .Y(_abc_19873_new_n1056_));
OAI21X1 OAI21X1_130 ( .A(core_siphash_word_54_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf53), .Y(_abc_19873_new_n1750_));
OAI21X1 OAI21X1_1300 ( .A(core_v2_reg_35_), .B(core__abc_21302_new_n5104__bF_buf6), .C(reset_n_bF_buf53), .Y(core__abc_21302_new_n5726_));
OAI21X1 OAI21X1_1301 ( .A(core__abc_21302_new_n5728_), .B(core__abc_21302_new_n2364__bF_buf0), .C(core__abc_21302_new_n5732_), .Y(core__abc_21302_new_n5733_));
OAI21X1 OAI21X1_1302 ( .A(core__abc_21302_new_n5734_), .B(core__abc_21302_new_n5731_), .C(reset_n_bF_buf52), .Y(core__abc_21302_new_n5735_));
OAI21X1 OAI21X1_1303 ( .A(core__abc_21302_new_n2673__bF_buf11), .B(core__abc_21302_new_n5739_), .C(core__abc_21302_new_n5740_), .Y(core__abc_21302_new_n5741_));
OAI21X1 OAI21X1_1304 ( .A(core__abc_21302_new_n5737_), .B(core__abc_21302_new_n5741_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n5742_));
OAI21X1 OAI21X1_1305 ( .A(core_v2_reg_37_), .B(core__abc_21302_new_n5104__bF_buf5), .C(reset_n_bF_buf51), .Y(core__abc_21302_new_n5743_));
OAI21X1 OAI21X1_1306 ( .A(core_key_38_), .B(core__abc_21302_new_n2640__bF_buf9), .C(core__abc_21302_new_n5747_), .Y(core__abc_21302_new_n5748_));
OAI21X1 OAI21X1_1307 ( .A(core_v2_reg_38_), .B(core__abc_21302_new_n5104__bF_buf3), .C(reset_n_bF_buf50), .Y(core__abc_21302_new_n5750_));
OAI21X1 OAI21X1_1308 ( .A(core__abc_21302_new_n5754_), .B(core__abc_21302_new_n5058_), .C(core__abc_21302_new_n5753_), .Y(core__abc_21302_new_n5755_));
OAI21X1 OAI21X1_1309 ( .A(core__abc_21302_new_n5758_), .B(core__abc_21302_new_n2640__bF_buf8), .C(core__abc_21302_new_n5759_), .Y(core__abc_21302_new_n5760_));
OAI21X1 OAI21X1_131 ( .A(core_siphash_word_55_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf52), .Y(_abc_19873_new_n1752_));
OAI21X1 OAI21X1_1310 ( .A(core_v2_reg_39_), .B(core__abc_21302_new_n5104__bF_buf2), .C(reset_n_bF_buf49), .Y(core__abc_21302_new_n5762_));
OAI21X1 OAI21X1_1311 ( .A(core__abc_21302_new_n5766_), .B(core__abc_21302_new_n2364__bF_buf5), .C(core__abc_21302_new_n5767_), .Y(core__abc_21302_new_n5768_));
OAI21X1 OAI21X1_1312 ( .A(core_v2_reg_40_), .B(core__abc_21302_new_n5104__bF_buf1), .C(reset_n_bF_buf48), .Y(core__abc_21302_new_n5770_));
OAI21X1 OAI21X1_1313 ( .A(core__abc_21302_new_n2673__bF_buf10), .B(core__abc_21302_new_n5776_), .C(core__abc_21302_new_n5777_), .Y(core__abc_21302_new_n5778_));
OAI21X1 OAI21X1_1314 ( .A(core__abc_21302_new_n5772_), .B(core__abc_21302_new_n5778_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n5779_));
OAI21X1 OAI21X1_1315 ( .A(core_v2_reg_41_), .B(core__abc_21302_new_n5104__bF_buf0), .C(reset_n_bF_buf47), .Y(core__abc_21302_new_n5780_));
OAI21X1 OAI21X1_1316 ( .A(core_key_42_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n5785_), .Y(core__abc_21302_new_n5786_));
OAI21X1 OAI21X1_1317 ( .A(core_v2_reg_42_), .B(core__abc_21302_new_n5104__bF_buf6), .C(reset_n_bF_buf46), .Y(core__abc_21302_new_n5788_));
OAI21X1 OAI21X1_1318 ( .A(core__abc_21302_new_n5008_), .B(core__abc_21302_new_n5782_), .C(core__abc_21302_new_n5002_), .Y(core__abc_21302_new_n5790_));
OAI21X1 OAI21X1_1319 ( .A(core_v2_reg_43_), .B(core__abc_21302_new_n5104__bF_buf4), .C(reset_n_bF_buf45), .Y(core__abc_21302_new_n5795_));
OAI21X1 OAI21X1_132 ( .A(core_siphash_word_56_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf51), .Y(_abc_19873_new_n1755_));
OAI21X1 OAI21X1_1320 ( .A(core__abc_21302_new_n5799_), .B(core__abc_21302_new_n5782_), .C(core__abc_21302_new_n5798_), .Y(core__abc_21302_new_n5800_));
OAI21X1 OAI21X1_1321 ( .A(core__abc_21302_new_n2702_), .B(core__abc_21302_new_n2364__bF_buf4), .C(core__abc_21302_new_n5806_), .Y(core__abc_21302_new_n5807_));
OAI21X1 OAI21X1_1322 ( .A(core_v2_reg_44_), .B(core__abc_21302_new_n5104__bF_buf3), .C(reset_n_bF_buf44), .Y(core__abc_21302_new_n5809_));
OAI21X1 OAI21X1_1323 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n5813_), .C(core__abc_21302_new_n5814_), .Y(core__abc_21302_new_n5815_));
OAI21X1 OAI21X1_1324 ( .A(core__abc_21302_new_n5811_), .B(core__abc_21302_new_n5815_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n5816_));
OAI21X1 OAI21X1_1325 ( .A(core_v2_reg_45_), .B(core__abc_21302_new_n5104__bF_buf2), .C(reset_n_bF_buf43), .Y(core__abc_21302_new_n5817_));
OAI21X1 OAI21X1_1326 ( .A(core__abc_21302_new_n4982_), .B(core__abc_21302_new_n5802_), .C(core__abc_21302_new_n4988_), .Y(core__abc_21302_new_n5819_));
OAI21X1 OAI21X1_1327 ( .A(core_key_46_), .B(core__abc_21302_new_n2640__bF_buf3), .C(core__abc_21302_new_n5822_), .Y(core__abc_21302_new_n5823_));
OAI21X1 OAI21X1_1328 ( .A(core_v2_reg_46_), .B(core__abc_21302_new_n5104__bF_buf0), .C(reset_n_bF_buf42), .Y(core__abc_21302_new_n5825_));
OAI21X1 OAI21X1_1329 ( .A(core__abc_21302_new_n5830_), .B(core__abc_21302_new_n5819_), .C(core__abc_21302_new_n4972_), .Y(core__abc_21302_new_n5831_));
OAI21X1 OAI21X1_133 ( .A(core_siphash_word_57_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf50), .Y(_abc_19873_new_n1758_));
OAI21X1 OAI21X1_1330 ( .A(core__abc_21302_new_n5828_), .B(core__abc_21302_new_n2364__bF_buf3), .C(core__abc_21302_new_n5833_), .Y(core__abc_21302_new_n5834_));
OAI21X1 OAI21X1_1331 ( .A(core__abc_21302_new_n5827_), .B(core__abc_21302_new_n5834_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n5835_));
OAI21X1 OAI21X1_1332 ( .A(core_v2_reg_47_), .B(core__abc_21302_new_n5104__bF_buf7), .C(reset_n_bF_buf41), .Y(core__abc_21302_new_n5836_));
OAI21X1 OAI21X1_1333 ( .A(core__abc_21302_new_n1753_), .B(core__abc_21302_new_n2364__bF_buf2), .C(core__abc_21302_new_n5844_), .Y(core__abc_21302_new_n5845_));
OAI21X1 OAI21X1_1334 ( .A(core_v2_reg_48_), .B(core__abc_21302_new_n5104__bF_buf5), .C(reset_n_bF_buf40), .Y(core__abc_21302_new_n5847_));
OAI21X1 OAI21X1_1335 ( .A(core__abc_21302_new_n5067_), .B(core__abc_21302_new_n5849_), .C(core__abc_21302_new_n4947_), .Y(core__abc_21302_new_n5850_));
OAI21X1 OAI21X1_1336 ( .A(core__abc_21302_new_n1763_), .B(core__abc_21302_new_n2364__bF_buf1), .C(core__abc_21302_new_n5852_), .Y(core__abc_21302_new_n5853_));
OAI21X1 OAI21X1_1337 ( .A(core__abc_21302_new_n2673__bF_buf8), .B(core__abc_21302_new_n5851_), .C(core__abc_21302_new_n5854_), .Y(core__abc_21302_new_n5855_));
OAI21X1 OAI21X1_1338 ( .A(core_v2_reg_49_), .B(core__abc_21302_new_n5104__bF_buf4), .C(core__abc_21302_new_n5855_), .Y(core__abc_21302_new_n5856_));
OAI21X1 OAI21X1_1339 ( .A(core__abc_21302_new_n4943_), .B(core__abc_21302_new_n4944_), .C(core__abc_21302_new_n5850_), .Y(core__abc_21302_new_n5858_));
OAI21X1 OAI21X1_134 ( .A(core_siphash_word_58_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf49), .Y(_abc_19873_new_n1760_));
OAI21X1 OAI21X1_1340 ( .A(core__abc_21302_new_n3340_), .B(core__abc_21302_new_n4945_), .C(core__abc_21302_new_n5858_), .Y(core__abc_21302_new_n5859_));
OAI21X1 OAI21X1_1341 ( .A(core__abc_21302_new_n5865_), .B(core__abc_21302_new_n2640__bF_buf1), .C(core__abc_21302_new_n5866_), .Y(core__abc_21302_new_n5867_));
OAI21X1 OAI21X1_1342 ( .A(core_v2_reg_50_), .B(core__abc_21302_new_n5104__bF_buf3), .C(reset_n_bF_buf39), .Y(core__abc_21302_new_n5869_));
OAI21X1 OAI21X1_1343 ( .A(core__abc_21302_new_n4929_), .B(core__abc_21302_new_n4951_), .C(core__abc_21302_new_n5860_), .Y(core__abc_21302_new_n5871_));
OAI21X1 OAI21X1_1344 ( .A(core_key_51_), .B(core__abc_21302_new_n2640__bF_buf0), .C(core__abc_21302_new_n5873_), .Y(core__abc_21302_new_n5874_));
OAI21X1 OAI21X1_1345 ( .A(core_v2_reg_51_), .B(core__abc_21302_new_n5104__bF_buf2), .C(reset_n_bF_buf38), .Y(core__abc_21302_new_n5876_));
OAI21X1 OAI21X1_1346 ( .A(core__abc_21302_new_n4955_), .B(core__abc_21302_new_n5878_), .C(core__abc_21302_new_n4926_), .Y(core__abc_21302_new_n5879_));
OAI21X1 OAI21X1_1347 ( .A(core_key_52_), .B(core__abc_21302_new_n2640__bF_buf11), .C(core__abc_21302_new_n5884_), .Y(core__abc_21302_new_n5885_));
OAI21X1 OAI21X1_1348 ( .A(core_v2_reg_52_), .B(core__abc_21302_new_n5104__bF_buf0), .C(reset_n_bF_buf37), .Y(core__abc_21302_new_n5887_));
OAI21X1 OAI21X1_1349 ( .A(core_key_53_), .B(core__abc_21302_new_n2640__bF_buf10), .C(core__abc_21302_new_n5894_), .Y(core__abc_21302_new_n5895_));
OAI21X1 OAI21X1_135 ( .A(core_siphash_word_59_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf48), .Y(_abc_19873_new_n1762_));
OAI21X1 OAI21X1_1350 ( .A(core_v2_reg_53_), .B(core__abc_21302_new_n5104__bF_buf6), .C(reset_n_bF_buf36), .Y(core__abc_21302_new_n5897_));
OAI21X1 OAI21X1_1351 ( .A(core__abc_21302_new_n4957_), .B(core__abc_21302_new_n5880_), .C(core__abc_21302_new_n4923_), .Y(core__abc_21302_new_n5900_));
OAI21X1 OAI21X1_1352 ( .A(core__abc_21302_new_n2673__bF_buf7), .B(core__abc_21302_new_n5903_), .C(core__abc_21302_new_n5905_), .Y(core__abc_21302_new_n5906_));
OAI21X1 OAI21X1_1353 ( .A(core_v2_reg_54_), .B(core__abc_21302_new_n5104__bF_buf4), .C(core__abc_21302_new_n5906_), .Y(core__abc_21302_new_n5907_));
OAI21X1 OAI21X1_1354 ( .A(core__abc_21302_new_n5899_), .B(core__abc_21302_new_n5900_), .C(core__abc_21302_new_n4910_), .Y(core__abc_21302_new_n5911_));
OAI21X1 OAI21X1_1355 ( .A(core__abc_21302_new_n2673__bF_buf6), .B(core__abc_21302_new_n5914_), .C(core__abc_21302_new_n5917_), .Y(core__abc_21302_new_n5918_));
OAI21X1 OAI21X1_1356 ( .A(core_v2_reg_55_), .B(core__abc_21302_new_n5104__bF_buf3), .C(core__abc_21302_new_n5918_), .Y(core__abc_21302_new_n5919_));
OAI21X1 OAI21X1_1357 ( .A(core_v2_reg_56_), .B(core__abc_21302_new_n5104__bF_buf1), .C(reset_n_bF_buf35), .Y(core__abc_21302_new_n5928_));
OAI21X1 OAI21X1_1358 ( .A(core__abc_21302_new_n4892_), .B(core__abc_21302_new_n5072_), .C(core__abc_21302_new_n4873_), .Y(core__abc_21302_new_n5930_));
OAI21X1 OAI21X1_1359 ( .A(core_v2_reg_57_), .B(core__abc_21302_new_n5104__bF_buf7), .C(reset_n_bF_buf34), .Y(core__abc_21302_new_n5935_));
OAI21X1 OAI21X1_136 ( .A(core_siphash_word_60_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf47), .Y(_abc_19873_new_n1765_));
OAI21X1 OAI21X1_1360 ( .A(core__abc_21302_new_n4890_), .B(core__abc_21302_new_n5922_), .C(core__abc_21302_new_n4875_), .Y(core__abc_21302_new_n5937_));
OAI21X1 OAI21X1_1361 ( .A(core_key_58_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n5939_), .Y(core__abc_21302_new_n5940_));
OAI21X1 OAI21X1_1362 ( .A(core_v2_reg_58_), .B(core__abc_21302_new_n5104__bF_buf6), .C(reset_n_bF_buf33), .Y(core__abc_21302_new_n5942_));
OAI21X1 OAI21X1_1363 ( .A(core__abc_21302_new_n2673__bF_buf5), .B(core__abc_21302_new_n5947_), .C(core__abc_21302_new_n5948_), .Y(core__abc_21302_new_n5949_));
OAI21X1 OAI21X1_1364 ( .A(core__abc_21302_new_n5944_), .B(core__abc_21302_new_n5949_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n5950_));
OAI21X1 OAI21X1_1365 ( .A(core_v2_reg_59_), .B(core__abc_21302_new_n5104__bF_buf4), .C(reset_n_bF_buf32), .Y(core__abc_21302_new_n5951_));
OAI21X1 OAI21X1_1366 ( .A(core__abc_21302_new_n4878_), .B(core__abc_21302_new_n5953_), .C(core__abc_21302_new_n4851_), .Y(core__abc_21302_new_n5954_));
OAI21X1 OAI21X1_1367 ( .A(core__abc_21302_new_n1902_), .B(core__abc_21302_new_n2364__bF_buf4), .C(core__abc_21302_new_n5960_), .Y(core__abc_21302_new_n5961_));
OAI21X1 OAI21X1_1368 ( .A(core_v2_reg_60_), .B(core__abc_21302_new_n5104__bF_buf2), .C(reset_n_bF_buf31), .Y(core__abc_21302_new_n5963_));
OAI21X1 OAI21X1_1369 ( .A(core__abc_21302_new_n4881_), .B(core__abc_21302_new_n5968_), .C(core__abc_21302_new_n5967_), .Y(core__abc_21302_new_n5969_));
OAI21X1 OAI21X1_137 ( .A(core_siphash_word_61_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf46), .Y(_abc_19873_new_n1767_));
OAI21X1 OAI21X1_1370 ( .A(core__abc_21302_new_n2673__bF_buf4), .B(core__abc_21302_new_n5970_), .C(core__abc_21302_new_n5972_), .Y(core__abc_21302_new_n5973_));
OAI21X1 OAI21X1_1371 ( .A(core_v2_reg_61_), .B(core__abc_21302_new_n5104__bF_buf1), .C(core__abc_21302_new_n5973_), .Y(core__abc_21302_new_n5974_));
OAI21X1 OAI21X1_1372 ( .A(core__abc_21302_new_n4852_), .B(core__abc_21302_new_n5955_), .C(core__abc_21302_new_n4882_), .Y(core__abc_21302_new_n5976_));
OAI21X1 OAI21X1_1373 ( .A(core__abc_21302_new_n2673__bF_buf3), .B(core__abc_21302_new_n5979_), .C(core__abc_21302_new_n5981_), .Y(core__abc_21302_new_n5982_));
OAI21X1 OAI21X1_1374 ( .A(core_v2_reg_62_), .B(core__abc_21302_new_n5104__bF_buf0), .C(core__abc_21302_new_n5982_), .Y(core__abc_21302_new_n5983_));
OAI21X1 OAI21X1_1375 ( .A(core__abc_21302_new_n2673__bF_buf2), .B(core__abc_21302_new_n5989_), .C(core__abc_21302_new_n5990_), .Y(core__abc_21302_new_n5991_));
OAI21X1 OAI21X1_1376 ( .A(core__abc_21302_new_n5986_), .B(core__abc_21302_new_n5991_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n5992_));
OAI21X1 OAI21X1_1377 ( .A(core_v2_reg_63_), .B(core__abc_21302_new_n5104__bF_buf7), .C(reset_n_bF_buf30), .Y(core__abc_21302_new_n5993_));
OAI21X1 OAI21X1_1378 ( .A(core__abc_21302_new_n1148_), .B(core__abc_21302_new_n2166_), .C(core__abc_21302_new_n2366_), .Y(core__abc_21302_new_n5995_));
OAI21X1 OAI21X1_1379 ( .A(core__abc_21302_new_n2363__bF_buf5), .B(core__abc_21302_new_n5995_), .C(core_v1_reg_0_), .Y(core__abc_21302_new_n5996_));
OAI21X1 OAI21X1_138 ( .A(core_siphash_word_62_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf45), .Y(_abc_19873_new_n1770_));
OAI21X1 OAI21X1_1380 ( .A(core_v1_reg_0_), .B(core__abc_21302_new_n5999__bF_buf5), .C(core__abc_21302_new_n5997_), .Y(core__abc_21302_new_n6000_));
OAI21X1 OAI21X1_1381 ( .A(core__abc_21302_new_n5373_), .B(core__abc_21302_new_n6001_), .C(core__abc_21302_new_n6002_), .Y(core__abc_21302_new_n6003_));
OAI21X1 OAI21X1_1382 ( .A(core__abc_21302_new_n6000_), .B(core__abc_21302_new_n6003_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n6004_));
OAI21X1 OAI21X1_1383 ( .A(core__abc_21302_new_n5405_), .B(core__abc_21302_new_n5710_), .C(core__abc_21302_new_n6006_), .Y(core__abc_21302_new_n6007_));
OAI21X1 OAI21X1_1384 ( .A(core__abc_21302_new_n4970_), .B(core__abc_21302_new_n5999__bF_buf4), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6010_));
OAI21X1 OAI21X1_1385 ( .A(core_v1_reg_1_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf29), .Y(core__abc_21302_new_n6012_));
OAI21X1 OAI21X1_1386 ( .A(core__abc_21302_new_n2363__bF_buf3), .B(core__abc_21302_new_n5995_), .C(core_v1_reg_2_), .Y(core__abc_21302_new_n6014_));
OAI21X1 OAI21X1_1387 ( .A(core__abc_21302_new_n5715_), .B(core__abc_21302_new_n5423_), .C(core__abc_21302_new_n6018_), .Y(core__abc_21302_new_n6019_));
OAI21X1 OAI21X1_1388 ( .A(core__abc_21302_new_n6016_), .B(core__abc_21302_new_n6019_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n6020_));
OAI21X1 OAI21X1_1389 ( .A(core__abc_21302_new_n2363__bF_buf2), .B(core__abc_21302_new_n5995_), .C(core_v1_reg_3_), .Y(core__abc_21302_new_n6022_));
OAI21X1 OAI21X1_139 ( .A(core_siphash_word_63_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf44), .Y(_abc_19873_new_n1772_));
OAI21X1 OAI21X1_1390 ( .A(core__abc_21302_new_n6027_), .B(core__abc_21302_new_n6025_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n6028_));
OAI21X1 OAI21X1_1391 ( .A(core__abc_21302_new_n2363__bF_buf1), .B(core__abc_21302_new_n5995_), .C(core_v1_reg_4_), .Y(core__abc_21302_new_n6030_));
OAI21X1 OAI21X1_1392 ( .A(core_v1_reg_4_), .B(core__abc_21302_new_n5999__bF_buf2), .C(core__abc_21302_new_n6032_), .Y(core__abc_21302_new_n6033_));
OAI21X1 OAI21X1_1393 ( .A(core__abc_21302_new_n5466_), .B(core__abc_21302_new_n6031_), .C(core__abc_21302_new_n6034_), .Y(core__abc_21302_new_n6035_));
OAI21X1 OAI21X1_1394 ( .A(core__abc_21302_new_n5479_), .B(core__abc_21302_new_n6038_), .C(core__abc_21302_new_n6039_), .Y(core__abc_21302_new_n6040_));
OAI21X1 OAI21X1_1395 ( .A(core__abc_21302_new_n1261_), .B(core__abc_21302_new_n5999__bF_buf1), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6042_));
OAI21X1 OAI21X1_1396 ( .A(core_v1_reg_5_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf28), .Y(core__abc_21302_new_n6044_));
OAI21X1 OAI21X1_1397 ( .A(core__abc_21302_new_n2363__bF_buf0), .B(core__abc_21302_new_n5995_), .C(core_v1_reg_6_), .Y(core__abc_21302_new_n6046_));
OAI21X1 OAI21X1_1398 ( .A(core__abc_21302_new_n6048_), .B(core__abc_21302_new_n6050_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n6051_));
OAI21X1 OAI21X1_1399 ( .A(core__abc_21302_new_n2363__bF_buf5), .B(core__abc_21302_new_n5995_), .C(core_v1_reg_7_), .Y(core__abc_21302_new_n6053_));
OAI21X1 OAI21X1_14 ( .A(_abc_19873_new_n1071_), .B(_abc_19873_new_n918_), .C(_abc_19873_new_n1072_), .Y(_abc_19873_new_n1073_));
OAI21X1 OAI21X1_140 ( .A(core_siphash_word_0_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf43), .Y(_abc_19873_new_n1775_));
OAI21X1 OAI21X1_1400 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n5756_), .C(core__abc_21302_new_n5509_), .Y(core__abc_21302_new_n6055_));
OAI21X1 OAI21X1_1401 ( .A(core__abc_21302_new_n6058_), .B(core__abc_21302_new_n6056_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n6059_));
OAI21X1 OAI21X1_1402 ( .A(core__abc_21302_new_n2673__bF_buf8), .B(core__abc_21302_new_n5764_), .C(core__abc_21302_new_n5530_), .Y(core__abc_21302_new_n6061_));
OAI21X1 OAI21X1_1403 ( .A(core__abc_21302_new_n2405_), .B(core__abc_21302_new_n5999__bF_buf4), .C(core__abc_21302_new_n6063_), .Y(core__abc_21302_new_n6064_));
OAI21X1 OAI21X1_1404 ( .A(core__abc_21302_new_n2915_), .B(core__abc_21302_new_n6064_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n6065_));
OAI21X1 OAI21X1_1405 ( .A(core_v1_reg_8_), .B(core__abc_21302_new_n6009__bF_buf5), .C(reset_n_bF_buf27), .Y(core__abc_21302_new_n6066_));
OAI21X1 OAI21X1_1406 ( .A(core__abc_21302_new_n5554_), .B(core__abc_21302_new_n5776_), .C(core__abc_21302_new_n2634__bF_buf2), .Y(core__abc_21302_new_n6069_));
OAI21X1 OAI21X1_1407 ( .A(core_key_73_), .B(core__abc_21302_new_n2640__bF_buf11), .C(core__abc_21302_new_n6071_), .Y(core__abc_21302_new_n6072_));
OAI21X1 OAI21X1_1408 ( .A(core__abc_21302_new_n6072_), .B(core__abc_21302_new_n6070_), .C(reset_n_bF_buf26), .Y(core__abc_21302_new_n6073_));
OAI21X1 OAI21X1_1409 ( .A(core__abc_21302_new_n5572_), .B(core__abc_21302_new_n5783_), .C(core__abc_21302_new_n2634__bF_buf1), .Y(core__abc_21302_new_n6076_));
OAI21X1 OAI21X1_141 ( .A(core_siphash_word_1_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf42), .Y(_abc_19873_new_n1778_));
OAI21X1 OAI21X1_1410 ( .A(core__abc_21302_new_n3000_), .B(core__abc_21302_new_n6077_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n6078_));
OAI21X1 OAI21X1_1411 ( .A(core_v1_reg_10_), .B(core__abc_21302_new_n6009__bF_buf2), .C(reset_n_bF_buf25), .Y(core__abc_21302_new_n6079_));
OAI21X1 OAI21X1_1412 ( .A(core__abc_21302_new_n6081_), .B(core__abc_21302_new_n5791_), .C(core__abc_21302_new_n2634__bF_buf0), .Y(core__abc_21302_new_n6082_));
OAI21X1 OAI21X1_1413 ( .A(core_key_75_), .B(core__abc_21302_new_n2640__bF_buf10), .C(core__abc_21302_new_n6084_), .Y(core__abc_21302_new_n6085_));
OAI21X1 OAI21X1_1414 ( .A(core__abc_21302_new_n6085_), .B(core__abc_21302_new_n6083_), .C(reset_n_bF_buf24), .Y(core__abc_21302_new_n6086_));
OAI21X1 OAI21X1_1415 ( .A(core__abc_21302_new_n5603_), .B(core__abc_21302_new_n5804_), .C(core__abc_21302_new_n2634__bF_buf8), .Y(core__abc_21302_new_n6089_));
OAI21X1 OAI21X1_1416 ( .A(core__abc_21302_new_n3082_), .B(core__abc_21302_new_n6090_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n6091_));
OAI21X1 OAI21X1_1417 ( .A(core_v1_reg_12_), .B(core__abc_21302_new_n6009__bF_buf0), .C(reset_n_bF_buf23), .Y(core__abc_21302_new_n6092_));
OAI21X1 OAI21X1_1418 ( .A(core__abc_21302_new_n5625_), .B(core__abc_21302_new_n5813_), .C(core__abc_21302_new_n2634__bF_buf7), .Y(core__abc_21302_new_n6094_));
OAI21X1 OAI21X1_1419 ( .A(core_key_77_), .B(core__abc_21302_new_n2640__bF_buf9), .C(core__abc_21302_new_n6096_), .Y(core__abc_21302_new_n6097_));
OAI21X1 OAI21X1_142 ( .A(core_siphash_word_2_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf41), .Y(_abc_19873_new_n1781_));
OAI21X1 OAI21X1_1420 ( .A(core__abc_21302_new_n6100_), .B(core__abc_21302_new_n5820_), .C(core__abc_21302_new_n6101_), .Y(core__abc_21302_new_n6102_));
OAI21X1 OAI21X1_1421 ( .A(core__abc_21302_new_n4360_), .B(core__abc_21302_new_n5999__bF_buf1), .C(core__abc_21302_new_n6102_), .Y(core__abc_21302_new_n6103_));
OAI21X1 OAI21X1_1422 ( .A(core__abc_21302_new_n3175_), .B(core__abc_21302_new_n6103_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n6104_));
OAI21X1 OAI21X1_1423 ( .A(core_v1_reg_14_), .B(core__abc_21302_new_n6009__bF_buf7), .C(reset_n_bF_buf22), .Y(core__abc_21302_new_n6105_));
OAI21X1 OAI21X1_1424 ( .A(core__abc_21302_new_n5670_), .B(core__abc_21302_new_n5832_), .C(core__abc_21302_new_n6107_), .Y(core__abc_21302_new_n6108_));
OAI21X1 OAI21X1_1425 ( .A(core__abc_21302_new_n4847_), .B(core__abc_21302_new_n5999__bF_buf0), .C(core__abc_21302_new_n6108_), .Y(core__abc_21302_new_n6109_));
OAI21X1 OAI21X1_1426 ( .A(core__abc_21302_new_n3259_), .B(core__abc_21302_new_n6109_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n6110_));
OAI21X1 OAI21X1_1427 ( .A(core_v1_reg_15_), .B(core__abc_21302_new_n6009__bF_buf5), .C(reset_n_bF_buf21), .Y(core__abc_21302_new_n6111_));
OAI21X1 OAI21X1_1428 ( .A(core__abc_21302_new_n5687_), .B(core__abc_21302_new_n5842_), .C(core__abc_21302_new_n2634__bF_buf6), .Y(core__abc_21302_new_n6114_));
OAI21X1 OAI21X1_1429 ( .A(core__abc_21302_new_n3266_), .B(core__abc_21302_new_n6115_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n6116_));
OAI21X1 OAI21X1_143 ( .A(core_siphash_word_3_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf40), .Y(_abc_19873_new_n1784_));
OAI21X1 OAI21X1_1430 ( .A(core_v1_reg_16_), .B(core__abc_21302_new_n6009__bF_buf3), .C(reset_n_bF_buf20), .Y(core__abc_21302_new_n6117_));
OAI21X1 OAI21X1_1431 ( .A(core__abc_21302_new_n5047_), .B(core__abc_21302_new_n5851_), .C(core__abc_21302_new_n6119_), .Y(core__abc_21302_new_n6120_));
OAI21X1 OAI21X1_1432 ( .A(core__abc_21302_new_n4833_), .B(core__abc_21302_new_n5999__bF_buf4), .C(core__abc_21302_new_n6120_), .Y(core__abc_21302_new_n6121_));
OAI21X1 OAI21X1_1433 ( .A(core__abc_21302_new_n3328_), .B(core__abc_21302_new_n6121_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n6122_));
OAI21X1 OAI21X1_1434 ( .A(core_v1_reg_17_), .B(core__abc_21302_new_n6009__bF_buf1), .C(reset_n_bF_buf19), .Y(core__abc_21302_new_n6123_));
OAI21X1 OAI21X1_1435 ( .A(core__abc_21302_new_n6125_), .B(core__abc_21302_new_n5863_), .C(core__abc_21302_new_n6126_), .Y(core__abc_21302_new_n6127_));
OAI21X1 OAI21X1_1436 ( .A(core__abc_21302_new_n4824_), .B(core__abc_21302_new_n5999__bF_buf3), .C(core__abc_21302_new_n6127_), .Y(core__abc_21302_new_n6128_));
OAI21X1 OAI21X1_1437 ( .A(core__abc_21302_new_n3368_), .B(core__abc_21302_new_n6128_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n6129_));
OAI21X1 OAI21X1_1438 ( .A(core_v1_reg_18_), .B(core__abc_21302_new_n6009__bF_buf9), .C(reset_n_bF_buf18), .Y(core__abc_21302_new_n6130_));
OAI21X1 OAI21X1_1439 ( .A(core__abc_21302_new_n6132_), .B(core__abc_21302_new_n5872_), .C(core__abc_21302_new_n6133_), .Y(core__abc_21302_new_n6134_));
OAI21X1 OAI21X1_144 ( .A(core_siphash_word_4_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf39), .Y(_abc_19873_new_n1787_));
OAI21X1 OAI21X1_1440 ( .A(core__abc_21302_new_n3452_), .B(core__abc_21302_new_n2640__bF_buf8), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6135_));
OAI21X1 OAI21X1_1441 ( .A(core_v1_reg_19_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf17), .Y(core__abc_21302_new_n6137_));
OAI21X1 OAI21X1_1442 ( .A(core__abc_21302_new_n6142_), .B(core__abc_21302_new_n5999__bF_buf2), .C(core__abc_21302_new_n6009__bF_buf5), .Y(core__abc_21302_new_n6143_));
OAI21X1 OAI21X1_1443 ( .A(core_v1_reg_20_), .B(core__abc_21302_new_n6009__bF_buf4), .C(reset_n_bF_buf16), .Y(core__abc_21302_new_n6145_));
OAI21X1 OAI21X1_1444 ( .A(core__abc_21302_new_n5035_), .B(core__abc_21302_new_n5892_), .C(core__abc_21302_new_n6147_), .Y(core__abc_21302_new_n6148_));
OAI21X1 OAI21X1_1445 ( .A(core__abc_21302_new_n5113_), .B(core__abc_21302_new_n5999__bF_buf1), .C(core__abc_21302_new_n6148_), .Y(core__abc_21302_new_n6149_));
OAI21X1 OAI21X1_1446 ( .A(core__abc_21302_new_n3499_), .B(core__abc_21302_new_n6149_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n6150_));
OAI21X1 OAI21X1_1447 ( .A(core_v1_reg_21_), .B(core__abc_21302_new_n6009__bF_buf3), .C(reset_n_bF_buf15), .Y(core__abc_21302_new_n6151_));
OAI21X1 OAI21X1_1448 ( .A(core__abc_21302_new_n6154_), .B(core__abc_21302_new_n6153_), .C(core__abc_21302_new_n2634__bF_buf4), .Y(core__abc_21302_new_n6155_));
OAI21X1 OAI21X1_1449 ( .A(core__abc_21302_new_n5136_), .B(core__abc_21302_new_n5999__bF_buf0), .C(core__abc_21302_new_n6155_), .Y(core__abc_21302_new_n6156_));
OAI21X1 OAI21X1_145 ( .A(core_siphash_word_5_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf38), .Y(_abc_19873_new_n1790_));
OAI21X1 OAI21X1_1450 ( .A(core__abc_21302_new_n3531_), .B(core__abc_21302_new_n6156_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n6157_));
OAI21X1 OAI21X1_1451 ( .A(core_v1_reg_22_), .B(core__abc_21302_new_n6009__bF_buf1), .C(reset_n_bF_buf14), .Y(core__abc_21302_new_n6158_));
OAI21X1 OAI21X1_1452 ( .A(core__abc_21302_new_n5025_), .B(core__abc_21302_new_n5914_), .C(core__abc_21302_new_n6160_), .Y(core__abc_21302_new_n6161_));
OAI21X1 OAI21X1_1453 ( .A(core__abc_21302_new_n6162_), .B(core__abc_21302_new_n5999__bF_buf5), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6163_));
OAI21X1 OAI21X1_1454 ( .A(core_v1_reg_23_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf13), .Y(core__abc_21302_new_n6165_));
OAI21X1 OAI21X1_1455 ( .A(core__abc_21302_new_n5017_), .B(core__abc_21302_new_n5018_), .C(core__abc_21302_new_n5923_), .Y(core__abc_21302_new_n6168_));
OAI21X1 OAI21X1_1456 ( .A(core__abc_21302_new_n2453_), .B(core__abc_21302_new_n5999__bF_buf4), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6170_));
OAI21X1 OAI21X1_1457 ( .A(core_v1_reg_24_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf12), .Y(core__abc_21302_new_n6172_));
OAI21X1 OAI21X1_1458 ( .A(core__abc_21302_new_n5012_), .B(core__abc_21302_new_n5931_), .C(core__abc_21302_new_n6174_), .Y(core__abc_21302_new_n6175_));
OAI21X1 OAI21X1_1459 ( .A(core__abc_21302_new_n6176_), .B(core__abc_21302_new_n5999__bF_buf3), .C(core__abc_21302_new_n6009__bF_buf5), .Y(core__abc_21302_new_n6177_));
OAI21X1 OAI21X1_146 ( .A(core_siphash_word_6_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf37), .Y(_abc_19873_new_n1793_));
OAI21X1 OAI21X1_1460 ( .A(core_v1_reg_25_), .B(core__abc_21302_new_n6009__bF_buf4), .C(reset_n_bF_buf11), .Y(core__abc_21302_new_n6179_));
OAI21X1 OAI21X1_1461 ( .A(core__abc_21302_new_n5010_), .B(core__abc_21302_new_n5938_), .C(core__abc_21302_new_n2634__bF_buf2), .Y(core__abc_21302_new_n6182_));
OAI21X1 OAI21X1_1462 ( .A(core__abc_21302_new_n5210_), .B(core__abc_21302_new_n5999__bF_buf2), .C(core__abc_21302_new_n6009__bF_buf3), .Y(core__abc_21302_new_n6183_));
OAI21X1 OAI21X1_1463 ( .A(core__abc_21302_new_n6181_), .B(core__abc_21302_new_n6182_), .C(core__abc_21302_new_n6184_), .Y(core__abc_21302_new_n6185_));
OAI21X1 OAI21X1_1464 ( .A(core_v1_reg_26_), .B(core__abc_21302_new_n6009__bF_buf2), .C(core__abc_21302_new_n6185_), .Y(core__abc_21302_new_n6186_));
OAI21X1 OAI21X1_1465 ( .A(core__abc_21302_new_n5001_), .B(core__abc_21302_new_n5947_), .C(core__abc_21302_new_n6188_), .Y(core__abc_21302_new_n6189_));
OAI21X1 OAI21X1_1466 ( .A(core_key_91_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n6009__bF_buf1), .Y(core__abc_21302_new_n6190_));
OAI21X1 OAI21X1_1467 ( .A(core_v1_reg_27_), .B(core__abc_21302_new_n6009__bF_buf0), .C(reset_n_bF_buf10), .Y(core__abc_21302_new_n6192_));
OAI21X1 OAI21X1_1468 ( .A(core__abc_21302_new_n5968_), .B(core__abc_21302_new_n5957_), .C(core__abc_21302_new_n5003_), .Y(core__abc_21302_new_n6195_));
OAI21X1 OAI21X1_1469 ( .A(core__abc_21302_new_n5248_), .B(core__abc_21302_new_n5999__bF_buf1), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6197_));
OAI21X1 OAI21X1_147 ( .A(core_siphash_word_7_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf36), .Y(_abc_19873_new_n1795_));
OAI21X1 OAI21X1_1470 ( .A(core_v1_reg_28_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf9), .Y(core__abc_21302_new_n6199_));
OAI21X1 OAI21X1_1471 ( .A(core__abc_21302_new_n4979_), .B(core__abc_21302_new_n5970_), .C(core__abc_21302_new_n6201_), .Y(core__abc_21302_new_n6202_));
OAI21X1 OAI21X1_1472 ( .A(core_key_93_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6203_));
OAI21X1 OAI21X1_1473 ( .A(core_v1_reg_29_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf8), .Y(core__abc_21302_new_n6205_));
OAI21X1 OAI21X1_1474 ( .A(core__abc_21302_new_n4977_), .B(core__abc_21302_new_n5979_), .C(core__abc_21302_new_n6208_), .Y(core__abc_21302_new_n6209_));
OAI21X1 OAI21X1_1475 ( .A(core__abc_21302_new_n6207_), .B(core__abc_21302_new_n5999__bF_buf0), .C(core__abc_21302_new_n6209_), .Y(core__abc_21302_new_n6210_));
OAI21X1 OAI21X1_1476 ( .A(core__abc_21302_new_n3830_), .B(core__abc_21302_new_n6210_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n6211_));
OAI21X1 OAI21X1_1477 ( .A(core_v1_reg_30_), .B(core__abc_21302_new_n6009__bF_buf5), .C(reset_n_bF_buf7), .Y(core__abc_21302_new_n6212_));
OAI21X1 OAI21X1_1478 ( .A(core__abc_21302_new_n4971_), .B(core__abc_21302_new_n5989_), .C(core__abc_21302_new_n6214_), .Y(core__abc_21302_new_n6215_));
OAI21X1 OAI21X1_1479 ( .A(core__abc_21302_new_n5311_), .B(core__abc_21302_new_n5999__bF_buf5), .C(core__abc_21302_new_n6009__bF_buf3), .Y(core__abc_21302_new_n6216_));
OAI21X1 OAI21X1_148 ( .A(core_siphash_word_8_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf35), .Y(_abc_19873_new_n1797_));
OAI21X1 OAI21X1_1480 ( .A(core_v1_reg_31_), .B(core__abc_21302_new_n6009__bF_buf2), .C(reset_n_bF_buf6), .Y(core__abc_21302_new_n6218_));
OAI21X1 OAI21X1_1481 ( .A(core__abc_21302_new_n5325_), .B(core__abc_21302_new_n5999__bF_buf4), .C(core__abc_21302_new_n6009__bF_buf1), .Y(core__abc_21302_new_n6223_));
OAI21X1 OAI21X1_1482 ( .A(core_v1_reg_32_), .B(core__abc_21302_new_n6009__bF_buf0), .C(reset_n_bF_buf5), .Y(core__abc_21302_new_n6225_));
OAI21X1 OAI21X1_1483 ( .A(core__abc_21302_new_n4946_), .B(core__abc_21302_new_n5097_), .C(core__abc_21302_new_n6227_), .Y(core__abc_21302_new_n6228_));
OAI21X1 OAI21X1_1484 ( .A(core__abc_21302_new_n1576_), .B(core__abc_21302_new_n5999__bF_buf3), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6229_));
OAI21X1 OAI21X1_1485 ( .A(core_v1_reg_33_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf4), .Y(core__abc_21302_new_n6231_));
OAI21X1 OAI21X1_1486 ( .A(core__abc_21302_new_n4945_), .B(core__abc_21302_new_n5124_), .C(core__abc_21302_new_n6233_), .Y(core__abc_21302_new_n6234_));
OAI21X1 OAI21X1_1487 ( .A(core__abc_21302_new_n1588_), .B(core__abc_21302_new_n5999__bF_buf2), .C(core__abc_21302_new_n6234_), .Y(core__abc_21302_new_n6235_));
OAI21X1 OAI21X1_1488 ( .A(core__abc_21302_new_n3970_), .B(core__abc_21302_new_n6235_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n6236_));
OAI21X1 OAI21X1_1489 ( .A(core_v1_reg_34_), .B(core__abc_21302_new_n6009__bF_buf7), .C(reset_n_bF_buf3), .Y(core__abc_21302_new_n6237_));
OAI21X1 OAI21X1_149 ( .A(core_siphash_word_9_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf34), .Y(_abc_19873_new_n1799_));
OAI21X1 OAI21X1_1490 ( .A(core__abc_21302_new_n4930_), .B(core__abc_21302_new_n5145_), .C(core__abc_21302_new_n6239_), .Y(core__abc_21302_new_n6240_));
OAI21X1 OAI21X1_1491 ( .A(core__abc_21302_new_n4025_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n6009__bF_buf5), .Y(core__abc_21302_new_n6241_));
OAI21X1 OAI21X1_1492 ( .A(core_v1_reg_35_), .B(core__abc_21302_new_n6009__bF_buf4), .C(reset_n_bF_buf2), .Y(core__abc_21302_new_n6243_));
OAI21X1 OAI21X1_1493 ( .A(core__abc_21302_new_n6245_), .B(core__abc_21302_new_n5168_), .C(core__abc_21302_new_n6246_), .Y(core__abc_21302_new_n6247_));
OAI21X1 OAI21X1_1494 ( .A(core__abc_21302_new_n5422_), .B(core__abc_21302_new_n5999__bF_buf1), .C(core__abc_21302_new_n6247_), .Y(core__abc_21302_new_n6248_));
OAI21X1 OAI21X1_1495 ( .A(core__abc_21302_new_n4031_), .B(core__abc_21302_new_n6248_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n6249_));
OAI21X1 OAI21X1_1496 ( .A(core_v1_reg_36_), .B(core__abc_21302_new_n6009__bF_buf3), .C(reset_n_bF_buf1), .Y(core__abc_21302_new_n6250_));
OAI21X1 OAI21X1_1497 ( .A(core__abc_21302_new_n4925_), .B(core__abc_21302_new_n5181_), .C(core__abc_21302_new_n6252_), .Y(core__abc_21302_new_n6253_));
OAI21X1 OAI21X1_1498 ( .A(core_key_101_), .B(core__abc_21302_new_n2640__bF_buf4), .C(core__abc_21302_new_n6009__bF_buf1), .Y(core__abc_21302_new_n6254_));
OAI21X1 OAI21X1_1499 ( .A(core_v1_reg_37_), .B(core__abc_21302_new_n6009__bF_buf0), .C(reset_n_bF_buf0), .Y(core__abc_21302_new_n6256_));
OAI21X1 OAI21X1_15 ( .A(_abc_19873_new_n1139_), .B(_abc_19873_new_n894__bF_buf0), .C(_abc_19873_new_n1140_), .Y(_abc_19873_new_n1141_));
OAI21X1 OAI21X1_150 ( .A(core_siphash_word_10_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf33), .Y(_abc_19873_new_n1801_));
OAI21X1 OAI21X1_1500 ( .A(core_key_102_), .B(core__abc_21302_new_n2640__bF_buf3), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6261_));
OAI21X1 OAI21X1_1501 ( .A(core_v1_reg_38_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf69), .Y(core__abc_21302_new_n6263_));
OAI21X1 OAI21X1_1502 ( .A(core__abc_21302_new_n5478_), .B(core__abc_21302_new_n5999__bF_buf0), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6270_));
OAI21X1 OAI21X1_1503 ( .A(core_v1_reg_39_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf68), .Y(core__abc_21302_new_n6272_));
OAI21X1 OAI21X1_1504 ( .A(core__abc_21302_new_n6274_), .B(core__abc_21302_new_n5242_), .C(core__abc_21302_new_n2634__bF_buf6), .Y(core__abc_21302_new_n6276_));
OAI21X1 OAI21X1_1505 ( .A(core__abc_21302_new_n6275_), .B(core__abc_21302_new_n6276_), .C(core__abc_21302_new_n6277_), .Y(core__abc_21302_new_n6278_));
OAI21X1 OAI21X1_1506 ( .A(core__abc_21302_new_n4154_), .B(core__abc_21302_new_n6278_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n6279_));
OAI21X1 OAI21X1_1507 ( .A(core_v1_reg_40_), .B(core__abc_21302_new_n6009__bF_buf5), .C(reset_n_bF_buf67), .Y(core__abc_21302_new_n6280_));
OAI21X1 OAI21X1_1508 ( .A(core__abc_21302_new_n6282_), .B(core__abc_21302_new_n5256_), .C(core__abc_21302_new_n6283_), .Y(core__abc_21302_new_n6284_));
OAI21X1 OAI21X1_1509 ( .A(core__abc_21302_new_n5507_), .B(core__abc_21302_new_n5999__bF_buf5), .C(core__abc_21302_new_n6009__bF_buf3), .Y(core__abc_21302_new_n6285_));
OAI21X1 OAI21X1_151 ( .A(core_siphash_word_11_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf32), .Y(_abc_19873_new_n1803_));
OAI21X1 OAI21X1_1510 ( .A(core_v1_reg_41_), .B(core__abc_21302_new_n6009__bF_buf2), .C(reset_n_bF_buf66), .Y(core__abc_21302_new_n6287_));
OAI21X1 OAI21X1_1511 ( .A(core__abc_21302_new_n4869_), .B(core__abc_21302_new_n5278_), .C(core__abc_21302_new_n6289_), .Y(core__abc_21302_new_n6290_));
OAI21X1 OAI21X1_1512 ( .A(core__abc_21302_new_n5528_), .B(core__abc_21302_new_n5999__bF_buf4), .C(core__abc_21302_new_n6009__bF_buf1), .Y(core__abc_21302_new_n6291_));
OAI21X1 OAI21X1_1513 ( .A(core_v1_reg_42_), .B(core__abc_21302_new_n6009__bF_buf0), .C(reset_n_bF_buf65), .Y(core__abc_21302_new_n6293_));
OAI21X1 OAI21X1_1514 ( .A(core__abc_21302_new_n4864_), .B(core__abc_21302_new_n5296_), .C(core__abc_21302_new_n6295_), .Y(core__abc_21302_new_n6296_));
OAI21X1 OAI21X1_1515 ( .A(core__abc_21302_new_n4268_), .B(core__abc_21302_new_n2640__bF_buf2), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6297_));
OAI21X1 OAI21X1_1516 ( .A(core_v1_reg_43_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf64), .Y(core__abc_21302_new_n6299_));
OAI21X1 OAI21X1_1517 ( .A(core__abc_21302_new_n6304_), .B(core__abc_21302_new_n5999__bF_buf3), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6305_));
OAI21X1 OAI21X1_1518 ( .A(core_v1_reg_44_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf63), .Y(core__abc_21302_new_n6307_));
OAI21X1 OAI21X1_1519 ( .A(core_key_109_), .B(core__abc_21302_new_n2640__bF_buf1), .C(core__abc_21302_new_n6009__bF_buf5), .Y(core__abc_21302_new_n6312_));
OAI21X1 OAI21X1_152 ( .A(core_siphash_word_12_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf31), .Y(_abc_19873_new_n1805_));
OAI21X1 OAI21X1_1520 ( .A(core_v1_reg_45_), .B(core__abc_21302_new_n6009__bF_buf4), .C(reset_n_bF_buf62), .Y(core__abc_21302_new_n6314_));
OAI21X1 OAI21X1_1521 ( .A(core__abc_21302_new_n6317_), .B(core__abc_21302_new_n5362_), .C(core__abc_21302_new_n6318_), .Y(core__abc_21302_new_n6319_));
OAI21X1 OAI21X1_1522 ( .A(core_key_110_), .B(core__abc_21302_new_n2640__bF_buf0), .C(core__abc_21302_new_n6009__bF_buf3), .Y(core__abc_21302_new_n6320_));
OAI21X1 OAI21X1_1523 ( .A(core_v1_reg_46_), .B(core__abc_21302_new_n6009__bF_buf2), .C(reset_n_bF_buf61), .Y(core__abc_21302_new_n6322_));
OAI21X1 OAI21X1_1524 ( .A(core__abc_21302_new_n4836_), .B(core__abc_21302_new_n5381_), .C(core__abc_21302_new_n6324_), .Y(core__abc_21302_new_n6325_));
OAI21X1 OAI21X1_1525 ( .A(core_v1_reg_47_), .B(core__abc_21302_new_n6009__bF_buf0), .C(reset_n_bF_buf60), .Y(core__abc_21302_new_n6328_));
OAI21X1 OAI21X1_1526 ( .A(core__abc_21302_new_n4828_), .B(core__abc_21302_new_n5409_), .C(core__abc_21302_new_n2634__bF_buf3), .Y(core__abc_21302_new_n6332_));
OAI21X1 OAI21X1_1527 ( .A(core__abc_21302_new_n4385_), .B(core__abc_21302_new_n6333_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n6334_));
OAI21X1 OAI21X1_1528 ( .A(core_v1_reg_48_), .B(core__abc_21302_new_n6009__bF_buf9), .C(reset_n_bF_buf59), .Y(core__abc_21302_new_n6335_));
OAI21X1 OAI21X1_1529 ( .A(core__abc_21302_new_n6337_), .B(core__abc_21302_new_n5427_), .C(core__abc_21302_new_n6338_), .Y(core__abc_21302_new_n6339_));
OAI21X1 OAI21X1_153 ( .A(core_siphash_word_13_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf30), .Y(_abc_19873_new_n1808_));
OAI21X1 OAI21X1_1530 ( .A(core__abc_21302_new_n3379_), .B(core__abc_21302_new_n5999__bF_buf1), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6340_));
OAI21X1 OAI21X1_1531 ( .A(core_v1_reg_49_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf58), .Y(core__abc_21302_new_n6342_));
OAI21X1 OAI21X1_1532 ( .A(core__abc_21302_new_n5447_), .B(core__abc_21302_new_n6345_), .C(core__abc_21302_new_n5107_), .Y(core__abc_21302_new_n6346_));
OAI21X1 OAI21X1_1533 ( .A(core_key_114_), .B(core__abc_21302_new_n2640__bF_buf11), .C(core__abc_21302_new_n6009__bF_buf5), .Y(core__abc_21302_new_n6348_));
OAI21X1 OAI21X1_1534 ( .A(core_v1_reg_50_), .B(core__abc_21302_new_n6009__bF_buf4), .C(reset_n_bF_buf57), .Y(core__abc_21302_new_n6350_));
OAI21X1 OAI21X1_1535 ( .A(core__abc_21302_new_n5133_), .B(core__abc_21302_new_n5459_), .C(core__abc_21302_new_n6352_), .Y(core__abc_21302_new_n6353_));
OAI21X1 OAI21X1_1536 ( .A(core__abc_21302_new_n6354_), .B(core__abc_21302_new_n5999__bF_buf0), .C(core__abc_21302_new_n6009__bF_buf3), .Y(core__abc_21302_new_n6355_));
OAI21X1 OAI21X1_1537 ( .A(core_v1_reg_51_), .B(core__abc_21302_new_n6009__bF_buf2), .C(reset_n_bF_buf56), .Y(core__abc_21302_new_n6357_));
OAI21X1 OAI21X1_1538 ( .A(core__abc_21302_new_n5155_), .B(core__abc_21302_new_n5485_), .C(core__abc_21302_new_n2634__bF_buf1), .Y(core__abc_21302_new_n6360_));
OAI21X1 OAI21X1_1539 ( .A(core__abc_21302_new_n1794_), .B(core__abc_21302_new_n5999__bF_buf5), .C(core__abc_21302_new_n6009__bF_buf1), .Y(core__abc_21302_new_n6361_));
OAI21X1 OAI21X1_154 ( .A(core_siphash_word_14_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf29), .Y(_abc_19873_new_n1810_));
OAI21X1 OAI21X1_1540 ( .A(core__abc_21302_new_n6359_), .B(core__abc_21302_new_n6360_), .C(core__abc_21302_new_n6362_), .Y(core__abc_21302_new_n6363_));
OAI21X1 OAI21X1_1541 ( .A(core_v1_reg_52_), .B(core__abc_21302_new_n6009__bF_buf0), .C(core__abc_21302_new_n6363_), .Y(core__abc_21302_new_n6364_));
OAI21X1 OAI21X1_1542 ( .A(core__abc_21302_new_n5151_), .B(core__abc_21302_new_n5501_), .C(core__abc_21302_new_n6366_), .Y(core__abc_21302_new_n6367_));
OAI21X1 OAI21X1_1543 ( .A(core_key_117_), .B(core__abc_21302_new_n2640__bF_buf10), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6368_));
OAI21X1 OAI21X1_1544 ( .A(core_v1_reg_53_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf55), .Y(core__abc_21302_new_n6370_));
OAI21X1 OAI21X1_1545 ( .A(core__abc_21302_new_n5176_), .B(core__abc_21302_new_n5522_), .C(core__abc_21302_new_n6372_), .Y(core__abc_21302_new_n6373_));
OAI21X1 OAI21X1_1546 ( .A(core_key_118_), .B(core__abc_21302_new_n2640__bF_buf9), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6374_));
OAI21X1 OAI21X1_1547 ( .A(core_v1_reg_54_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf54), .Y(core__abc_21302_new_n6376_));
OAI21X1 OAI21X1_1548 ( .A(core__abc_21302_new_n5536_), .B(core__abc_21302_new_n5519_), .C(core__abc_21302_new_n5534_), .Y(core__abc_21302_new_n6379_));
OAI21X1 OAI21X1_1549 ( .A(core__abc_21302_new_n5034_), .B(core__abc_21302_new_n5999__bF_buf4), .C(core__abc_21302_new_n6009__bF_buf5), .Y(core__abc_21302_new_n6383_));
OAI21X1 OAI21X1_155 ( .A(core_siphash_word_15_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf28), .Y(_abc_19873_new_n1812_));
OAI21X1 OAI21X1_1550 ( .A(core_v1_reg_55_), .B(core__abc_21302_new_n6009__bF_buf4), .C(reset_n_bF_buf53), .Y(core__abc_21302_new_n6385_));
OAI21X1 OAI21X1_1551 ( .A(core__abc_21302_new_n5231_), .B(core__abc_21302_new_n5563_), .C(core__abc_21302_new_n6387_), .Y(core__abc_21302_new_n6388_));
OAI21X1 OAI21X1_1552 ( .A(core__abc_21302_new_n1845_), .B(core__abc_21302_new_n5999__bF_buf3), .C(core__abc_21302_new_n6009__bF_buf3), .Y(core__abc_21302_new_n6389_));
OAI21X1 OAI21X1_1553 ( .A(core_v1_reg_56_), .B(core__abc_21302_new_n6009__bF_buf2), .C(reset_n_bF_buf52), .Y(core__abc_21302_new_n6391_));
OAI21X1 OAI21X1_1554 ( .A(core__abc_21302_new_n5024_), .B(core__abc_21302_new_n5999__bF_buf2), .C(core__abc_21302_new_n6009__bF_buf1), .Y(core__abc_21302_new_n6398_));
OAI21X1 OAI21X1_1555 ( .A(core_v1_reg_57_), .B(core__abc_21302_new_n6009__bF_buf0), .C(reset_n_bF_buf51), .Y(core__abc_21302_new_n6400_));
OAI21X1 OAI21X1_1556 ( .A(core__abc_21302_new_n5252_), .B(core__abc_21302_new_n5595_), .C(core__abc_21302_new_n6402_), .Y(core__abc_21302_new_n6403_));
OAI21X1 OAI21X1_1557 ( .A(core_key_122_), .B(core__abc_21302_new_n2640__bF_buf8), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6404_));
OAI21X1 OAI21X1_1558 ( .A(core_v1_reg_58_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf50), .Y(core__abc_21302_new_n6406_));
OAI21X1 OAI21X1_1559 ( .A(core__abc_21302_new_n5609_), .B(core__abc_21302_new_n5592_), .C(core__abc_21302_new_n5607_), .Y(core__abc_21302_new_n6409_));
OAI21X1 OAI21X1_156 ( .A(core_siphash_word_16_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf27), .Y(_abc_19873_new_n1814_));
OAI21X1 OAI21X1_1560 ( .A(core__abc_21302_new_n4692_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n6009__bF_buf7), .Y(core__abc_21302_new_n6414_));
OAI21X1 OAI21X1_1561 ( .A(core_v1_reg_59_), .B(core__abc_21302_new_n6009__bF_buf6), .C(reset_n_bF_buf49), .Y(core__abc_21302_new_n6416_));
OAI21X1 OAI21X1_1562 ( .A(core__abc_21302_new_n6419_), .B(core__abc_21302_new_n5638_), .C(core__abc_21302_new_n6420_), .Y(core__abc_21302_new_n6421_));
OAI21X1 OAI21X1_1563 ( .A(core__abc_21302_new_n6422_), .B(core__abc_21302_new_n2139_), .C(core__abc_21302_new_n6009__bF_buf5), .Y(core__abc_21302_new_n6423_));
OAI21X1 OAI21X1_1564 ( .A(core_v1_reg_60_), .B(core__abc_21302_new_n6009__bF_buf4), .C(reset_n_bF_buf48), .Y(core__abc_21302_new_n6425_));
OAI21X1 OAI21X1_1565 ( .A(core__abc_21302_new_n5312_), .B(core__abc_21302_new_n5657_), .C(core__abc_21302_new_n6427_), .Y(core__abc_21302_new_n6428_));
OAI21X1 OAI21X1_1566 ( .A(core_key_125_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n6009__bF_buf3), .Y(core__abc_21302_new_n6429_));
OAI21X1 OAI21X1_1567 ( .A(core_v1_reg_61_), .B(core__abc_21302_new_n6009__bF_buf2), .C(reset_n_bF_buf47), .Y(core__abc_21302_new_n6431_));
OAI21X1 OAI21X1_1568 ( .A(core__abc_21302_new_n5328_), .B(core__abc_21302_new_n5677_), .C(core__abc_21302_new_n6433_), .Y(core__abc_21302_new_n6434_));
OAI21X1 OAI21X1_1569 ( .A(core_key_126_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n6009__bF_buf1), .Y(core__abc_21302_new_n6435_));
OAI21X1 OAI21X1_157 ( .A(core_siphash_word_17_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf26), .Y(_abc_19873_new_n1816_));
OAI21X1 OAI21X1_1570 ( .A(core_v1_reg_62_), .B(core__abc_21302_new_n6009__bF_buf0), .C(reset_n_bF_buf46), .Y(core__abc_21302_new_n6437_));
OAI21X1 OAI21X1_1571 ( .A(core__abc_21302_new_n5683_), .B(core__abc_21302_new_n5691_), .C(core__abc_21302_new_n5689_), .Y(core__abc_21302_new_n6440_));
OAI21X1 OAI21X1_1572 ( .A(core__abc_21302_new_n4978_), .B(core__abc_21302_new_n5999__bF_buf1), .C(core__abc_21302_new_n6009__bF_buf9), .Y(core__abc_21302_new_n6444_));
OAI21X1 OAI21X1_1573 ( .A(core_v1_reg_63_), .B(core__abc_21302_new_n6009__bF_buf8), .C(reset_n_bF_buf45), .Y(core__abc_21302_new_n6446_));
OAI21X1 OAI21X1_1574 ( .A(core__abc_21302_new_n1148_), .B(core__abc_21302_new_n1157_), .C(core__abc_21302_new_n2138_), .Y(core__abc_21302_new_n6448_));
OAI21X1 OAI21X1_1575 ( .A(core__abc_21302_new_n6449__bF_buf7), .B(core__abc_21302_new_n5084_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n6450_));
OAI21X1 OAI21X1_1576 ( .A(core__abc_21302_new_n2673__bF_buf11), .B(core__abc_21302_new_n2512_), .C(core__abc_21302_new_n6453_), .Y(core__abc_21302_new_n6454_));
OAI21X1 OAI21X1_1577 ( .A(core__abc_21302_new_n4822_), .B(core__abc_21302_new_n6454_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n6455_));
OAI21X1 OAI21X1_1578 ( .A(core__abc_21302_new_n6460_), .B(core__abc_21302_new_n6457_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n6461_));
OAI21X1 OAI21X1_1579 ( .A(core_key_2_), .B(core__abc_21302_new_n2640__bF_buf4), .C(core__abc_21302_new_n6467_), .Y(core__abc_21302_new_n6468_));
OAI21X1 OAI21X1_158 ( .A(core_siphash_word_18_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf25), .Y(_abc_19873_new_n1818_));
OAI21X1 OAI21X1_1580 ( .A(core__abc_21302_new_n6468_), .B(core__abc_21302_new_n6465_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n6469_));
OAI21X1 OAI21X1_1581 ( .A(core__abc_21302_new_n5131_), .B(core__abc_21302_new_n2640__bF_buf3), .C(core__abc_21302_new_n6474_), .Y(core__abc_21302_new_n6475_));
OAI21X1 OAI21X1_1582 ( .A(core__abc_21302_new_n6475_), .B(core__abc_21302_new_n2754_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n6476_));
OAI21X1 OAI21X1_1583 ( .A(core_key_4_), .B(core__abc_21302_new_n2640__bF_buf2), .C(core__abc_21302_new_n6480_), .Y(core__abc_21302_new_n6481_));
OAI21X1 OAI21X1_1584 ( .A(core__abc_21302_new_n6481_), .B(core__abc_21302_new_n6478_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n6482_));
OAI21X1 OAI21X1_1585 ( .A(core_key_5_), .B(core__abc_21302_new_n2640__bF_buf1), .C(core__abc_21302_new_n6487_), .Y(core__abc_21302_new_n6488_));
OAI21X1 OAI21X1_1586 ( .A(core__abc_21302_new_n6488_), .B(core__abc_21302_new_n6485_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n6489_));
OAI21X1 OAI21X1_1587 ( .A(core__abc_21302_new_n2673__bF_buf8), .B(core__abc_21302_new_n6492_), .C(core__abc_21302_new_n6494_), .Y(core__abc_21302_new_n6495_));
OAI21X1 OAI21X1_1588 ( .A(core__abc_21302_new_n5187_), .B(core__abc_21302_new_n6495_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n6496_));
OAI21X1 OAI21X1_1589 ( .A(core__abc_21302_new_n5221_), .B(core__abc_21302_new_n2640__bF_buf0), .C(core__abc_21302_new_n6501_), .Y(core__abc_21302_new_n6502_));
OAI21X1 OAI21X1_159 ( .A(core_siphash_word_19_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf24), .Y(_abc_19873_new_n1820_));
OAI21X1 OAI21X1_1590 ( .A(core__abc_21302_new_n6502_), .B(core__abc_21302_new_n6499_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n6503_));
OAI21X1 OAI21X1_1591 ( .A(core_key_8_), .B(core__abc_21302_new_n2640__bF_buf11), .C(core__abc_21302_new_n6508_), .Y(core__abc_21302_new_n6509_));
OAI21X1 OAI21X1_1592 ( .A(core__abc_21302_new_n6509_), .B(core__abc_21302_new_n6506_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n6510_));
OAI21X1 OAI21X1_1593 ( .A(core__abc_21302_new_n6514_), .B(core__abc_21302_new_n2640__bF_buf10), .C(core__abc_21302_new_n6516_), .Y(core__abc_21302_new_n6517_));
OAI21X1 OAI21X1_1594 ( .A(core__abc_21302_new_n6517_), .B(core__abc_21302_new_n6513_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n6518_));
OAI21X1 OAI21X1_1595 ( .A(core_key_10_), .B(core__abc_21302_new_n2640__bF_buf9), .C(core__abc_21302_new_n6523_), .Y(core__abc_21302_new_n6524_));
OAI21X1 OAI21X1_1596 ( .A(core__abc_21302_new_n6524_), .B(core__abc_21302_new_n6521_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n6525_));
OAI21X1 OAI21X1_1597 ( .A(core__abc_21302_new_n5297_), .B(core__abc_21302_new_n2640__bF_buf8), .C(core__abc_21302_new_n6530_), .Y(core__abc_21302_new_n6531_));
OAI21X1 OAI21X1_1598 ( .A(core__abc_21302_new_n6531_), .B(core__abc_21302_new_n6528_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n6532_));
OAI21X1 OAI21X1_1599 ( .A(core__abc_21302_new_n6536_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n6538_), .Y(core__abc_21302_new_n6539_));
OAI21X1 OAI21X1_16 ( .A(_abc_19873_new_n1147_), .B(_abc_19873_new_n960__bF_buf0), .C(_abc_19873_new_n1148_), .Y(_abc_19873_new_n1149_));
OAI21X1 OAI21X1_160 ( .A(core_siphash_word_20_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf23), .Y(_abc_19873_new_n1822_));
OAI21X1 OAI21X1_1600 ( .A(core__abc_21302_new_n6539_), .B(core__abc_21302_new_n6535_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n6540_));
OAI21X1 OAI21X1_1601 ( .A(core_key_13_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n6545_), .Y(core__abc_21302_new_n6546_));
OAI21X1 OAI21X1_1602 ( .A(core__abc_21302_new_n6546_), .B(core__abc_21302_new_n6543_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n6547_));
OAI21X1 OAI21X1_1603 ( .A(core_key_14_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n6552_), .Y(core__abc_21302_new_n6553_));
OAI21X1 OAI21X1_1604 ( .A(core__abc_21302_new_n6553_), .B(core__abc_21302_new_n6550_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n6554_));
OAI21X1 OAI21X1_1605 ( .A(core__abc_21302_new_n5382_), .B(core__abc_21302_new_n2640__bF_buf4), .C(core__abc_21302_new_n6559_), .Y(core__abc_21302_new_n6560_));
OAI21X1 OAI21X1_1606 ( .A(core__abc_21302_new_n6560_), .B(core__abc_21302_new_n6557_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n6561_));
OAI21X1 OAI21X1_1607 ( .A(core_key_16_), .B(core__abc_21302_new_n2640__bF_buf3), .C(core__abc_21302_new_n6566_), .Y(core__abc_21302_new_n6567_));
OAI21X1 OAI21X1_1608 ( .A(core__abc_21302_new_n6567_), .B(core__abc_21302_new_n6564_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n6568_));
OAI21X1 OAI21X1_1609 ( .A(core_key_17_), .B(core__abc_21302_new_n2640__bF_buf2), .C(core__abc_21302_new_n6573_), .Y(core__abc_21302_new_n6574_));
OAI21X1 OAI21X1_161 ( .A(core_siphash_word_21_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf22), .Y(_abc_19873_new_n1825_));
OAI21X1 OAI21X1_1610 ( .A(core__abc_21302_new_n6574_), .B(core__abc_21302_new_n6571_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n6575_));
OAI21X1 OAI21X1_1611 ( .A(core__abc_21302_new_n6579_), .B(core__abc_21302_new_n2640__bF_buf1), .C(core__abc_21302_new_n6581_), .Y(core__abc_21302_new_n6582_));
OAI21X1 OAI21X1_1612 ( .A(core__abc_21302_new_n6582_), .B(core__abc_21302_new_n6578_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n6583_));
OAI21X1 OAI21X1_1613 ( .A(core__abc_21302_new_n5460_), .B(core__abc_21302_new_n2640__bF_buf0), .C(core__abc_21302_new_n6588_), .Y(core__abc_21302_new_n6589_));
OAI21X1 OAI21X1_1614 ( .A(core__abc_21302_new_n6589_), .B(core__abc_21302_new_n6586_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n6590_));
OAI21X1 OAI21X1_1615 ( .A(core_key_20_), .B(core__abc_21302_new_n2640__bF_buf11), .C(core__abc_21302_new_n6595_), .Y(core__abc_21302_new_n6596_));
OAI21X1 OAI21X1_1616 ( .A(core__abc_21302_new_n6596_), .B(core__abc_21302_new_n6593_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n6597_));
OAI21X1 OAI21X1_1617 ( .A(core_key_21_), .B(core__abc_21302_new_n2640__bF_buf10), .C(core__abc_21302_new_n6602_), .Y(core__abc_21302_new_n6603_));
OAI21X1 OAI21X1_1618 ( .A(core__abc_21302_new_n6603_), .B(core__abc_21302_new_n6600_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n6604_));
OAI21X1 OAI21X1_1619 ( .A(core_key_22_), .B(core__abc_21302_new_n2640__bF_buf9), .C(core__abc_21302_new_n6609_), .Y(core__abc_21302_new_n6610_));
OAI21X1 OAI21X1_162 ( .A(core_siphash_word_22_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf21), .Y(_abc_19873_new_n1827_));
OAI21X1 OAI21X1_1620 ( .A(core__abc_21302_new_n6610_), .B(core__abc_21302_new_n6607_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n6611_));
OAI21X1 OAI21X1_1621 ( .A(core__abc_21302_new_n5540_), .B(core__abc_21302_new_n2640__bF_buf8), .C(core__abc_21302_new_n6616_), .Y(core__abc_21302_new_n6617_));
OAI21X1 OAI21X1_1622 ( .A(core__abc_21302_new_n6617_), .B(core__abc_21302_new_n6614_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n6618_));
OAI21X1 OAI21X1_1623 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n6623_), .C(core__abc_21302_new_n5564_), .Y(core__abc_21302_new_n6624_));
OAI21X1 OAI21X1_1624 ( .A(core__abc_21302_new_n6622_), .B(core__abc_21302_new_n6624_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n6625_));
OAI21X1 OAI21X1_1625 ( .A(core__abc_21302_new_n6629_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n6631_), .Y(core__abc_21302_new_n6632_));
OAI21X1 OAI21X1_1626 ( .A(core__abc_21302_new_n6632_), .B(core__abc_21302_new_n6628_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n6633_));
OAI21X1 OAI21X1_1627 ( .A(core__abc_21302_new_n6637_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n6639_), .Y(core__abc_21302_new_n6640_));
OAI21X1 OAI21X1_1628 ( .A(core__abc_21302_new_n6640_), .B(core__abc_21302_new_n6636_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n6641_));
OAI21X1 OAI21X1_1629 ( .A(core__abc_21302_new_n6645_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n6647_), .Y(core__abc_21302_new_n6648_));
OAI21X1 OAI21X1_163 ( .A(core_siphash_word_23_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf20), .Y(_abc_19873_new_n1829_));
OAI21X1 OAI21X1_1630 ( .A(core__abc_21302_new_n6648_), .B(core__abc_21302_new_n6644_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n6649_));
OAI21X1 OAI21X1_1631 ( .A(core_key_28_), .B(core__abc_21302_new_n2640__bF_buf4), .C(core__abc_21302_new_n6654_), .Y(core__abc_21302_new_n6655_));
OAI21X1 OAI21X1_1632 ( .A(core__abc_21302_new_n6655_), .B(core__abc_21302_new_n6652_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n6656_));
OAI21X1 OAI21X1_1633 ( .A(core_key_29_), .B(core__abc_21302_new_n2640__bF_buf3), .C(core__abc_21302_new_n6661_), .Y(core__abc_21302_new_n6662_));
OAI21X1 OAI21X1_1634 ( .A(core__abc_21302_new_n6662_), .B(core__abc_21302_new_n6659_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n6663_));
OAI21X1 OAI21X1_1635 ( .A(core_key_30_), .B(core__abc_21302_new_n2640__bF_buf2), .C(core__abc_21302_new_n6668_), .Y(core__abc_21302_new_n6669_));
OAI21X1 OAI21X1_1636 ( .A(core__abc_21302_new_n6669_), .B(core__abc_21302_new_n6666_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n6670_));
OAI21X1 OAI21X1_1637 ( .A(core__abc_21302_new_n5694_), .B(core__abc_21302_new_n2640__bF_buf1), .C(core__abc_21302_new_n6675_), .Y(core__abc_21302_new_n6676_));
OAI21X1 OAI21X1_1638 ( .A(core__abc_21302_new_n6676_), .B(core__abc_21302_new_n6673_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n6677_));
OAI21X1 OAI21X1_1639 ( .A(core__abc_21302_new_n2673__bF_buf4), .B(core__abc_21302_new_n3933_), .C(core__abc_21302_new_n6681_), .Y(core__abc_21302_new_n6682_));
OAI21X1 OAI21X1_164 ( .A(core_siphash_word_24_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf19), .Y(_abc_19873_new_n1831_));
OAI21X1 OAI21X1_1640 ( .A(core__abc_21302_new_n5699_), .B(core__abc_21302_new_n6682_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n6683_));
OAI21X1 OAI21X1_1641 ( .A(core__abc_21302_new_n2673__bF_buf3), .B(core__abc_21302_new_n3962_), .C(core__abc_21302_new_n6687_), .Y(core__abc_21302_new_n6688_));
OAI21X1 OAI21X1_1642 ( .A(core__abc_21302_new_n5707_), .B(core__abc_21302_new_n6688_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n6689_));
OAI21X1 OAI21X1_1643 ( .A(core_key_34_), .B(core__abc_21302_new_n2640__bF_buf0), .C(core__abc_21302_new_n6694_), .Y(core__abc_21302_new_n6695_));
OAI21X1 OAI21X1_1644 ( .A(core__abc_21302_new_n6695_), .B(core__abc_21302_new_n6692_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n6696_));
OAI21X1 OAI21X1_1645 ( .A(core__abc_21302_new_n5723_), .B(core__abc_21302_new_n2640__bF_buf11), .C(core__abc_21302_new_n6701_), .Y(core__abc_21302_new_n6702_));
OAI21X1 OAI21X1_1646 ( .A(core__abc_21302_new_n6702_), .B(core__abc_21302_new_n6699_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n6703_));
OAI21X1 OAI21X1_1647 ( .A(core__abc_21302_new_n6709_), .B(core__abc_21302_new_n6706_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n6710_));
OAI21X1 OAI21X1_1648 ( .A(core__abc_21302_new_n2673__bF_buf1), .B(core__abc_21302_new_n4083_), .C(core__abc_21302_new_n6714_), .Y(core__abc_21302_new_n6715_));
OAI21X1 OAI21X1_1649 ( .A(core__abc_21302_new_n5737_), .B(core__abc_21302_new_n6715_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n6716_));
OAI21X1 OAI21X1_165 ( .A(core_siphash_word_25_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf18), .Y(_abc_19873_new_n1833_));
OAI21X1 OAI21X1_1650 ( .A(core_key_38_), .B(core__abc_21302_new_n2640__bF_buf10), .C(core__abc_21302_new_n6721_), .Y(core__abc_21302_new_n6722_));
OAI21X1 OAI21X1_1651 ( .A(core__abc_21302_new_n6722_), .B(core__abc_21302_new_n6719_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n6723_));
OAI21X1 OAI21X1_1652 ( .A(core__abc_21302_new_n5758_), .B(core__abc_21302_new_n2640__bF_buf9), .C(core__abc_21302_new_n6728_), .Y(core__abc_21302_new_n6729_));
OAI21X1 OAI21X1_1653 ( .A(core__abc_21302_new_n6729_), .B(core__abc_21302_new_n6726_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n6730_));
OAI21X1 OAI21X1_1654 ( .A(core__abc_21302_new_n2673__bF_buf10), .B(core__abc_21302_new_n4184_), .C(core__abc_21302_new_n5767_), .Y(core__abc_21302_new_n6735_));
OAI21X1 OAI21X1_1655 ( .A(core__abc_21302_new_n6734_), .B(core__abc_21302_new_n6735_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n6736_));
OAI21X1 OAI21X1_1656 ( .A(core__abc_21302_new_n6740_), .B(core__abc_21302_new_n2640__bF_buf8), .C(core__abc_21302_new_n6742_), .Y(core__abc_21302_new_n6743_));
OAI21X1 OAI21X1_1657 ( .A(core__abc_21302_new_n6743_), .B(core__abc_21302_new_n6739_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n6744_));
OAI21X1 OAI21X1_1658 ( .A(core_key_42_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n6749_), .Y(core__abc_21302_new_n6750_));
OAI21X1 OAI21X1_1659 ( .A(core__abc_21302_new_n6750_), .B(core__abc_21302_new_n6747_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n6751_));
OAI21X1 OAI21X1_166 ( .A(core_siphash_word_26_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf17), .Y(_abc_19873_new_n1835_));
OAI21X1 OAI21X1_1660 ( .A(core_key_43_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n6756_), .Y(core__abc_21302_new_n6757_));
OAI21X1 OAI21X1_1661 ( .A(core__abc_21302_new_n6757_), .B(core__abc_21302_new_n6754_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n6758_));
OAI21X1 OAI21X1_1662 ( .A(core__abc_21302_new_n6764_), .B(core__abc_21302_new_n6761_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n6765_));
OAI21X1 OAI21X1_1663 ( .A(core__abc_21302_new_n2673__bF_buf7), .B(core__abc_21302_new_n6768_), .C(core__abc_21302_new_n6770_), .Y(core__abc_21302_new_n6771_));
OAI21X1 OAI21X1_1664 ( .A(core__abc_21302_new_n5811_), .B(core__abc_21302_new_n6771_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n6772_));
OAI21X1 OAI21X1_1665 ( .A(core_key_46_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n6777_), .Y(core__abc_21302_new_n6778_));
OAI21X1 OAI21X1_1666 ( .A(core__abc_21302_new_n6778_), .B(core__abc_21302_new_n6775_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n6779_));
OAI21X1 OAI21X1_1667 ( .A(core__abc_21302_new_n2673__bF_buf5), .B(core__abc_21302_new_n6782_), .C(core__abc_21302_new_n6784_), .Y(core__abc_21302_new_n6785_));
OAI21X1 OAI21X1_1668 ( .A(core__abc_21302_new_n5827_), .B(core__abc_21302_new_n6785_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n6786_));
OAI21X1 OAI21X1_1669 ( .A(core__abc_21302_new_n2673__bF_buf4), .B(core__abc_21302_new_n4404_), .C(core__abc_21302_new_n5844_), .Y(core__abc_21302_new_n6791_));
OAI21X1 OAI21X1_167 ( .A(core_siphash_word_27_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf16), .Y(_abc_19873_new_n1837_));
OAI21X1 OAI21X1_1670 ( .A(core__abc_21302_new_n6790_), .B(core__abc_21302_new_n6791_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n6792_));
OAI21X1 OAI21X1_1671 ( .A(core_key_49_), .B(core__abc_21302_new_n2640__bF_buf4), .C(core__abc_21302_new_n6797_), .Y(core__abc_21302_new_n6798_));
OAI21X1 OAI21X1_1672 ( .A(core__abc_21302_new_n6798_), .B(core__abc_21302_new_n6795_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n6799_));
OAI21X1 OAI21X1_1673 ( .A(core_key_50_), .B(core__abc_21302_new_n2640__bF_buf3), .C(core__abc_21302_new_n6804_), .Y(core__abc_21302_new_n6805_));
OAI21X1 OAI21X1_1674 ( .A(core__abc_21302_new_n6805_), .B(core__abc_21302_new_n6802_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n6806_));
OAI21X1 OAI21X1_1675 ( .A(core_key_51_), .B(core__abc_21302_new_n2640__bF_buf2), .C(core__abc_21302_new_n6811_), .Y(core__abc_21302_new_n6812_));
OAI21X1 OAI21X1_1676 ( .A(core__abc_21302_new_n6812_), .B(core__abc_21302_new_n6809_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n6813_));
OAI21X1 OAI21X1_1677 ( .A(core__abc_21302_new_n6817_), .B(core__abc_21302_new_n2640__bF_buf1), .C(core__abc_21302_new_n6819_), .Y(core__abc_21302_new_n6820_));
OAI21X1 OAI21X1_1678 ( .A(core__abc_21302_new_n6820_), .B(core__abc_21302_new_n6816_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n6821_));
OAI21X1 OAI21X1_1679 ( .A(core_key_53_), .B(core__abc_21302_new_n2640__bF_buf0), .C(core__abc_21302_new_n6826_), .Y(core__abc_21302_new_n6827_));
OAI21X1 OAI21X1_168 ( .A(core_siphash_word_28_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf15), .Y(_abc_19873_new_n1839_));
OAI21X1 OAI21X1_1680 ( .A(core__abc_21302_new_n6827_), .B(core__abc_21302_new_n6824_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n6828_));
OAI21X1 OAI21X1_1681 ( .A(core_key_54_), .B(core__abc_21302_new_n2640__bF_buf11), .C(core__abc_21302_new_n6833_), .Y(core__abc_21302_new_n6834_));
OAI21X1 OAI21X1_1682 ( .A(core__abc_21302_new_n6834_), .B(core__abc_21302_new_n6831_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n6835_));
OAI21X1 OAI21X1_1683 ( .A(core__abc_21302_new_n5915_), .B(core__abc_21302_new_n2640__bF_buf10), .C(core__abc_21302_new_n6840_), .Y(core__abc_21302_new_n6841_));
OAI21X1 OAI21X1_1684 ( .A(core__abc_21302_new_n6841_), .B(core__abc_21302_new_n6838_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n6842_));
OAI21X1 OAI21X1_1685 ( .A(core_key_56_), .B(core__abc_21302_new_n2640__bF_buf9), .C(core__abc_21302_new_n6847_), .Y(core__abc_21302_new_n6848_));
OAI21X1 OAI21X1_1686 ( .A(core__abc_21302_new_n6848_), .B(core__abc_21302_new_n6845_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n6849_));
OAI21X1 OAI21X1_1687 ( .A(core_key_57_), .B(core__abc_21302_new_n2640__bF_buf8), .C(core__abc_21302_new_n6855_), .Y(core__abc_21302_new_n6856_));
OAI21X1 OAI21X1_1688 ( .A(core__abc_21302_new_n6856_), .B(core__abc_21302_new_n6853_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n6857_));
OAI21X1 OAI21X1_1689 ( .A(core__abc_21302_new_n6861_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n6863_), .Y(core__abc_21302_new_n6864_));
OAI21X1 OAI21X1_169 ( .A(core_siphash_word_29_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf14), .Y(_abc_19873_new_n1841_));
OAI21X1 OAI21X1_1690 ( .A(core__abc_21302_new_n6864_), .B(core__abc_21302_new_n6860_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n6865_));
OAI21X1 OAI21X1_1691 ( .A(core__abc_21302_new_n6869_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n6871_), .Y(core__abc_21302_new_n6872_));
OAI21X1 OAI21X1_1692 ( .A(core__abc_21302_new_n6872_), .B(core__abc_21302_new_n6868_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n6873_));
OAI21X1 OAI21X1_1693 ( .A(core_key_60_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n6878_), .Y(core__abc_21302_new_n6879_));
OAI21X1 OAI21X1_1694 ( .A(core__abc_21302_new_n6879_), .B(core__abc_21302_new_n6876_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n6880_));
OAI21X1 OAI21X1_1695 ( .A(core_key_61_), .B(core__abc_21302_new_n2640__bF_buf4), .C(core__abc_21302_new_n6885_), .Y(core__abc_21302_new_n6886_));
OAI21X1 OAI21X1_1696 ( .A(core__abc_21302_new_n6886_), .B(core__abc_21302_new_n6883_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n6887_));
OAI21X1 OAI21X1_1697 ( .A(core_key_62_), .B(core__abc_21302_new_n2640__bF_buf3), .C(core__abc_21302_new_n6893_), .Y(core__abc_21302_new_n6894_));
OAI21X1 OAI21X1_1698 ( .A(core__abc_21302_new_n6894_), .B(core__abc_21302_new_n6891_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n6895_));
OAI21X1 OAI21X1_1699 ( .A(core__abc_21302_new_n5985_), .B(core__abc_21302_new_n2640__bF_buf2), .C(core__abc_21302_new_n6900_), .Y(core__abc_21302_new_n6901_));
OAI21X1 OAI21X1_17 ( .A(_abc_19873_new_n905__bF_buf2), .B(_abc_19873_new_n893__bF_buf1), .C(_abc_19873_new_n877_), .Y(_abc_19873_new_n1159_));
OAI21X1 OAI21X1_170 ( .A(core_siphash_word_30_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf13), .Y(_abc_19873_new_n1843_));
OAI21X1 OAI21X1_1700 ( .A(core__abc_21302_new_n6901_), .B(core__abc_21302_new_n6898_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n6902_));
OAI21X1 OAI21X1_1701 ( .A(core__abc_21302_new_n1147_), .B(core__abc_21302_new_n2166_), .C(core_siphash_valid_reg), .Y(core__abc_21302_new_n6912_));
OAI21X1 OAI21X1_171 ( .A(core_siphash_word_31_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf12), .Y(_abc_19873_new_n1845_));
OAI21X1 OAI21X1_172 ( .A(\write_data[0] ), .B(_abc_19873_new_n1849__bF_buf7), .C(reset_n_bF_buf11), .Y(_abc_19873_new_n1850_));
OAI21X1 OAI21X1_173 ( .A(\write_data[1] ), .B(_abc_19873_new_n1849__bF_buf5), .C(reset_n_bF_buf10), .Y(_abc_19873_new_n1853_));
OAI21X1 OAI21X1_174 ( .A(\write_data[2] ), .B(_abc_19873_new_n1849__bF_buf3), .C(reset_n_bF_buf9), .Y(_abc_19873_new_n1855_));
OAI21X1 OAI21X1_175 ( .A(\write_data[3] ), .B(_abc_19873_new_n1849__bF_buf1), .C(reset_n_bF_buf8), .Y(_abc_19873_new_n1857_));
OAI21X1 OAI21X1_176 ( .A(\write_data[4] ), .B(_abc_19873_new_n1849__bF_buf7), .C(reset_n_bF_buf7), .Y(_abc_19873_new_n1859_));
OAI21X1 OAI21X1_177 ( .A(\write_data[5] ), .B(_abc_19873_new_n1849__bF_buf5), .C(reset_n_bF_buf6), .Y(_abc_19873_new_n1862_));
OAI21X1 OAI21X1_178 ( .A(\write_data[6] ), .B(_abc_19873_new_n1849__bF_buf3), .C(reset_n_bF_buf5), .Y(_abc_19873_new_n1864_));
OAI21X1 OAI21X1_179 ( .A(\write_data[7] ), .B(_abc_19873_new_n1849__bF_buf1), .C(reset_n_bF_buf4), .Y(_abc_19873_new_n1866_));
OAI21X1 OAI21X1_18 ( .A(_abc_19873_new_n1158_), .B(_abc_19873_new_n894__bF_buf4), .C(_abc_19873_new_n1159_), .Y(_abc_19873_new_n1160_));
OAI21X1 OAI21X1_180 ( .A(\write_data[8] ), .B(_abc_19873_new_n1849__bF_buf7), .C(reset_n_bF_buf3), .Y(_abc_19873_new_n1868_));
OAI21X1 OAI21X1_181 ( .A(\write_data[9] ), .B(_abc_19873_new_n1849__bF_buf5), .C(reset_n_bF_buf2), .Y(_abc_19873_new_n1870_));
OAI21X1 OAI21X1_182 ( .A(\write_data[10] ), .B(_abc_19873_new_n1849__bF_buf3), .C(reset_n_bF_buf1), .Y(_abc_19873_new_n1872_));
OAI21X1 OAI21X1_183 ( .A(\write_data[11] ), .B(_abc_19873_new_n1849__bF_buf1), .C(reset_n_bF_buf0), .Y(_abc_19873_new_n1874_));
OAI21X1 OAI21X1_184 ( .A(\write_data[12] ), .B(_abc_19873_new_n1849__bF_buf7), .C(reset_n_bF_buf69), .Y(_abc_19873_new_n1876_));
OAI21X1 OAI21X1_185 ( .A(\write_data[13] ), .B(_abc_19873_new_n1849__bF_buf5), .C(reset_n_bF_buf68), .Y(_abc_19873_new_n1878_));
OAI21X1 OAI21X1_186 ( .A(\write_data[14] ), .B(_abc_19873_new_n1849__bF_buf3), .C(reset_n_bF_buf67), .Y(_abc_19873_new_n1881_));
OAI21X1 OAI21X1_187 ( .A(\write_data[15] ), .B(_abc_19873_new_n1849__bF_buf1), .C(reset_n_bF_buf66), .Y(_abc_19873_new_n1883_));
OAI21X1 OAI21X1_188 ( .A(\write_data[16] ), .B(_abc_19873_new_n1849__bF_buf7), .C(reset_n_bF_buf65), .Y(_abc_19873_new_n1886_));
OAI21X1 OAI21X1_189 ( .A(\write_data[17] ), .B(_abc_19873_new_n1849__bF_buf5), .C(reset_n_bF_buf64), .Y(_abc_19873_new_n1888_));
OAI21X1 OAI21X1_19 ( .A(_abc_19873_new_n1166_), .B(_abc_19873_new_n960__bF_buf4), .C(_abc_19873_new_n1167_), .Y(_abc_19873_new_n1168_));
OAI21X1 OAI21X1_190 ( .A(\write_data[18] ), .B(_abc_19873_new_n1849__bF_buf3), .C(reset_n_bF_buf63), .Y(_abc_19873_new_n1890_));
OAI21X1 OAI21X1_191 ( .A(\write_data[19] ), .B(_abc_19873_new_n1849__bF_buf1), .C(reset_n_bF_buf62), .Y(_abc_19873_new_n1893_));
OAI21X1 OAI21X1_192 ( .A(\write_data[20] ), .B(_abc_19873_new_n1849__bF_buf7), .C(reset_n_bF_buf61), .Y(_abc_19873_new_n1895_));
OAI21X1 OAI21X1_193 ( .A(\write_data[21] ), .B(_abc_19873_new_n1849__bF_buf5), .C(reset_n_bF_buf60), .Y(_abc_19873_new_n1897_));
OAI21X1 OAI21X1_194 ( .A(\write_data[22] ), .B(_abc_19873_new_n1849__bF_buf3), .C(reset_n_bF_buf59), .Y(_abc_19873_new_n1900_));
OAI21X1 OAI21X1_195 ( .A(\write_data[23] ), .B(_abc_19873_new_n1849__bF_buf1), .C(reset_n_bF_buf58), .Y(_abc_19873_new_n1902_));
OAI21X1 OAI21X1_196 ( .A(\write_data[24] ), .B(_abc_19873_new_n1849__bF_buf7), .C(reset_n_bF_buf57), .Y(_abc_19873_new_n1905_));
OAI21X1 OAI21X1_197 ( .A(\write_data[25] ), .B(_abc_19873_new_n1849__bF_buf5), .C(reset_n_bF_buf56), .Y(_abc_19873_new_n1908_));
OAI21X1 OAI21X1_198 ( .A(\write_data[26] ), .B(_abc_19873_new_n1849__bF_buf3), .C(reset_n_bF_buf55), .Y(_abc_19873_new_n1910_));
OAI21X1 OAI21X1_199 ( .A(\write_data[27] ), .B(_abc_19873_new_n1849__bF_buf1), .C(reset_n_bF_buf54), .Y(_abc_19873_new_n1912_));
OAI21X1 OAI21X1_2 ( .A(_abc_19873_new_n916_), .B(_abc_19873_new_n918_), .C(_abc_19873_new_n919_), .Y(_abc_19873_new_n920_));
OAI21X1 OAI21X1_20 ( .A(_abc_19873_new_n1195_), .B(_abc_19873_new_n894__bF_buf2), .C(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1196_));
OAI21X1 OAI21X1_200 ( .A(\write_data[28] ), .B(_abc_19873_new_n1849__bF_buf7), .C(reset_n_bF_buf53), .Y(_abc_19873_new_n1915_));
OAI21X1 OAI21X1_201 ( .A(\write_data[29] ), .B(_abc_19873_new_n1849__bF_buf5), .C(reset_n_bF_buf52), .Y(_abc_19873_new_n1918_));
OAI21X1 OAI21X1_202 ( .A(\write_data[30] ), .B(_abc_19873_new_n1849__bF_buf3), .C(reset_n_bF_buf51), .Y(_abc_19873_new_n1921_));
OAI21X1 OAI21X1_203 ( .A(\write_data[31] ), .B(_abc_19873_new_n1849__bF_buf1), .C(reset_n_bF_buf50), .Y(_abc_19873_new_n1923_));
OAI21X1 OAI21X1_204 ( .A(\write_data[0] ), .B(_abc_19873_new_n1925__bF_buf7), .C(reset_n_bF_buf49), .Y(_abc_19873_new_n1926_));
OAI21X1 OAI21X1_205 ( .A(\write_data[1] ), .B(_abc_19873_new_n1925__bF_buf5), .C(reset_n_bF_buf48), .Y(_abc_19873_new_n1928_));
OAI21X1 OAI21X1_206 ( .A(\write_data[2] ), .B(_abc_19873_new_n1925__bF_buf3), .C(reset_n_bF_buf47), .Y(_abc_19873_new_n1930_));
OAI21X1 OAI21X1_207 ( .A(\write_data[3] ), .B(_abc_19873_new_n1925__bF_buf1), .C(reset_n_bF_buf46), .Y(_abc_19873_new_n1932_));
OAI21X1 OAI21X1_208 ( .A(\write_data[4] ), .B(_abc_19873_new_n1925__bF_buf7), .C(reset_n_bF_buf45), .Y(_abc_19873_new_n1934_));
OAI21X1 OAI21X1_209 ( .A(\write_data[5] ), .B(_abc_19873_new_n1925__bF_buf5), .C(reset_n_bF_buf44), .Y(_abc_19873_new_n1936_));
OAI21X1 OAI21X1_21 ( .A(_abc_19873_new_n1198_), .B(_abc_19873_new_n1064__bF_buf1), .C(_abc_19873_new_n1199_), .Y(_abc_19873_new_n1200_));
OAI21X1 OAI21X1_210 ( .A(\write_data[6] ), .B(_abc_19873_new_n1925__bF_buf3), .C(reset_n_bF_buf43), .Y(_abc_19873_new_n1938_));
OAI21X1 OAI21X1_211 ( .A(\write_data[7] ), .B(_abc_19873_new_n1925__bF_buf1), .C(reset_n_bF_buf42), .Y(_abc_19873_new_n1940_));
OAI21X1 OAI21X1_212 ( .A(\write_data[8] ), .B(_abc_19873_new_n1925__bF_buf7), .C(reset_n_bF_buf41), .Y(_abc_19873_new_n1942_));
OAI21X1 OAI21X1_213 ( .A(\write_data[9] ), .B(_abc_19873_new_n1925__bF_buf5), .C(reset_n_bF_buf40), .Y(_abc_19873_new_n1944_));
OAI21X1 OAI21X1_214 ( .A(\write_data[10] ), .B(_abc_19873_new_n1925__bF_buf3), .C(reset_n_bF_buf39), .Y(_abc_19873_new_n1946_));
OAI21X1 OAI21X1_215 ( .A(\write_data[11] ), .B(_abc_19873_new_n1925__bF_buf1), .C(reset_n_bF_buf38), .Y(_abc_19873_new_n1948_));
OAI21X1 OAI21X1_216 ( .A(\write_data[12] ), .B(_abc_19873_new_n1925__bF_buf7), .C(reset_n_bF_buf37), .Y(_abc_19873_new_n1950_));
OAI21X1 OAI21X1_217 ( .A(\write_data[13] ), .B(_abc_19873_new_n1925__bF_buf5), .C(reset_n_bF_buf36), .Y(_abc_19873_new_n1952_));
OAI21X1 OAI21X1_218 ( .A(\write_data[14] ), .B(_abc_19873_new_n1925__bF_buf3), .C(reset_n_bF_buf35), .Y(_abc_19873_new_n1954_));
OAI21X1 OAI21X1_219 ( .A(\write_data[15] ), .B(_abc_19873_new_n1925__bF_buf1), .C(reset_n_bF_buf34), .Y(_abc_19873_new_n1956_));
OAI21X1 OAI21X1_22 ( .A(_abc_19873_new_n1232_), .B(_abc_19873_new_n894__bF_buf0), .C(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1233_));
OAI21X1 OAI21X1_220 ( .A(\write_data[16] ), .B(_abc_19873_new_n1925__bF_buf7), .C(reset_n_bF_buf33), .Y(_abc_19873_new_n1958_));
OAI21X1 OAI21X1_221 ( .A(\write_data[17] ), .B(_abc_19873_new_n1925__bF_buf5), .C(reset_n_bF_buf32), .Y(_abc_19873_new_n1961_));
OAI21X1 OAI21X1_222 ( .A(\write_data[18] ), .B(_abc_19873_new_n1925__bF_buf3), .C(reset_n_bF_buf31), .Y(_abc_19873_new_n1963_));
OAI21X1 OAI21X1_223 ( .A(\write_data[19] ), .B(_abc_19873_new_n1925__bF_buf1), .C(reset_n_bF_buf30), .Y(_abc_19873_new_n1965_));
OAI21X1 OAI21X1_224 ( .A(\write_data[20] ), .B(_abc_19873_new_n1925__bF_buf7), .C(reset_n_bF_buf29), .Y(_abc_19873_new_n1967_));
OAI21X1 OAI21X1_225 ( .A(\write_data[21] ), .B(_abc_19873_new_n1925__bF_buf5), .C(reset_n_bF_buf28), .Y(_abc_19873_new_n1969_));
OAI21X1 OAI21X1_226 ( .A(\write_data[22] ), .B(_abc_19873_new_n1925__bF_buf3), .C(reset_n_bF_buf27), .Y(_abc_19873_new_n1971_));
OAI21X1 OAI21X1_227 ( .A(\write_data[23] ), .B(_abc_19873_new_n1925__bF_buf1), .C(reset_n_bF_buf26), .Y(_abc_19873_new_n1973_));
OAI21X1 OAI21X1_228 ( .A(\write_data[24] ), .B(_abc_19873_new_n1925__bF_buf7), .C(reset_n_bF_buf25), .Y(_abc_19873_new_n1975_));
OAI21X1 OAI21X1_229 ( .A(\write_data[25] ), .B(_abc_19873_new_n1925__bF_buf5), .C(reset_n_bF_buf24), .Y(_abc_19873_new_n1977_));
OAI21X1 OAI21X1_23 ( .A(_abc_19873_new_n1235_), .B(_abc_19873_new_n1064__bF_buf3), .C(_abc_19873_new_n1236_), .Y(_abc_19873_new_n1237_));
OAI21X1 OAI21X1_230 ( .A(\write_data[26] ), .B(_abc_19873_new_n1925__bF_buf3), .C(reset_n_bF_buf23), .Y(_abc_19873_new_n1979_));
OAI21X1 OAI21X1_231 ( .A(\write_data[27] ), .B(_abc_19873_new_n1925__bF_buf1), .C(reset_n_bF_buf22), .Y(_abc_19873_new_n1981_));
OAI21X1 OAI21X1_232 ( .A(\write_data[28] ), .B(_abc_19873_new_n1925__bF_buf7), .C(reset_n_bF_buf21), .Y(_abc_19873_new_n1983_));
OAI21X1 OAI21X1_233 ( .A(\write_data[29] ), .B(_abc_19873_new_n1925__bF_buf5), .C(reset_n_bF_buf20), .Y(_abc_19873_new_n1986_));
OAI21X1 OAI21X1_234 ( .A(\write_data[30] ), .B(_abc_19873_new_n1925__bF_buf3), .C(reset_n_bF_buf19), .Y(_abc_19873_new_n1988_));
OAI21X1 OAI21X1_235 ( .A(\write_data[31] ), .B(_abc_19873_new_n1925__bF_buf1), .C(reset_n_bF_buf18), .Y(_abc_19873_new_n1990_));
OAI21X1 OAI21X1_236 ( .A(\write_data[0] ), .B(_abc_19873_new_n1992__bF_buf7), .C(reset_n_bF_buf17), .Y(_abc_19873_new_n1993_));
OAI21X1 OAI21X1_237 ( .A(\write_data[1] ), .B(_abc_19873_new_n1992__bF_buf5), .C(reset_n_bF_buf16), .Y(_abc_19873_new_n1995_));
OAI21X1 OAI21X1_238 ( .A(\write_data[2] ), .B(_abc_19873_new_n1992__bF_buf3), .C(reset_n_bF_buf15), .Y(_abc_19873_new_n1997_));
OAI21X1 OAI21X1_239 ( .A(\write_data[3] ), .B(_abc_19873_new_n1992__bF_buf1), .C(reset_n_bF_buf14), .Y(_abc_19873_new_n1999_));
OAI21X1 OAI21X1_24 ( .A(_abc_19873_new_n895__bF_buf0), .B(_abc_19873_new_n893__bF_buf2), .C(_abc_19873_new_n877_), .Y(_abc_19873_new_n1248_));
OAI21X1 OAI21X1_240 ( .A(\write_data[4] ), .B(_abc_19873_new_n1992__bF_buf7), .C(reset_n_bF_buf13), .Y(_abc_19873_new_n2001_));
OAI21X1 OAI21X1_241 ( .A(\write_data[5] ), .B(_abc_19873_new_n1992__bF_buf5), .C(reset_n_bF_buf12), .Y(_abc_19873_new_n2003_));
OAI21X1 OAI21X1_242 ( .A(\write_data[6] ), .B(_abc_19873_new_n1992__bF_buf3), .C(reset_n_bF_buf11), .Y(_abc_19873_new_n2005_));
OAI21X1 OAI21X1_243 ( .A(\write_data[7] ), .B(_abc_19873_new_n1992__bF_buf1), .C(reset_n_bF_buf10), .Y(_abc_19873_new_n2007_));
OAI21X1 OAI21X1_244 ( .A(\write_data[8] ), .B(_abc_19873_new_n1992__bF_buf7), .C(reset_n_bF_buf9), .Y(_abc_19873_new_n2009_));
OAI21X1 OAI21X1_245 ( .A(\write_data[9] ), .B(_abc_19873_new_n1992__bF_buf5), .C(reset_n_bF_buf8), .Y(_abc_19873_new_n2011_));
OAI21X1 OAI21X1_246 ( .A(\write_data[10] ), .B(_abc_19873_new_n1992__bF_buf3), .C(reset_n_bF_buf7), .Y(_abc_19873_new_n2013_));
OAI21X1 OAI21X1_247 ( .A(\write_data[11] ), .B(_abc_19873_new_n1992__bF_buf1), .C(reset_n_bF_buf6), .Y(_abc_19873_new_n2015_));
OAI21X1 OAI21X1_248 ( .A(\write_data[12] ), .B(_abc_19873_new_n1992__bF_buf7), .C(reset_n_bF_buf5), .Y(_abc_19873_new_n2017_));
OAI21X1 OAI21X1_249 ( .A(\write_data[13] ), .B(_abc_19873_new_n1992__bF_buf5), .C(reset_n_bF_buf4), .Y(_abc_19873_new_n2019_));
OAI21X1 OAI21X1_25 ( .A(_abc_19873_new_n1247_), .B(_abc_19873_new_n960__bF_buf4), .C(_abc_19873_new_n1248_), .Y(_abc_19873_new_n1249_));
OAI21X1 OAI21X1_250 ( .A(\write_data[14] ), .B(_abc_19873_new_n1992__bF_buf3), .C(reset_n_bF_buf3), .Y(_abc_19873_new_n2021_));
OAI21X1 OAI21X1_251 ( .A(\write_data[15] ), .B(_abc_19873_new_n1992__bF_buf1), .C(reset_n_bF_buf2), .Y(_abc_19873_new_n2023_));
OAI21X1 OAI21X1_252 ( .A(\write_data[16] ), .B(_abc_19873_new_n1992__bF_buf7), .C(reset_n_bF_buf1), .Y(_abc_19873_new_n2025_));
OAI21X1 OAI21X1_253 ( .A(\write_data[17] ), .B(_abc_19873_new_n1992__bF_buf5), .C(reset_n_bF_buf0), .Y(_abc_19873_new_n2027_));
OAI21X1 OAI21X1_254 ( .A(\write_data[18] ), .B(_abc_19873_new_n1992__bF_buf3), .C(reset_n_bF_buf69), .Y(_abc_19873_new_n2029_));
OAI21X1 OAI21X1_255 ( .A(\write_data[19] ), .B(_abc_19873_new_n1992__bF_buf1), .C(reset_n_bF_buf68), .Y(_abc_19873_new_n2031_));
OAI21X1 OAI21X1_256 ( .A(\write_data[20] ), .B(_abc_19873_new_n1992__bF_buf7), .C(reset_n_bF_buf67), .Y(_abc_19873_new_n2033_));
OAI21X1 OAI21X1_257 ( .A(\write_data[21] ), .B(_abc_19873_new_n1992__bF_buf5), .C(reset_n_bF_buf66), .Y(_abc_19873_new_n2035_));
OAI21X1 OAI21X1_258 ( .A(\write_data[22] ), .B(_abc_19873_new_n1992__bF_buf3), .C(reset_n_bF_buf65), .Y(_abc_19873_new_n2037_));
OAI21X1 OAI21X1_259 ( .A(\write_data[23] ), .B(_abc_19873_new_n1992__bF_buf1), .C(reset_n_bF_buf64), .Y(_abc_19873_new_n2039_));
OAI21X1 OAI21X1_26 ( .A(_abc_19873_new_n1261_), .B(_abc_19873_new_n913__bF_buf2), .C(_abc_19873_new_n1262_), .Y(_abc_19873_new_n1263_));
OAI21X1 OAI21X1_260 ( .A(\write_data[24] ), .B(_abc_19873_new_n1992__bF_buf7), .C(reset_n_bF_buf63), .Y(_abc_19873_new_n2041_));
OAI21X1 OAI21X1_261 ( .A(\write_data[25] ), .B(_abc_19873_new_n1992__bF_buf5), .C(reset_n_bF_buf62), .Y(_abc_19873_new_n2043_));
OAI21X1 OAI21X1_262 ( .A(\write_data[26] ), .B(_abc_19873_new_n1992__bF_buf3), .C(reset_n_bF_buf61), .Y(_abc_19873_new_n2045_));
OAI21X1 OAI21X1_263 ( .A(\write_data[27] ), .B(_abc_19873_new_n1992__bF_buf1), .C(reset_n_bF_buf60), .Y(_abc_19873_new_n2047_));
OAI21X1 OAI21X1_264 ( .A(\write_data[28] ), .B(_abc_19873_new_n1992__bF_buf7), .C(reset_n_bF_buf59), .Y(_abc_19873_new_n2049_));
OAI21X1 OAI21X1_265 ( .A(\write_data[29] ), .B(_abc_19873_new_n1992__bF_buf5), .C(reset_n_bF_buf58), .Y(_abc_19873_new_n2052_));
OAI21X1 OAI21X1_266 ( .A(\write_data[30] ), .B(_abc_19873_new_n1992__bF_buf3), .C(reset_n_bF_buf57), .Y(_abc_19873_new_n2054_));
OAI21X1 OAI21X1_267 ( .A(\write_data[31] ), .B(_abc_19873_new_n1992__bF_buf1), .C(reset_n_bF_buf56), .Y(_abc_19873_new_n2056_));
OAI21X1 OAI21X1_268 ( .A(\write_data[0] ), .B(_abc_19873_new_n2058__bF_buf7), .C(reset_n_bF_buf55), .Y(_abc_19873_new_n2059_));
OAI21X1 OAI21X1_269 ( .A(\write_data[1] ), .B(_abc_19873_new_n2058__bF_buf5), .C(reset_n_bF_buf54), .Y(_abc_19873_new_n2061_));
OAI21X1 OAI21X1_27 ( .A(_abc_19873_new_n1269_), .B(_abc_19873_new_n894__bF_buf3), .C(_abc_19873_new_n1003_), .Y(_abc_19873_new_n1270_));
OAI21X1 OAI21X1_270 ( .A(\write_data[2] ), .B(_abc_19873_new_n2058__bF_buf3), .C(reset_n_bF_buf53), .Y(_abc_19873_new_n2063_));
OAI21X1 OAI21X1_271 ( .A(\write_data[3] ), .B(_abc_19873_new_n2058__bF_buf1), .C(reset_n_bF_buf52), .Y(_abc_19873_new_n2065_));
OAI21X1 OAI21X1_272 ( .A(\write_data[4] ), .B(_abc_19873_new_n2058__bF_buf7), .C(reset_n_bF_buf51), .Y(_abc_19873_new_n2067_));
OAI21X1 OAI21X1_273 ( .A(\write_data[5] ), .B(_abc_19873_new_n2058__bF_buf5), .C(reset_n_bF_buf50), .Y(_abc_19873_new_n2069_));
OAI21X1 OAI21X1_274 ( .A(\write_data[6] ), .B(_abc_19873_new_n2058__bF_buf3), .C(reset_n_bF_buf49), .Y(_abc_19873_new_n2072_));
OAI21X1 OAI21X1_275 ( .A(\write_data[7] ), .B(_abc_19873_new_n2058__bF_buf1), .C(reset_n_bF_buf48), .Y(_abc_19873_new_n2075_));
OAI21X1 OAI21X1_276 ( .A(\write_data[8] ), .B(_abc_19873_new_n2058__bF_buf7), .C(reset_n_bF_buf47), .Y(_abc_19873_new_n2077_));
OAI21X1 OAI21X1_277 ( .A(\write_data[9] ), .B(_abc_19873_new_n2058__bF_buf5), .C(reset_n_bF_buf46), .Y(_abc_19873_new_n2079_));
OAI21X1 OAI21X1_278 ( .A(\write_data[10] ), .B(_abc_19873_new_n2058__bF_buf3), .C(reset_n_bF_buf45), .Y(_abc_19873_new_n2081_));
OAI21X1 OAI21X1_279 ( .A(\write_data[11] ), .B(_abc_19873_new_n2058__bF_buf1), .C(reset_n_bF_buf44), .Y(_abc_19873_new_n2083_));
OAI21X1 OAI21X1_28 ( .A(_abc_19873_new_n1276_), .B(_abc_19873_new_n960__bF_buf3), .C(_abc_19873_new_n1277_), .Y(_abc_19873_new_n1278_));
OAI21X1 OAI21X1_280 ( .A(\write_data[12] ), .B(_abc_19873_new_n2058__bF_buf7), .C(reset_n_bF_buf43), .Y(_abc_19873_new_n2085_));
OAI21X1 OAI21X1_281 ( .A(\write_data[13] ), .B(_abc_19873_new_n2058__bF_buf5), .C(reset_n_bF_buf42), .Y(_abc_19873_new_n2087_));
OAI21X1 OAI21X1_282 ( .A(\write_data[14] ), .B(_abc_19873_new_n2058__bF_buf3), .C(reset_n_bF_buf41), .Y(_abc_19873_new_n2089_));
OAI21X1 OAI21X1_283 ( .A(\write_data[15] ), .B(_abc_19873_new_n2058__bF_buf1), .C(reset_n_bF_buf40), .Y(_abc_19873_new_n2091_));
OAI21X1 OAI21X1_284 ( .A(\write_data[16] ), .B(_abc_19873_new_n2058__bF_buf7), .C(reset_n_bF_buf39), .Y(_abc_19873_new_n2093_));
OAI21X1 OAI21X1_285 ( .A(\write_data[17] ), .B(_abc_19873_new_n2058__bF_buf5), .C(reset_n_bF_buf38), .Y(_abc_19873_new_n2095_));
OAI21X1 OAI21X1_286 ( .A(\write_data[18] ), .B(_abc_19873_new_n2058__bF_buf3), .C(reset_n_bF_buf37), .Y(_abc_19873_new_n2097_));
OAI21X1 OAI21X1_287 ( .A(\write_data[19] ), .B(_abc_19873_new_n2058__bF_buf1), .C(reset_n_bF_buf36), .Y(_abc_19873_new_n2099_));
OAI21X1 OAI21X1_288 ( .A(\write_data[20] ), .B(_abc_19873_new_n2058__bF_buf7), .C(reset_n_bF_buf35), .Y(_abc_19873_new_n2101_));
OAI21X1 OAI21X1_289 ( .A(\write_data[21] ), .B(_abc_19873_new_n2058__bF_buf5), .C(reset_n_bF_buf34), .Y(_abc_19873_new_n2103_));
OAI21X1 OAI21X1_29 ( .A(_abc_19873_new_n1287_), .B(_abc_19873_new_n894__bF_buf2), .C(_abc_19873_new_n1159_), .Y(_abc_19873_new_n1288_));
OAI21X1 OAI21X1_290 ( .A(\write_data[22] ), .B(_abc_19873_new_n2058__bF_buf3), .C(reset_n_bF_buf33), .Y(_abc_19873_new_n2105_));
OAI21X1 OAI21X1_291 ( .A(\write_data[23] ), .B(_abc_19873_new_n2058__bF_buf1), .C(reset_n_bF_buf32), .Y(_abc_19873_new_n2107_));
OAI21X1 OAI21X1_292 ( .A(\write_data[24] ), .B(_abc_19873_new_n2058__bF_buf7), .C(reset_n_bF_buf31), .Y(_abc_19873_new_n2109_));
OAI21X1 OAI21X1_293 ( .A(\write_data[25] ), .B(_abc_19873_new_n2058__bF_buf5), .C(reset_n_bF_buf30), .Y(_abc_19873_new_n2111_));
OAI21X1 OAI21X1_294 ( .A(\write_data[26] ), .B(_abc_19873_new_n2058__bF_buf3), .C(reset_n_bF_buf29), .Y(_abc_19873_new_n2113_));
OAI21X1 OAI21X1_295 ( .A(\write_data[27] ), .B(_abc_19873_new_n2058__bF_buf1), .C(reset_n_bF_buf28), .Y(_abc_19873_new_n2115_));
OAI21X1 OAI21X1_296 ( .A(\write_data[28] ), .B(_abc_19873_new_n2058__bF_buf7), .C(reset_n_bF_buf27), .Y(_abc_19873_new_n2117_));
OAI21X1 OAI21X1_297 ( .A(\write_data[29] ), .B(_abc_19873_new_n2058__bF_buf5), .C(reset_n_bF_buf26), .Y(_abc_19873_new_n2119_));
OAI21X1 OAI21X1_298 ( .A(\write_data[30] ), .B(_abc_19873_new_n2058__bF_buf3), .C(reset_n_bF_buf25), .Y(_abc_19873_new_n2121_));
OAI21X1 OAI21X1_299 ( .A(\write_data[31] ), .B(_abc_19873_new_n2058__bF_buf1), .C(reset_n_bF_buf24), .Y(_abc_19873_new_n2123_));
OAI21X1 OAI21X1_3 ( .A(_abc_19873_new_n930_), .B(_abc_19873_new_n878_), .C(_abc_19873_new_n931_), .Y(_abc_19873_new_n932_));
OAI21X1 OAI21X1_30 ( .A(_abc_19873_new_n1290_), .B(_abc_19873_new_n1064__bF_buf0), .C(_abc_19873_new_n1291_), .Y(_abc_19873_new_n1292_));
OAI21X1 OAI21X1_300 ( .A(\write_data[0] ), .B(_abc_19873_new_n2125__bF_buf7), .C(reset_n_bF_buf23), .Y(_abc_19873_new_n2126_));
OAI21X1 OAI21X1_301 ( .A(\write_data[1] ), .B(_abc_19873_new_n2125__bF_buf5), .C(reset_n_bF_buf22), .Y(_abc_19873_new_n2128_));
OAI21X1 OAI21X1_302 ( .A(\write_data[2] ), .B(_abc_19873_new_n2125__bF_buf3), .C(reset_n_bF_buf21), .Y(_abc_19873_new_n2130_));
OAI21X1 OAI21X1_303 ( .A(\write_data[3] ), .B(_abc_19873_new_n2125__bF_buf1), .C(reset_n_bF_buf20), .Y(_abc_19873_new_n2133_));
OAI21X1 OAI21X1_304 ( .A(\write_data[4] ), .B(_abc_19873_new_n2125__bF_buf7), .C(reset_n_bF_buf19), .Y(_abc_19873_new_n2136_));
OAI21X1 OAI21X1_305 ( .A(\write_data[5] ), .B(_abc_19873_new_n2125__bF_buf5), .C(reset_n_bF_buf18), .Y(_abc_19873_new_n2139_));
OAI21X1 OAI21X1_306 ( .A(\write_data[6] ), .B(_abc_19873_new_n2125__bF_buf3), .C(reset_n_bF_buf17), .Y(_abc_19873_new_n2141_));
OAI21X1 OAI21X1_307 ( .A(\write_data[7] ), .B(_abc_19873_new_n2125__bF_buf1), .C(reset_n_bF_buf16), .Y(_abc_19873_new_n2143_));
OAI21X1 OAI21X1_308 ( .A(\write_data[8] ), .B(_abc_19873_new_n2125__bF_buf7), .C(reset_n_bF_buf15), .Y(_abc_19873_new_n2145_));
OAI21X1 OAI21X1_309 ( .A(\write_data[9] ), .B(_abc_19873_new_n2125__bF_buf5), .C(reset_n_bF_buf14), .Y(_abc_19873_new_n2147_));
OAI21X1 OAI21X1_31 ( .A(_abc_19873_new_n1305_), .B(_abc_19873_new_n894__bF_buf1), .C(_abc_19873_new_n1140_), .Y(_abc_19873_new_n1306_));
OAI21X1 OAI21X1_310 ( .A(\write_data[10] ), .B(_abc_19873_new_n2125__bF_buf3), .C(reset_n_bF_buf13), .Y(_abc_19873_new_n2149_));
OAI21X1 OAI21X1_311 ( .A(\write_data[11] ), .B(_abc_19873_new_n2125__bF_buf1), .C(reset_n_bF_buf12), .Y(_abc_19873_new_n2152_));
OAI21X1 OAI21X1_312 ( .A(\write_data[12] ), .B(_abc_19873_new_n2125__bF_buf7), .C(reset_n_bF_buf11), .Y(_abc_19873_new_n2155_));
OAI21X1 OAI21X1_313 ( .A(\write_data[13] ), .B(_abc_19873_new_n2125__bF_buf5), .C(reset_n_bF_buf10), .Y(_abc_19873_new_n2157_));
OAI21X1 OAI21X1_314 ( .A(\write_data[14] ), .B(_abc_19873_new_n2125__bF_buf3), .C(reset_n_bF_buf9), .Y(_abc_19873_new_n2159_));
OAI21X1 OAI21X1_315 ( .A(\write_data[15] ), .B(_abc_19873_new_n2125__bF_buf1), .C(reset_n_bF_buf8), .Y(_abc_19873_new_n2161_));
OAI21X1 OAI21X1_316 ( .A(\write_data[16] ), .B(_abc_19873_new_n2125__bF_buf7), .C(reset_n_bF_buf7), .Y(_abc_19873_new_n2163_));
OAI21X1 OAI21X1_317 ( .A(\write_data[17] ), .B(_abc_19873_new_n2125__bF_buf5), .C(reset_n_bF_buf6), .Y(_abc_19873_new_n2165_));
OAI21X1 OAI21X1_318 ( .A(\write_data[18] ), .B(_abc_19873_new_n2125__bF_buf3), .C(reset_n_bF_buf5), .Y(_abc_19873_new_n2168_));
OAI21X1 OAI21X1_319 ( .A(\write_data[19] ), .B(_abc_19873_new_n2125__bF_buf1), .C(reset_n_bF_buf4), .Y(_abc_19873_new_n2170_));
OAI21X1 OAI21X1_32 ( .A(_abc_19873_new_n1312_), .B(_abc_19873_new_n960__bF_buf1), .C(_abc_19873_new_n1313_), .Y(_abc_19873_new_n1314_));
OAI21X1 OAI21X1_320 ( .A(\write_data[20] ), .B(_abc_19873_new_n2125__bF_buf7), .C(reset_n_bF_buf3), .Y(_abc_19873_new_n2173_));
OAI21X1 OAI21X1_321 ( .A(\write_data[21] ), .B(_abc_19873_new_n2125__bF_buf5), .C(reset_n_bF_buf2), .Y(_abc_19873_new_n2175_));
OAI21X1 OAI21X1_322 ( .A(\write_data[22] ), .B(_abc_19873_new_n2125__bF_buf3), .C(reset_n_bF_buf1), .Y(_abc_19873_new_n2177_));
OAI21X1 OAI21X1_323 ( .A(\write_data[23] ), .B(_abc_19873_new_n2125__bF_buf1), .C(reset_n_bF_buf0), .Y(_abc_19873_new_n2179_));
OAI21X1 OAI21X1_324 ( .A(\write_data[24] ), .B(_abc_19873_new_n2125__bF_buf7), .C(reset_n_bF_buf69), .Y(_abc_19873_new_n2181_));
OAI21X1 OAI21X1_325 ( .A(\write_data[25] ), .B(_abc_19873_new_n2125__bF_buf5), .C(reset_n_bF_buf68), .Y(_abc_19873_new_n2183_));
OAI21X1 OAI21X1_326 ( .A(\write_data[26] ), .B(_abc_19873_new_n2125__bF_buf3), .C(reset_n_bF_buf67), .Y(_abc_19873_new_n2185_));
OAI21X1 OAI21X1_327 ( .A(\write_data[27] ), .B(_abc_19873_new_n2125__bF_buf1), .C(reset_n_bF_buf66), .Y(_abc_19873_new_n2187_));
OAI21X1 OAI21X1_328 ( .A(\write_data[28] ), .B(_abc_19873_new_n2125__bF_buf7), .C(reset_n_bF_buf65), .Y(_abc_19873_new_n2189_));
OAI21X1 OAI21X1_329 ( .A(\write_data[29] ), .B(_abc_19873_new_n2125__bF_buf5), .C(reset_n_bF_buf64), .Y(_abc_19873_new_n2191_));
OAI21X1 OAI21X1_33 ( .A(_abc_19873_new_n1341_), .B(_abc_19873_new_n894__bF_buf4), .C(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1342_));
OAI21X1 OAI21X1_330 ( .A(\write_data[30] ), .B(_abc_19873_new_n2125__bF_buf3), .C(reset_n_bF_buf63), .Y(_abc_19873_new_n2193_));
OAI21X1 OAI21X1_331 ( .A(\write_data[31] ), .B(_abc_19873_new_n2125__bF_buf1), .C(reset_n_bF_buf62), .Y(_abc_19873_new_n2195_));
OAI21X1 OAI21X1_332 ( .A(\write_data[0] ), .B(_abc_19873_new_n2198__bF_buf7), .C(reset_n_bF_buf61), .Y(_abc_19873_new_n2199_));
OAI21X1 OAI21X1_333 ( .A(\write_data[1] ), .B(_abc_19873_new_n2198__bF_buf5), .C(reset_n_bF_buf60), .Y(_abc_19873_new_n2202_));
OAI21X1 OAI21X1_334 ( .A(\write_data[2] ), .B(_abc_19873_new_n2198__bF_buf3), .C(reset_n_bF_buf59), .Y(_abc_19873_new_n2204_));
OAI21X1 OAI21X1_335 ( .A(\write_data[3] ), .B(_abc_19873_new_n2198__bF_buf1), .C(reset_n_bF_buf58), .Y(_abc_19873_new_n2206_));
OAI21X1 OAI21X1_336 ( .A(\write_data[4] ), .B(_abc_19873_new_n2198__bF_buf7), .C(reset_n_bF_buf57), .Y(_abc_19873_new_n2208_));
OAI21X1 OAI21X1_337 ( .A(\write_data[5] ), .B(_abc_19873_new_n2198__bF_buf5), .C(reset_n_bF_buf56), .Y(_abc_19873_new_n2210_));
OAI21X1 OAI21X1_338 ( .A(\write_data[6] ), .B(_abc_19873_new_n2198__bF_buf3), .C(reset_n_bF_buf55), .Y(_abc_19873_new_n2212_));
OAI21X1 OAI21X1_339 ( .A(\write_data[7] ), .B(_abc_19873_new_n2198__bF_buf1), .C(reset_n_bF_buf54), .Y(_abc_19873_new_n2214_));
OAI21X1 OAI21X1_34 ( .A(_abc_19873_new_n1344_), .B(_abc_19873_new_n1064__bF_buf2), .C(_abc_19873_new_n1345_), .Y(_abc_19873_new_n1346_));
OAI21X1 OAI21X1_340 ( .A(\write_data[8] ), .B(_abc_19873_new_n2198__bF_buf7), .C(reset_n_bF_buf53), .Y(_abc_19873_new_n2216_));
OAI21X1 OAI21X1_341 ( .A(\write_data[9] ), .B(_abc_19873_new_n2198__bF_buf5), .C(reset_n_bF_buf52), .Y(_abc_19873_new_n2218_));
OAI21X1 OAI21X1_342 ( .A(\write_data[10] ), .B(_abc_19873_new_n2198__bF_buf3), .C(reset_n_bF_buf51), .Y(_abc_19873_new_n2220_));
OAI21X1 OAI21X1_343 ( .A(\write_data[11] ), .B(_abc_19873_new_n2198__bF_buf1), .C(reset_n_bF_buf50), .Y(_abc_19873_new_n2222_));
OAI21X1 OAI21X1_344 ( .A(\write_data[12] ), .B(_abc_19873_new_n2198__bF_buf7), .C(reset_n_bF_buf49), .Y(_abc_19873_new_n2224_));
OAI21X1 OAI21X1_345 ( .A(\write_data[13] ), .B(_abc_19873_new_n2198__bF_buf5), .C(reset_n_bF_buf48), .Y(_abc_19873_new_n2226_));
OAI21X1 OAI21X1_346 ( .A(\write_data[14] ), .B(_abc_19873_new_n2198__bF_buf3), .C(reset_n_bF_buf47), .Y(_abc_19873_new_n2228_));
OAI21X1 OAI21X1_347 ( .A(\write_data[15] ), .B(_abc_19873_new_n2198__bF_buf1), .C(reset_n_bF_buf46), .Y(_abc_19873_new_n2230_));
OAI21X1 OAI21X1_348 ( .A(\write_data[16] ), .B(_abc_19873_new_n2198__bF_buf7), .C(reset_n_bF_buf45), .Y(_abc_19873_new_n2232_));
OAI21X1 OAI21X1_349 ( .A(\write_data[17] ), .B(_abc_19873_new_n2198__bF_buf5), .C(reset_n_bF_buf44), .Y(_abc_19873_new_n2234_));
OAI21X1 OAI21X1_35 ( .A(_abc_19873_new_n1378_), .B(_abc_19873_new_n894__bF_buf2), .C(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1379_));
OAI21X1 OAI21X1_350 ( .A(\write_data[18] ), .B(_abc_19873_new_n2198__bF_buf3), .C(reset_n_bF_buf43), .Y(_abc_19873_new_n2236_));
OAI21X1 OAI21X1_351 ( .A(\write_data[19] ), .B(_abc_19873_new_n2198__bF_buf1), .C(reset_n_bF_buf42), .Y(_abc_19873_new_n2238_));
OAI21X1 OAI21X1_352 ( .A(\write_data[20] ), .B(_abc_19873_new_n2198__bF_buf7), .C(reset_n_bF_buf41), .Y(_abc_19873_new_n2240_));
OAI21X1 OAI21X1_353 ( .A(\write_data[21] ), .B(_abc_19873_new_n2198__bF_buf5), .C(reset_n_bF_buf40), .Y(_abc_19873_new_n2242_));
OAI21X1 OAI21X1_354 ( .A(\write_data[22] ), .B(_abc_19873_new_n2198__bF_buf3), .C(reset_n_bF_buf39), .Y(_abc_19873_new_n2244_));
OAI21X1 OAI21X1_355 ( .A(\write_data[23] ), .B(_abc_19873_new_n2198__bF_buf1), .C(reset_n_bF_buf38), .Y(_abc_19873_new_n2246_));
OAI21X1 OAI21X1_356 ( .A(\write_data[24] ), .B(_abc_19873_new_n2198__bF_buf7), .C(reset_n_bF_buf37), .Y(_abc_19873_new_n2248_));
OAI21X1 OAI21X1_357 ( .A(\write_data[25] ), .B(_abc_19873_new_n2198__bF_buf5), .C(reset_n_bF_buf36), .Y(_abc_19873_new_n2250_));
OAI21X1 OAI21X1_358 ( .A(\write_data[26] ), .B(_abc_19873_new_n2198__bF_buf3), .C(reset_n_bF_buf35), .Y(_abc_19873_new_n2252_));
OAI21X1 OAI21X1_359 ( .A(\write_data[27] ), .B(_abc_19873_new_n2198__bF_buf1), .C(reset_n_bF_buf34), .Y(_abc_19873_new_n2254_));
OAI21X1 OAI21X1_36 ( .A(_abc_19873_new_n1381_), .B(_abc_19873_new_n1064__bF_buf0), .C(_abc_19873_new_n1382_), .Y(_abc_19873_new_n1383_));
OAI21X1 OAI21X1_360 ( .A(\write_data[28] ), .B(_abc_19873_new_n2198__bF_buf7), .C(reset_n_bF_buf33), .Y(_abc_19873_new_n2256_));
OAI21X1 OAI21X1_361 ( .A(\write_data[29] ), .B(_abc_19873_new_n2198__bF_buf5), .C(reset_n_bF_buf32), .Y(_abc_19873_new_n2259_));
OAI21X1 OAI21X1_362 ( .A(\write_data[30] ), .B(_abc_19873_new_n2198__bF_buf3), .C(reset_n_bF_buf31), .Y(_abc_19873_new_n2261_));
OAI21X1 OAI21X1_363 ( .A(\write_data[31] ), .B(_abc_19873_new_n2198__bF_buf1), .C(reset_n_bF_buf30), .Y(_abc_19873_new_n2263_));
OAI21X1 OAI21X1_364 ( .A(\write_data[0] ), .B(_abc_19873_new_n2266_), .C(reset_n_bF_buf29), .Y(_abc_19873_new_n2267_));
OAI21X1 OAI21X1_365 ( .A(_abc_19873_new_n944_), .B(_abc_19873_new_n2265_), .C(_abc_19873_new_n2270_), .Y(_0param_reg_7_0__1_));
OAI21X1 OAI21X1_366 ( .A(\write_data[2] ), .B(_abc_19873_new_n2266_), .C(reset_n_bF_buf27), .Y(_abc_19873_new_n2272_));
OAI21X1 OAI21X1_367 ( .A(\write_data[3] ), .B(_abc_19873_new_n2266_), .C(reset_n_bF_buf26), .Y(_abc_19873_new_n2274_));
OAI21X1 OAI21X1_368 ( .A(\write_data[4] ), .B(_abc_19873_new_n2266_), .C(reset_n_bF_buf25), .Y(_abc_19873_new_n2276_));
OAI21X1 OAI21X1_369 ( .A(\write_data[5] ), .B(_abc_19873_new_n2266_), .C(reset_n_bF_buf24), .Y(_abc_19873_new_n2278_));
OAI21X1 OAI21X1_37 ( .A(_abc_19873_new_n1396_), .B(_abc_19873_new_n894__bF_buf1), .C(_abc_19873_new_n1159_), .Y(_abc_19873_new_n1397_));
OAI21X1 OAI21X1_370 ( .A(_abc_19873_new_n1045_), .B(_abc_19873_new_n2265_), .C(_abc_19873_new_n2280_), .Y(_0param_reg_7_0__6_));
OAI21X1 OAI21X1_371 ( .A(\write_data[7] ), .B(_abc_19873_new_n2266_), .C(reset_n_bF_buf23), .Y(_abc_19873_new_n2282_));
OAI21X1 OAI21X1_372 ( .A(\write_data[0] ), .B(_abc_19873_new_n2295_), .C(reset_n_bF_buf21), .Y(_abc_19873_new_n2296_));
OAI21X1 OAI21X1_373 ( .A(core_loop_ctr_reg_3_), .B(core__abc_21302_new_n1133_), .C(core__abc_21302_new_n1143_), .Y(core__abc_21302_new_n1144_));
OAI21X1 OAI21X1_374 ( .A(core_finalize), .B(core_compress), .C(core__abc_21302_new_n1147_), .Y(core__abc_21302_new_n1148_));
OAI21X1 OAI21X1_375 ( .A(core_final_rounds_1_), .B(core_final_rounds_0_), .C(core_final_rounds_2_), .Y(core__abc_21302_new_n1166_));
OAI21X1 OAI21X1_376 ( .A(core__abc_21302_new_n1183_), .B(core__abc_21302_new_n1180_), .C(core__abc_21302_new_n1186_), .Y(core__abc_21302_new_n1187_));
OAI21X1 OAI21X1_377 ( .A(core__abc_21302_new_n1189_), .B(core__abc_21302_new_n1190_), .C(core__abc_21302_new_n1179_), .Y(core__abc_21302_new_n1191_));
OAI21X1 OAI21X1_378 ( .A(core__abc_21302_new_n1203_), .B(core__abc_21302_new_n1196_), .C(core__abc_21302_new_n1206_), .Y(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_6_));
OAI21X1 OAI21X1_379 ( .A(core_siphash_word1_we_bF_buf9), .B(core_siphash_word_64_), .C(reset_n_bF_buf18), .Y(core__abc_21302_new_n1218_));
OAI21X1 OAI21X1_38 ( .A(_abc_19873_new_n1399_), .B(_abc_19873_new_n1064__bF_buf3), .C(_abc_19873_new_n1400_), .Y(_abc_19873_new_n1401_));
OAI21X1 OAI21X1_380 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_65_), .C(reset_n_bF_buf17), .Y(core__abc_21302_new_n1230_));
OAI21X1 OAI21X1_381 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_66_), .C(reset_n_bF_buf16), .Y(core__abc_21302_new_n1239_));
OAI21X1 OAI21X1_382 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_67_), .C(reset_n_bF_buf15), .Y(core__abc_21302_new_n1249_));
OAI21X1 OAI21X1_383 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_68_), .C(reset_n_bF_buf14), .Y(core__abc_21302_new_n1259_));
OAI21X1 OAI21X1_384 ( .A(core_siphash_word1_we_bF_buf10), .B(core_siphash_word_69_), .C(reset_n_bF_buf13), .Y(core__abc_21302_new_n1271_));
OAI21X1 OAI21X1_385 ( .A(core_siphash_word1_we_bF_buf8), .B(core_siphash_word_70_), .C(reset_n_bF_buf12), .Y(core__abc_21302_new_n1281_));
OAI21X1 OAI21X1_386 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_71_), .C(reset_n_bF_buf11), .Y(core__abc_21302_new_n1291_));
OAI21X1 OAI21X1_387 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_72_), .C(reset_n_bF_buf10), .Y(core__abc_21302_new_n1299_));
OAI21X1 OAI21X1_388 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_73_), .C(reset_n_bF_buf9), .Y(core__abc_21302_new_n1310_));
OAI21X1 OAI21X1_389 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_74_), .C(reset_n_bF_buf8), .Y(core__abc_21302_new_n1322_));
OAI21X1 OAI21X1_39 ( .A(_abc_19873_new_n1452_), .B(_abc_19873_new_n894__bF_buf3), .C(_abc_19873_new_n1159_), .Y(_abc_19873_new_n1453_));
OAI21X1 OAI21X1_390 ( .A(core_siphash_word1_we_bF_buf9), .B(core_siphash_word_75_), .C(reset_n_bF_buf7), .Y(core__abc_21302_new_n1334_));
OAI21X1 OAI21X1_391 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_76_), .C(reset_n_bF_buf6), .Y(core__abc_21302_new_n1344_));
OAI21X1 OAI21X1_392 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_77_), .C(reset_n_bF_buf5), .Y(core__abc_21302_new_n1356_));
OAI21X1 OAI21X1_393 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_78_), .C(reset_n_bF_buf4), .Y(core__abc_21302_new_n1368_));
OAI21X1 OAI21X1_394 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_79_), .C(reset_n_bF_buf3), .Y(core__abc_21302_new_n1380_));
OAI21X1 OAI21X1_395 ( .A(core_siphash_word1_we_bF_buf10), .B(core_siphash_word_80_), .C(reset_n_bF_buf2), .Y(core__abc_21302_new_n1391_));
OAI21X1 OAI21X1_396 ( .A(core_siphash_word1_we_bF_buf8), .B(core_siphash_word_81_), .C(reset_n_bF_buf1), .Y(core__abc_21302_new_n1403_));
OAI21X1 OAI21X1_397 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_82_), .C(reset_n_bF_buf0), .Y(core__abc_21302_new_n1415_));
OAI21X1 OAI21X1_398 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_83_), .C(reset_n_bF_buf69), .Y(core__abc_21302_new_n1427_));
OAI21X1 OAI21X1_399 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_84_), .C(reset_n_bF_buf68), .Y(core__abc_21302_new_n1439_));
OAI21X1 OAI21X1_4 ( .A(_abc_19873_new_n944_), .B(_abc_19873_new_n918_), .C(_abc_19873_new_n945_), .Y(_abc_19873_new_n946_));
OAI21X1 OAI21X1_40 ( .A(_abc_19873_new_n1455_), .B(_abc_19873_new_n1064__bF_buf0), .C(_abc_19873_new_n1456_), .Y(_abc_19873_new_n1457_));
OAI21X1 OAI21X1_400 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_85_), .C(reset_n_bF_buf67), .Y(core__abc_21302_new_n1451_));
OAI21X1 OAI21X1_401 ( .A(core_siphash_word1_we_bF_buf9), .B(core_siphash_word_86_), .C(reset_n_bF_buf66), .Y(core__abc_21302_new_n1463_));
OAI21X1 OAI21X1_402 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_87_), .C(reset_n_bF_buf65), .Y(core__abc_21302_new_n1471_));
OAI21X1 OAI21X1_403 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_88_), .C(reset_n_bF_buf64), .Y(core__abc_21302_new_n1483_));
OAI21X1 OAI21X1_404 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_89_), .C(reset_n_bF_buf63), .Y(core__abc_21302_new_n1493_));
OAI21X1 OAI21X1_405 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_90_), .C(reset_n_bF_buf62), .Y(core__abc_21302_new_n1505_));
OAI21X1 OAI21X1_406 ( .A(core_siphash_word1_we_bF_buf10), .B(core_siphash_word_91_), .C(reset_n_bF_buf61), .Y(core__abc_21302_new_n1517_));
OAI21X1 OAI21X1_407 ( .A(core_siphash_word1_we_bF_buf8), .B(core_siphash_word_92_), .C(reset_n_bF_buf60), .Y(core__abc_21302_new_n1529_));
OAI21X1 OAI21X1_408 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_93_), .C(reset_n_bF_buf59), .Y(core__abc_21302_new_n1542_));
OAI21X1 OAI21X1_409 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_94_), .C(reset_n_bF_buf58), .Y(core__abc_21302_new_n1554_));
OAI21X1 OAI21X1_41 ( .A(_abc_19873_new_n893__bF_buf3), .B(_abc_19873_new_n1480_), .C(_abc_19873_new_n877_), .Y(_abc_19873_new_n1481_));
OAI21X1 OAI21X1_410 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_95_), .C(reset_n_bF_buf57), .Y(core__abc_21302_new_n1562_));
OAI21X1 OAI21X1_411 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_96_), .C(reset_n_bF_buf56), .Y(core__abc_21302_new_n1574_));
OAI21X1 OAI21X1_412 ( .A(core_siphash_word1_we_bF_buf9), .B(core_siphash_word_97_), .C(reset_n_bF_buf55), .Y(core__abc_21302_new_n1586_));
OAI21X1 OAI21X1_413 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_98_), .C(reset_n_bF_buf54), .Y(core__abc_21302_new_n1600_));
OAI21X1 OAI21X1_414 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_99_), .C(reset_n_bF_buf53), .Y(core__abc_21302_new_n1612_));
OAI21X1 OAI21X1_415 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_100_), .C(reset_n_bF_buf52), .Y(core__abc_21302_new_n1623_));
OAI21X1 OAI21X1_416 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_101_), .C(reset_n_bF_buf51), .Y(core__abc_21302_new_n1636_));
OAI21X1 OAI21X1_417 ( .A(core_siphash_word1_we_bF_buf10), .B(core_siphash_word_102_), .C(reset_n_bF_buf50), .Y(core__abc_21302_new_n1645_));
OAI21X1 OAI21X1_418 ( .A(core_siphash_word1_we_bF_buf8), .B(core_siphash_word_103_), .C(reset_n_bF_buf49), .Y(core__abc_21302_new_n1656_));
OAI21X1 OAI21X1_419 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_104_), .C(reset_n_bF_buf48), .Y(core__abc_21302_new_n1667_));
OAI21X1 OAI21X1_42 ( .A(_abc_19873_new_n1490_), .B(_abc_19873_new_n894__bF_buf1), .C(_abc_19873_new_n1018_), .Y(_abc_19873_new_n1491_));
OAI21X1 OAI21X1_420 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_105_), .C(reset_n_bF_buf47), .Y(core__abc_21302_new_n1678_));
OAI21X1 OAI21X1_421 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_106_), .C(reset_n_bF_buf46), .Y(core__abc_21302_new_n1689_));
OAI21X1 OAI21X1_422 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_107_), .C(reset_n_bF_buf45), .Y(core__abc_21302_new_n1700_));
OAI21X1 OAI21X1_423 ( .A(core_siphash_word1_we_bF_buf9), .B(core_siphash_word_108_), .C(reset_n_bF_buf44), .Y(core__abc_21302_new_n1712_));
OAI21X1 OAI21X1_424 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_109_), .C(reset_n_bF_buf43), .Y(core__abc_21302_new_n1723_));
OAI21X1 OAI21X1_425 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_110_), .C(reset_n_bF_buf42), .Y(core__abc_21302_new_n1735_));
OAI21X1 OAI21X1_426 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_111_), .C(reset_n_bF_buf41), .Y(core__abc_21302_new_n1746_));
OAI21X1 OAI21X1_427 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_112_), .C(reset_n_bF_buf40), .Y(core__abc_21302_new_n1759_));
OAI21X1 OAI21X1_428 ( .A(core_siphash_word1_we_bF_buf10), .B(core_siphash_word_113_), .C(reset_n_bF_buf39), .Y(core__abc_21302_new_n1768_));
OAI21X1 OAI21X1_429 ( .A(core_siphash_word1_we_bF_buf8), .B(core_siphash_word_114_), .C(reset_n_bF_buf38), .Y(core__abc_21302_new_n1780_));
OAI21X1 OAI21X1_43 ( .A(_abc_19873_new_n1493_), .B(_abc_19873_new_n1064__bF_buf2), .C(_abc_19873_new_n1494_), .Y(_abc_19873_new_n1495_));
OAI21X1 OAI21X1_430 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_115_), .C(reset_n_bF_buf37), .Y(core__abc_21302_new_n1791_));
OAI21X1 OAI21X1_431 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_116_), .C(reset_n_bF_buf36), .Y(core__abc_21302_new_n1805_));
OAI21X1 OAI21X1_432 ( .A(core_siphash_word1_we_bF_buf2), .B(core_siphash_word_117_), .C(reset_n_bF_buf35), .Y(core__abc_21302_new_n1816_));
OAI21X1 OAI21X1_433 ( .A(core_siphash_word1_we_bF_buf0), .B(core_siphash_word_118_), .C(reset_n_bF_buf34), .Y(core__abc_21302_new_n1829_));
OAI21X1 OAI21X1_434 ( .A(core_siphash_word1_we_bF_buf9), .B(core_siphash_word_119_), .C(reset_n_bF_buf33), .Y(core__abc_21302_new_n1842_));
OAI21X1 OAI21X1_435 ( .A(core_siphash_word1_we_bF_buf7), .B(core_siphash_word_120_), .C(reset_n_bF_buf32), .Y(core__abc_21302_new_n1856_));
OAI21X1 OAI21X1_436 ( .A(core_siphash_word1_we_bF_buf5), .B(core_siphash_word_121_), .C(reset_n_bF_buf31), .Y(core__abc_21302_new_n1868_));
OAI21X1 OAI21X1_437 ( .A(core_siphash_word1_we_bF_buf3), .B(core_siphash_word_122_), .C(reset_n_bF_buf30), .Y(core__abc_21302_new_n1882_));
OAI21X1 OAI21X1_438 ( .A(core_siphash_word1_we_bF_buf1), .B(core_siphash_word_123_), .C(reset_n_bF_buf29), .Y(core__abc_21302_new_n1894_));
OAI21X1 OAI21X1_439 ( .A(core_siphash_word1_we_bF_buf10), .B(core_siphash_word_124_), .C(reset_n_bF_buf28), .Y(core__abc_21302_new_n1908_));
OAI21X1 OAI21X1_44 ( .A(core_siphash_word_96_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf69), .Y(_abc_19873_new_n1525_));
OAI21X1 OAI21X1_440 ( .A(core_siphash_word1_we_bF_buf8), .B(core_siphash_word_125_), .C(reset_n_bF_buf27), .Y(core__abc_21302_new_n1922_));
OAI21X1 OAI21X1_441 ( .A(core_siphash_word1_we_bF_buf6), .B(core_siphash_word_126_), .C(reset_n_bF_buf26), .Y(core__abc_21302_new_n1935_));
OAI21X1 OAI21X1_442 ( .A(core_siphash_word1_we_bF_buf4), .B(core_siphash_word_127_), .C(reset_n_bF_buf25), .Y(core__abc_21302_new_n1941_));
OAI21X1 OAI21X1_443 ( .A(core_siphash_word_0_), .B(core__abc_21302_new_n1945__bF_buf9), .C(core__abc_21302_new_n1946_), .Y(core__abc_21302_new_n1947_));
OAI21X1 OAI21X1_444 ( .A(core_siphash_word_1_), .B(core__abc_21302_new_n1945__bF_buf7), .C(core__abc_21302_new_n1949_), .Y(core__abc_21302_new_n1950_));
OAI21X1 OAI21X1_445 ( .A(core_siphash_word_2_), .B(core__abc_21302_new_n1945__bF_buf5), .C(core__abc_21302_new_n1952_), .Y(core__abc_21302_new_n1953_));
OAI21X1 OAI21X1_446 ( .A(core_siphash_word_3_), .B(core__abc_21302_new_n1945__bF_buf3), .C(core__abc_21302_new_n1955_), .Y(core__abc_21302_new_n1956_));
OAI21X1 OAI21X1_447 ( .A(core_siphash_word_4_), .B(core__abc_21302_new_n1945__bF_buf1), .C(core__abc_21302_new_n1958_), .Y(core__abc_21302_new_n1959_));
OAI21X1 OAI21X1_448 ( .A(core_siphash_word_5_), .B(core__abc_21302_new_n1945__bF_buf10), .C(core__abc_21302_new_n1961_), .Y(core__abc_21302_new_n1962_));
OAI21X1 OAI21X1_449 ( .A(core_siphash_word_6_), .B(core__abc_21302_new_n1945__bF_buf8), .C(core__abc_21302_new_n1964_), .Y(core__abc_21302_new_n1965_));
OAI21X1 OAI21X1_45 ( .A(core_siphash_word_97_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf68), .Y(_abc_19873_new_n1527_));
OAI21X1 OAI21X1_450 ( .A(core_siphash_word_7_), .B(core__abc_21302_new_n1945__bF_buf6), .C(core__abc_21302_new_n1967_), .Y(core__abc_21302_new_n1968_));
OAI21X1 OAI21X1_451 ( .A(core_siphash_word_8_), .B(core__abc_21302_new_n1945__bF_buf4), .C(core__abc_21302_new_n1970_), .Y(core__abc_21302_new_n1971_));
OAI21X1 OAI21X1_452 ( .A(core_siphash_word_9_), .B(core__abc_21302_new_n1945__bF_buf2), .C(core__abc_21302_new_n1973_), .Y(core__abc_21302_new_n1974_));
OAI21X1 OAI21X1_453 ( .A(core_siphash_word_10_), .B(core__abc_21302_new_n1945__bF_buf0), .C(core__abc_21302_new_n1976_), .Y(core__abc_21302_new_n1977_));
OAI21X1 OAI21X1_454 ( .A(core_siphash_word_11_), .B(core__abc_21302_new_n1945__bF_buf9), .C(core__abc_21302_new_n1979_), .Y(core__abc_21302_new_n1980_));
OAI21X1 OAI21X1_455 ( .A(core_siphash_word_12_), .B(core__abc_21302_new_n1945__bF_buf7), .C(core__abc_21302_new_n1982_), .Y(core__abc_21302_new_n1983_));
OAI21X1 OAI21X1_456 ( .A(core_siphash_word_13_), .B(core__abc_21302_new_n1945__bF_buf5), .C(core__abc_21302_new_n1985_), .Y(core__abc_21302_new_n1986_));
OAI21X1 OAI21X1_457 ( .A(core_siphash_word_14_), .B(core__abc_21302_new_n1945__bF_buf3), .C(core__abc_21302_new_n1988_), .Y(core__abc_21302_new_n1989_));
OAI21X1 OAI21X1_458 ( .A(core_siphash_word_15_), .B(core__abc_21302_new_n1945__bF_buf1), .C(core__abc_21302_new_n1991_), .Y(core__abc_21302_new_n1992_));
OAI21X1 OAI21X1_459 ( .A(core_siphash_word_16_), .B(core__abc_21302_new_n1945__bF_buf10), .C(core__abc_21302_new_n1994_), .Y(core__abc_21302_new_n1995_));
OAI21X1 OAI21X1_46 ( .A(core_siphash_word_98_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf67), .Y(_abc_19873_new_n1530_));
OAI21X1 OAI21X1_460 ( .A(core_siphash_word_17_), .B(core__abc_21302_new_n1945__bF_buf8), .C(core__abc_21302_new_n1997_), .Y(core__abc_21302_new_n1998_));
OAI21X1 OAI21X1_461 ( .A(core_siphash_word_18_), .B(core__abc_21302_new_n1945__bF_buf6), .C(core__abc_21302_new_n2000_), .Y(core__abc_21302_new_n2001_));
OAI21X1 OAI21X1_462 ( .A(core_siphash_word_19_), .B(core__abc_21302_new_n1945__bF_buf4), .C(core__abc_21302_new_n2003_), .Y(core__abc_21302_new_n2004_));
OAI21X1 OAI21X1_463 ( .A(core_siphash_word_20_), .B(core__abc_21302_new_n1945__bF_buf2), .C(core__abc_21302_new_n2006_), .Y(core__abc_21302_new_n2007_));
OAI21X1 OAI21X1_464 ( .A(core_siphash_word_21_), .B(core__abc_21302_new_n1945__bF_buf0), .C(core__abc_21302_new_n2009_), .Y(core__abc_21302_new_n2010_));
OAI21X1 OAI21X1_465 ( .A(core_siphash_word_22_), .B(core__abc_21302_new_n1945__bF_buf9), .C(core__abc_21302_new_n2012_), .Y(core__abc_21302_new_n2013_));
OAI21X1 OAI21X1_466 ( .A(core_siphash_word_23_), .B(core__abc_21302_new_n1945__bF_buf7), .C(core__abc_21302_new_n2015_), .Y(core__abc_21302_new_n2016_));
OAI21X1 OAI21X1_467 ( .A(core_siphash_word_24_), .B(core__abc_21302_new_n1945__bF_buf5), .C(core__abc_21302_new_n2018_), .Y(core__abc_21302_new_n2019_));
OAI21X1 OAI21X1_468 ( .A(core_siphash_word_25_), .B(core__abc_21302_new_n1945__bF_buf3), .C(core__abc_21302_new_n2021_), .Y(core__abc_21302_new_n2022_));
OAI21X1 OAI21X1_469 ( .A(core_siphash_word_26_), .B(core__abc_21302_new_n1945__bF_buf1), .C(core__abc_21302_new_n2024_), .Y(core__abc_21302_new_n2025_));
OAI21X1 OAI21X1_47 ( .A(core_siphash_word_99_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf66), .Y(_abc_19873_new_n1532_));
OAI21X1 OAI21X1_470 ( .A(core_siphash_word_27_), .B(core__abc_21302_new_n1945__bF_buf10), .C(core__abc_21302_new_n2027_), .Y(core__abc_21302_new_n2028_));
OAI21X1 OAI21X1_471 ( .A(core_siphash_word_28_), .B(core__abc_21302_new_n1945__bF_buf8), .C(core__abc_21302_new_n2030_), .Y(core__abc_21302_new_n2031_));
OAI21X1 OAI21X1_472 ( .A(core_siphash_word_29_), .B(core__abc_21302_new_n1945__bF_buf6), .C(core__abc_21302_new_n2033_), .Y(core__abc_21302_new_n2034_));
OAI21X1 OAI21X1_473 ( .A(core_siphash_word_30_), .B(core__abc_21302_new_n1945__bF_buf4), .C(core__abc_21302_new_n2036_), .Y(core__abc_21302_new_n2037_));
OAI21X1 OAI21X1_474 ( .A(core_siphash_word_31_), .B(core__abc_21302_new_n1945__bF_buf2), .C(core__abc_21302_new_n2039_), .Y(core__abc_21302_new_n2040_));
OAI21X1 OAI21X1_475 ( .A(core_siphash_word_32_), .B(core__abc_21302_new_n1945__bF_buf0), .C(core__abc_21302_new_n2042_), .Y(core__abc_21302_new_n2043_));
OAI21X1 OAI21X1_476 ( .A(core_siphash_word_33_), .B(core__abc_21302_new_n1945__bF_buf9), .C(core__abc_21302_new_n2045_), .Y(core__abc_21302_new_n2046_));
OAI21X1 OAI21X1_477 ( .A(core_siphash_word_34_), .B(core__abc_21302_new_n1945__bF_buf7), .C(core__abc_21302_new_n2048_), .Y(core__abc_21302_new_n2049_));
OAI21X1 OAI21X1_478 ( .A(core_siphash_word_35_), .B(core__abc_21302_new_n1945__bF_buf5), .C(core__abc_21302_new_n2051_), .Y(core__abc_21302_new_n2052_));
OAI21X1 OAI21X1_479 ( .A(core_siphash_word_36_), .B(core__abc_21302_new_n1945__bF_buf3), .C(core__abc_21302_new_n2054_), .Y(core__abc_21302_new_n2055_));
OAI21X1 OAI21X1_48 ( .A(core_siphash_word_100_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf65), .Y(_abc_19873_new_n1534_));
OAI21X1 OAI21X1_480 ( .A(core_siphash_word_37_), .B(core__abc_21302_new_n1945__bF_buf1), .C(core__abc_21302_new_n2057_), .Y(core__abc_21302_new_n2058_));
OAI21X1 OAI21X1_481 ( .A(core_siphash_word_38_), .B(core__abc_21302_new_n1945__bF_buf10), .C(core__abc_21302_new_n2060_), .Y(core__abc_21302_new_n2061_));
OAI21X1 OAI21X1_482 ( .A(core_siphash_word_39_), .B(core__abc_21302_new_n1945__bF_buf8), .C(core__abc_21302_new_n2063_), .Y(core__abc_21302_new_n2064_));
OAI21X1 OAI21X1_483 ( .A(core_siphash_word_40_), .B(core__abc_21302_new_n1945__bF_buf6), .C(core__abc_21302_new_n2066_), .Y(core__abc_21302_new_n2067_));
OAI21X1 OAI21X1_484 ( .A(core_siphash_word_41_), .B(core__abc_21302_new_n1945__bF_buf4), .C(core__abc_21302_new_n2069_), .Y(core__abc_21302_new_n2070_));
OAI21X1 OAI21X1_485 ( .A(core_siphash_word_42_), .B(core__abc_21302_new_n1945__bF_buf2), .C(core__abc_21302_new_n2072_), .Y(core__abc_21302_new_n2073_));
OAI21X1 OAI21X1_486 ( .A(core_siphash_word_43_), .B(core__abc_21302_new_n1945__bF_buf0), .C(core__abc_21302_new_n2075_), .Y(core__abc_21302_new_n2076_));
OAI21X1 OAI21X1_487 ( .A(core_siphash_word_44_), .B(core__abc_21302_new_n1945__bF_buf9), .C(core__abc_21302_new_n2078_), .Y(core__abc_21302_new_n2079_));
OAI21X1 OAI21X1_488 ( .A(core_siphash_word_45_), .B(core__abc_21302_new_n1945__bF_buf7), .C(core__abc_21302_new_n2081_), .Y(core__abc_21302_new_n2082_));
OAI21X1 OAI21X1_489 ( .A(core_siphash_word_46_), .B(core__abc_21302_new_n1945__bF_buf5), .C(core__abc_21302_new_n2084_), .Y(core__abc_21302_new_n2085_));
OAI21X1 OAI21X1_49 ( .A(core_siphash_word_101_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf64), .Y(_abc_19873_new_n1536_));
OAI21X1 OAI21X1_490 ( .A(core_siphash_word_47_), .B(core__abc_21302_new_n1945__bF_buf3), .C(core__abc_21302_new_n2087_), .Y(core__abc_21302_new_n2088_));
OAI21X1 OAI21X1_491 ( .A(core_siphash_word_48_), .B(core__abc_21302_new_n1945__bF_buf1), .C(core__abc_21302_new_n2090_), .Y(core__abc_21302_new_n2091_));
OAI21X1 OAI21X1_492 ( .A(core_siphash_word_49_), .B(core__abc_21302_new_n1945__bF_buf10), .C(core__abc_21302_new_n2093_), .Y(core__abc_21302_new_n2094_));
OAI21X1 OAI21X1_493 ( .A(core_siphash_word_50_), .B(core__abc_21302_new_n1945__bF_buf8), .C(core__abc_21302_new_n2096_), .Y(core__abc_21302_new_n2097_));
OAI21X1 OAI21X1_494 ( .A(core_siphash_word_51_), .B(core__abc_21302_new_n1945__bF_buf6), .C(core__abc_21302_new_n2099_), .Y(core__abc_21302_new_n2100_));
OAI21X1 OAI21X1_495 ( .A(core_siphash_word_52_), .B(core__abc_21302_new_n1945__bF_buf4), .C(core__abc_21302_new_n2102_), .Y(core__abc_21302_new_n2103_));
OAI21X1 OAI21X1_496 ( .A(core_siphash_word_53_), .B(core__abc_21302_new_n1945__bF_buf2), .C(core__abc_21302_new_n2105_), .Y(core__abc_21302_new_n2106_));
OAI21X1 OAI21X1_497 ( .A(core_siphash_word_54_), .B(core__abc_21302_new_n1945__bF_buf0), .C(core__abc_21302_new_n2108_), .Y(core__abc_21302_new_n2109_));
OAI21X1 OAI21X1_498 ( .A(core_siphash_word_55_), .B(core__abc_21302_new_n1945__bF_buf9), .C(core__abc_21302_new_n2111_), .Y(core__abc_21302_new_n2112_));
OAI21X1 OAI21X1_499 ( .A(core_siphash_word_56_), .B(core__abc_21302_new_n1945__bF_buf7), .C(core__abc_21302_new_n2114_), .Y(core__abc_21302_new_n2115_));
OAI21X1 OAI21X1_5 ( .A(_abc_19873_new_n971_), .B(_abc_19873_new_n918_), .C(_abc_19873_new_n972_), .Y(_abc_19873_new_n973_));
OAI21X1 OAI21X1_50 ( .A(core_siphash_word_102_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf63), .Y(_abc_19873_new_n1538_));
OAI21X1 OAI21X1_500 ( .A(core_siphash_word_57_), .B(core__abc_21302_new_n1945__bF_buf5), .C(core__abc_21302_new_n2117_), .Y(core__abc_21302_new_n2118_));
OAI21X1 OAI21X1_501 ( .A(core_siphash_word_58_), .B(core__abc_21302_new_n1945__bF_buf3), .C(core__abc_21302_new_n2120_), .Y(core__abc_21302_new_n2121_));
OAI21X1 OAI21X1_502 ( .A(core_siphash_word_59_), .B(core__abc_21302_new_n1945__bF_buf1), .C(core__abc_21302_new_n2123_), .Y(core__abc_21302_new_n2124_));
OAI21X1 OAI21X1_503 ( .A(core_siphash_word_60_), .B(core__abc_21302_new_n1945__bF_buf10), .C(core__abc_21302_new_n2126_), .Y(core__abc_21302_new_n2127_));
OAI21X1 OAI21X1_504 ( .A(core_siphash_word_61_), .B(core__abc_21302_new_n1945__bF_buf8), .C(core__abc_21302_new_n2129_), .Y(core__abc_21302_new_n2130_));
OAI21X1 OAI21X1_505 ( .A(core_siphash_word_62_), .B(core__abc_21302_new_n1945__bF_buf6), .C(core__abc_21302_new_n2132_), .Y(core__abc_21302_new_n2133_));
OAI21X1 OAI21X1_506 ( .A(core_siphash_word_63_), .B(core__abc_21302_new_n1945__bF_buf4), .C(core__abc_21302_new_n2135_), .Y(core__abc_21302_new_n2136_));
OAI21X1 OAI21X1_507 ( .A(core__abc_21302_new_n1148_), .B(core__abc_21302_new_n2139_), .C(core_ready), .Y(core__abc_21302_new_n2140_));
OAI21X1 OAI21X1_508 ( .A(core__abc_21302_new_n1148_), .B(core__abc_21302_new_n1157_), .C(core__abc_21302_new_n1194_), .Y(core__abc_21302_new_n2144_));
OAI21X1 OAI21X1_509 ( .A(core_loop_ctr_reg_0_), .B(core__abc_21302_new_n2143_), .C(reset_n_bF_buf24), .Y(core__abc_21302_new_n2147_));
OAI21X1 OAI21X1_51 ( .A(core_siphash_word_103_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf62), .Y(_abc_19873_new_n1541_));
OAI21X1 OAI21X1_510 ( .A(core_loop_ctr_reg_1_), .B(core__abc_21302_new_n2146_), .C(reset_n_bF_buf23), .Y(core__abc_21302_new_n2152_));
OAI21X1 OAI21X1_511 ( .A(core_loop_ctr_reg_3_), .B(core__abc_21302_new_n2157_), .C(reset_n_bF_buf21), .Y(core__abc_21302_new_n2162_));
OAI21X1 OAI21X1_512 ( .A(core_mi_0_), .B(core__abc_21302_new_n2168__bF_buf12), .C(reset_n_bF_buf20), .Y(core__abc_21302_new_n2169_));
OAI21X1 OAI21X1_513 ( .A(core_mi_1_), .B(core__abc_21302_new_n2168__bF_buf10), .C(reset_n_bF_buf19), .Y(core__abc_21302_new_n2172_));
OAI21X1 OAI21X1_514 ( .A(core_mi_2_), .B(core__abc_21302_new_n2168__bF_buf8), .C(reset_n_bF_buf18), .Y(core__abc_21302_new_n2175_));
OAI21X1 OAI21X1_515 ( .A(core_mi_3_), .B(core__abc_21302_new_n2168__bF_buf6), .C(reset_n_bF_buf17), .Y(core__abc_21302_new_n2178_));
OAI21X1 OAI21X1_516 ( .A(core_mi_4_), .B(core__abc_21302_new_n2168__bF_buf4), .C(reset_n_bF_buf16), .Y(core__abc_21302_new_n2181_));
OAI21X1 OAI21X1_517 ( .A(core_mi_5_), .B(core__abc_21302_new_n2168__bF_buf2), .C(reset_n_bF_buf15), .Y(core__abc_21302_new_n2184_));
OAI21X1 OAI21X1_518 ( .A(core_mi_6_), .B(core__abc_21302_new_n2168__bF_buf0), .C(reset_n_bF_buf14), .Y(core__abc_21302_new_n2187_));
OAI21X1 OAI21X1_519 ( .A(core_mi_7_), .B(core__abc_21302_new_n2168__bF_buf11), .C(reset_n_bF_buf13), .Y(core__abc_21302_new_n2190_));
OAI21X1 OAI21X1_52 ( .A(core_siphash_word_104_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf61), .Y(_abc_19873_new_n1543_));
OAI21X1 OAI21X1_520 ( .A(core_mi_8_), .B(core__abc_21302_new_n2168__bF_buf9), .C(reset_n_bF_buf12), .Y(core__abc_21302_new_n2193_));
OAI21X1 OAI21X1_521 ( .A(core_mi_9_), .B(core__abc_21302_new_n2168__bF_buf7), .C(reset_n_bF_buf11), .Y(core__abc_21302_new_n2196_));
OAI21X1 OAI21X1_522 ( .A(core_mi_10_), .B(core__abc_21302_new_n2168__bF_buf5), .C(reset_n_bF_buf10), .Y(core__abc_21302_new_n2199_));
OAI21X1 OAI21X1_523 ( .A(core_mi_11_), .B(core__abc_21302_new_n2168__bF_buf3), .C(reset_n_bF_buf9), .Y(core__abc_21302_new_n2202_));
OAI21X1 OAI21X1_524 ( .A(core_mi_12_), .B(core__abc_21302_new_n2168__bF_buf1), .C(reset_n_bF_buf8), .Y(core__abc_21302_new_n2205_));
OAI21X1 OAI21X1_525 ( .A(core_mi_13_), .B(core__abc_21302_new_n2168__bF_buf12), .C(reset_n_bF_buf7), .Y(core__abc_21302_new_n2208_));
OAI21X1 OAI21X1_526 ( .A(core_mi_14_), .B(core__abc_21302_new_n2168__bF_buf10), .C(reset_n_bF_buf6), .Y(core__abc_21302_new_n2211_));
OAI21X1 OAI21X1_527 ( .A(core_mi_15_), .B(core__abc_21302_new_n2168__bF_buf8), .C(reset_n_bF_buf5), .Y(core__abc_21302_new_n2214_));
OAI21X1 OAI21X1_528 ( .A(core_mi_16_), .B(core__abc_21302_new_n2168__bF_buf6), .C(reset_n_bF_buf4), .Y(core__abc_21302_new_n2217_));
OAI21X1 OAI21X1_529 ( .A(core_mi_17_), .B(core__abc_21302_new_n2168__bF_buf4), .C(reset_n_bF_buf3), .Y(core__abc_21302_new_n2220_));
OAI21X1 OAI21X1_53 ( .A(core_siphash_word_105_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf60), .Y(_abc_19873_new_n1545_));
OAI21X1 OAI21X1_530 ( .A(core_mi_18_), .B(core__abc_21302_new_n2168__bF_buf2), .C(reset_n_bF_buf2), .Y(core__abc_21302_new_n2223_));
OAI21X1 OAI21X1_531 ( .A(core_mi_19_), .B(core__abc_21302_new_n2168__bF_buf0), .C(reset_n_bF_buf1), .Y(core__abc_21302_new_n2226_));
OAI21X1 OAI21X1_532 ( .A(core_mi_20_), .B(core__abc_21302_new_n2168__bF_buf11), .C(reset_n_bF_buf0), .Y(core__abc_21302_new_n2229_));
OAI21X1 OAI21X1_533 ( .A(core_mi_21_), .B(core__abc_21302_new_n2168__bF_buf9), .C(reset_n_bF_buf69), .Y(core__abc_21302_new_n2232_));
OAI21X1 OAI21X1_534 ( .A(core_mi_22_), .B(core__abc_21302_new_n2168__bF_buf7), .C(reset_n_bF_buf68), .Y(core__abc_21302_new_n2235_));
OAI21X1 OAI21X1_535 ( .A(core_mi_23_), .B(core__abc_21302_new_n2168__bF_buf5), .C(reset_n_bF_buf67), .Y(core__abc_21302_new_n2238_));
OAI21X1 OAI21X1_536 ( .A(core_mi_24_), .B(core__abc_21302_new_n2168__bF_buf3), .C(reset_n_bF_buf66), .Y(core__abc_21302_new_n2241_));
OAI21X1 OAI21X1_537 ( .A(core_mi_25_), .B(core__abc_21302_new_n2168__bF_buf1), .C(reset_n_bF_buf65), .Y(core__abc_21302_new_n2244_));
OAI21X1 OAI21X1_538 ( .A(core_mi_26_), .B(core__abc_21302_new_n2168__bF_buf12), .C(reset_n_bF_buf64), .Y(core__abc_21302_new_n2247_));
OAI21X1 OAI21X1_539 ( .A(core_mi_27_), .B(core__abc_21302_new_n2168__bF_buf10), .C(reset_n_bF_buf63), .Y(core__abc_21302_new_n2250_));
OAI21X1 OAI21X1_54 ( .A(core_siphash_word_106_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf59), .Y(_abc_19873_new_n1547_));
OAI21X1 OAI21X1_540 ( .A(core_mi_28_), .B(core__abc_21302_new_n2168__bF_buf8), .C(reset_n_bF_buf62), .Y(core__abc_21302_new_n2253_));
OAI21X1 OAI21X1_541 ( .A(core_mi_29_), .B(core__abc_21302_new_n2168__bF_buf6), .C(reset_n_bF_buf61), .Y(core__abc_21302_new_n2256_));
OAI21X1 OAI21X1_542 ( .A(core_mi_30_), .B(core__abc_21302_new_n2168__bF_buf4), .C(reset_n_bF_buf60), .Y(core__abc_21302_new_n2259_));
OAI21X1 OAI21X1_543 ( .A(core_mi_31_), .B(core__abc_21302_new_n2168__bF_buf2), .C(reset_n_bF_buf59), .Y(core__abc_21302_new_n2262_));
OAI21X1 OAI21X1_544 ( .A(core_mi_32_), .B(core__abc_21302_new_n2168__bF_buf0), .C(reset_n_bF_buf58), .Y(core__abc_21302_new_n2265_));
OAI21X1 OAI21X1_545 ( .A(core_mi_33_), .B(core__abc_21302_new_n2168__bF_buf11), .C(reset_n_bF_buf57), .Y(core__abc_21302_new_n2268_));
OAI21X1 OAI21X1_546 ( .A(core_mi_34_), .B(core__abc_21302_new_n2168__bF_buf9), .C(reset_n_bF_buf56), .Y(core__abc_21302_new_n2271_));
OAI21X1 OAI21X1_547 ( .A(core_mi_35_), .B(core__abc_21302_new_n2168__bF_buf7), .C(reset_n_bF_buf55), .Y(core__abc_21302_new_n2274_));
OAI21X1 OAI21X1_548 ( .A(core_mi_36_), .B(core__abc_21302_new_n2168__bF_buf5), .C(reset_n_bF_buf54), .Y(core__abc_21302_new_n2277_));
OAI21X1 OAI21X1_549 ( .A(core_mi_37_), .B(core__abc_21302_new_n2168__bF_buf3), .C(reset_n_bF_buf53), .Y(core__abc_21302_new_n2280_));
OAI21X1 OAI21X1_55 ( .A(core_siphash_word_107_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf58), .Y(_abc_19873_new_n1550_));
OAI21X1 OAI21X1_550 ( .A(core_mi_38_), .B(core__abc_21302_new_n2168__bF_buf1), .C(reset_n_bF_buf52), .Y(core__abc_21302_new_n2283_));
OAI21X1 OAI21X1_551 ( .A(core_mi_39_), .B(core__abc_21302_new_n2168__bF_buf12), .C(reset_n_bF_buf51), .Y(core__abc_21302_new_n2286_));
OAI21X1 OAI21X1_552 ( .A(core_mi_40_), .B(core__abc_21302_new_n2168__bF_buf10), .C(reset_n_bF_buf50), .Y(core__abc_21302_new_n2289_));
OAI21X1 OAI21X1_553 ( .A(core_mi_41_), .B(core__abc_21302_new_n2168__bF_buf8), .C(reset_n_bF_buf49), .Y(core__abc_21302_new_n2292_));
OAI21X1 OAI21X1_554 ( .A(core_mi_42_), .B(core__abc_21302_new_n2168__bF_buf6), .C(reset_n_bF_buf48), .Y(core__abc_21302_new_n2295_));
OAI21X1 OAI21X1_555 ( .A(core_mi_43_), .B(core__abc_21302_new_n2168__bF_buf4), .C(reset_n_bF_buf47), .Y(core__abc_21302_new_n2298_));
OAI21X1 OAI21X1_556 ( .A(core_mi_44_), .B(core__abc_21302_new_n2168__bF_buf2), .C(reset_n_bF_buf46), .Y(core__abc_21302_new_n2301_));
OAI21X1 OAI21X1_557 ( .A(core_mi_45_), .B(core__abc_21302_new_n2168__bF_buf0), .C(reset_n_bF_buf45), .Y(core__abc_21302_new_n2304_));
OAI21X1 OAI21X1_558 ( .A(core_mi_46_), .B(core__abc_21302_new_n2168__bF_buf11), .C(reset_n_bF_buf44), .Y(core__abc_21302_new_n2307_));
OAI21X1 OAI21X1_559 ( .A(core_mi_47_), .B(core__abc_21302_new_n2168__bF_buf9), .C(reset_n_bF_buf43), .Y(core__abc_21302_new_n2310_));
OAI21X1 OAI21X1_56 ( .A(core_siphash_word_108_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf57), .Y(_abc_19873_new_n1553_));
OAI21X1 OAI21X1_560 ( .A(core_mi_48_), .B(core__abc_21302_new_n2168__bF_buf7), .C(reset_n_bF_buf42), .Y(core__abc_21302_new_n2313_));
OAI21X1 OAI21X1_561 ( .A(core_mi_49_), .B(core__abc_21302_new_n2168__bF_buf5), .C(reset_n_bF_buf41), .Y(core__abc_21302_new_n2316_));
OAI21X1 OAI21X1_562 ( .A(core_mi_50_), .B(core__abc_21302_new_n2168__bF_buf3), .C(reset_n_bF_buf40), .Y(core__abc_21302_new_n2319_));
OAI21X1 OAI21X1_563 ( .A(core_mi_51_), .B(core__abc_21302_new_n2168__bF_buf1), .C(reset_n_bF_buf39), .Y(core__abc_21302_new_n2322_));
OAI21X1 OAI21X1_564 ( .A(core_mi_52_), .B(core__abc_21302_new_n2168__bF_buf12), .C(reset_n_bF_buf38), .Y(core__abc_21302_new_n2325_));
OAI21X1 OAI21X1_565 ( .A(core_mi_53_), .B(core__abc_21302_new_n2168__bF_buf10), .C(reset_n_bF_buf37), .Y(core__abc_21302_new_n2328_));
OAI21X1 OAI21X1_566 ( .A(core_mi_54_), .B(core__abc_21302_new_n2168__bF_buf8), .C(reset_n_bF_buf36), .Y(core__abc_21302_new_n2331_));
OAI21X1 OAI21X1_567 ( .A(core_mi_55_), .B(core__abc_21302_new_n2168__bF_buf6), .C(reset_n_bF_buf35), .Y(core__abc_21302_new_n2334_));
OAI21X1 OAI21X1_568 ( .A(core_mi_56_), .B(core__abc_21302_new_n2168__bF_buf4), .C(reset_n_bF_buf34), .Y(core__abc_21302_new_n2337_));
OAI21X1 OAI21X1_569 ( .A(core_mi_57_), .B(core__abc_21302_new_n2168__bF_buf2), .C(reset_n_bF_buf33), .Y(core__abc_21302_new_n2340_));
OAI21X1 OAI21X1_57 ( .A(core_siphash_word_109_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf56), .Y(_abc_19873_new_n1556_));
OAI21X1 OAI21X1_570 ( .A(core_mi_58_), .B(core__abc_21302_new_n2168__bF_buf0), .C(reset_n_bF_buf32), .Y(core__abc_21302_new_n2343_));
OAI21X1 OAI21X1_571 ( .A(core_mi_59_), .B(core__abc_21302_new_n2168__bF_buf11), .C(reset_n_bF_buf31), .Y(core__abc_21302_new_n2346_));
OAI21X1 OAI21X1_572 ( .A(core_mi_60_), .B(core__abc_21302_new_n2168__bF_buf9), .C(reset_n_bF_buf30), .Y(core__abc_21302_new_n2349_));
OAI21X1 OAI21X1_573 ( .A(core_mi_61_), .B(core__abc_21302_new_n2168__bF_buf7), .C(reset_n_bF_buf29), .Y(core__abc_21302_new_n2352_));
OAI21X1 OAI21X1_574 ( .A(core_mi_62_), .B(core__abc_21302_new_n2168__bF_buf5), .C(reset_n_bF_buf28), .Y(core__abc_21302_new_n2355_));
OAI21X1 OAI21X1_575 ( .A(core_mi_63_), .B(core__abc_21302_new_n2168__bF_buf3), .C(reset_n_bF_buf27), .Y(core__abc_21302_new_n2358_));
OAI21X1 OAI21X1_576 ( .A(core__abc_21302_new_n1148_), .B(core__abc_21302_new_n1177_), .C(core__abc_21302_new_n1154_), .Y(core__abc_21302_new_n2367_));
OAI21X1 OAI21X1_577 ( .A(core__abc_21302_new_n2138_), .B(core__abc_21302_new_n2367_), .C(core__abc_21302_new_n2366_), .Y(core__abc_21302_new_n2368_));
OAI21X1 OAI21X1_578 ( .A(core__abc_21302_new_n1209_), .B(core__abc_21302_new_n1220_), .C(core__abc_21302_new_n1221_), .Y(core__abc_21302_new_n2375_));
OAI21X1 OAI21X1_579 ( .A(core__abc_21302_new_n1252_), .B(core__abc_21302_new_n2387_), .C(core__abc_21302_new_n1264_), .Y(core__abc_21302_new_n2392_));
OAI21X1 OAI21X1_58 ( .A(core_siphash_word_110_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf55), .Y(_abc_19873_new_n1559_));
OAI21X1 OAI21X1_580 ( .A(core__abc_21302_new_n1274_), .B(core__abc_21302_new_n2382_), .C(core__abc_21302_new_n1284_), .Y(core__abc_21302_new_n2394_));
OAI21X1 OAI21X1_581 ( .A(core__abc_21302_new_n2393_), .B(core__abc_21302_new_n2385_), .C(core__abc_21302_new_n2395_), .Y(core__abc_21302_new_n2396_));
OAI21X1 OAI21X1_582 ( .A(core__abc_21302_new_n2405_), .B(core__abc_21302_new_n2406_), .C(core__abc_21302_new_n2407_), .Y(core__abc_21302_new_n2408_));
OAI21X1 OAI21X1_583 ( .A(core_v1_reg_9_), .B(core_v0_reg_9_), .C(core__abc_21302_new_n2408_), .Y(core__abc_21302_new_n2409_));
OAI21X1 OAI21X1_584 ( .A(core__abc_21302_new_n1313_), .B(core__abc_21302_new_n1325_), .C(core__abc_21302_new_n2410_), .Y(core__abc_21302_new_n2411_));
OAI21X1 OAI21X1_585 ( .A(core__abc_21302_new_n2409_), .B(core__abc_21302_new_n2402_), .C(core__abc_21302_new_n2411_), .Y(core__abc_21302_new_n2412_));
OAI21X1 OAI21X1_586 ( .A(core__abc_21302_new_n2413_), .B(core__abc_21302_new_n1346_), .C(core__abc_21302_new_n2414_), .Y(core__abc_21302_new_n2415_));
OAI21X1 OAI21X1_587 ( .A(core__abc_21302_new_n2404_), .B(core__abc_21302_new_n2397_), .C(core__abc_21302_new_n2419_), .Y(core__abc_21302_new_n2420_));
OAI21X1 OAI21X1_588 ( .A(core__abc_21302_new_n2436_), .B(core__abc_21302_new_n2437_), .C(core__abc_21302_new_n2438_), .Y(core__abc_21302_new_n2439_));
OAI21X1 OAI21X1_589 ( .A(core_v1_reg_17_), .B(core_v0_reg_17_), .C(core__abc_21302_new_n2439_), .Y(core__abc_21302_new_n2440_));
OAI21X1 OAI21X1_59 ( .A(core_siphash_word_111_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf54), .Y(_abc_19873_new_n1561_));
OAI21X1 OAI21X1_590 ( .A(core__abc_21302_new_n2441_), .B(core__abc_21302_new_n1417_), .C(core__abc_21302_new_n2442_), .Y(core__abc_21302_new_n2443_));
OAI21X1 OAI21X1_591 ( .A(core__abc_21302_new_n2440_), .B(core__abc_21302_new_n2435_), .C(core__abc_21302_new_n2444_), .Y(core__abc_21302_new_n2445_));
OAI21X1 OAI21X1_592 ( .A(core__abc_21302_new_n2446_), .B(core__abc_21302_new_n1441_), .C(core__abc_21302_new_n2447_), .Y(core__abc_21302_new_n2448_));
OAI21X1 OAI21X1_593 ( .A(core__abc_21302_new_n2428_), .B(core__abc_21302_new_n2449_), .C(core__abc_21302_new_n2450_), .Y(core__abc_21302_new_n2451_));
OAI21X1 OAI21X1_594 ( .A(core__abc_21302_new_n2453_), .B(core__abc_21302_new_n2454_), .C(core__abc_21302_new_n2455_), .Y(core__abc_21302_new_n2456_));
OAI21X1 OAI21X1_595 ( .A(core_v1_reg_25_), .B(core_v0_reg_25_), .C(core__abc_21302_new_n2456_), .Y(core__abc_21302_new_n2457_));
OAI21X1 OAI21X1_596 ( .A(core__abc_21302_new_n2425_), .B(core__abc_21302_new_n2457_), .C(core__abc_21302_new_n2458_), .Y(core__abc_21302_new_n2459_));
OAI21X1 OAI21X1_597 ( .A(core__abc_21302_new_n2461_), .B(core__abc_21302_new_n1531_), .C(core__abc_21302_new_n1532_), .Y(core__abc_21302_new_n2462_));
OAI21X1 OAI21X1_598 ( .A(core__abc_21302_new_n2427_), .B(core__abc_21302_new_n2452_), .C(core__abc_21302_new_n2465_), .Y(core__abc_21302_new_n2466_));
OAI21X1 OAI21X1_599 ( .A(core__abc_21302_new_n2478_), .B(core__abc_21302_new_n2475_), .C(core__abc_21302_new_n2479_), .Y(core__abc_21302_new_n2480_));
OAI21X1 OAI21X1_6 ( .A(_abc_19873_new_n981_), .B(_abc_19873_new_n918_), .C(_abc_19873_new_n982_), .Y(_abc_19873_new_n983_));
OAI21X1 OAI21X1_60 ( .A(core_siphash_word_112_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf53), .Y(_abc_19873_new_n1564_));
OAI21X1 OAI21X1_600 ( .A(core__abc_21302_new_n2483_), .B(core__abc_21302_new_n2489_), .C(core__abc_21302_new_n2490_), .Y(core__abc_21302_new_n2491_));
OAI21X1 OAI21X1_601 ( .A(core__abc_21302_new_n2497_), .B(core__abc_21302_new_n2492_), .C(core__abc_21302_new_n2504_), .Y(core__abc_21302_new_n2505_));
OAI21X1 OAI21X1_602 ( .A(core__abc_21302_new_n2468_), .B(core__abc_21302_new_n2506_), .C(core__abc_21302_new_n2507_), .Y(core__abc_21302_new_n2508_));
OAI21X1 OAI21X1_603 ( .A(core__abc_21302_new_n1661_), .B(core__abc_21302_new_n1674_), .C(core__abc_21302_new_n1672_), .Y(core__abc_21302_new_n2514_));
OAI21X1 OAI21X1_604 ( .A(core__abc_21302_new_n1213_), .B(core__abc_21302_new_n1226_), .C(core__abc_21302_new_n1224_), .Y(core__abc_21302_new_n2517_));
OAI21X1 OAI21X1_605 ( .A(core__abc_21302_new_n2520_), .B(core__abc_21302_new_n2523_), .C(core__abc_21302_new_n2524_), .Y(core__abc_21302_new_n2525_));
OAI21X1 OAI21X1_606 ( .A(core__abc_21302_new_n1294_), .B(core__abc_21302_new_n1305_), .C(core__abc_21302_new_n1304_), .Y(core__abc_21302_new_n2537_));
OAI21X1 OAI21X1_607 ( .A(core__abc_21302_new_n2538_), .B(core__abc_21302_new_n2536_), .C(core__abc_21302_new_n2540_), .Y(core__abc_21302_new_n2541_));
OAI21X1 OAI21X1_608 ( .A(core__abc_21302_new_n1350_), .B(core__abc_21302_new_n1351_), .C(core__abc_21302_new_n1337_), .Y(core__abc_21302_new_n2542_));
OAI21X1 OAI21X1_609 ( .A(core_v2_reg_13_), .B(core_v3_reg_13_), .C(core__abc_21302_new_n2542_), .Y(core__abc_21302_new_n2543_));
OAI21X1 OAI21X1_61 ( .A(core_siphash_word_113_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf52), .Y(_abc_19873_new_n1567_));
OAI21X1 OAI21X1_610 ( .A(core__abc_21302_new_n2543_), .B(core__abc_21302_new_n2527_), .C(core__abc_21302_new_n2545_), .Y(core__abc_21302_new_n2546_));
OAI21X1 OAI21X1_611 ( .A(core__abc_21302_new_n2526_), .B(core__abc_21302_new_n2533_), .C(core__abc_21302_new_n2547_), .Y(core__abc_21302_new_n2548_));
OAI21X1 OAI21X1_612 ( .A(core__abc_21302_new_n1385_), .B(core__abc_21302_new_n1400_), .C(core__abc_21302_new_n1396_), .Y(core__abc_21302_new_n2571_));
OAI21X1 OAI21X1_613 ( .A(core__abc_21302_new_n1408_), .B(core__abc_21302_new_n1424_), .C(core__abc_21302_new_n1420_), .Y(core__abc_21302_new_n2572_));
OAI21X1 OAI21X1_614 ( .A(core__abc_21302_new_n1432_), .B(core__abc_21302_new_n1448_), .C(core__abc_21302_new_n1444_), .Y(core__abc_21302_new_n2578_));
OAI21X1 OAI21X1_615 ( .A(core__abc_21302_new_n2577_), .B(core__abc_21302_new_n2579_), .C(core__abc_21302_new_n2584_), .Y(core__abc_21302_new_n2585_));
OAI21X1 OAI21X1_616 ( .A(core_v2_reg_31_), .B(core_v3_reg_31_), .C(core__abc_21302_new_n2589_), .Y(core__abc_21302_new_n2590_));
OAI21X1 OAI21X1_617 ( .A(core__abc_21302_new_n2587_), .B(core__abc_21302_new_n2588_), .C(core__abc_21302_new_n2590_), .Y(core__abc_21302_new_n2591_));
OAI21X1 OAI21X1_618 ( .A(core_v2_reg_25_), .B(core_v3_reg_25_), .C(core__abc_21302_new_n1478_), .Y(core__abc_21302_new_n2594_));
OAI21X1 OAI21X1_619 ( .A(core__abc_21302_new_n1487_), .B(core__abc_21302_new_n1488_), .C(core__abc_21302_new_n2594_), .Y(core__abc_21302_new_n2595_));
OAI21X1 OAI21X1_62 ( .A(core_siphash_word_114_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf51), .Y(_abc_19873_new_n1570_));
OAI21X1 OAI21X1_620 ( .A(core__abc_21302_new_n1498_), .B(core__abc_21302_new_n1514_), .C(core__abc_21302_new_n1510_), .Y(core__abc_21302_new_n2596_));
OAI21X1 OAI21X1_621 ( .A(core__abc_21302_new_n1522_), .B(core__abc_21302_new_n1539_), .C(core__abc_21302_new_n1535_), .Y(core__abc_21302_new_n2598_));
OAI21X1 OAI21X1_622 ( .A(core__abc_21302_new_n2592_), .B(core__abc_21302_new_n2597_), .C(core__abc_21302_new_n2599_), .Y(core__abc_21302_new_n2600_));
OAI21X1 OAI21X1_623 ( .A(core__abc_21302_new_n2556_), .B(core__abc_21302_new_n2586_), .C(core__abc_21302_new_n2601_), .Y(core__abc_21302_new_n2602_));
OAI21X1 OAI21X1_624 ( .A(core__abc_21302_new_n2602_), .B(core__abc_21302_new_n2568_), .C(core__abc_21302_new_n2609_), .Y(core__abc_21302_new_n2610_));
OAI21X1 OAI21X1_625 ( .A(core__abc_21302_new_n1568_), .B(core__abc_21302_new_n1583_), .C(core__abc_21302_new_n1581_), .Y(core__abc_21302_new_n2611_));
OAI21X1 OAI21X1_626 ( .A(core__abc_21302_new_n1596_), .B(core__abc_21302_new_n1609_), .C(core__abc_21302_new_n1605_), .Y(core__abc_21302_new_n2612_));
OAI21X1 OAI21X1_627 ( .A(core__abc_21302_new_n1618_), .B(core__abc_21302_new_n1632_), .C(core__abc_21302_new_n1630_), .Y(core__abc_21302_new_n2617_));
OAI21X1 OAI21X1_628 ( .A(core__abc_21302_new_n2514_), .B(core__abc_21302_new_n2623_), .C(core__abc_21302_new_n1686_), .Y(core__abc_21302_new_n2624_));
OAI21X1 OAI21X1_629 ( .A(core__abc_21302_new_n1684_), .B(core__abc_21302_new_n2626_), .C(core__abc_21302_new_n1697_), .Y(core__abc_21302_new_n2627_));
OAI21X1 OAI21X1_63 ( .A(core_siphash_word_115_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf50), .Y(_abc_19873_new_n1573_));
OAI21X1 OAI21X1_630 ( .A(core__abc_21302_new_n1684_), .B(core__abc_21302_new_n2626_), .C(core__abc_21302_new_n2513_), .Y(core__abc_21302_new_n2630_));
OAI21X1 OAI21X1_631 ( .A(core__abc_21302_new_n2512_), .B(core__abc_21302_new_n2632_), .C(core__abc_21302_new_n2634__bF_buf8), .Y(core__abc_21302_new_n2635_));
OAI21X1 OAI21X1_632 ( .A(core__abc_21302_new_n2168__bF_buf1), .B(core__abc_21302_new_n2642_), .C(core__abc_21302_new_n2369__bF_buf6), .Y(core__abc_21302_new_n2643_));
OAI21X1 OAI21X1_633 ( .A(core__abc_21302_new_n2644_), .B(core__abc_21302_new_n2636_), .C(reset_n_bF_buf26), .Y(core__abc_21302_new_n2645_));
OAI21X1 OAI21X1_634 ( .A(core__abc_21302_new_n2371_), .B(core__abc_21302_new_n2467_), .C(core__abc_21302_new_n2648_), .Y(core__abc_21302_new_n2649_));
OAI21X1 OAI21X1_635 ( .A(core__abc_21302_new_n1566_), .B(core__abc_21302_new_n2468_), .C(core__abc_21302_new_n2647_), .Y(core__abc_21302_new_n2650_));
OAI21X1 OAI21X1_636 ( .A(core__abc_21302_new_n2659_), .B(core__abc_21302_new_n2660_), .C(core__abc_21302_new_n2661_), .Y(core__abc_21302_new_n2662_));
OAI21X1 OAI21X1_637 ( .A(core__abc_21302_new_n1706_), .B(core__abc_21302_new_n1708_), .C(core__abc_21302_new_n2665_), .Y(core__abc_21302_new_n2666_));
OAI21X1 OAI21X1_638 ( .A(core__abc_21302_new_n2662_), .B(core__abc_21302_new_n2664_), .C(core__abc_21302_new_n1709_), .Y(core__abc_21302_new_n2667_));
OAI21X1 OAI21X1_639 ( .A(core__abc_21302_new_n2658_), .B(core__abc_21302_new_n2672_), .C(core__abc_21302_new_n2674_), .Y(core__abc_21302_new_n2675_));
OAI21X1 OAI21X1_64 ( .A(core_siphash_word_116_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf49), .Y(_abc_19873_new_n1576_));
OAI21X1 OAI21X1_640 ( .A(core_v3_reg_1_), .B(core__abc_21302_new_n2369__bF_buf5), .C(reset_n_bF_buf25), .Y(core__abc_21302_new_n2679_));
OAI21X1 OAI21X1_641 ( .A(core__abc_21302_new_n2511_), .B(core__abc_21302_new_n2654_), .C(core__abc_21302_new_n2655_), .Y(core__abc_21302_new_n2681_));
OAI21X1 OAI21X1_642 ( .A(core__abc_21302_new_n1565_), .B(core__abc_21302_new_n1580_), .C(core__abc_21302_new_n1579_), .Y(core__abc_21302_new_n2684_));
OAI21X1 OAI21X1_643 ( .A(core__abc_21302_new_n2683_), .B(core__abc_21302_new_n2467_), .C(core__abc_21302_new_n2685_), .Y(core__abc_21302_new_n2686_));
OAI21X1 OAI21X1_644 ( .A(core__abc_21302_new_n2689_), .B(core__abc_21302_new_n2688_), .C(core__abc_21302_new_n2693_), .Y(core__abc_21302_new_n2694_));
OAI21X1 OAI21X1_645 ( .A(core__abc_21302_new_n2702_), .B(core__abc_21302_new_n2703_), .C(core__abc_21302_new_n2667_), .Y(core__abc_21302_new_n2704_));
OAI21X1 OAI21X1_646 ( .A(core__abc_21302_new_n2700_), .B(core__abc_21302_new_n2710_), .C(core__abc_21302_new_n2711_), .Y(core__abc_21302_new_n2712_));
OAI21X1 OAI21X1_647 ( .A(core__abc_21302_new_n2714_), .B(core__abc_21302_new_n2640__bF_buf9), .C(core__abc_21302_new_n2369__bF_buf4), .Y(core__abc_21302_new_n2715_));
OAI21X1 OAI21X1_648 ( .A(core_v3_reg_2_), .B(core__abc_21302_new_n2369__bF_buf3), .C(reset_n_bF_buf24), .Y(core__abc_21302_new_n2717_));
OAI21X1 OAI21X1_649 ( .A(core__abc_21302_new_n2662_), .B(core__abc_21302_new_n2664_), .C(core__abc_21302_new_n2720_), .Y(core__abc_21302_new_n2721_));
OAI21X1 OAI21X1_65 ( .A(core_siphash_word_117_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf48), .Y(_abc_19873_new_n1579_));
OAI21X1 OAI21X1_650 ( .A(core__abc_21302_new_n1707_), .B(core__abc_21302_new_n1717_), .C(core__abc_21302_new_n1718_), .Y(core__abc_21302_new_n2722_));
OAI21X1 OAI21X1_651 ( .A(core__abc_21302_new_n2719_), .B(core__abc_21302_new_n2665_), .C(core__abc_21302_new_n2723_), .Y(core__abc_21302_new_n2726_));
OAI21X1 OAI21X1_652 ( .A(core__abc_21302_new_n2724_), .B(core__abc_21302_new_n2727_), .C(core__abc_21302_new_n1549_), .Y(core__abc_21302_new_n2728_));
OAI21X1 OAI21X1_653 ( .A(core__abc_21302_new_n2736_), .B(core__abc_21302_new_n2688_), .C(core__abc_21302_new_n2737_), .Y(core__abc_21302_new_n2738_));
OAI21X1 OAI21X1_654 ( .A(core__abc_21302_new_n2741_), .B(core__abc_21302_new_n2742_), .C(core__abc_21302_new_n2690_), .Y(core__abc_21302_new_n2743_));
OAI21X1 OAI21X1_655 ( .A(core__abc_21302_new_n2673__bF_buf9), .B(core__abc_21302_new_n2752_), .C(core__abc_21302_new_n2733_), .Y(core__abc_21302_new_n2753_));
OAI21X1 OAI21X1_656 ( .A(core__abc_21302_new_n2733_), .B(core__abc_21302_new_n2754_), .C(core__abc_21302_new_n2753_), .Y(core__abc_21302_new_n2755_));
OAI21X1 OAI21X1_657 ( .A(core__abc_21302_new_n2757_), .B(core__abc_21302_new_n2640__bF_buf8), .C(core__abc_21302_new_n2369__bF_buf2), .Y(core__abc_21302_new_n2758_));
OAI21X1 OAI21X1_658 ( .A(core_v3_reg_3_), .B(core__abc_21302_new_n2369__bF_buf1), .C(reset_n_bF_buf23), .Y(core__abc_21302_new_n2760_));
OAI21X1 OAI21X1_659 ( .A(core__abc_21302_new_n2766_), .B(core__abc_21302_new_n2467_), .C(core__abc_21302_new_n2764_), .Y(core__abc_21302_new_n2767_));
OAI21X1 OAI21X1_66 ( .A(core_siphash_word_118_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf47), .Y(_abc_19873_new_n1582_));
OAI21X1 OAI21X1_660 ( .A(core__abc_21302_new_n1254_), .B(core__abc_21302_new_n1255_), .C(core__abc_21302_new_n2770_), .Y(core__abc_21302_new_n2771_));
OAI21X1 OAI21X1_661 ( .A(core__abc_21302_new_n2769_), .B(core__abc_21302_new_n2768_), .C(core__abc_21302_new_n2775_), .Y(core__abc_21302_new_n2776_));
OAI21X1 OAI21X1_662 ( .A(core__abc_21302_new_n2748_), .B(core__abc_21302_new_n2734_), .C(core__abc_21302_new_n2747_), .Y(core__abc_21302_new_n2780_));
OAI21X1 OAI21X1_663 ( .A(core__abc_21302_new_n1731_), .B(core__abc_21302_new_n2724_), .C(core__abc_21302_new_n2783_), .Y(core__abc_21302_new_n2784_));
OAI21X1 OAI21X1_664 ( .A(core__abc_21302_new_n1731_), .B(core__abc_21302_new_n2724_), .C(core__abc_21302_new_n1743_), .Y(core__abc_21302_new_n2787_));
OAI21X1 OAI21X1_665 ( .A(core__abc_21302_new_n2781_), .B(core__abc_21302_new_n2789_), .C(core__abc_21302_new_n2634__bF_buf6), .Y(core__abc_21302_new_n2791_));
OAI21X1 OAI21X1_666 ( .A(core_key_68_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n2369__bF_buf0), .Y(core__abc_21302_new_n2793_));
OAI21X1 OAI21X1_667 ( .A(core__abc_21302_new_n2790_), .B(core__abc_21302_new_n2791_), .C(core__abc_21302_new_n2794_), .Y(core__abc_21302_new_n2795_));
OAI21X1 OAI21X1_668 ( .A(core_v3_reg_4_), .B(core__abc_21302_new_n2369__bF_buf7), .C(core__abc_21302_new_n2795_), .Y(core__abc_21302_new_n2796_));
OAI21X1 OAI21X1_669 ( .A(core__abc_21302_new_n2779_), .B(core__abc_21302_new_n2798_), .C(core__abc_21302_new_n2778_), .Y(core__abc_21302_new_n2799_));
OAI21X1 OAI21X1_67 ( .A(core_siphash_word_119_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf46), .Y(_abc_19873_new_n1584_));
OAI21X1 OAI21X1_670 ( .A(core__abc_21302_new_n1615_), .B(core__abc_21302_new_n2768_), .C(core__abc_21302_new_n1629_), .Y(core__abc_21302_new_n2803_));
OAI21X1 OAI21X1_671 ( .A(core__abc_21302_new_n2602_), .B(core__abc_21302_new_n2568_), .C(core__abc_21302_new_n2817_), .Y(core__abc_21302_new_n2818_));
OAI21X1 OAI21X1_672 ( .A(core__abc_21302_new_n1730_), .B(core__abc_21302_new_n1740_), .C(core__abc_21302_new_n1741_), .Y(core__abc_21302_new_n2820_));
OAI21X1 OAI21X1_673 ( .A(core__abc_21302_new_n2619_), .B(core__abc_21302_new_n2614_), .C(core__abc_21302_new_n2816_), .Y(core__abc_21302_new_n2823_));
OAI21X1 OAI21X1_674 ( .A(core__abc_21302_new_n2830_), .B(core__abc_21302_new_n2813_), .C(core__abc_21302_new_n2634__bF_buf5), .Y(core__abc_21302_new_n2832_));
OAI21X1 OAI21X1_675 ( .A(core_key_69_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n2369__bF_buf6), .Y(core__abc_21302_new_n2834_));
OAI21X1 OAI21X1_676 ( .A(core__abc_21302_new_n2831_), .B(core__abc_21302_new_n2832_), .C(core__abc_21302_new_n2835_), .Y(core__abc_21302_new_n2836_));
OAI21X1 OAI21X1_677 ( .A(core_v3_reg_5_), .B(core__abc_21302_new_n2369__bF_buf5), .C(core__abc_21302_new_n2836_), .Y(core__abc_21302_new_n2837_));
OAI21X1 OAI21X1_678 ( .A(core_v1_reg_37_), .B(core_v0_reg_37_), .C(core__abc_21302_new_n1615_), .Y(core__abc_21302_new_n2839_));
OAI21X1 OAI21X1_679 ( .A(core__abc_21302_new_n1625_), .B(core__abc_21302_new_n1626_), .C(core__abc_21302_new_n2839_), .Y(core__abc_21302_new_n2840_));
OAI21X1 OAI21X1_68 ( .A(core_siphash_word_120_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf45), .Y(_abc_19873_new_n1587_));
OAI21X1 OAI21X1_680 ( .A(core__abc_21302_new_n2846_), .B(core__abc_21302_new_n2845_), .C(core__abc_21302_new_n1278_), .Y(core__abc_21302_new_n2847_));
OAI21X1 OAI21X1_681 ( .A(core__abc_21302_new_n1276_), .B(core__abc_21302_new_n1277_), .C(core__abc_21302_new_n2848_), .Y(core__abc_21302_new_n2849_));
OAI21X1 OAI21X1_682 ( .A(core__abc_21302_new_n2843_), .B(core__abc_21302_new_n2844_), .C(core__abc_21302_new_n2851_), .Y(core__abc_21302_new_n2852_));
OAI21X1 OAI21X1_683 ( .A(core__abc_21302_new_n2778_), .B(core__abc_21302_new_n2859_), .C(core__abc_21302_new_n2858_), .Y(core__abc_21302_new_n2860_));
OAI21X1 OAI21X1_684 ( .A(core__abc_21302_new_n1762_), .B(core__abc_21302_new_n1765_), .C(core__abc_21302_new_n2864_), .Y(core__abc_21302_new_n2865_));
OAI21X1 OAI21X1_685 ( .A(core__abc_21302_new_n1755_), .B(core__abc_21302_new_n2828_), .C(core__abc_21302_new_n1766_), .Y(core__abc_21302_new_n2866_));
OAI21X1 OAI21X1_686 ( .A(core__abc_21302_new_n2828_), .B(core__abc_21302_new_n2865_), .C(core__abc_21302_new_n2866_), .Y(core__abc_21302_new_n2867_));
OAI21X1 OAI21X1_687 ( .A(core__abc_21302_new_n2863_), .B(core__abc_21302_new_n2871_), .C(core__abc_21302_new_n2872_), .Y(core__abc_21302_new_n2873_));
OAI21X1 OAI21X1_688 ( .A(core_key_70_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n2369__bF_buf4), .Y(core__abc_21302_new_n2875_));
OAI21X1 OAI21X1_689 ( .A(core_v3_reg_6_), .B(core__abc_21302_new_n2369__bF_buf3), .C(reset_n_bF_buf22), .Y(core__abc_21302_new_n2877_));
OAI21X1 OAI21X1_69 ( .A(core_siphash_word_121_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf44), .Y(_abc_19873_new_n1590_));
OAI21X1 OAI21X1_690 ( .A(core__abc_21302_new_n2882_), .B(core__abc_21302_new_n2883_), .C(core__abc_21302_new_n2847_), .Y(core__abc_21302_new_n2884_));
OAI21X1 OAI21X1_691 ( .A(core__abc_21302_new_n2856_), .B(core__abc_21302_new_n2862_), .C(core__abc_21302_new_n2855_), .Y(core__abc_21302_new_n2893_));
OAI21X1 OAI21X1_692 ( .A(core__abc_21302_new_n2902_), .B(core__abc_21302_new_n2901_), .C(core__abc_21302_new_n1594_), .Y(core__abc_21302_new_n2903_));
OAI21X1 OAI21X1_693 ( .A(core__abc_21302_new_n2906_), .B(core__abc_21302_new_n2894_), .C(core__abc_21302_new_n2634__bF_buf4), .Y(core__abc_21302_new_n2908_));
OAI21X1 OAI21X1_694 ( .A(core__abc_21302_new_n2168__bF_buf12), .B(core__abc_21302_new_n2909_), .C(core__abc_21302_new_n2369__bF_buf2), .Y(core__abc_21302_new_n2910_));
OAI21X1 OAI21X1_695 ( .A(core__abc_21302_new_n2907_), .B(core__abc_21302_new_n2908_), .C(core__abc_21302_new_n2911_), .Y(core__abc_21302_new_n2912_));
OAI21X1 OAI21X1_696 ( .A(core_v3_reg_7_), .B(core__abc_21302_new_n2369__bF_buf1), .C(core__abc_21302_new_n2912_), .Y(core__abc_21302_new_n2913_));
OAI21X1 OAI21X1_697 ( .A(core__abc_21302_new_n2916_), .B(core__abc_21302_new_n2862_), .C(core__abc_21302_new_n2918_), .Y(core__abc_21302_new_n2919_));
OAI21X1 OAI21X1_698 ( .A(core__abc_21302_new_n2922_), .B(core__abc_21302_new_n2764_), .C(core__abc_21302_new_n2925_), .Y(core__abc_21302_new_n2926_));
OAI21X1 OAI21X1_699 ( .A(core__abc_21302_new_n2765_), .B(core__abc_21302_new_n2685_), .C(core__abc_21302_new_n2763_), .Y(core__abc_21302_new_n2930_));
OAI21X1 OAI21X1_7 ( .A(_abc_19873_new_n989_), .B(_abc_19873_new_n960__bF_buf3), .C(_abc_19873_new_n990_), .Y(_abc_19873_new_n991_));
OAI21X1 OAI21X1_70 ( .A(core_siphash_word_122_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf43), .Y(_abc_19873_new_n1592_));
OAI21X1 OAI21X1_700 ( .A(core__abc_21302_new_n2934_), .B(core__abc_21302_new_n2467_), .C(core__abc_21302_new_n2933_), .Y(core__abc_21302_new_n2935_));
OAI21X1 OAI21X1_701 ( .A(core__abc_21302_new_n2936_), .B(core__abc_21302_new_n2929_), .C(core__abc_21302_new_n2940_), .Y(core__abc_21302_new_n2943_));
OAI21X1 OAI21X1_702 ( .A(core__abc_21302_new_n2895_), .B(core__abc_21302_new_n2900_), .C(core__abc_21302_new_n1775_), .Y(core__abc_21302_new_n2949_));
OAI21X1 OAI21X1_703 ( .A(core__abc_21302_new_n1786_), .B(core__abc_21302_new_n1787_), .C(core__abc_21302_new_n2949_), .Y(core__abc_21302_new_n2951_));
OAI21X1 OAI21X1_704 ( .A(core__abc_21302_new_n2947_), .B(core__abc_21302_new_n2956_), .C(core__abc_21302_new_n2957_), .Y(core__abc_21302_new_n2958_));
OAI21X1 OAI21X1_705 ( .A(core__abc_21302_new_n2168__bF_buf11), .B(core__abc_21302_new_n2959_), .C(core__abc_21302_new_n2958_), .Y(core__abc_21302_new_n2960_));
OAI21X1 OAI21X1_706 ( .A(core__abc_21302_new_n2915_), .B(core__abc_21302_new_n2960_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n2961_));
OAI21X1 OAI21X1_707 ( .A(core_v3_reg_8_), .B(core__abc_21302_new_n2369__bF_buf0), .C(reset_n_bF_buf21), .Y(core__abc_21302_new_n2962_));
OAI21X1 OAI21X1_708 ( .A(core__abc_21302_new_n1659_), .B(core__abc_21302_new_n2929_), .C(core__abc_21302_new_n2966_), .Y(core__abc_21302_new_n2967_));
OAI21X1 OAI21X1_709 ( .A(core__abc_21302_new_n1296_), .B(core__abc_21302_new_n2526_), .C(core__abc_21302_new_n1294_), .Y(core__abc_21302_new_n2969_));
OAI21X1 OAI21X1_71 ( .A(core_siphash_word_123_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf42), .Y(_abc_19873_new_n1594_));
OAI21X1 OAI21X1_710 ( .A(core__abc_21302_new_n1765_), .B(core__abc_21302_new_n2898_), .C(core__abc_21302_new_n2981_), .Y(core__abc_21302_new_n2984_));
OAI21X1 OAI21X1_711 ( .A(core__abc_21302_new_n1798_), .B(core__abc_21302_new_n1801_), .C(core__abc_21302_new_n2987_), .Y(core__abc_21302_new_n2988_));
OAI21X1 OAI21X1_712 ( .A(core__abc_21302_new_n2986_), .B(core__abc_21302_new_n2983_), .C(core__abc_21302_new_n1802_), .Y(core__abc_21302_new_n2989_));
OAI21X1 OAI21X1_713 ( .A(core__abc_21302_new_n2991_), .B(core__abc_21302_new_n2979_), .C(core__abc_21302_new_n2634__bF_buf3), .Y(core__abc_21302_new_n2993_));
OAI21X1 OAI21X1_714 ( .A(core__abc_21302_new_n2168__bF_buf10), .B(core__abc_21302_new_n2994_), .C(core__abc_21302_new_n2369__bF_buf6), .Y(core__abc_21302_new_n2995_));
OAI21X1 OAI21X1_715 ( .A(core__abc_21302_new_n2992_), .B(core__abc_21302_new_n2993_), .C(core__abc_21302_new_n2996_), .Y(core__abc_21302_new_n2997_));
OAI21X1 OAI21X1_716 ( .A(core_v3_reg_9_), .B(core__abc_21302_new_n2369__bF_buf5), .C(core__abc_21302_new_n2997_), .Y(core__abc_21302_new_n2998_));
OAI21X1 OAI21X1_717 ( .A(core__abc_21302_new_n3002_), .B(core__abc_21302_new_n3001_), .C(core__abc_21302_new_n3004_), .Y(core__abc_21302_new_n3005_));
OAI21X1 OAI21X1_718 ( .A(core__abc_21302_new_n2525_), .B(core__abc_21302_new_n3015_), .C(core__abc_21302_new_n2530_), .Y(core__abc_21302_new_n3016_));
OAI21X1 OAI21X1_719 ( .A(core__abc_21302_new_n3013_), .B(core__abc_21302_new_n3014_), .C(core__abc_21302_new_n3019_), .Y(core__abc_21302_new_n3020_));
OAI21X1 OAI21X1_72 ( .A(core_siphash_word_124_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf41), .Y(_abc_19873_new_n1597_));
OAI21X1 OAI21X1_720 ( .A(core__abc_21302_new_n1799_), .B(core__abc_21302_new_n1800_), .C(core__abc_21302_new_n2989_), .Y(core__abc_21302_new_n3026_));
OAI21X1 OAI21X1_721 ( .A(core__abc_21302_new_n3025_), .B(core__abc_21302_new_n3034_), .C(core__abc_21302_new_n3035_), .Y(core__abc_21302_new_n3036_));
OAI21X1 OAI21X1_722 ( .A(core__abc_21302_new_n2168__bF_buf9), .B(core__abc_21302_new_n3037_), .C(core__abc_21302_new_n3036_), .Y(core__abc_21302_new_n3038_));
OAI21X1 OAI21X1_723 ( .A(core__abc_21302_new_n3000_), .B(core__abc_21302_new_n3038_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n3039_));
OAI21X1 OAI21X1_724 ( .A(core_v3_reg_10_), .B(core__abc_21302_new_n2369__bF_buf4), .C(reset_n_bF_buf20), .Y(core__abc_21302_new_n3040_));
OAI21X1 OAI21X1_725 ( .A(core__abc_21302_new_n3042_), .B(core__abc_21302_new_n3019_), .C(core__abc_21302_new_n3043_), .Y(core__abc_21302_new_n3044_));
OAI21X1 OAI21X1_726 ( .A(core__abc_21302_new_n1681_), .B(core__abc_21302_new_n3013_), .C(core__abc_21302_new_n3047_), .Y(core__abc_21302_new_n3048_));
OAI21X1 OAI21X1_727 ( .A(core__abc_21302_new_n1316_), .B(core__abc_21302_new_n1317_), .C(core__abc_21302_new_n3049_), .Y(core__abc_21302_new_n3050_));
OAI21X1 OAI21X1_728 ( .A(core__abc_21302_new_n3064_), .B(core__abc_21302_new_n2987_), .C(core__abc_21302_new_n3065_), .Y(core__abc_21302_new_n3066_));
OAI21X1 OAI21X1_729 ( .A(core__abc_21302_new_n3069_), .B(core__abc_21302_new_n3068_), .C(core__abc_21302_new_n3063_), .Y(core__abc_21302_new_n3070_));
OAI21X1 OAI21X1_73 ( .A(core_siphash_word_125_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf40), .Y(_abc_19873_new_n1599_));
OAI21X1 OAI21X1_730 ( .A(core__abc_21302_new_n3062_), .B(core__abc_21302_new_n3074_), .C(core__abc_21302_new_n3075_), .Y(core__abc_21302_new_n3076_));
OAI21X1 OAI21X1_731 ( .A(core__abc_21302_new_n2168__bF_buf8), .B(core__abc_21302_new_n3077_), .C(core__abc_21302_new_n2369__bF_buf2), .Y(core__abc_21302_new_n3078_));
OAI21X1 OAI21X1_732 ( .A(core_v3_reg_11_), .B(core__abc_21302_new_n2369__bF_buf1), .C(reset_n_bF_buf19), .Y(core__abc_21302_new_n3080_));
OAI21X1 OAI21X1_733 ( .A(core__abc_21302_new_n3042_), .B(core__abc_21302_new_n3019_), .C(core__abc_21302_new_n3060_), .Y(core__abc_21302_new_n3084_));
OAI21X1 OAI21X1_734 ( .A(core__abc_21302_new_n3004_), .B(core__abc_21302_new_n3083_), .C(core__abc_21302_new_n3085_), .Y(core__abc_21302_new_n3086_));
OAI21X1 OAI21X1_735 ( .A(core__abc_21302_new_n3089_), .B(core__abc_21302_new_n3001_), .C(core__abc_21302_new_n3087_), .Y(core__abc_21302_new_n3090_));
OAI21X1 OAI21X1_736 ( .A(core__abc_21302_new_n3010_), .B(core__abc_21302_new_n3091_), .C(core__abc_21302_new_n3092_), .Y(core__abc_21302_new_n3093_));
OAI21X1 OAI21X1_737 ( .A(core__abc_21302_new_n3096_), .B(core__abc_21302_new_n2928_), .C(core__abc_21302_new_n3094_), .Y(core__abc_21302_new_n3097_));
OAI21X1 OAI21X1_738 ( .A(core__abc_21302_new_n1702_), .B(core__abc_21302_new_n1704_), .C(core__abc_21302_new_n3099_), .Y(core__abc_21302_new_n3100_));
OAI21X1 OAI21X1_739 ( .A(core__abc_21302_new_n2536_), .B(core__abc_21302_new_n3016_), .C(core__abc_21302_new_n3102_), .Y(core__abc_21302_new_n3103_));
OAI21X1 OAI21X1_74 ( .A(core_siphash_word_126_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf39), .Y(_abc_19873_new_n1602_));
OAI21X1 OAI21X1_740 ( .A(core__abc_21302_new_n1825_), .B(core__abc_21302_new_n3068_), .C(core__abc_21302_new_n3114_), .Y(core__abc_21302_new_n3115_));
OAI21X1 OAI21X1_741 ( .A(core__abc_21302_new_n3110_), .B(core__abc_21302_new_n3121_), .C(core__abc_21302_new_n3122_), .Y(core__abc_21302_new_n3123_));
OAI21X1 OAI21X1_742 ( .A(core__abc_21302_new_n2168__bF_buf7), .B(core__abc_21302_new_n3124_), .C(core__abc_21302_new_n3123_), .Y(core__abc_21302_new_n3125_));
OAI21X1 OAI21X1_743 ( .A(core__abc_21302_new_n3082_), .B(core__abc_21302_new_n3125_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n3126_));
OAI21X1 OAI21X1_744 ( .A(core_v3_reg_12_), .B(core__abc_21302_new_n2369__bF_buf0), .C(reset_n_bF_buf18), .Y(core__abc_21302_new_n3127_));
OAI21X1 OAI21X1_745 ( .A(core__abc_21302_new_n1704_), .B(core__abc_21302_new_n3131_), .C(core__abc_21302_new_n3134_), .Y(core__abc_21302_new_n3135_));
OAI21X1 OAI21X1_746 ( .A(core__abc_21302_new_n1338_), .B(core__abc_21302_new_n1339_), .C(core__abc_21302_new_n3104_), .Y(core__abc_21302_new_n3138_));
OAI21X1 OAI21X1_747 ( .A(core__abc_21302_new_n3101_), .B(core__abc_21302_new_n3108_), .C(core__abc_21302_new_n3150_), .Y(core__abc_21302_new_n3151_));
OAI21X1 OAI21X1_748 ( .A(core__abc_21302_new_n1835_), .B(core__abc_21302_new_n3112_), .C(core__abc_21302_new_n3156_), .Y(core__abc_21302_new_n3157_));
OAI21X1 OAI21X1_749 ( .A(core__abc_21302_new_n3154_), .B(core__abc_21302_new_n3167_), .C(core__abc_21302_new_n3168_), .Y(core__abc_21302_new_n3169_));
OAI21X1 OAI21X1_75 ( .A(core_siphash_word_127_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf38), .Y(_abc_19873_new_n1604_));
OAI21X1 OAI21X1_750 ( .A(core__abc_21302_new_n2168__bF_buf6), .B(core__abc_21302_new_n3170_), .C(core__abc_21302_new_n3169_), .Y(core__abc_21302_new_n3171_));
OAI21X1 OAI21X1_751 ( .A(core__abc_21302_new_n3129_), .B(core__abc_21302_new_n3171_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n3172_));
OAI21X1 OAI21X1_752 ( .A(core_v3_reg_13_), .B(core__abc_21302_new_n2369__bF_buf6), .C(reset_n_bF_buf17), .Y(core__abc_21302_new_n3173_));
OAI21X1 OAI21X1_753 ( .A(core__abc_21302_new_n1703_), .B(core__abc_21302_new_n1716_), .C(core__abc_21302_new_n1715_), .Y(core__abc_21302_new_n3178_));
OAI21X1 OAI21X1_754 ( .A(core__abc_21302_new_n3179_), .B(core__abc_21302_new_n3099_), .C(core__abc_21302_new_n3183_), .Y(core__abc_21302_new_n3184_));
OAI21X1 OAI21X1_755 ( .A(core__abc_21302_new_n2525_), .B(core__abc_21302_new_n3015_), .C(core__abc_21302_new_n2532_), .Y(core__abc_21302_new_n3188_));
OAI21X1 OAI21X1_756 ( .A(core__abc_21302_new_n3187_), .B(core__abc_21302_new_n3189_), .C(core__abc_21302_new_n1365_), .Y(core__abc_21302_new_n3192_));
OAI21X1 OAI21X1_757 ( .A(core__abc_21302_new_n3193_), .B(core__abc_21302_new_n3191_), .C(core__abc_21302_new_n1930_), .Y(core__abc_21302_new_n3194_));
OAI21X1 OAI21X1_758 ( .A(core__abc_21302_new_n3185_), .B(core__abc_21302_new_n3182_), .C(core__abc_21302_new_n3197_), .Y(core__abc_21302_new_n3198_));
OAI21X1 OAI21X1_759 ( .A(core__abc_21302_new_n1725_), .B(core__abc_21302_new_n1727_), .C(core__abc_21302_new_n3181_), .Y(core__abc_21302_new_n3200_));
OAI21X1 OAI21X1_76 ( .A(core_siphash_word_64_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf37), .Y(_abc_19873_new_n1607_));
OAI21X1 OAI21X1_760 ( .A(core__abc_21302_new_n1850_), .B(core__abc_21302_new_n1851_), .C(core__abc_21302_new_n3162_), .Y(core__abc_21302_new_n3206_));
OAI21X1 OAI21X1_761 ( .A(core__abc_21302_new_n1865_), .B(core__abc_21302_new_n3206_), .C(core__abc_21302_new_n3208_), .Y(core__abc_21302_new_n3209_));
OAI21X1 OAI21X1_762 ( .A(core__abc_21302_new_n3205_), .B(core__abc_21302_new_n3215_), .C(core__abc_21302_new_n3216_), .Y(core__abc_21302_new_n3217_));
OAI21X1 OAI21X1_763 ( .A(core__abc_21302_new_n2168__bF_buf5), .B(core__abc_21302_new_n3218_), .C(core__abc_21302_new_n3217_), .Y(core__abc_21302_new_n3219_));
OAI21X1 OAI21X1_764 ( .A(core__abc_21302_new_n3175_), .B(core__abc_21302_new_n3219_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n3220_));
OAI21X1 OAI21X1_765 ( .A(core_v3_reg_14_), .B(core__abc_21302_new_n2369__bF_buf4), .C(reset_n_bF_buf16), .Y(core__abc_21302_new_n3221_));
OAI21X1 OAI21X1_766 ( .A(core__abc_21302_new_n3204_), .B(core__abc_21302_new_n3176_), .C(core__abc_21302_new_n3202_), .Y(core__abc_21302_new_n3223_));
OAI21X1 OAI21X1_767 ( .A(core__abc_21302_new_n3177_), .B(core__abc_21302_new_n3181_), .C(core__abc_21302_new_n1726_), .Y(core__abc_21302_new_n3225_));
OAI21X1 OAI21X1_768 ( .A(core__abc_21302_new_n1737_), .B(core__abc_21302_new_n1738_), .C(core__abc_21302_new_n3225_), .Y(core__abc_21302_new_n3226_));
OAI21X1 OAI21X1_769 ( .A(core__abc_21302_new_n1362_), .B(core__abc_21302_new_n1363_), .C(core__abc_21302_new_n3192_), .Y(core__abc_21302_new_n3228_));
OAI21X1 OAI21X1_77 ( .A(core_siphash_word_65_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf36), .Y(_abc_19873_new_n1610_));
OAI21X1 OAI21X1_770 ( .A(core__abc_21302_new_n1375_), .B(core__abc_21302_new_n1376_), .C(core__abc_21302_new_n3228_), .Y(core__abc_21302_new_n3229_));
OAI21X1 OAI21X1_771 ( .A(core__abc_21302_new_n3239_), .B(core__abc_21302_new_n3238_), .C(core__abc_21302_new_n3240_), .Y(core__abc_21302_new_n3241_));
OAI21X1 OAI21X1_772 ( .A(core__abc_21302_new_n3249_), .B(core__abc_21302_new_n3250_), .C(core__abc_21302_new_n3246_), .Y(core__abc_21302_new_n3251_));
OAI21X1 OAI21X1_773 ( .A(core__abc_21302_new_n3245_), .B(core__abc_21302_new_n3256_), .C(core__abc_21302_new_n3257_), .Y(core__abc_21302_new_n3258_));
OAI21X1 OAI21X1_774 ( .A(core__abc_21302_new_n2168__bF_buf4), .B(core__abc_21302_new_n3260_), .C(core__abc_21302_new_n2369__bF_buf2), .Y(core__abc_21302_new_n3261_));
OAI21X1 OAI21X1_775 ( .A(core_v3_reg_15_), .B(core__abc_21302_new_n2369__bF_buf1), .C(reset_n_bF_buf15), .Y(core__abc_21302_new_n3263_));
OAI21X1 OAI21X1_776 ( .A(core__abc_21302_new_n2363__bF_buf4), .B(core__abc_21302_new_n2368__bF_buf3), .C(core_v3_reg_16_), .Y(core__abc_21302_new_n3265_));
OAI21X1 OAI21X1_777 ( .A(core__abc_21302_new_n1704_), .B(core__abc_21302_new_n3131_), .C(core__abc_21302_new_n1716_), .Y(core__abc_21302_new_n3268_));
OAI21X1 OAI21X1_778 ( .A(core__abc_21302_new_n3280_), .B(core__abc_21302_new_n3240_), .C(core__abc_21302_new_n3281_), .Y(core__abc_21302_new_n3282_));
OAI21X1 OAI21X1_779 ( .A(core__abc_21302_new_n3279_), .B(core__abc_21302_new_n3273_), .C(core__abc_21302_new_n3282_), .Y(core__abc_21302_new_n3283_));
OAI21X1 OAI21X1_78 ( .A(core_siphash_word_66_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf35), .Y(_abc_19873_new_n1612_));
OAI21X1 OAI21X1_780 ( .A(core__abc_21302_new_n3286_), .B(core__abc_21302_new_n3183_), .C(core__abc_21302_new_n3290_), .Y(core__abc_21302_new_n3291_));
OAI21X1 OAI21X1_781 ( .A(core__abc_21302_new_n3295_), .B(core__abc_21302_new_n2467_), .C(core__abc_21302_new_n3294_), .Y(core__abc_21302_new_n3296_));
OAI21X1 OAI21X1_782 ( .A(core__abc_21302_new_n3297_), .B(core__abc_21302_new_n3298_), .C(core__abc_21302_new_n3301_), .Y(core__abc_21302_new_n3302_));
OAI21X1 OAI21X1_783 ( .A(core__abc_21302_new_n1878_), .B(core__abc_21302_new_n3250_), .C(core__abc_21302_new_n1891_), .Y(core__abc_21302_new_n3315_));
OAI21X1 OAI21X1_784 ( .A(core__abc_21302_new_n1888_), .B(core__abc_21302_new_n1890_), .C(core__abc_21302_new_n3312_), .Y(core__abc_21302_new_n3317_));
OAI21X1 OAI21X1_785 ( .A(core__abc_21302_new_n3266_), .B(core__abc_21302_new_n3325_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n3326_));
OAI21X1 OAI21X1_786 ( .A(core__abc_21302_new_n3288_), .B(core__abc_21302_new_n2933_), .C(core__abc_21302_new_n3292_), .Y(core__abc_21302_new_n3329_));
OAI21X1 OAI21X1_787 ( .A(core__abc_21302_new_n1748_), .B(core__abc_21302_new_n3331_), .C(core__abc_21302_new_n1749_), .Y(core__abc_21302_new_n3332_));
OAI21X1 OAI21X1_788 ( .A(core__abc_21302_new_n3335_), .B(core__abc_21302_new_n3331_), .C(core__abc_21302_new_n3334_), .Y(core__abc_21302_new_n3336_));
OAI21X1 OAI21X1_789 ( .A(core__abc_21302_new_n3333_), .B(core__abc_21302_new_n3336_), .C(core__abc_21302_new_n3343_), .Y(core__abc_21302_new_n3344_));
OAI21X1 OAI21X1_79 ( .A(core_siphash_word_67_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf34), .Y(_abc_19873_new_n1615_));
OAI21X1 OAI21X1_790 ( .A(core__abc_21302_new_n3313_), .B(core__abc_21302_new_n3253_), .C(core__abc_21302_new_n3352_), .Y(core__abc_21302_new_n3353_));
OAI21X1 OAI21X1_791 ( .A(core__abc_21302_new_n3355_), .B(core__abc_21302_new_n3354_), .C(core__abc_21302_new_n2703_), .Y(core__abc_21302_new_n3356_));
OAI21X1 OAI21X1_792 ( .A(core__abc_21302_new_n3351_), .B(core__abc_21302_new_n3360_), .C(core__abc_21302_new_n3361_), .Y(core__abc_21302_new_n3362_));
OAI21X1 OAI21X1_793 ( .A(core__abc_21302_new_n2168__bF_buf2), .B(core__abc_21302_new_n3363_), .C(core__abc_21302_new_n3362_), .Y(core__abc_21302_new_n3364_));
OAI21X1 OAI21X1_794 ( .A(core__abc_21302_new_n3328_), .B(core__abc_21302_new_n3364_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n3365_));
OAI21X1 OAI21X1_795 ( .A(core_v3_reg_17_), .B(core__abc_21302_new_n2369__bF_buf0), .C(reset_n_bF_buf14), .Y(core__abc_21302_new_n3366_));
OAI21X1 OAI21X1_796 ( .A(core__abc_21302_new_n3333_), .B(core__abc_21302_new_n3336_), .C(core__abc_21302_new_n3341_), .Y(core__abc_21302_new_n3373_));
OAI21X1 OAI21X1_797 ( .A(core__abc_21302_new_n3379_), .B(core__abc_21302_new_n3380_), .C(core__abc_21302_new_n3334_), .Y(core__abc_21302_new_n3381_));
OAI21X1 OAI21X1_798 ( .A(core__abc_21302_new_n1770_), .B(core__abc_21302_new_n1772_), .C(core__abc_21302_new_n3382_), .Y(core__abc_21302_new_n3384_));
OAI21X1 OAI21X1_799 ( .A(core__abc_21302_new_n3390_), .B(core__abc_21302_new_n3391_), .C(core__abc_21302_new_n3392_), .Y(core__abc_21302_new_n3393_));
OAI21X1 OAI21X1_8 ( .A(_abc_19873_new_n1002_), .B(_abc_19873_new_n918_), .C(_abc_19873_new_n1003_), .Y(_abc_19873_new_n1004_));
OAI21X1 OAI21X1_80 ( .A(core_siphash_word_68_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf33), .Y(_abc_19873_new_n1618_));
OAI21X1 OAI21X1_800 ( .A(core__abc_21302_new_n1904_), .B(core__abc_21302_new_n3354_), .C(core__abc_21302_new_n1919_), .Y(core__abc_21302_new_n3397_));
OAI21X1 OAI21X1_801 ( .A(core__abc_21302_new_n1904_), .B(core__abc_21302_new_n3354_), .C(core__abc_21302_new_n3399_), .Y(core__abc_21302_new_n3404_));
OAI21X1 OAI21X1_802 ( .A(core__abc_21302_new_n3396_), .B(core__abc_21302_new_n3407_), .C(core__abc_21302_new_n3408_), .Y(core__abc_21302_new_n3409_));
OAI21X1 OAI21X1_803 ( .A(core__abc_21302_new_n2168__bF_buf1), .B(core__abc_21302_new_n3410_), .C(core__abc_21302_new_n3409_), .Y(core__abc_21302_new_n3411_));
OAI21X1 OAI21X1_804 ( .A(core__abc_21302_new_n3368_), .B(core__abc_21302_new_n3411_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n3412_));
OAI21X1 OAI21X1_805 ( .A(core_v3_reg_18_), .B(core__abc_21302_new_n2369__bF_buf6), .C(reset_n_bF_buf13), .Y(core__abc_21302_new_n3413_));
OAI21X1 OAI21X1_806 ( .A(core__abc_21302_new_n3415_), .B(core__abc_21302_new_n3376_), .C(core__abc_21302_new_n3389_), .Y(core__abc_21302_new_n3416_));
OAI21X1 OAI21X1_807 ( .A(core__abc_21302_new_n1772_), .B(core__abc_21302_new_n3390_), .C(core__abc_21302_new_n3418_), .Y(core__abc_21302_new_n3419_));
OAI21X1 OAI21X1_808 ( .A(core__abc_21302_new_n1412_), .B(core__abc_21302_new_n3386_), .C(core__abc_21302_new_n1408_), .Y(core__abc_21302_new_n3420_));
OAI21X1 OAI21X1_809 ( .A(core__abc_21302_new_n3425_), .B(core__abc_21302_new_n3426_), .C(core__abc_21302_new_n3424_), .Y(core__abc_21302_new_n3427_));
OAI21X1 OAI21X1_81 ( .A(core_siphash_word_69_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf32), .Y(_abc_19873_new_n1621_));
OAI21X1 OAI21X1_810 ( .A(core__abc_21302_new_n1772_), .B(core__abc_21302_new_n3390_), .C(core__abc_21302_new_n1785_), .Y(core__abc_21302_new_n3431_));
OAI21X1 OAI21X1_811 ( .A(core__abc_21302_new_n1915_), .B(core__abc_21302_new_n3398_), .C(core__abc_21302_new_n3439_), .Y(core__abc_21302_new_n3440_));
OAI21X1 OAI21X1_812 ( .A(core__abc_21302_new_n1928_), .B(core__abc_21302_new_n1931_), .C(core__abc_21302_new_n3443_), .Y(core__abc_21302_new_n3444_));
OAI21X1 OAI21X1_813 ( .A(core__abc_21302_new_n3440_), .B(core__abc_21302_new_n3442_), .C(core__abc_21302_new_n1932_), .Y(core__abc_21302_new_n3445_));
OAI21X1 OAI21X1_814 ( .A(core__abc_21302_new_n3452_), .B(core__abc_21302_new_n2640__bF_buf11), .C(core__abc_21302_new_n2369__bF_buf4), .Y(core__abc_21302_new_n3453_));
OAI21X1 OAI21X1_815 ( .A(core__abc_21302_new_n2673__bF_buf8), .B(core__abc_21302_new_n3450_), .C(core__abc_21302_new_n3454_), .Y(core__abc_21302_new_n3455_));
OAI21X1 OAI21X1_816 ( .A(core_v3_reg_19_), .B(core__abc_21302_new_n2369__bF_buf3), .C(core__abc_21302_new_n3455_), .Y(core__abc_21302_new_n3456_));
OAI21X1 OAI21X1_817 ( .A(core__abc_21302_new_n3429_), .B(core__abc_21302_new_n3433_), .C(core__abc_21302_new_n3394_), .Y(core__abc_21302_new_n3460_));
OAI21X1 OAI21X1_818 ( .A(core__abc_21302_new_n1929_), .B(core__abc_21302_new_n1930_), .C(core__abc_21302_new_n3445_), .Y(core__abc_21302_new_n3489_));
OAI21X1 OAI21X1_819 ( .A(core__abc_21302_new_n3488_), .B(core__abc_21302_new_n3491_), .C(core__abc_21302_new_n3492_), .Y(core__abc_21302_new_n3493_));
OAI21X1 OAI21X1_82 ( .A(core_siphash_word_70_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf31), .Y(_abc_19873_new_n1624_));
OAI21X1 OAI21X1_820 ( .A(core_v3_reg_20_), .B(core__abc_21302_new_n2369__bF_buf2), .C(reset_n_bF_buf12), .Y(core__abc_21302_new_n3497_));
OAI21X1 OAI21X1_821 ( .A(core__abc_21302_new_n3473_), .B(core__abc_21302_new_n3331_), .C(core__abc_21302_new_n3500_), .Y(core__abc_21302_new_n3501_));
OAI21X1 OAI21X1_822 ( .A(core__abc_21302_new_n1809_), .B(core__abc_21302_new_n1810_), .C(core__abc_21302_new_n3502_), .Y(core__abc_21302_new_n3503_));
OAI21X1 OAI21X1_823 ( .A(core__abc_21302_new_n1793_), .B(core__abc_21302_new_n3475_), .C(core__abc_21302_new_n3504_), .Y(core__abc_21302_new_n3505_));
OAI21X1 OAI21X1_824 ( .A(core__abc_21302_new_n1436_), .B(core__abc_21302_new_n3478_), .C(core__abc_21302_new_n1432_), .Y(core__abc_21302_new_n3508_));
OAI21X1 OAI21X1_825 ( .A(core__abc_21302_new_n3485_), .B(core__abc_21302_new_n3468_), .C(core__abc_21302_new_n3483_), .Y(core__abc_21302_new_n3521_));
OAI21X1 OAI21X1_826 ( .A(core__abc_21302_new_n2510_), .B(core__abc_21302_new_n3523_), .C(core__abc_21302_new_n3524_), .Y(core__abc_21302_new_n3525_));
OAI21X1 OAI21X1_827 ( .A(core__abc_21302_new_n2168__bF_buf12), .B(core__abc_21302_new_n3526_), .C(core__abc_21302_new_n3525_), .Y(core__abc_21302_new_n3527_));
OAI21X1 OAI21X1_828 ( .A(core__abc_21302_new_n3499_), .B(core__abc_21302_new_n3527_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n3528_));
OAI21X1 OAI21X1_829 ( .A(core_v3_reg_21_), .B(core__abc_21302_new_n2369__bF_buf1), .C(reset_n_bF_buf11), .Y(core__abc_21302_new_n3529_));
OAI21X1 OAI21X1_83 ( .A(core_siphash_word_71_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf30), .Y(_abc_19873_new_n1627_));
OAI21X1 OAI21X1_830 ( .A(core__abc_21302_new_n3532_), .B(core__abc_21302_new_n3468_), .C(core__abc_21302_new_n3535_), .Y(core__abc_21302_new_n3536_));
OAI21X1 OAI21X1_831 ( .A(core__abc_21302_new_n1807_), .B(core__abc_21302_new_n1808_), .C(core__abc_21302_new_n3504_), .Y(core__abc_21302_new_n3541_));
OAI21X1 OAI21X1_832 ( .A(core__abc_21302_new_n3539_), .B(core__abc_21302_new_n3475_), .C(core__abc_21302_new_n3545_), .Y(core__abc_21302_new_n3546_));
OAI21X1 OAI21X1_833 ( .A(core__abc_21302_new_n3548_), .B(core__abc_21302_new_n3478_), .C(core__abc_21302_new_n2579_), .Y(core__abc_21302_new_n3549_));
OAI21X1 OAI21X1_834 ( .A(core__abc_21302_new_n3551_), .B(core__abc_21302_new_n3550_), .C(core_v3_reg_6_), .Y(core__abc_21302_new_n3552_));
OAI21X1 OAI21X1_835 ( .A(core__abc_21302_new_n3547_), .B(core__abc_21302_new_n3543_), .C(core__abc_21302_new_n3556_), .Y(core__abc_21302_new_n3557_));
OAI21X1 OAI21X1_836 ( .A(core__abc_21302_new_n1818_), .B(core__abc_21302_new_n1820_), .C(core__abc_21302_new_n3542_), .Y(core__abc_21302_new_n3559_));
OAI21X1 OAI21X1_837 ( .A(core__abc_21302_new_n2653_), .B(core__abc_21302_new_n3565_), .C(core__abc_21302_new_n3566_), .Y(core__abc_21302_new_n3567_));
OAI21X1 OAI21X1_838 ( .A(core__abc_21302_new_n2168__bF_buf11), .B(core__abc_21302_new_n3568_), .C(core__abc_21302_new_n3567_), .Y(core__abc_21302_new_n3569_));
OAI21X1 OAI21X1_839 ( .A(core__abc_21302_new_n3531_), .B(core__abc_21302_new_n3569_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n3570_));
OAI21X1 OAI21X1_84 ( .A(core_siphash_word_72_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf29), .Y(_abc_19873_new_n1629_));
OAI21X1 OAI21X1_840 ( .A(core_v3_reg_22_), .B(core__abc_21302_new_n2369__bF_buf7), .C(reset_n_bF_buf10), .Y(core__abc_21302_new_n3571_));
OAI21X1 OAI21X1_841 ( .A(core__abc_21302_new_n3537_), .B(core__abc_21302_new_n3542_), .C(core__abc_21302_new_n1819_), .Y(core__abc_21302_new_n3578_));
OAI21X1 OAI21X1_842 ( .A(core__abc_21302_new_n2580_), .B(core__abc_21302_new_n3550_), .C(core__abc_21302_new_n1468_), .Y(core__abc_21302_new_n3581_));
OAI21X1 OAI21X1_843 ( .A(core__abc_21302_new_n2580_), .B(core__abc_21302_new_n3550_), .C(core__abc_21302_new_n2576_), .Y(core__abc_21302_new_n3585_));
OAI21X1 OAI21X1_844 ( .A(core__abc_21302_new_n3573_), .B(core__abc_21302_new_n3595_), .C(core__abc_21302_new_n3596_), .Y(core__abc_21302_new_n3597_));
OAI21X1 OAI21X1_845 ( .A(core__abc_21302_new_n2168__bF_buf10), .B(core__abc_21302_new_n3599_), .C(core__abc_21302_new_n2369__bF_buf5), .Y(core__abc_21302_new_n3600_));
OAI21X1 OAI21X1_846 ( .A(core_v3_reg_23_), .B(core__abc_21302_new_n2369__bF_buf4), .C(reset_n_bF_buf9), .Y(core__abc_21302_new_n3602_));
OAI21X1 OAI21X1_847 ( .A(core__abc_21302_new_n3618_), .B(core__abc_21302_new_n3545_), .C(core__abc_21302_new_n3623_), .Y(core__abc_21302_new_n3624_));
OAI21X1 OAI21X1_848 ( .A(core__abc_21302_new_n3628_), .B(core__abc_21302_new_n3331_), .C(core__abc_21302_new_n3629_), .Y(core__abc_21302_new_n3630_));
OAI21X1 OAI21X1_849 ( .A(core__abc_21302_new_n3632_), .B(core__abc_21302_new_n3634_), .C(core__abc_21302_new_n1480_), .Y(core__abc_21302_new_n3635_));
OAI21X1 OAI21X1_85 ( .A(core_siphash_word_73_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf28), .Y(_abc_19873_new_n1631_));
OAI21X1 OAI21X1_850 ( .A(core__abc_21302_new_n1478_), .B(core__abc_21302_new_n1479_), .C(core__abc_21302_new_n3636_), .Y(core__abc_21302_new_n3637_));
OAI21X1 OAI21X1_851 ( .A(core__abc_21302_new_n3627_), .B(core__abc_21302_new_n3631_), .C(core__abc_21302_new_n3640_), .Y(core__abc_21302_new_n3641_));
OAI21X1 OAI21X1_852 ( .A(core__abc_21302_new_n2745_), .B(core__abc_21302_new_n3646_), .C(core__abc_21302_new_n2634__bF_buf2), .Y(core__abc_21302_new_n3648_));
OAI21X1 OAI21X1_853 ( .A(core_key_88_), .B(core__abc_21302_new_n2640__bF_buf7), .C(core__abc_21302_new_n2369__bF_buf3), .Y(core__abc_21302_new_n3650_));
OAI21X1 OAI21X1_854 ( .A(core__abc_21302_new_n3647_), .B(core__abc_21302_new_n3648_), .C(core__abc_21302_new_n3651_), .Y(core__abc_21302_new_n3652_));
OAI21X1 OAI21X1_855 ( .A(core_v3_reg_24_), .B(core__abc_21302_new_n2369__bF_buf2), .C(core__abc_21302_new_n3652_), .Y(core__abc_21302_new_n3653_));
OAI21X1 OAI21X1_856 ( .A(core__abc_21302_new_n1844_), .B(core__abc_21302_new_n3626_), .C(core__abc_21302_new_n3655_), .Y(core__abc_21302_new_n3656_));
OAI21X1 OAI21X1_857 ( .A(core__abc_21302_new_n1858_), .B(core__abc_21302_new_n1860_), .C(core__abc_21302_new_n3657_), .Y(core__abc_21302_new_n3658_));
OAI21X1 OAI21X1_858 ( .A(core__abc_21302_new_n1847_), .B(core__abc_21302_new_n3627_), .C(core__abc_21302_new_n1861_), .Y(core__abc_21302_new_n3659_));
OAI21X1 OAI21X1_859 ( .A(core__abc_21302_new_n1479_), .B(core__abc_21302_new_n3636_), .C(core__abc_21302_new_n3662_), .Y(core__abc_21302_new_n3663_));
OAI21X1 OAI21X1_86 ( .A(core_siphash_word_74_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf27), .Y(_abc_19873_new_n1633_));
OAI21X1 OAI21X1_860 ( .A(core__abc_21302_new_n3644_), .B(core__abc_21302_new_n3616_), .C(core__abc_21302_new_n3643_), .Y(core__abc_21302_new_n3677_));
OAI21X1 OAI21X1_861 ( .A(core__abc_21302_new_n2775_), .B(core__abc_21302_new_n3678_), .C(core__abc_21302_new_n3679_), .Y(core__abc_21302_new_n3680_));
OAI21X1 OAI21X1_862 ( .A(core__abc_21302_new_n3682_), .B(core__abc_21302_new_n2640__bF_buf6), .C(core__abc_21302_new_n2369__bF_buf1), .Y(core__abc_21302_new_n3683_));
OAI21X1 OAI21X1_863 ( .A(core_v3_reg_25_), .B(core__abc_21302_new_n2369__bF_buf0), .C(reset_n_bF_buf8), .Y(core__abc_21302_new_n3685_));
OAI21X1 OAI21X1_864 ( .A(core__abc_21302_new_n3660_), .B(core__abc_21302_new_n3672_), .C(core__abc_21302_new_n3643_), .Y(core__abc_21302_new_n3692_));
OAI21X1 OAI21X1_865 ( .A(core__abc_21302_new_n3655_), .B(core__abc_21302_new_n3694_), .C(core__abc_21302_new_n1859_), .Y(core__abc_21302_new_n3697_));
OAI21X1 OAI21X1_866 ( .A(core__abc_21302_new_n3696_), .B(core__abc_21302_new_n3626_), .C(core__abc_21302_new_n3698_), .Y(core__abc_21302_new_n3699_));
OAI21X1 OAI21X1_867 ( .A(core__abc_21302_new_n2554_), .B(core__abc_21302_new_n3636_), .C(core__abc_21302_new_n3703_), .Y(core__abc_21302_new_n3704_));
OAI21X1 OAI21X1_868 ( .A(core__abc_21302_new_n3705_), .B(core__abc_21302_new_n3706_), .C(core__abc_21302_new_n1317_), .Y(core__abc_21302_new_n3707_));
OAI21X1 OAI21X1_869 ( .A(core__abc_21302_new_n3702_), .B(core__abc_21302_new_n3701_), .C(core__abc_21302_new_n3710_), .Y(core__abc_21302_new_n3711_));
OAI21X1 OAI21X1_87 ( .A(core_siphash_word_75_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf26), .Y(_abc_19873_new_n1636_));
OAI21X1 OAI21X1_870 ( .A(core__abc_21302_new_n1870_), .B(core__abc_21302_new_n1873_), .C(core__abc_21302_new_n3712_), .Y(core__abc_21302_new_n3713_));
OAI21X1 OAI21X1_871 ( .A(core__abc_21302_new_n2807_), .B(core__abc_21302_new_n3717_), .C(core__abc_21302_new_n2634__bF_buf1), .Y(core__abc_21302_new_n3719_));
OAI21X1 OAI21X1_872 ( .A(core__abc_21302_new_n3688_), .B(core__abc_21302_new_n3721_), .C(core__abc_21302_new_n2362__bF_buf0), .Y(core__abc_21302_new_n3722_));
OAI21X1 OAI21X1_873 ( .A(core_v3_reg_26_), .B(core__abc_21302_new_n2369__bF_buf7), .C(reset_n_bF_buf7), .Y(core__abc_21302_new_n3723_));
OAI21X1 OAI21X1_874 ( .A(core__abc_21302_new_n1870_), .B(core__abc_21302_new_n3712_), .C(core__abc_21302_new_n3730_), .Y(core__abc_21302_new_n3732_));
OAI21X1 OAI21X1_875 ( .A(core__abc_21302_new_n1884_), .B(core__abc_21302_new_n1886_), .C(core__abc_21302_new_n3732_), .Y(core__abc_21302_new_n3733_));
OAI21X1 OAI21X1_876 ( .A(core__abc_21302_new_n3736_), .B(core__abc_21302_new_n3706_), .C(core__abc_21302_new_n1514_), .Y(core__abc_21302_new_n3737_));
OAI21X1 OAI21X1_877 ( .A(core__abc_21302_new_n3736_), .B(core__abc_21302_new_n3706_), .C(core__abc_21302_new_n2552_), .Y(core__abc_21302_new_n3740_));
OAI21X1 OAI21X1_878 ( .A(core__abc_21302_new_n3745_), .B(core__abc_21302_new_n3744_), .C(core__abc_21302_new_n3746_), .Y(core__abc_21302_new_n3747_));
OAI21X1 OAI21X1_879 ( .A(core__abc_21302_new_n2854_), .B(core__abc_21302_new_n3751_), .C(core__abc_21302_new_n3752_), .Y(core__abc_21302_new_n3753_));
OAI21X1 OAI21X1_88 ( .A(core_siphash_word_76_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf25), .Y(_abc_19873_new_n1639_));
OAI21X1 OAI21X1_880 ( .A(core_key_91_), .B(core__abc_21302_new_n2640__bF_buf4), .C(core__abc_21302_new_n2369__bF_buf5), .Y(core__abc_21302_new_n3755_));
OAI21X1 OAI21X1_881 ( .A(core_v3_reg_27_), .B(core__abc_21302_new_n2369__bF_buf4), .C(reset_n_bF_buf6), .Y(core__abc_21302_new_n3757_));
OAI21X1 OAI21X1_882 ( .A(core__abc_21302_new_n2363__bF_buf3), .B(core__abc_21302_new_n2368__bF_buf2), .C(core_v3_reg_28_), .Y(core__abc_21302_new_n3759_));
OAI21X1 OAI21X1_883 ( .A(core__abc_21302_new_n3674_), .B(core__abc_21302_new_n3671_), .C(core__abc_21302_new_n3692_), .Y(core__abc_21302_new_n3760_));
OAI21X1 OAI21X1_884 ( .A(core__abc_21302_new_n3761_), .B(core__abc_21302_new_n3760_), .C(core__abc_21302_new_n3763_), .Y(core__abc_21302_new_n3764_));
OAI21X1 OAI21X1_885 ( .A(core__abc_21302_new_n3766_), .B(core__abc_21302_new_n3616_), .C(core__abc_21302_new_n3765_), .Y(core__abc_21302_new_n3767_));
OAI21X1 OAI21X1_886 ( .A(core__abc_21302_new_n1884_), .B(core__abc_21302_new_n3730_), .C(core__abc_21302_new_n1885_), .Y(core__abc_21302_new_n3771_));
OAI21X1 OAI21X1_887 ( .A(core__abc_21302_new_n3770_), .B(core__abc_21302_new_n3626_), .C(core__abc_21302_new_n3772_), .Y(core__abc_21302_new_n3773_));
OAI21X1 OAI21X1_888 ( .A(core__abc_21302_new_n3775_), .B(core__abc_21302_new_n3636_), .C(core__abc_21302_new_n2597_), .Y(core__abc_21302_new_n3776_));
OAI21X1 OAI21X1_889 ( .A(core__abc_21302_new_n3781_), .B(core__abc_21302_new_n3780_), .C(core__abc_21302_new_n2886_), .Y(core__abc_21302_new_n3784_));
OAI21X1 OAI21X1_89 ( .A(core_siphash_word_77_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf24), .Y(_abc_19873_new_n1641_));
OAI21X1 OAI21X1_890 ( .A(core__abc_21302_new_n3787_), .B(core__abc_21302_new_n3785_), .C(core__abc_21302_new_n2362__bF_buf11), .Y(core__abc_21302_new_n3788_));
OAI21X1 OAI21X1_891 ( .A(core__abc_21302_new_n2396_), .B(core__abc_21302_new_n3794_), .C(core__abc_21302_new_n2486_), .Y(core__abc_21302_new_n3795_));
OAI21X1 OAI21X1_892 ( .A(core__abc_21302_new_n2466_), .B(core__abc_21302_new_n3796_), .C(core__abc_21302_new_n3330_), .Y(core__abc_21302_new_n3797_));
OAI21X1 OAI21X1_893 ( .A(core__abc_21302_new_n3625_), .B(core__abc_21302_new_n3798_), .C(core__abc_21302_new_n3799_), .Y(core__abc_21302_new_n3800_));
OAI21X1 OAI21X1_894 ( .A(core__abc_21302_new_n1523_), .B(core__abc_21302_new_n1524_), .C(core__abc_21302_new_n3808_), .Y(core__abc_21302_new_n3810_));
OAI21X1 OAI21X1_895 ( .A(core__abc_21302_new_n3814_), .B(core__abc_21302_new_n3813_), .C(core__abc_21302_new_n1351_), .Y(core__abc_21302_new_n3815_));
OAI21X1 OAI21X1_896 ( .A(core__abc_21302_new_n2940_), .B(core__abc_21302_new_n3821_), .C(core__abc_21302_new_n2634__bF_buf0), .Y(core__abc_21302_new_n3823_));
OAI21X1 OAI21X1_897 ( .A(core_key_93_), .B(core__abc_21302_new_n2640__bF_buf2), .C(core__abc_21302_new_n2369__bF_buf3), .Y(core__abc_21302_new_n3825_));
OAI21X1 OAI21X1_898 ( .A(core__abc_21302_new_n3822_), .B(core__abc_21302_new_n3823_), .C(core__abc_21302_new_n3826_), .Y(core__abc_21302_new_n3827_));
OAI21X1 OAI21X1_899 ( .A(core_v3_reg_29_), .B(core__abc_21302_new_n2369__bF_buf2), .C(core__abc_21302_new_n3827_), .Y(core__abc_21302_new_n3828_));
OAI21X1 OAI21X1_9 ( .A(_abc_19873_new_n1010_), .B(_abc_19873_new_n960__bF_buf2), .C(_abc_19873_new_n1011_), .Y(_abc_19873_new_n1012_));
OAI21X1 OAI21X1_90 ( .A(core_siphash_word_78_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf23), .Y(_abc_19873_new_n1644_));
OAI21X1 OAI21X1_900 ( .A(core__abc_21302_new_n1911_), .B(core__abc_21302_new_n1912_), .C(core__abc_21302_new_n3791_), .Y(core__abc_21302_new_n3832_));
OAI21X1 OAI21X1_901 ( .A(core__abc_21302_new_n1536_), .B(core__abc_21302_new_n1537_), .C(core__abc_21302_new_n1522_), .Y(core__abc_21302_new_n3836_));
OAI21X1 OAI21X1_902 ( .A(core__abc_21302_new_n3838_), .B(core__abc_21302_new_n3839_), .C(core_v3_reg_14_), .Y(core__abc_21302_new_n3840_));
OAI21X1 OAI21X1_903 ( .A(core__abc_21302_new_n3632_), .B(core__abc_21302_new_n3634_), .C(core__abc_21302_new_n2555_), .Y(core__abc_21302_new_n3843_));
OAI21X1 OAI21X1_904 ( .A(core__abc_21302_new_n2598_), .B(core__abc_21302_new_n3844_), .C(core__abc_21302_new_n3841_), .Y(core__abc_21302_new_n3845_));
OAI21X1 OAI21X1_905 ( .A(core__abc_21302_new_n3834_), .B(core__abc_21302_new_n3835_), .C(core__abc_21302_new_n3848_), .Y(core__abc_21302_new_n3849_));
OAI21X1 OAI21X1_906 ( .A(core__abc_21302_new_n3832_), .B(core__abc_21302_new_n3804_), .C(core__abc_21302_new_n1927_), .Y(core__abc_21302_new_n3850_));
OAI21X1 OAI21X1_907 ( .A(core__abc_21302_new_n1924_), .B(core__abc_21302_new_n1926_), .C(core__abc_21302_new_n3833_), .Y(core__abc_21302_new_n3851_));
OAI21X1 OAI21X1_908 ( .A(core__abc_21302_new_n3855_), .B(core__abc_21302_new_n3817_), .C(core__abc_21302_new_n3818_), .Y(core__abc_21302_new_n3856_));
OAI21X1 OAI21X1_909 ( .A(core__abc_21302_new_n3858_), .B(core__abc_21302_new_n3801_), .C(core__abc_21302_new_n3805_), .Y(core__abc_21302_new_n3859_));
OAI21X1 OAI21X1_91 ( .A(core_siphash_word_79_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf22), .Y(_abc_19873_new_n1646_));
OAI21X1 OAI21X1_910 ( .A(core__abc_21302_new_n2971_), .B(core__abc_21302_new_n3869_), .C(core__abc_21302_new_n2634__bF_buf8), .Y(core__abc_21302_new_n3871_));
OAI21X1 OAI21X1_911 ( .A(core__abc_21302_new_n3830_), .B(core__abc_21302_new_n3873_), .C(core__abc_21302_new_n2362__bF_buf10), .Y(core__abc_21302_new_n3874_));
OAI21X1 OAI21X1_912 ( .A(core_v3_reg_30_), .B(core__abc_21302_new_n2369__bF_buf1), .C(reset_n_bF_buf5), .Y(core__abc_21302_new_n3875_));
OAI21X1 OAI21X1_913 ( .A(core__abc_21302_new_n3831_), .B(core__abc_21302_new_n3833_), .C(core__abc_21302_new_n1925_), .Y(core__abc_21302_new_n3881_));
OAI21X1 OAI21X1_914 ( .A(core__abc_21302_new_n2589_), .B(core__abc_21302_new_n3838_), .C(core__abc_21302_new_n1559_), .Y(core__abc_21302_new_n3885_));
OAI21X1 OAI21X1_915 ( .A(core__abc_21302_new_n2589_), .B(core__abc_21302_new_n3838_), .C(core__abc_21302_new_n3883_), .Y(core__abc_21302_new_n3888_));
OAI21X1 OAI21X1_916 ( .A(core__abc_21302_new_n3877_), .B(core__abc_21302_new_n3865_), .C(core__abc_21302_new_n3897_), .Y(core__abc_21302_new_n3898_));
OAI21X1 OAI21X1_917 ( .A(core__abc_21302_new_n3022_), .B(core__abc_21302_new_n3899_), .C(core__abc_21302_new_n3900_), .Y(core__abc_21302_new_n3901_));
OAI21X1 OAI21X1_918 ( .A(core__abc_21302_new_n2168__bF_buf6), .B(core__abc_21302_new_n3903_), .C(core__abc_21302_new_n2369__bF_buf7), .Y(core__abc_21302_new_n3904_));
OAI21X1 OAI21X1_919 ( .A(core_v3_reg_31_), .B(core__abc_21302_new_n2369__bF_buf6), .C(reset_n_bF_buf4), .Y(core__abc_21302_new_n3906_));
OAI21X1 OAI21X1_92 ( .A(core_siphash_word_80_), .B(_abc_19873_new_n1524__bF_buf15), .C(reset_n_bF_buf21), .Y(_abc_19873_new_n1649_));
OAI21X1 OAI21X1_920 ( .A(core__abc_21302_new_n2363__bF_buf2), .B(core__abc_21302_new_n2368__bF_buf1), .C(core_v3_reg_32_), .Y(core__abc_21302_new_n3908_));
OAI21X1 OAI21X1_921 ( .A(core__abc_21302_new_n3857_), .B(core__abc_21302_new_n3915_), .C(core__abc_21302_new_n3917_), .Y(core__abc_21302_new_n3918_));
OAI21X1 OAI21X1_922 ( .A(core__abc_21302_new_n1569_), .B(core__abc_21302_new_n1570_), .C(core__abc_21302_new_n3921_), .Y(core__abc_21302_new_n3922_));
OAI21X1 OAI21X1_923 ( .A(core__abc_21302_new_n2602_), .B(core__abc_21302_new_n2568_), .C(core__abc_21302_new_n3923_), .Y(core__abc_21302_new_n3924_));
OAI21X1 OAI21X1_924 ( .A(core__abc_21302_new_n3913_), .B(core__abc_21302_new_n3920_), .C(core__abc_21302_new_n3929_), .Y(core__abc_21302_new_n3930_));
OAI21X1 OAI21X1_925 ( .A(core__abc_21302_new_n3927_), .B(core__abc_21302_new_n3928_), .C(core__abc_21302_new_n3931_), .Y(core__abc_21302_new_n3932_));
OAI21X1 OAI21X1_926 ( .A(core__abc_21302_new_n3939_), .B(core__abc_21302_new_n3936_), .C(core__abc_21302_new_n2362__bF_buf9), .Y(core__abc_21302_new_n3940_));
OAI21X1 OAI21X1_927 ( .A(core__abc_21302_new_n2363__bF_buf1), .B(core__abc_21302_new_n2368__bF_buf0), .C(core_v3_reg_33_), .Y(core__abc_21302_new_n3942_));
OAI21X1 OAI21X1_928 ( .A(core__abc_21302_new_n3928_), .B(core__abc_21302_new_n3931_), .C(core__abc_21302_new_n3943_), .Y(core__abc_21302_new_n3944_));
OAI21X1 OAI21X1_929 ( .A(core__abc_21302_new_n1220_), .B(core__abc_21302_new_n1222_), .C(core__abc_21302_new_n1209_), .Y(core__abc_21302_new_n3946_));
OAI21X1 OAI21X1_93 ( .A(core_siphash_word_81_), .B(_abc_19873_new_n1524__bF_buf13), .C(reset_n_bF_buf20), .Y(_abc_19873_new_n1652_));
OAI21X1 OAI21X1_930 ( .A(core__abc_21302_new_n1570_), .B(core__abc_21302_new_n3921_), .C(core__abc_21302_new_n1568_), .Y(core__abc_21302_new_n3952_));
OAI21X1 OAI21X1_931 ( .A(core__abc_21302_new_n3955_), .B(core__abc_21302_new_n3957_), .C(core__abc_21302_new_n3948_), .Y(core__abc_21302_new_n3958_));
OAI21X1 OAI21X1_932 ( .A(core__abc_21302_new_n3966_), .B(core__abc_21302_new_n3964_), .C(core__abc_21302_new_n2362__bF_buf8), .Y(core__abc_21302_new_n3967_));
OAI21X1 OAI21X1_933 ( .A(core__abc_21302_new_n2363__bF_buf0), .B(core__abc_21302_new_n2368__bF_buf4), .C(core_v3_reg_34_), .Y(core__abc_21302_new_n3969_));
OAI21X1 OAI21X1_934 ( .A(core__abc_21302_new_n3947_), .B(core__abc_21302_new_n3959_), .C(core__abc_21302_new_n3943_), .Y(core__abc_21302_new_n3972_));
OAI21X1 OAI21X1_935 ( .A(core__abc_21302_new_n3948_), .B(core__abc_21302_new_n3971_), .C(core__abc_21302_new_n3972_), .Y(core__abc_21302_new_n3973_));
OAI21X1 OAI21X1_936 ( .A(core__abc_21302_new_n3974_), .B(core__abc_21302_new_n3931_), .C(core__abc_21302_new_n3973_), .Y(core__abc_21302_new_n3975_));
OAI21X1 OAI21X1_937 ( .A(core__abc_21302_new_n3981_), .B(core__abc_21302_new_n3921_), .C(core__abc_21302_new_n3982_), .Y(core__abc_21302_new_n3983_));
OAI21X1 OAI21X1_938 ( .A(core__abc_21302_new_n3986_), .B(core__abc_21302_new_n3985_), .C(core__abc_21302_new_n1410_), .Y(core__abc_21302_new_n3987_));
OAI21X1 OAI21X1_939 ( .A(core__abc_21302_new_n3986_), .B(core__abc_21302_new_n3985_), .C(core_v3_reg_18_), .Y(core__abc_21302_new_n3991_));
OAI21X1 OAI21X1_94 ( .A(core_siphash_word_82_), .B(_abc_19873_new_n1524__bF_buf11), .C(reset_n_bF_buf19), .Y(_abc_19873_new_n1655_));
OAI21X1 OAI21X1_940 ( .A(core__abc_21302_new_n3970_), .B(core__abc_21302_new_n3998_), .C(core__abc_21302_new_n2362__bF_buf7), .Y(core__abc_21302_new_n3999_));
OAI21X1 OAI21X1_941 ( .A(core__abc_21302_new_n3978_), .B(core__abc_21302_new_n4001_), .C(core__abc_21302_new_n4002_), .Y(core__abc_21302_new_n4003_));
OAI21X1 OAI21X1_942 ( .A(core__abc_21302_new_n2471_), .B(core__abc_21302_new_n2469_), .C(core__abc_21302_new_n3976_), .Y(core__abc_21302_new_n4004_));
OAI21X1 OAI21X1_943 ( .A(core__abc_21302_new_n1593_), .B(core__abc_21302_new_n1594_), .C(core__abc_21302_new_n3984_), .Y(core__abc_21302_new_n4008_));
OAI21X1 OAI21X1_944 ( .A(core__abc_21302_new_n3201_), .B(core__abc_21302_new_n4021_), .C(core__abc_21302_new_n4022_), .Y(core__abc_21302_new_n4023_));
OAI21X1 OAI21X1_945 ( .A(core__abc_21302_new_n4025_), .B(core__abc_21302_new_n2640__bF_buf10), .C(core__abc_21302_new_n2369__bF_buf5), .Y(core__abc_21302_new_n4026_));
OAI21X1 OAI21X1_946 ( .A(core_v3_reg_35_), .B(core__abc_21302_new_n2369__bF_buf4), .C(reset_n_bF_buf3), .Y(core__abc_21302_new_n4028_));
OAI21X1 OAI21X1_947 ( .A(core__abc_21302_new_n2363__bF_buf5), .B(core__abc_21302_new_n2368__bF_buf3), .C(core_v3_reg_36_), .Y(core__abc_21302_new_n4030_));
OAI21X1 OAI21X1_948 ( .A(core__abc_21302_new_n3973_), .B(core__abc_21302_new_n4032_), .C(core__abc_21302_new_n4035_), .Y(core__abc_21302_new_n4036_));
OAI21X1 OAI21X1_949 ( .A(core__abc_21302_new_n2608_), .B(core__abc_21302_new_n3921_), .C(core__abc_21302_new_n2613_), .Y(core__abc_21302_new_n4045_));
OAI21X1 OAI21X1_95 ( .A(core_siphash_word_83_), .B(_abc_19873_new_n1524__bF_buf9), .C(reset_n_bF_buf18), .Y(_abc_19873_new_n1658_));
OAI21X1 OAI21X1_950 ( .A(core__abc_21302_new_n4031_), .B(core__abc_21302_new_n4059_), .C(core__abc_21302_new_n2362__bF_buf6), .Y(core__abc_21302_new_n4060_));
OAI21X1 OAI21X1_951 ( .A(core__abc_21302_new_n2363__bF_buf4), .B(core__abc_21302_new_n2368__bF_buf2), .C(core_v3_reg_37_), .Y(core__abc_21302_new_n4062_));
OAI21X1 OAI21X1_952 ( .A(core__abc_21302_new_n1253_), .B(core__abc_21302_new_n2475_), .C(core__abc_21302_new_n1252_), .Y(core__abc_21302_new_n4063_));
OAI21X1 OAI21X1_953 ( .A(core__abc_21302_new_n1631_), .B(core__abc_21302_new_n1632_), .C(core__abc_21302_new_n4069_), .Y(core__abc_21302_new_n4070_));
OAI21X1 OAI21X1_954 ( .A(core__abc_21302_new_n1631_), .B(core__abc_21302_new_n1632_), .C(core__abc_21302_new_n4067_), .Y(core__abc_21302_new_n4072_));
OAI21X1 OAI21X1_955 ( .A(core__abc_21302_new_n4054_), .B(core__abc_21302_new_n4040_), .C(core__abc_21302_new_n4051_), .Y(core__abc_21302_new_n4079_));
OAI21X1 OAI21X1_956 ( .A(core__abc_21302_new_n4087_), .B(core__abc_21302_new_n4085_), .C(core__abc_21302_new_n2362__bF_buf5), .Y(core__abc_21302_new_n4088_));
OAI21X1 OAI21X1_957 ( .A(core__abc_21302_new_n2363__bF_buf3), .B(core__abc_21302_new_n2368__bF_buf1), .C(core_v3_reg_38_), .Y(core__abc_21302_new_n4090_));
OAI21X1 OAI21X1_958 ( .A(core__abc_21302_new_n4036_), .B(core__abc_21302_new_n4039_), .C(core__abc_21302_new_n4091_), .Y(core__abc_21302_new_n4092_));
OAI21X1 OAI21X1_959 ( .A(core__abc_21302_new_n4051_), .B(core__abc_21302_new_n4076_), .C(core__abc_21302_new_n4094_), .Y(core__abc_21302_new_n4095_));
OAI21X1 OAI21X1_96 ( .A(core_siphash_word_84_), .B(_abc_19873_new_n1524__bF_buf7), .C(reset_n_bF_buf17), .Y(_abc_19873_new_n1661_));
OAI21X1 OAI21X1_960 ( .A(core__abc_21302_new_n2379_), .B(core__abc_21302_new_n2380_), .C(core__abc_21302_new_n4096_), .Y(core__abc_21302_new_n4098_));
OAI21X1 OAI21X1_961 ( .A(core__abc_21302_new_n1639_), .B(core__abc_21302_new_n1641_), .C(core__abc_21302_new_n4100_), .Y(core__abc_21302_new_n4101_));
OAI21X1 OAI21X1_962 ( .A(core__abc_21302_new_n4095_), .B(core__abc_21302_new_n4093_), .C(core__abc_21302_new_n4113_), .Y(core__abc_21302_new_n4114_));
OAI21X1 OAI21X1_963 ( .A(core__abc_21302_new_n4122_), .B(core__abc_21302_new_n4120_), .C(core__abc_21302_new_n2362__bF_buf4), .Y(core__abc_21302_new_n4123_));
OAI21X1 OAI21X1_964 ( .A(core__abc_21302_new_n2379_), .B(core__abc_21302_new_n4096_), .C(core__abc_21302_new_n1274_), .Y(core__abc_21302_new_n4125_));
OAI21X1 OAI21X1_965 ( .A(core__abc_21302_new_n1642_), .B(core__abc_21302_new_n4100_), .C(core__abc_21302_new_n1640_), .Y(core__abc_21302_new_n4127_));
OAI21X1 OAI21X1_966 ( .A(core__abc_21302_new_n1651_), .B(core__abc_21302_new_n1652_), .C(core__abc_21302_new_n4127_), .Y(core__abc_21302_new_n4129_));
OAI21X1 OAI21X1_967 ( .A(core__abc_21302_new_n4136_), .B(core__abc_21302_new_n4137_), .C(core__abc_21302_new_n4135_), .Y(core__abc_21302_new_n4138_));
OAI21X1 OAI21X1_968 ( .A(core__abc_21302_new_n4141_), .B(core__abc_21302_new_n4144_), .C(core__abc_21302_new_n3388_), .Y(core__abc_21302_new_n4145_));
OAI21X1 OAI21X1_969 ( .A(core__abc_21302_new_n2168__bF_buf12), .B(core__abc_21302_new_n4148_), .C(core__abc_21302_new_n4147_), .Y(core__abc_21302_new_n4149_));
OAI21X1 OAI21X1_97 ( .A(core_siphash_word_85_), .B(_abc_19873_new_n1524__bF_buf5), .C(reset_n_bF_buf16), .Y(_abc_19873_new_n1663_));
OAI21X1 OAI21X1_970 ( .A(core_v3_reg_39_), .B(core__abc_21302_new_n2369__bF_buf3), .C(reset_n_bF_buf2), .Y(core__abc_21302_new_n4151_));
OAI21X1 OAI21X1_971 ( .A(core__abc_21302_new_n2363__bF_buf2), .B(core__abc_21302_new_n2368__bF_buf0), .C(core_v3_reg_40_), .Y(core__abc_21302_new_n4153_));
OAI21X1 OAI21X1_972 ( .A(core__abc_21302_new_n4135_), .B(core__abc_21302_new_n4157_), .C(core__abc_21302_new_n4111_), .Y(core__abc_21302_new_n4159_));
OAI21X1 OAI21X1_973 ( .A(core__abc_21302_new_n4161_), .B(core__abc_21302_new_n4172_), .C(core__abc_21302_new_n4179_), .Y(core__abc_21302_new_n4180_));
OAI21X1 OAI21X1_974 ( .A(core__abc_21302_new_n4154_), .B(core__abc_21302_new_n4187_), .C(core__abc_21302_new_n2362__bF_buf3), .Y(core__abc_21302_new_n4188_));
OAI21X1 OAI21X1_975 ( .A(core__abc_21302_new_n2363__bF_buf1), .B(core__abc_21302_new_n2368__bF_buf4), .C(core_v3_reg_41_), .Y(core__abc_21302_new_n4190_));
OAI21X1 OAI21X1_976 ( .A(core__abc_21302_new_n4173_), .B(core__abc_21302_new_n4176_), .C(core__abc_21302_new_n4180_), .Y(core__abc_21302_new_n4191_));
OAI21X1 OAI21X1_977 ( .A(core__abc_21302_new_n2396_), .B(core__abc_21302_new_n3794_), .C(core__abc_21302_new_n1293_), .Y(core__abc_21302_new_n4192_));
OAI21X1 OAI21X1_978 ( .A(core__abc_21302_new_n2405_), .B(core__abc_21302_new_n2406_), .C(core__abc_21302_new_n4192_), .Y(core__abc_21302_new_n4193_));
OAI21X1 OAI21X1_979 ( .A(core__abc_21302_new_n4205_), .B(core__abc_21302_new_n4204_), .C(core__abc_21302_new_n4194_), .Y(core__abc_21302_new_n4206_));
OAI21X1 OAI21X1_98 ( .A(core_siphash_word_86_), .B(_abc_19873_new_n1524__bF_buf3), .C(reset_n_bF_buf15), .Y(_abc_19873_new_n1666_));
OAI21X1 OAI21X1_980 ( .A(core__abc_21302_new_n4214_), .B(core__abc_21302_new_n4211_), .C(core__abc_21302_new_n2362__bF_buf2), .Y(core__abc_21302_new_n4215_));
OAI21X1 OAI21X1_981 ( .A(core__abc_21302_new_n2363__bF_buf0), .B(core__abc_21302_new_n2368__bF_buf3), .C(core_v3_reg_42_), .Y(core__abc_21302_new_n4217_));
OAI21X1 OAI21X1_982 ( .A(core__abc_21302_new_n2401_), .B(core__abc_21302_new_n2397_), .C(core__abc_21302_new_n2409_), .Y(core__abc_21302_new_n4218_));
OAI21X1 OAI21X1_983 ( .A(core__abc_21302_new_n2626_), .B(core__abc_21302_new_n4223_), .C(core__abc_21302_new_n1500_), .Y(core__abc_21302_new_n4224_));
OAI21X1 OAI21X1_984 ( .A(core__abc_21302_new_n1684_), .B(core__abc_21302_new_n1685_), .C(core__abc_21302_new_n4222_), .Y(core__abc_21302_new_n4225_));
OAI21X1 OAI21X1_985 ( .A(core__abc_21302_new_n2626_), .B(core__abc_21302_new_n4223_), .C(core_v3_reg_26_), .Y(core__abc_21302_new_n4228_));
OAI21X1 OAI21X1_986 ( .A(core__abc_21302_new_n4173_), .B(core__abc_21302_new_n4176_), .C(core__abc_21302_new_n4203_), .Y(core__abc_21302_new_n4233_));
OAI21X1 OAI21X1_987 ( .A(core__abc_21302_new_n4195_), .B(core__abc_21302_new_n4232_), .C(core__abc_21302_new_n4233_), .Y(core__abc_21302_new_n4234_));
OAI21X1 OAI21X1_988 ( .A(core__abc_21302_new_n4235_), .B(core__abc_21302_new_n4181_), .C(core__abc_21302_new_n4234_), .Y(core__abc_21302_new_n4236_));
OAI21X1 OAI21X1_989 ( .A(core__abc_21302_new_n4239_), .B(core__abc_21302_new_n4238_), .C(core__abc_21302_new_n3516_), .Y(core__abc_21302_new_n4240_));
OAI21X1 OAI21X1_99 ( .A(core_siphash_word_87_), .B(_abc_19873_new_n1524__bF_buf1), .C(reset_n_bF_buf14), .Y(_abc_19873_new_n1668_));
OAI21X1 OAI21X1_990 ( .A(core__abc_21302_new_n4245_), .B(core__abc_21302_new_n4243_), .C(core__abc_21302_new_n2362__bF_buf1), .Y(core__abc_21302_new_n4246_));
OAI21X1 OAI21X1_991 ( .A(core__abc_21302_new_n4248_), .B(core__abc_21302_new_n4249_), .C(core__abc_21302_new_n4250_), .Y(core__abc_21302_new_n4251_));
OAI21X1 OAI21X1_992 ( .A(core__abc_21302_new_n2631_), .B(core__abc_21302_new_n2628_), .C(core__abc_21302_new_n4252_), .Y(core__abc_21302_new_n4253_));
OAI21X1 OAI21X1_993 ( .A(core__abc_21302_new_n4262_), .B(core__abc_21302_new_n4238_), .C(core__abc_21302_new_n4259_), .Y(core__abc_21302_new_n4263_));
OAI21X1 OAI21X1_994 ( .A(core__abc_21302_new_n3560_), .B(core__abc_21302_new_n4264_), .C(core__abc_21302_new_n4265_), .Y(core__abc_21302_new_n4266_));
OAI21X1 OAI21X1_995 ( .A(core__abc_21302_new_n4268_), .B(core__abc_21302_new_n2640__bF_buf5), .C(core__abc_21302_new_n2369__bF_buf2), .Y(core__abc_21302_new_n4269_));
OAI21X1 OAI21X1_996 ( .A(core_v3_reg_43_), .B(core__abc_21302_new_n2369__bF_buf1), .C(reset_n_bF_buf1), .Y(core__abc_21302_new_n4271_));
OAI21X1 OAI21X1_997 ( .A(core__abc_21302_new_n2363__bF_buf5), .B(core__abc_21302_new_n2368__bF_buf2), .C(core_v3_reg_44_), .Y(core__abc_21302_new_n4273_));
OAI21X1 OAI21X1_998 ( .A(core__abc_21302_new_n4234_), .B(core__abc_21302_new_n4274_), .C(core__abc_21302_new_n4276_), .Y(core__abc_21302_new_n4277_));
OAI21X1 OAI21X1_999 ( .A(core__abc_21302_new_n3913_), .B(core__abc_21302_new_n3920_), .C(core__abc_21302_new_n4279_), .Y(core__abc_21302_new_n4280_));
OAI22X1 OAI22X1_1 ( .A(_abc_19873_new_n884_), .B(_abc_19873_new_n894__bF_buf4), .C(_abc_19873_new_n885_), .D(_abc_19873_new_n896__bF_buf4), .Y(_abc_19873_new_n897_));
OAI22X1 OAI22X1_10 ( .A(_abc_19873_new_n979_), .B(_abc_19873_new_n914__bF_buf1), .C(_abc_19873_new_n978_), .D(_abc_19873_new_n969__bF_buf2), .Y(_abc_19873_new_n980_));
OAI22X1 OAI22X1_100 ( .A(core__abc_21302_new_n2168__bF_buf4), .B(core__abc_21302_new_n3965_), .C(core_key_97_), .D(core__abc_21302_new_n2640__bF_buf11), .Y(core__abc_21302_new_n3966_));
OAI22X1 OAI22X1_101 ( .A(core__abc_21302_new_n2168__bF_buf3), .B(core__abc_21302_new_n3997_), .C(core__abc_21302_new_n2673__bF_buf9), .D(core__abc_21302_new_n3996_), .Y(core__abc_21302_new_n3998_));
OAI22X1 OAI22X1_102 ( .A(core__abc_21302_new_n2168__bF_buf2), .B(core__abc_21302_new_n4058_), .C(core__abc_21302_new_n2673__bF_buf7), .D(core__abc_21302_new_n4057_), .Y(core__abc_21302_new_n4059_));
OAI22X1 OAI22X1_103 ( .A(core__abc_21302_new_n2168__bF_buf1), .B(core__abc_21302_new_n4086_), .C(core_key_101_), .D(core__abc_21302_new_n2640__bF_buf9), .Y(core__abc_21302_new_n4087_));
OAI22X1 OAI22X1_104 ( .A(core__abc_21302_new_n2168__bF_buf0), .B(core__abc_21302_new_n4121_), .C(core_key_102_), .D(core__abc_21302_new_n2640__bF_buf8), .Y(core__abc_21302_new_n4122_));
OAI22X1 OAI22X1_105 ( .A(core__abc_21302_new_n2168__bF_buf11), .B(core__abc_21302_new_n4186_), .C(core__abc_21302_new_n2673__bF_buf4), .D(core__abc_21302_new_n4185_), .Y(core__abc_21302_new_n4187_));
OAI22X1 OAI22X1_106 ( .A(core__abc_21302_new_n2168__bF_buf10), .B(core__abc_21302_new_n4213_), .C(core__abc_21302_new_n4212_), .D(core__abc_21302_new_n2640__bF_buf7), .Y(core__abc_21302_new_n4214_));
OAI22X1 OAI22X1_107 ( .A(core__abc_21302_new_n2168__bF_buf9), .B(core__abc_21302_new_n4244_), .C(core_key_106_), .D(core__abc_21302_new_n2640__bF_buf6), .Y(core__abc_21302_new_n4245_));
OAI22X1 OAI22X1_108 ( .A(core__abc_21302_new_n2168__bF_buf8), .B(core__abc_21302_new_n4295_), .C(core__abc_21302_new_n4294_), .D(core__abc_21302_new_n2640__bF_buf4), .Y(core__abc_21302_new_n4296_));
OAI22X1 OAI22X1_109 ( .A(core__abc_21302_new_n2168__bF_buf7), .B(core__abc_21302_new_n4318_), .C(core_key_109_), .D(core__abc_21302_new_n2640__bF_buf3), .Y(core__abc_21302_new_n4319_));
OAI22X1 OAI22X1_11 ( .A(_abc_19873_new_n992_), .B(_abc_19873_new_n913__bF_buf1), .C(_abc_19873_new_n993_), .D(_abc_19873_new_n894__bF_buf1), .Y(_abc_19873_new_n994_));
OAI22X1 OAI22X1_110 ( .A(core__abc_21302_new_n2168__bF_buf6), .B(core__abc_21302_new_n4353_), .C(core_key_110_), .D(core__abc_21302_new_n2640__bF_buf2), .Y(core__abc_21302_new_n4354_));
OAI22X1 OAI22X1_111 ( .A(core__abc_21302_new_n2168__bF_buf4), .B(core__abc_21302_new_n4406_), .C(core__abc_21302_new_n2673__bF_buf8), .D(core__abc_21302_new_n4405_), .Y(core__abc_21302_new_n4407_));
OAI22X1 OAI22X1_112 ( .A(core__abc_21302_new_n2168__bF_buf3), .B(core__abc_21302_new_n4438_), .C(core__abc_21302_new_n4437_), .D(core__abc_21302_new_n2640__bF_buf0), .Y(core__abc_21302_new_n4439_));
OAI22X1 OAI22X1_113 ( .A(core__abc_21302_new_n2168__bF_buf2), .B(core__abc_21302_new_n4465_), .C(core_key_114_), .D(core__abc_21302_new_n2640__bF_buf11), .Y(core__abc_21302_new_n4466_));
OAI22X1 OAI22X1_114 ( .A(core__abc_21302_new_n2168__bF_buf1), .B(core__abc_21302_new_n4487_), .C(core__abc_21302_new_n4486_), .D(core__abc_21302_new_n2640__bF_buf10), .Y(core__abc_21302_new_n4488_));
OAI22X1 OAI22X1_115 ( .A(core__abc_21302_new_n2168__bF_buf0), .B(core__abc_21302_new_n4510_), .C(core__abc_21302_new_n2673__bF_buf4), .D(core__abc_21302_new_n4509_), .Y(core__abc_21302_new_n4511_));
OAI22X1 OAI22X1_116 ( .A(core__abc_21302_new_n2168__bF_buf12), .B(core__abc_21302_new_n4534_), .C(core_key_117_), .D(core__abc_21302_new_n2640__bF_buf9), .Y(core__abc_21302_new_n4535_));
OAI22X1 OAI22X1_117 ( .A(core__abc_21302_new_n2168__bF_buf11), .B(core__abc_21302_new_n4559_), .C(core_key_118_), .D(core__abc_21302_new_n2640__bF_buf8), .Y(core__abc_21302_new_n4560_));
OAI22X1 OAI22X1_118 ( .A(core__abc_21302_new_n2168__bF_buf9), .B(core__abc_21302_new_n4612_), .C(core__abc_21302_new_n2673__bF_buf0), .D(core__abc_21302_new_n4611_), .Y(core__abc_21302_new_n4613_));
OAI22X1 OAI22X1_119 ( .A(core__abc_21302_new_n2168__bF_buf7), .B(core__abc_21302_new_n4667_), .C(core_key_122_), .D(core__abc_21302_new_n2640__bF_buf7), .Y(core__abc_21302_new_n4668_));
OAI22X1 OAI22X1_12 ( .A(_abc_19873_new_n1000_), .B(_abc_19873_new_n914__bF_buf0), .C(_abc_19873_new_n999_), .D(_abc_19873_new_n969__bF_buf1), .Y(_abc_19873_new_n1001_));
OAI22X1 OAI22X1_120 ( .A(core__abc_21302_new_n4136_), .B(core__abc_21302_new_n4137_), .C(core__abc_21302_new_n4719_), .D(core__abc_21302_new_n4721_), .Y(core__abc_21302_new_n4722_));
OAI22X1 OAI22X1_121 ( .A(core__abc_21302_new_n2168__bF_buf6), .B(core__abc_21302_new_n4726_), .C(core_key_124_), .D(core__abc_21302_new_n2640__bF_buf5), .Y(core__abc_21302_new_n4727_));
OAI22X1 OAI22X1_122 ( .A(core__abc_21302_new_n2168__bF_buf5), .B(core__abc_21302_new_n4758_), .C(core_key_125_), .D(core__abc_21302_new_n2640__bF_buf4), .Y(core__abc_21302_new_n4759_));
OAI22X1 OAI22X1_123 ( .A(core__abc_21302_new_n2168__bF_buf4), .B(core__abc_21302_new_n4791_), .C(core_key_126_), .D(core__abc_21302_new_n2640__bF_buf3), .Y(core__abc_21302_new_n4792_));
OAI22X1 OAI22X1_124 ( .A(core_v2_reg_5_), .B(core__abc_21302_new_n2364__bF_buf0), .C(core_key_5_), .D(core__abc_21302_new_n2640__bF_buf10), .Y(core__abc_21302_new_n5183_));
OAI22X1 OAI22X1_125 ( .A(core_v2_reg_7_), .B(core__abc_21302_new_n2364__bF_buf4), .C(core__abc_21302_new_n5221_), .D(core__abc_21302_new_n2640__bF_buf8), .Y(core__abc_21302_new_n5222_));
OAI22X1 OAI22X1_126 ( .A(core__abc_21302_new_n1328_), .B(core__abc_21302_new_n2364__bF_buf3), .C(core__abc_21302_new_n5297_), .D(core__abc_21302_new_n2640__bF_buf6), .Y(core__abc_21302_new_n5298_));
OAI22X1 OAI22X1_127 ( .A(core__abc_21302_new_n1350_), .B(core__abc_21302_new_n2364__bF_buf2), .C(core_key_13_), .D(core__abc_21302_new_n2640__bF_buf4), .Y(core__abc_21302_new_n5338_));
OAI22X1 OAI22X1_128 ( .A(core__abc_21302_new_n1362_), .B(core__abc_21302_new_n2364__bF_buf1), .C(core_key_14_), .D(core__abc_21302_new_n2640__bF_buf3), .Y(core__abc_21302_new_n5363_));
OAI22X1 OAI22X1_129 ( .A(core__abc_21302_new_n1373_), .B(core__abc_21302_new_n2364__bF_buf0), .C(core__abc_21302_new_n5382_), .D(core__abc_21302_new_n2640__bF_buf2), .Y(core__abc_21302_new_n5383_));
OAI22X1 OAI22X1_13 ( .A(_abc_19873_new_n1013_), .B(_abc_19873_new_n913__bF_buf0), .C(_abc_19873_new_n1014_), .D(_abc_19873_new_n894__bF_buf0), .Y(_abc_19873_new_n1015_));
OAI22X1 OAI22X1_130 ( .A(core__abc_21302_new_n1409_), .B(core__abc_21302_new_n2364__bF_buf4), .C(core_key_18_), .D(core__abc_21302_new_n2640__bF_buf0), .Y(core__abc_21302_new_n5450_));
OAI22X1 OAI22X1_131 ( .A(core__abc_21302_new_n1421_), .B(core__abc_21302_new_n2364__bF_buf3), .C(core__abc_21302_new_n5460_), .D(core__abc_21302_new_n2640__bF_buf11), .Y(core__abc_21302_new_n5461_));
OAI22X1 OAI22X1_132 ( .A(core__abc_21302_new_n1445_), .B(core__abc_21302_new_n2364__bF_buf1), .C(core_key_21_), .D(core__abc_21302_new_n2640__bF_buf10), .Y(core__abc_21302_new_n5502_));
OAI22X1 OAI22X1_133 ( .A(core__abc_21302_new_n1457_), .B(core__abc_21302_new_n2364__bF_buf0), .C(core_key_22_), .D(core__abc_21302_new_n2640__bF_buf9), .Y(core__abc_21302_new_n5523_));
OAI22X1 OAI22X1_134 ( .A(core__abc_21302_new_n2581_), .B(core__abc_21302_new_n2364__bF_buf5), .C(core__abc_21302_new_n5540_), .D(core__abc_21302_new_n2640__bF_buf8), .Y(core__abc_21302_new_n5541_));
OAI22X1 OAI22X1_135 ( .A(core__abc_21302_new_n1487_), .B(core__abc_21302_new_n2364__bF_buf3), .C(core_key_25_), .D(core__abc_21302_new_n2640__bF_buf7), .Y(core__abc_21302_new_n5579_));
OAI22X1 OAI22X1_136 ( .A(core__abc_21302_new_n1499_), .B(core__abc_21302_new_n2364__bF_buf2), .C(core_key_26_), .D(core__abc_21302_new_n2640__bF_buf6), .Y(core__abc_21302_new_n5596_));
OAI22X1 OAI22X1_137 ( .A(core__abc_21302_new_n1511_), .B(core__abc_21302_new_n2364__bF_buf1), .C(core_key_27_), .D(core__abc_21302_new_n2640__bF_buf5), .Y(core__abc_21302_new_n5613_));
OAI22X1 OAI22X1_138 ( .A(core__abc_21302_new_n1536_), .B(core__abc_21302_new_n2364__bF_buf5), .C(core_key_29_), .D(core__abc_21302_new_n2640__bF_buf4), .Y(core__abc_21302_new_n5658_));
OAI22X1 OAI22X1_139 ( .A(core__abc_21302_new_n1548_), .B(core__abc_21302_new_n2364__bF_buf4), .C(core_key_30_), .D(core__abc_21302_new_n2640__bF_buf3), .Y(core__abc_21302_new_n5678_));
OAI22X1 OAI22X1_14 ( .A(_abc_19873_new_n1021_), .B(_abc_19873_new_n918_), .C(_abc_19873_new_n1020_), .D(_abc_19873_new_n894__bF_buf4), .Y(_abc_19873_new_n1022_));
OAI22X1 OAI22X1_140 ( .A(core__abc_21302_new_n2587_), .B(core__abc_21302_new_n2364__bF_buf3), .C(core__abc_21302_new_n5694_), .D(core__abc_21302_new_n2640__bF_buf2), .Y(core__abc_21302_new_n5695_));
OAI22X1 OAI22X1_141 ( .A(core__abc_21302_new_n1593_), .B(core__abc_21302_new_n2364__bF_buf2), .C(core_key_34_), .D(core__abc_21302_new_n2640__bF_buf0), .Y(core__abc_21302_new_n5716_));
OAI22X1 OAI22X1_142 ( .A(core__abc_21302_new_n1606_), .B(core__abc_21302_new_n2364__bF_buf1), .C(core__abc_21302_new_n5723_), .D(core__abc_21302_new_n2640__bF_buf11), .Y(core__abc_21302_new_n5724_));
OAI22X1 OAI22X1_143 ( .A(core__abc_21302_new_n1823_), .B(core__abc_21302_new_n2364__bF_buf0), .C(core_key_54_), .D(core__abc_21302_new_n2640__bF_buf9), .Y(core__abc_21302_new_n5904_));
OAI22X1 OAI22X1_144 ( .A(core__abc_21302_new_n1836_), .B(core__abc_21302_new_n2364__bF_buf5), .C(core__abc_21302_new_n5915_), .D(core__abc_21302_new_n2640__bF_buf8), .Y(core__abc_21302_new_n5916_));
OAI22X1 OAI22X1_145 ( .A(core__abc_21302_new_n1916_), .B(core__abc_21302_new_n2364__bF_buf3), .C(core_key_61_), .D(core__abc_21302_new_n2640__bF_buf5), .Y(core__abc_21302_new_n5971_));
OAI22X1 OAI22X1_146 ( .A(core__abc_21302_new_n1929_), .B(core__abc_21302_new_n2364__bF_buf2), .C(core_key_62_), .D(core__abc_21302_new_n2640__bF_buf4), .Y(core__abc_21302_new_n5980_));
OAI22X1 OAI22X1_147 ( .A(core_v1_reg_3_), .B(core__abc_21302_new_n5999__bF_buf3), .C(core__abc_21302_new_n2640__bF_buf2), .D(core__abc_21302_new_n6026_), .Y(core__abc_21302_new_n6027_));
OAI22X1 OAI22X1_148 ( .A(core_v1_reg_6_), .B(core__abc_21302_new_n5999__bF_buf0), .C(core__abc_21302_new_n2673__bF_buf10), .D(core__abc_21302_new_n6049_), .Y(core__abc_21302_new_n6050_));
OAI22X1 OAI22X1_149 ( .A(core_v1_reg_7_), .B(core__abc_21302_new_n5999__bF_buf5), .C(core__abc_21302_new_n2640__bF_buf0), .D(core__abc_21302_new_n6057_), .Y(core__abc_21302_new_n6058_));
OAI22X1 OAI22X1_15 ( .A(_abc_19873_new_n1032_), .B(_abc_19873_new_n913__bF_buf4), .C(_abc_19873_new_n1031_), .D(_abc_19873_new_n914__bF_buf4), .Y(_abc_19873_new_n1033_));
OAI22X1 OAI22X1_150 ( .A(core__abc_21302_new_n4248_), .B(core__abc_21302_new_n5999__bF_buf3), .C(core__abc_21302_new_n6075_), .D(core__abc_21302_new_n6076_), .Y(core__abc_21302_new_n6077_));
OAI22X1 OAI22X1_151 ( .A(core__abc_21302_new_n4868_), .B(core__abc_21302_new_n5999__bF_buf2), .C(core__abc_21302_new_n6088_), .D(core__abc_21302_new_n6089_), .Y(core__abc_21302_new_n6090_));
OAI22X1 OAI22X1_152 ( .A(core_v1_reg_13_), .B(core__abc_21302_new_n6009__bF_buf8), .C(core__abc_21302_new_n6097_), .D(core__abc_21302_new_n6095_), .Y(core__abc_21302_new_n6098_));
OAI22X1 OAI22X1_153 ( .A(core__abc_21302_new_n2436_), .B(core__abc_21302_new_n5999__bF_buf5), .C(core__abc_21302_new_n6113_), .D(core__abc_21302_new_n6114_), .Y(core__abc_21302_new_n6115_));
OAI22X1 OAI22X1_154 ( .A(core__abc_21302_new_n5646_), .B(core__abc_21302_new_n5999__bF_buf2), .C(core__abc_21302_new_n6332_), .D(core__abc_21302_new_n6331_), .Y(core__abc_21302_new_n6333_));
OAI22X1 OAI22X1_16 ( .A(_abc_19873_new_n1034_), .B(_abc_19873_new_n924_), .C(_abc_19873_new_n1035_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1036_));
OAI22X1 OAI22X1_17 ( .A(_abc_19873_new_n1042_), .B(_abc_19873_new_n914__bF_buf3), .C(_abc_19873_new_n1041_), .D(_abc_19873_new_n969__bF_buf0), .Y(_abc_19873_new_n1043_));
OAI22X1 OAI22X1_18 ( .A(_abc_19873_new_n1045_), .B(_abc_19873_new_n918_), .C(_abc_19873_new_n1044_), .D(_abc_19873_new_n960__bF_buf0), .Y(_abc_19873_new_n1046_));
OAI22X1 OAI22X1_19 ( .A(_abc_19873_new_n1059_), .B(_abc_19873_new_n960__bF_buf4), .C(_abc_19873_new_n1060_), .D(_abc_19873_new_n896__bF_buf0), .Y(_abc_19873_new_n1061_));
OAI22X1 OAI22X1_2 ( .A(_abc_19873_new_n910_), .B(_abc_19873_new_n913__bF_buf4), .C(_abc_19873_new_n909_), .D(_abc_19873_new_n914__bF_buf4), .Y(_abc_19873_new_n915_));
OAI22X1 OAI22X1_20 ( .A(_abc_19873_new_n1062_), .B(_abc_19873_new_n1064__bF_buf3), .C(_abc_19873_new_n1063_), .D(_abc_19873_new_n969__bF_buf3), .Y(_abc_19873_new_n1065_));
OAI22X1 OAI22X1_21 ( .A(_abc_19873_new_n1075_), .B(_abc_19873_new_n913__bF_buf2), .C(_abc_19873_new_n1074_), .D(_abc_19873_new_n914__bF_buf2), .Y(_abc_19873_new_n1076_));
OAI22X1 OAI22X1_22 ( .A(_abc_19873_new_n1081_), .B(_abc_19873_new_n913__bF_buf1), .C(_abc_19873_new_n1082_), .D(_abc_19873_new_n894__bF_buf3), .Y(_abc_19873_new_n1083_));
OAI22X1 OAI22X1_23 ( .A(_abc_19873_new_n1085_), .B(_abc_19873_new_n1064__bF_buf2), .C(_abc_19873_new_n1084_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1086_));
OAI22X1 OAI22X1_24 ( .A(_abc_19873_new_n1091_), .B(_abc_19873_new_n960__bF_buf3), .C(_abc_19873_new_n1090_), .D(_abc_19873_new_n896__bF_buf4), .Y(_abc_19873_new_n1092_));
OAI22X1 OAI22X1_25 ( .A(_abc_19873_new_n1094_), .B(_abc_19873_new_n914__bF_buf1), .C(_abc_19873_new_n1093_), .D(_abc_19873_new_n969__bF_buf2), .Y(_abc_19873_new_n1095_));
OAI22X1 OAI22X1_26 ( .A(_abc_19873_new_n1100_), .B(_abc_19873_new_n913__bF_buf0), .C(_abc_19873_new_n1101_), .D(_abc_19873_new_n894__bF_buf2), .Y(_abc_19873_new_n1102_));
OAI22X1 OAI22X1_27 ( .A(_abc_19873_new_n1104_), .B(_abc_19873_new_n1064__bF_buf1), .C(_abc_19873_new_n1103_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1105_));
OAI22X1 OAI22X1_28 ( .A(_abc_19873_new_n1110_), .B(_abc_19873_new_n960__bF_buf2), .C(_abc_19873_new_n1109_), .D(_abc_19873_new_n896__bF_buf3), .Y(_abc_19873_new_n1111_));
OAI22X1 OAI22X1_29 ( .A(_abc_19873_new_n1113_), .B(_abc_19873_new_n914__bF_buf0), .C(_abc_19873_new_n1112_), .D(_abc_19873_new_n969__bF_buf1), .Y(_abc_19873_new_n1114_));
OAI22X1 OAI22X1_3 ( .A(_abc_19873_new_n921_), .B(_abc_19873_new_n924_), .C(_abc_19873_new_n922_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n925_));
OAI22X1 OAI22X1_30 ( .A(_abc_19873_new_n1119_), .B(_abc_19873_new_n913__bF_buf4), .C(_abc_19873_new_n1120_), .D(_abc_19873_new_n894__bF_buf1), .Y(_abc_19873_new_n1121_));
OAI22X1 OAI22X1_31 ( .A(_abc_19873_new_n1123_), .B(_abc_19873_new_n1064__bF_buf0), .C(_abc_19873_new_n1122_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1124_));
OAI22X1 OAI22X1_32 ( .A(_abc_19873_new_n1129_), .B(_abc_19873_new_n960__bF_buf1), .C(_abc_19873_new_n1128_), .D(_abc_19873_new_n896__bF_buf2), .Y(_abc_19873_new_n1130_));
OAI22X1 OAI22X1_33 ( .A(_abc_19873_new_n1132_), .B(_abc_19873_new_n914__bF_buf4), .C(_abc_19873_new_n1131_), .D(_abc_19873_new_n969__bF_buf0), .Y(_abc_19873_new_n1133_));
OAI22X1 OAI22X1_34 ( .A(_abc_19873_new_n1137_), .B(_abc_19873_new_n913__bF_buf3), .C(_abc_19873_new_n1136_), .D(_abc_19873_new_n914__bF_buf3), .Y(_abc_19873_new_n1138_));
OAI22X1 OAI22X1_35 ( .A(_abc_19873_new_n1150_), .B(_abc_19873_new_n1064__bF_buf3), .C(_abc_19873_new_n1151_), .D(_abc_19873_new_n969__bF_buf3), .Y(_abc_19873_new_n1152_));
OAI22X1 OAI22X1_36 ( .A(_abc_19873_new_n1156_), .B(_abc_19873_new_n913__bF_buf2), .C(_abc_19873_new_n1155_), .D(_abc_19873_new_n914__bF_buf2), .Y(_abc_19873_new_n1157_));
OAI22X1 OAI22X1_37 ( .A(_abc_19873_new_n1169_), .B(_abc_19873_new_n1064__bF_buf2), .C(_abc_19873_new_n1170_), .D(_abc_19873_new_n969__bF_buf2), .Y(_abc_19873_new_n1171_));
OAI22X1 OAI22X1_38 ( .A(_abc_19873_new_n1175_), .B(_abc_19873_new_n960__bF_buf3), .C(_abc_19873_new_n1174_), .D(_abc_19873_new_n896__bF_buf1), .Y(_abc_19873_new_n1176_));
OAI22X1 OAI22X1_39 ( .A(_abc_19873_new_n1179_), .B(_abc_19873_new_n913__bF_buf1), .C(_abc_19873_new_n1180_), .D(_abc_19873_new_n894__bF_buf3), .Y(_abc_19873_new_n1181_));
OAI22X1 OAI22X1_4 ( .A(_abc_19873_new_n933_), .B(_abc_19873_new_n894__bF_buf3), .C(_abc_19873_new_n934_), .D(_abc_19873_new_n896__bF_buf3), .Y(_abc_19873_new_n935_));
OAI22X1 OAI22X1_40 ( .A(_abc_19873_new_n1184_), .B(_abc_19873_new_n914__bF_buf1), .C(_abc_19873_new_n1183_), .D(_abc_19873_new_n969__bF_buf1), .Y(_abc_19873_new_n1185_));
OAI22X1 OAI22X1_41 ( .A(_abc_19873_new_n1193_), .B(_abc_19873_new_n913__bF_buf0), .C(_abc_19873_new_n1192_), .D(_abc_19873_new_n914__bF_buf0), .Y(_abc_19873_new_n1194_));
OAI22X1 OAI22X1_42 ( .A(_abc_19873_new_n1206_), .B(_abc_19873_new_n960__bF_buf2), .C(_abc_19873_new_n1205_), .D(_abc_19873_new_n896__bF_buf0), .Y(_abc_19873_new_n1207_));
OAI22X1 OAI22X1_43 ( .A(_abc_19873_new_n1212_), .B(_abc_19873_new_n913__bF_buf4), .C(_abc_19873_new_n1213_), .D(_abc_19873_new_n894__bF_buf1), .Y(_abc_19873_new_n1214_));
OAI22X1 OAI22X1_44 ( .A(_abc_19873_new_n1216_), .B(_abc_19873_new_n1064__bF_buf0), .C(_abc_19873_new_n1215_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1217_));
OAI22X1 OAI22X1_45 ( .A(_abc_19873_new_n1222_), .B(_abc_19873_new_n960__bF_buf1), .C(_abc_19873_new_n1221_), .D(_abc_19873_new_n896__bF_buf4), .Y(_abc_19873_new_n1223_));
OAI22X1 OAI22X1_46 ( .A(_abc_19873_new_n1225_), .B(_abc_19873_new_n914__bF_buf4), .C(_abc_19873_new_n1224_), .D(_abc_19873_new_n969__bF_buf0), .Y(_abc_19873_new_n1226_));
OAI22X1 OAI22X1_47 ( .A(_abc_19873_new_n1230_), .B(_abc_19873_new_n913__bF_buf3), .C(_abc_19873_new_n1229_), .D(_abc_19873_new_n914__bF_buf3), .Y(_abc_19873_new_n1231_));
OAI22X1 OAI22X1_48 ( .A(_abc_19873_new_n1243_), .B(_abc_19873_new_n960__bF_buf0), .C(_abc_19873_new_n1242_), .D(_abc_19873_new_n896__bF_buf3), .Y(_abc_19873_new_n1244_));
OAI22X1 OAI22X1_49 ( .A(_abc_19873_new_n1250_), .B(_abc_19873_new_n1064__bF_buf2), .C(_abc_19873_new_n1251_), .D(_abc_19873_new_n969__bF_buf3), .Y(_abc_19873_new_n1252_));
OAI22X1 OAI22X1_5 ( .A(_abc_19873_new_n942_), .B(_abc_19873_new_n913__bF_buf3), .C(_abc_19873_new_n941_), .D(_abc_19873_new_n914__bF_buf3), .Y(_abc_19873_new_n943_));
OAI22X1 OAI22X1_50 ( .A(_abc_19873_new_n1254_), .B(_abc_19873_new_n894__bF_buf4), .C(_abc_19873_new_n1255_), .D(_abc_19873_new_n896__bF_buf2), .Y(_abc_19873_new_n1256_));
OAI22X1 OAI22X1_51 ( .A(_abc_19873_new_n1267_), .B(_abc_19873_new_n913__bF_buf1), .C(_abc_19873_new_n1266_), .D(_abc_19873_new_n914__bF_buf2), .Y(_abc_19873_new_n1268_));
OAI22X1 OAI22X1_52 ( .A(_abc_19873_new_n1279_), .B(_abc_19873_new_n1064__bF_buf1), .C(_abc_19873_new_n1280_), .D(_abc_19873_new_n969__bF_buf2), .Y(_abc_19873_new_n1281_));
OAI22X1 OAI22X1_53 ( .A(_abc_19873_new_n1285_), .B(_abc_19873_new_n913__bF_buf0), .C(_abc_19873_new_n1284_), .D(_abc_19873_new_n914__bF_buf1), .Y(_abc_19873_new_n1286_));
OAI22X1 OAI22X1_54 ( .A(_abc_19873_new_n1298_), .B(_abc_19873_new_n960__bF_buf2), .C(_abc_19873_new_n1297_), .D(_abc_19873_new_n896__bF_buf1), .Y(_abc_19873_new_n1299_));
OAI22X1 OAI22X1_55 ( .A(_abc_19873_new_n1303_), .B(_abc_19873_new_n913__bF_buf4), .C(_abc_19873_new_n1302_), .D(_abc_19873_new_n914__bF_buf0), .Y(_abc_19873_new_n1304_));
OAI22X1 OAI22X1_56 ( .A(_abc_19873_new_n1315_), .B(_abc_19873_new_n1064__bF_buf3), .C(_abc_19873_new_n1316_), .D(_abc_19873_new_n969__bF_buf1), .Y(_abc_19873_new_n1317_));
OAI22X1 OAI22X1_57 ( .A(_abc_19873_new_n1323_), .B(_abc_19873_new_n960__bF_buf0), .C(_abc_19873_new_n1322_), .D(_abc_19873_new_n896__bF_buf0), .Y(_abc_19873_new_n1324_));
OAI22X1 OAI22X1_58 ( .A(_abc_19873_new_n1325_), .B(_abc_19873_new_n913__bF_buf3), .C(_abc_19873_new_n1326_), .D(_abc_19873_new_n894__bF_buf0), .Y(_abc_19873_new_n1327_));
OAI22X1 OAI22X1_59 ( .A(_abc_19873_new_n1330_), .B(_abc_19873_new_n914__bF_buf4), .C(_abc_19873_new_n1329_), .D(_abc_19873_new_n969__bF_buf0), .Y(_abc_19873_new_n1331_));
OAI22X1 OAI22X1_6 ( .A(_abc_19873_new_n947_), .B(_abc_19873_new_n924_), .C(_abc_19873_new_n948_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n949_));
OAI22X1 OAI22X1_60 ( .A(_abc_19873_new_n1339_), .B(_abc_19873_new_n913__bF_buf2), .C(_abc_19873_new_n1338_), .D(_abc_19873_new_n914__bF_buf3), .Y(_abc_19873_new_n1340_));
OAI22X1 OAI22X1_61 ( .A(_abc_19873_new_n1352_), .B(_abc_19873_new_n960__bF_buf4), .C(_abc_19873_new_n1351_), .D(_abc_19873_new_n896__bF_buf4), .Y(_abc_19873_new_n1353_));
OAI22X1 OAI22X1_62 ( .A(_abc_19873_new_n1358_), .B(_abc_19873_new_n913__bF_buf1), .C(_abc_19873_new_n1359_), .D(_abc_19873_new_n894__bF_buf3), .Y(_abc_19873_new_n1360_));
OAI22X1 OAI22X1_63 ( .A(_abc_19873_new_n1362_), .B(_abc_19873_new_n1064__bF_buf1), .C(_abc_19873_new_n1361_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1363_));
OAI22X1 OAI22X1_64 ( .A(_abc_19873_new_n1368_), .B(_abc_19873_new_n960__bF_buf3), .C(_abc_19873_new_n1367_), .D(_abc_19873_new_n896__bF_buf3), .Y(_abc_19873_new_n1369_));
OAI22X1 OAI22X1_65 ( .A(_abc_19873_new_n1371_), .B(_abc_19873_new_n914__bF_buf2), .C(_abc_19873_new_n1370_), .D(_abc_19873_new_n969__bF_buf3), .Y(_abc_19873_new_n1372_));
OAI22X1 OAI22X1_66 ( .A(_abc_19873_new_n1376_), .B(_abc_19873_new_n913__bF_buf0), .C(_abc_19873_new_n1375_), .D(_abc_19873_new_n914__bF_buf1), .Y(_abc_19873_new_n1377_));
OAI22X1 OAI22X1_67 ( .A(_abc_19873_new_n1389_), .B(_abc_19873_new_n960__bF_buf2), .C(_abc_19873_new_n1388_), .D(_abc_19873_new_n896__bF_buf2), .Y(_abc_19873_new_n1390_));
OAI22X1 OAI22X1_68 ( .A(_abc_19873_new_n1394_), .B(_abc_19873_new_n913__bF_buf4), .C(_abc_19873_new_n1393_), .D(_abc_19873_new_n914__bF_buf0), .Y(_abc_19873_new_n1395_));
OAI22X1 OAI22X1_69 ( .A(_abc_19873_new_n1407_), .B(_abc_19873_new_n960__bF_buf1), .C(_abc_19873_new_n1406_), .D(_abc_19873_new_n896__bF_buf1), .Y(_abc_19873_new_n1408_));
OAI22X1 OAI22X1_7 ( .A(_abc_19873_new_n955_), .B(_abc_19873_new_n913__bF_buf2), .C(_abc_19873_new_n956_), .D(_abc_19873_new_n894__bF_buf2), .Y(_abc_19873_new_n957_));
OAI22X1 OAI22X1_70 ( .A(_abc_19873_new_n1413_), .B(_abc_19873_new_n913__bF_buf3), .C(_abc_19873_new_n1414_), .D(_abc_19873_new_n894__bF_buf0), .Y(_abc_19873_new_n1415_));
OAI22X1 OAI22X1_71 ( .A(_abc_19873_new_n1417_), .B(_abc_19873_new_n1064__bF_buf2), .C(_abc_19873_new_n1416_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1418_));
OAI22X1 OAI22X1_72 ( .A(_abc_19873_new_n1423_), .B(_abc_19873_new_n960__bF_buf0), .C(_abc_19873_new_n1422_), .D(_abc_19873_new_n896__bF_buf0), .Y(_abc_19873_new_n1424_));
OAI22X1 OAI22X1_73 ( .A(_abc_19873_new_n1426_), .B(_abc_19873_new_n914__bF_buf4), .C(_abc_19873_new_n1425_), .D(_abc_19873_new_n969__bF_buf2), .Y(_abc_19873_new_n1427_));
OAI22X1 OAI22X1_74 ( .A(_abc_19873_new_n1432_), .B(_abc_19873_new_n913__bF_buf2), .C(_abc_19873_new_n1433_), .D(_abc_19873_new_n894__bF_buf4), .Y(_abc_19873_new_n1434_));
OAI22X1 OAI22X1_75 ( .A(_abc_19873_new_n1436_), .B(_abc_19873_new_n1064__bF_buf1), .C(_abc_19873_new_n1435_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1437_));
OAI22X1 OAI22X1_76 ( .A(_abc_19873_new_n1442_), .B(_abc_19873_new_n960__bF_buf4), .C(_abc_19873_new_n1441_), .D(_abc_19873_new_n896__bF_buf4), .Y(_abc_19873_new_n1443_));
OAI22X1 OAI22X1_77 ( .A(_abc_19873_new_n1445_), .B(_abc_19873_new_n914__bF_buf3), .C(_abc_19873_new_n1444_), .D(_abc_19873_new_n969__bF_buf1), .Y(_abc_19873_new_n1446_));
OAI22X1 OAI22X1_78 ( .A(_abc_19873_new_n1450_), .B(_abc_19873_new_n913__bF_buf1), .C(_abc_19873_new_n1449_), .D(_abc_19873_new_n914__bF_buf2), .Y(_abc_19873_new_n1451_));
OAI22X1 OAI22X1_79 ( .A(_abc_19873_new_n1463_), .B(_abc_19873_new_n960__bF_buf3), .C(_abc_19873_new_n1462_), .D(_abc_19873_new_n896__bF_buf3), .Y(_abc_19873_new_n1464_));
OAI22X1 OAI22X1_8 ( .A(_abc_19873_new_n959_), .B(_abc_19873_new_n960__bF_buf4), .C(_abc_19873_new_n958_), .D(_abc_19873_new_n896__bF_buf2), .Y(_abc_19873_new_n961_));
OAI22X1 OAI22X1_80 ( .A(_abc_19873_new_n1468_), .B(_abc_19873_new_n1064__bF_buf3), .C(_abc_19873_new_n1467_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1469_));
OAI22X1 OAI22X1_81 ( .A(_abc_19873_new_n1470_), .B(_abc_19873_new_n924_), .C(_abc_19873_new_n1471_), .D(_abc_19873_new_n953_), .Y(_abc_19873_new_n1472_));
OAI22X1 OAI22X1_82 ( .A(_abc_19873_new_n1477_), .B(_abc_19873_new_n894__bF_buf2), .C(_abc_19873_new_n1478_), .D(_abc_19873_new_n896__bF_buf2), .Y(_abc_19873_new_n1479_));
OAI22X1 OAI22X1_83 ( .A(_abc_19873_new_n1488_), .B(_abc_19873_new_n913__bF_buf0), .C(_abc_19873_new_n1487_), .D(_abc_19873_new_n914__bF_buf1), .Y(_abc_19873_new_n1489_));
OAI22X1 OAI22X1_84 ( .A(_abc_19873_new_n1501_), .B(_abc_19873_new_n960__bF_buf2), .C(_abc_19873_new_n1500_), .D(_abc_19873_new_n896__bF_buf1), .Y(_abc_19873_new_n1502_));
OAI22X1 OAI22X1_85 ( .A(_abc_19873_new_n1507_), .B(_abc_19873_new_n913__bF_buf4), .C(_abc_19873_new_n1508_), .D(_abc_19873_new_n894__bF_buf0), .Y(_abc_19873_new_n1509_));
OAI22X1 OAI22X1_86 ( .A(_abc_19873_new_n1511_), .B(_abc_19873_new_n1064__bF_buf1), .C(_abc_19873_new_n1510_), .D(_abc_19873_new_n923_), .Y(_abc_19873_new_n1512_));
OAI22X1 OAI22X1_87 ( .A(_abc_19873_new_n1517_), .B(_abc_19873_new_n960__bF_buf1), .C(_abc_19873_new_n1516_), .D(_abc_19873_new_n896__bF_buf0), .Y(_abc_19873_new_n1518_));
OAI22X1 OAI22X1_88 ( .A(_abc_19873_new_n1520_), .B(_abc_19873_new_n914__bF_buf0), .C(_abc_19873_new_n1519_), .D(_abc_19873_new_n969__bF_buf0), .Y(_abc_19873_new_n1521_));
OAI22X1 OAI22X1_89 ( .A(core__abc_21302_new_n1184_), .B(core__abc_21302_new_n1147_), .C(core__abc_21302_new_n1152_), .D(core__abc_21302_new_n1175_), .Y(core__abc_21302_new_n1190_));
OAI22X1 OAI22X1_9 ( .A(_abc_19873_new_n968_), .B(_abc_19873_new_n914__bF_buf2), .C(_abc_19873_new_n967_), .D(_abc_19873_new_n969__bF_buf3), .Y(_abc_19873_new_n970_));
OAI22X1 OAI22X1_90 ( .A(core__abc_21302_new_n1194_), .B(core__abc_21302_new_n1185__bF_buf11), .C(core__abc_21302_new_n1195_), .D(core__abc_21302_new_n1196_), .Y(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_3_));
OAI22X1 OAI22X1_91 ( .A(core__abc_21302_new_n1200_), .B(core__abc_21302_new_n1201_), .C(core__abc_21302_new_n1188_), .D(core__abc_21302_new_n1196_), .Y(core__abc_15204_auto_fsm_map_cc_170_map_fsm_1439_4_));
OAI22X1 OAI22X1_92 ( .A(core__abc_21302_new_n2168__bF_buf0), .B(core__abc_21302_new_n2676_), .C(core_key_65_), .D(core__abc_21302_new_n2640__bF_buf10), .Y(core__abc_21302_new_n2677_));
OAI22X1 OAI22X1_93 ( .A(core__abc_21302_new_n2168__bF_buf3), .B(core__abc_21302_new_n3324_), .C(core__abc_21302_new_n2673__bF_buf11), .D(core__abc_21302_new_n3323_), .Y(core__abc_21302_new_n3325_));
OAI22X1 OAI22X1_94 ( .A(core__abc_21302_new_n3459_), .B(core__abc_21302_new_n3463_), .C(core__abc_21302_new_n3374_), .D(core__abc_21302_new_n3460_), .Y(core__abc_21302_new_n3464_));
OAI22X1 OAI22X1_95 ( .A(core__abc_21302_new_n2168__bF_buf0), .B(core__abc_21302_new_n3494_), .C(core_key_84_), .D(core__abc_21302_new_n2640__bF_buf10), .Y(core__abc_21302_new_n3495_));
OAI22X1 OAI22X1_96 ( .A(core__abc_21302_new_n2168__bF_buf9), .B(core__abc_21302_new_n3720_), .C(core__abc_21302_new_n3718_), .D(core__abc_21302_new_n3719_), .Y(core__abc_21302_new_n3721_));
OAI22X1 OAI22X1_97 ( .A(core__abc_21302_new_n2168__bF_buf8), .B(core__abc_21302_new_n3786_), .C(core_key_92_), .D(core__abc_21302_new_n2640__bF_buf3), .Y(core__abc_21302_new_n3787_));
OAI22X1 OAI22X1_98 ( .A(core__abc_21302_new_n2168__bF_buf7), .B(core__abc_21302_new_n3872_), .C(core__abc_21302_new_n3870_), .D(core__abc_21302_new_n3871_), .Y(core__abc_21302_new_n3873_));
OAI22X1 OAI22X1_99 ( .A(core__abc_21302_new_n2168__bF_buf5), .B(core__abc_21302_new_n3938_), .C(core__abc_21302_new_n3937_), .D(core__abc_21302_new_n2640__bF_buf0), .Y(core__abc_21302_new_n3939_));
OR2X2 OR2X2_1 ( .A(\addr[0] ), .B(\addr[1] ), .Y(_abc_19873_new_n871_));
OR2X2 OR2X2_10 ( .A(core_v1_reg_3_), .B(core_v0_reg_3_), .Y(core__abc_21302_new_n1241_));
OR2X2 OR2X2_100 ( .A(core__abc_21302_new_n5151_), .B(core__abc_21302_new_n4049_), .Y(core__abc_21302_new_n5153_));
OR2X2 OR2X2_101 ( .A(core__abc_21302_new_n5167_), .B(core__abc_21302_new_n5163_), .Y(core__abc_21302_new_n5168_));
OR2X2 OR2X2_102 ( .A(core__abc_21302_new_n5254_), .B(core__abc_21302_new_n5241_), .Y(core__abc_21302_new_n5262_));
OR2X2 OR2X2_103 ( .A(core__abc_21302_new_n5271_), .B(core__abc_21302_new_n5267_), .Y(core__abc_21302_new_n5272_));
OR2X2 OR2X2_104 ( .A(core__abc_21302_new_n5276_), .B(core__abc_21302_new_n5274_), .Y(core__abc_21302_new_n5277_));
OR2X2 OR2X2_105 ( .A(core__abc_21302_new_n5285_), .B(core__abc_21302_new_n5293_), .Y(core__abc_21302_new_n5294_));
OR2X2 OR2X2_106 ( .A(core__abc_21302_new_n5262_), .B(core__abc_21302_new_n5303_), .Y(core__abc_21302_new_n5309_));
OR2X2 OR2X2_107 ( .A(core__abc_21302_new_n5312_), .B(core__abc_21302_new_n2668_), .Y(core__abc_21302_new_n5313_));
OR2X2 OR2X2_108 ( .A(core__abc_21302_new_n5324_), .B(core__abc_21302_new_n5333_), .Y(core__abc_21302_new_n5335_));
OR2X2 OR2X2_109 ( .A(core__abc_21302_new_n5423_), .B(core__abc_21302_new_n2868_), .Y(core__abc_21302_new_n5425_));
OR2X2 OR2X2_11 ( .A(core_v1_reg_4_), .B(core_v0_reg_4_), .Y(core__abc_21302_new_n1251_));
OR2X2 OR2X2_110 ( .A(core__abc_21302_new_n5454_), .B(core__abc_21302_new_n5456_), .Y(core__abc_21302_new_n5457_));
OR2X2 OR2X2_111 ( .A(core__abc_21302_new_n3030_), .B(core__abc_21302_new_n5493_), .Y(core__abc_21302_new_n5495_));
OR2X2 OR2X2_112 ( .A(core__abc_21302_new_n5534_), .B(core__abc_21302_new_n5513_), .Y(core__abc_21302_new_n5545_));
OR2X2 OR2X2_113 ( .A(core__abc_21302_new_n5547_), .B(core__abc_21302_new_n5550_), .Y(core__abc_21302_new_n5551_));
OR2X2 OR2X2_114 ( .A(core__abc_21302_new_n5583_), .B(core__abc_21302_new_n5584_), .Y(core__abc_21302_new_n5585_));
OR2X2 OR2X2_115 ( .A(core__abc_21302_new_n5622_), .B(core__abc_21302_new_n5623_), .Y(core__abc_21302_new_n5635_));
OR2X2 OR2X2_116 ( .A(core__abc_21302_new_n5645_), .B(core__abc_21302_new_n5647_), .Y(core__abc_21302_new_n5648_));
OR2X2 OR2X2_117 ( .A(core__abc_21302_new_n5667_), .B(core__abc_21302_new_n5670_), .Y(core__abc_21302_new_n5671_));
OR2X2 OR2X2_118 ( .A(core__abc_21302_new_n5085__bF_buf4), .B(core__abc_21302_new_n5733_), .Y(core__abc_21302_new_n5734_));
OR2X2 OR2X2_119 ( .A(core__abc_21302_new_n2640__bF_buf7), .B(core_key_40_), .Y(core__abc_21302_new_n5767_));
OR2X2 OR2X2_12 ( .A(core_v1_reg_6_), .B(core_v0_reg_6_), .Y(core__abc_21302_new_n1273_));
OR2X2 OR2X2_120 ( .A(core__abc_21302_new_n5005_), .B(core__abc_21302_new_n5008_), .Y(core__abc_21302_new_n5799_));
OR2X2 OR2X2_121 ( .A(core__abc_21302_new_n2640__bF_buf2), .B(core_key_48_), .Y(core__abc_21302_new_n5844_));
OR2X2 OR2X2_122 ( .A(core__abc_21302_new_n5878_), .B(core__abc_21302_new_n4955_), .Y(core__abc_21302_new_n5881_));
OR2X2 OR2X2_123 ( .A(core__abc_21302_new_n4925_), .B(core__abc_21302_new_n3481_), .Y(core__abc_21302_new_n5890_));
OR2X2 OR2X2_124 ( .A(core__abc_21302_new_n5900_), .B(core__abc_21302_new_n5899_), .Y(core__abc_21302_new_n5901_));
OR2X2 OR2X2_125 ( .A(core__abc_21302_new_n5911_), .B(core__abc_21302_new_n5910_), .Y(core__abc_21302_new_n5912_));
OR2X2 OR2X2_126 ( .A(core__abc_21302_new_n5072_), .B(core__abc_21302_new_n4892_), .Y(core__abc_21302_new_n5922_));
OR2X2 OR2X2_127 ( .A(core__abc_21302_new_n5976_), .B(core__abc_21302_new_n4837_), .Y(core__abc_21302_new_n5978_));
OR2X2 OR2X2_128 ( .A(core__abc_21302_new_n5883_), .B(core__abc_21302_new_n5037_), .Y(core__abc_21302_new_n6140_));
OR2X2 OR2X2_129 ( .A(core__abc_21302_new_n5079_), .B(core__abc_21302_new_n4984_), .Y(core__abc_21302_new_n6221_));
OR2X2 OR2X2_13 ( .A(core_v1_reg_7_), .B(core_v0_reg_7_), .Y(core__abc_21302_new_n1283_));
OR2X2 OR2X2_130 ( .A(core__abc_21302_new_n5199_), .B(core__abc_21302_new_n4956_), .Y(core__abc_21302_new_n6259_));
OR2X2 OR2X2_131 ( .A(core__abc_21302_new_n5316_), .B(core__abc_21302_new_n4857_), .Y(core__abc_21302_new_n6302_));
OR2X2 OR2X2_132 ( .A(core__abc_21302_new_n6906_), .B(core__abc_21302_new_n1203_), .Y(core__abc_21302_new_n6907_));
OR2X2 OR2X2_14 ( .A(core_v2_reg_8_), .B(core_v3_reg_8_), .Y(core__abc_21302_new_n1295_));
OR2X2 OR2X2_15 ( .A(core__abc_21302_new_n1383_), .B(core__abc_21302_new_n1382_), .Y(core__abc_21302_new_n1384_));
OR2X2 OR2X2_16 ( .A(core__abc_21302_new_n1394_), .B(core__abc_21302_new_n1393_), .Y(core__abc_21302_new_n1395_));
OR2X2 OR2X2_17 ( .A(core__abc_21302_new_n1569_), .B(core__abc_21302_new_n1570_), .Y(core__abc_21302_new_n1571_));
OR2X2 OR2X2_18 ( .A(core_v2_reg_33_), .B(core_v3_reg_33_), .Y(core__abc_21302_new_n1582_));
OR2X2 OR2X2_19 ( .A(core__abc_21302_new_n1603_), .B(core__abc_21302_new_n1602_), .Y(core__abc_21302_new_n1604_));
OR2X2 OR2X2_2 ( .A(\addr[7] ), .B(\addr[6] ), .Y(_abc_19873_new_n886_));
OR2X2 OR2X2_20 ( .A(core__abc_21302_new_n1619_), .B(core__abc_21302_new_n1617_), .Y(core__abc_21302_new_n1620_));
OR2X2 OR2X2_21 ( .A(core__abc_21302_new_n1631_), .B(core__abc_21302_new_n1632_), .Y(core__abc_21302_new_n1633_));
OR2X2 OR2X2_22 ( .A(core__abc_21302_new_n1641_), .B(core__abc_21302_new_n1639_), .Y(core__abc_21302_new_n1642_));
OR2X2 OR2X2_23 ( .A(core__abc_21302_new_n1648_), .B(core__abc_21302_new_n1647_), .Y(core__abc_21302_new_n1649_));
OR2X2 OR2X2_24 ( .A(core__abc_21302_new_n1651_), .B(core__abc_21302_new_n1652_), .Y(core__abc_21302_new_n1653_));
OR2X2 OR2X2_25 ( .A(core__abc_21302_new_n1662_), .B(core__abc_21302_new_n1663_), .Y(core__abc_21302_new_n1664_));
OR2X2 OR2X2_26 ( .A(core__abc_21302_new_n1673_), .B(core__abc_21302_new_n1674_), .Y(core__abc_21302_new_n1675_));
OR2X2 OR2X2_27 ( .A(core_v1_reg_45_), .B(core_v0_reg_45_), .Y(core__abc_21302_new_n1714_));
OR2X2 OR2X2_28 ( .A(core__abc_21302_new_n1731_), .B(core__abc_21302_new_n1729_), .Y(core__abc_21302_new_n1732_));
OR2X2 OR2X2_29 ( .A(core__abc_21302_new_n1742_), .B(core__abc_21302_new_n1740_), .Y(core__abc_21302_new_n1743_));
OR2X2 OR2X2_3 ( .A(\addr[3] ), .B(\addr[2] ), .Y(_abc_19873_new_n890_));
OR2X2 OR2X2_30 ( .A(core__abc_21302_new_n1313_), .B(core__abc_21302_new_n1325_), .Y(core__abc_21302_new_n2488_));
OR2X2 OR2X2_31 ( .A(core__abc_21302_new_n2428_), .B(core__abc_21302_new_n2429_), .Y(core__abc_21302_new_n2494_));
OR2X2 OR2X2_32 ( .A(core__abc_21302_new_n2641_), .B(core__abc_21302_new_n2643_), .Y(core__abc_21302_new_n2644_));
OR2X2 OR2X2_33 ( .A(core__abc_21302_new_n2622_), .B(core__abc_21302_new_n2660_), .Y(core__abc_21302_new_n2663_));
OR2X2 OR2X2_34 ( .A(core__abc_21302_new_n2517_), .B(core__abc_21302_new_n1237_), .Y(core__abc_21302_new_n2691_));
OR2X2 OR2X2_35 ( .A(core__abc_21302_new_n1719_), .B(core__abc_21302_new_n1717_), .Y(core__abc_21302_new_n2701_));
OR2X2 OR2X2_36 ( .A(core__abc_21302_new_n2726_), .B(core__abc_21302_new_n2725_), .Y(core__abc_21302_new_n2730_));
OR2X2 OR2X2_37 ( .A(core__abc_21302_new_n2739_), .B(core__abc_21302_new_n2746_), .Y(core__abc_21302_new_n2747_));
OR2X2 OR2X2_38 ( .A(core__abc_21302_new_n2765_), .B(core__abc_21302_new_n2683_), .Y(core__abc_21302_new_n2766_));
OR2X2 OR2X2_39 ( .A(core__abc_21302_new_n2898_), .B(core__abc_21302_new_n1765_), .Y(core__abc_21302_new_n2899_));
OR2X2 OR2X2_4 ( .A(_abc_19873_new_n969__bF_buf3), .B(_abc_19873_new_n1848_), .Y(_abc_19873_new_n1849_));
OR2X2 OR2X2_40 ( .A(core__abc_21302_new_n2766_), .B(core__abc_21302_new_n2922_), .Y(core__abc_21302_new_n2934_));
OR2X2 OR2X2_41 ( .A(core__abc_21302_new_n2949_), .B(core__abc_21302_new_n2948_), .Y(core__abc_21302_new_n2950_));
OR2X2 OR2X2_42 ( .A(core__abc_21302_new_n3026_), .B(core__abc_21302_new_n1814_), .Y(core__abc_21302_new_n3027_));
OR2X2 OR2X2_43 ( .A(core__abc_21302_new_n3030_), .B(core_v3_reg_37_), .Y(core__abc_21302_new_n3031_));
OR2X2 OR2X2_44 ( .A(core__abc_21302_new_n3050_), .B(core__abc_21302_new_n1331_), .Y(core__abc_21302_new_n3051_));
OR2X2 OR2X2_45 ( .A(core__abc_21302_new_n3053_), .B(core_v3_reg_59_), .Y(core__abc_21302_new_n3055_));
OR2X2 OR2X2_46 ( .A(core__abc_21302_new_n3138_), .B(core__abc_21302_new_n3137_), .Y(core__abc_21302_new_n3139_));
OR2X2 OR2X2_47 ( .A(core__abc_21302_new_n2987_), .B(core__abc_21302_new_n3064_), .Y(core__abc_21302_new_n3155_));
OR2X2 OR2X2_48 ( .A(core__abc_21302_new_n3161_), .B(core__abc_21302_new_n1853_), .Y(core__abc_21302_new_n3163_));
OR2X2 OR2X2_49 ( .A(core__abc_21302_new_n3164_), .B(core_v3_reg_40_), .Y(core__abc_21302_new_n3166_));
OR2X2 OR2X2_5 ( .A(_abc_19873_new_n914__bF_buf4), .B(_abc_19873_new_n1848_), .Y(_abc_19873_new_n1925_));
OR2X2 OR2X2_50 ( .A(core__abc_21302_new_n3223_), .B(core__abc_21302_new_n3242_), .Y(core__abc_21302_new_n3243_));
OR2X2 OR2X2_51 ( .A(core__abc_21302_new_n3248_), .B(core__abc_21302_new_n1879_), .Y(core__abc_21302_new_n3252_));
OR2X2 OR2X2_52 ( .A(core__abc_21302_new_n3108_), .B(core__abc_21302_new_n3101_), .Y(core__abc_21302_new_n3277_));
OR2X2 OR2X2_53 ( .A(core__abc_21302_new_n3333_), .B(core__abc_21302_new_n3336_), .Y(core__abc_21302_new_n3371_));
OR2X2 OR2X2_54 ( .A(core__abc_21302_new_n3382_), .B(core__abc_21302_new_n3377_), .Y(core__abc_21302_new_n3383_));
OR2X2 OR2X2_55 ( .A(core__abc_21302_new_n3420_), .B(core__abc_21302_new_n1424_), .Y(core__abc_21302_new_n3421_));
OR2X2 OR2X2_56 ( .A(core__abc_21302_new_n3433_), .B(core__abc_21302_new_n3429_), .Y(core__abc_21302_new_n3434_));
OR2X2 OR2X2_57 ( .A(core__abc_21302_new_n3416_), .B(core__abc_21302_new_n3435_), .Y(core__abc_21302_new_n3436_));
OR2X2 OR2X2_58 ( .A(core__abc_21302_new_n3478_), .B(core__abc_21302_new_n1436_), .Y(core__abc_21302_new_n3479_));
OR2X2 OR2X2_59 ( .A(core__abc_21302_new_n3482_), .B(core__abc_21302_new_n3476_), .Y(core__abc_21302_new_n3484_));
OR2X2 OR2X2_6 ( .A(_abc_19873_new_n913__bF_buf3), .B(_abc_19873_new_n1848_), .Y(_abc_19873_new_n1992_));
OR2X2 OR2X2_60 ( .A(core__abc_21302_new_n3549_), .B(core__abc_21302_new_n2575_), .Y(core__abc_21302_new_n3554_));
OR2X2 OR2X2_61 ( .A(core__abc_21302_new_n3575_), .B(core__abc_21302_new_n3592_), .Y(core__abc_21302_new_n3594_));
OR2X2 OR2X2_62 ( .A(core__abc_21302_new_n3622_), .B(core__abc_21302_new_n3624_), .Y(core__abc_21302_new_n3625_));
OR2X2 OR2X2_63 ( .A(core__abc_21302_new_n2574_), .B(core__abc_21302_new_n2585_), .Y(core__abc_21302_new_n3632_));
OR2X2 OR2X2_64 ( .A(core__abc_21302_new_n3729_), .B(core__abc_21302_new_n3748_), .Y(core__abc_21302_new_n3750_));
OR2X2 OR2X2_65 ( .A(core__abc_21302_new_n3690_), .B(core__abc_21302_new_n3761_), .Y(core__abc_21302_new_n3766_));
OR2X2 OR2X2_66 ( .A(core__abc_21302_new_n3933_), .B(core__abc_21302_new_n3059_), .Y(core__abc_21302_new_n3935_));
OR2X2 OR2X2_67 ( .A(core__abc_21302_new_n2375_), .B(core__abc_21302_new_n1234_), .Y(core__abc_21302_new_n3977_));
OR2X2 OR2X2_68 ( .A(core__abc_21302_new_n4003_), .B(core__abc_21302_new_n4018_), .Y(core__abc_21302_new_n4019_));
OR2X2 OR2X2_69 ( .A(core__abc_21302_new_n4079_), .B(core__abc_21302_new_n4078_), .Y(core__abc_21302_new_n4080_));
OR2X2 OR2X2_7 ( .A(_abc_19873_new_n894__bF_buf4), .B(_abc_19873_new_n1848_), .Y(_abc_19873_new_n2058_));
OR2X2 OR2X2_70 ( .A(core__abc_21302_new_n4096_), .B(core__abc_21302_new_n1275_), .Y(core__abc_21302_new_n4097_));
OR2X2 OR2X2_71 ( .A(core__abc_21302_new_n4100_), .B(core__abc_21302_new_n1642_), .Y(core__abc_21302_new_n4102_));
OR2X2 OR2X2_72 ( .A(core__abc_21302_new_n4117_), .B(core__abc_21302_new_n3343_), .Y(core__abc_21302_new_n4119_));
OR2X2 OR2X2_73 ( .A(core__abc_21302_new_n4127_), .B(core__abc_21302_new_n1653_), .Y(core__abc_21302_new_n4128_));
OR2X2 OR2X2_74 ( .A(core__abc_21302_new_n4176_), .B(core__abc_21302_new_n4173_), .Y(core__abc_21302_new_n4177_));
OR2X2 OR2X2_75 ( .A(core__abc_21302_new_n4208_), .B(core__abc_21302_new_n3482_), .Y(core__abc_21302_new_n4210_));
OR2X2 OR2X2_76 ( .A(core__abc_21302_new_n4235_), .B(core__abc_21302_new_n4274_), .Y(core__abc_21302_new_n4281_));
OR2X2 OR2X2_77 ( .A(core__abc_21302_new_n4300_), .B(core__abc_21302_new_n4309_), .Y(core__abc_21302_new_n4310_));
OR2X2 OR2X2_78 ( .A(core__abc_21302_new_n4300_), .B(core__abc_21302_new_n4313_), .Y(core__abc_21302_new_n4314_));
OR2X2 OR2X2_79 ( .A(core__abc_21302_new_n4330_), .B(core__abc_21302_new_n4342_), .Y(core__abc_21302_new_n4350_));
OR2X2 OR2X2_8 ( .A(_abc_19873_new_n896__bF_buf4), .B(_abc_19873_new_n1848_), .Y(_abc_19873_new_n2125_));
OR2X2 OR2X2_80 ( .A(core__abc_21302_new_n4424_), .B(core__abc_21302_new_n4432_), .Y(core__abc_21302_new_n4434_));
OR2X2 OR2X2_81 ( .A(core__abc_21302_new_n4434_), .B(core__abc_21302_new_n3778_), .Y(core__abc_21302_new_n4435_));
OR2X2 OR2X2_82 ( .A(core__abc_21302_new_n4493_), .B(core__abc_21302_new_n4497_), .Y(core__abc_21302_new_n4498_));
OR2X2 OR2X2_83 ( .A(core__abc_21302_new_n2991_), .B(core__abc_21302_new_n4504_), .Y(core__abc_21302_new_n4505_));
OR2X2 OR2X2_84 ( .A(core__abc_21302_new_n4700_), .B(core__abc_21302_new_n4647_), .Y(core__abc_21302_new_n4735_));
OR2X2 OR2X2_85 ( .A(core__abc_21302_new_n4872_), .B(core__abc_21302_new_n3638_), .Y(core__abc_21302_new_n4873_));
OR2X2 OR2X2_86 ( .A(core__abc_21302_new_n4946_), .B(core__abc_21302_new_n3299_), .Y(core__abc_21302_new_n4947_));
OR2X2 OR2X2_87 ( .A(core__abc_21302_new_n3191_), .B(core__abc_21302_new_n3193_), .Y(core__abc_21302_new_n4969_));
OR2X2 OR2X2_88 ( .A(core__abc_21302_new_n4971_), .B(core__abc_21302_new_n4969_), .Y(core__abc_21302_new_n4972_));
OR2X2 OR2X2_89 ( .A(core__abc_21302_new_n4990_), .B(core__abc_21302_new_n4992_), .Y(core__abc_21302_new_n4993_));
OR2X2 OR2X2_9 ( .A(_abc_19873_new_n960__bF_buf0), .B(_abc_19873_new_n1848_), .Y(_abc_19873_new_n2198_));
OR2X2 OR2X2_90 ( .A(core__abc_21302_new_n4975_), .B(core__abc_21302_new_n4993_), .Y(core__abc_21302_new_n4994_));
OR2X2 OR2X2_91 ( .A(core__abc_21302_new_n5001_), .B(core__abc_21302_new_n3018_), .Y(core__abc_21302_new_n5002_));
OR2X2 OR2X2_92 ( .A(core__abc_21302_new_n5030_), .B(core__abc_21302_new_n2806_), .Y(core__abc_21302_new_n5031_));
OR2X2 OR2X2_93 ( .A(core__abc_21302_new_n5035_), .B(core__abc_21302_new_n2773_), .Y(core__abc_21302_new_n5036_));
OR2X2 OR2X2_94 ( .A(core__abc_21302_new_n5037_), .B(core__abc_21302_new_n2744_), .Y(core__abc_21302_new_n5040_));
OR2X2 OR2X2_95 ( .A(core__abc_21302_new_n5041_), .B(core__abc_21302_new_n2692_), .Y(core__abc_21302_new_n5042_));
OR2X2 OR2X2_96 ( .A(core__abc_21302_new_n5012_), .B(core__abc_21302_new_n2939_), .Y(core__abc_21302_new_n5060_));
OR2X2 OR2X2_97 ( .A(core__abc_21302_new_n5074_), .B(core__abc_21302_new_n3925_), .Y(core__abc_21302_new_n5075_));
OR2X2 OR2X2_98 ( .A(core__abc_21302_new_n5122_), .B(core__abc_21302_new_n5120_), .Y(core__abc_21302_new_n5123_));
OR2X2 OR2X2_99 ( .A(core__abc_21302_new_n2739_), .B(core__abc_21302_new_n5136_), .Y(core__abc_21302_new_n5138_));
XNOR2X1 XNOR2X1_1 ( .A(core__abc_21302_new_n1132_), .B(core_compression_rounds_3_), .Y(core__abc_21302_new_n1133_));
XNOR2X1 XNOR2X1_10 ( .A(core__abc_21302_new_n1253_), .B(core__abc_21302_new_n1256_), .Y(core__abc_21302_new_n1257_));
XNOR2X1 XNOR2X1_100 ( .A(core__abc_21302_new_n3468_), .B(core__abc_21302_new_n3486_), .Y(core__abc_21302_new_n3487_));
XNOR2X1 XNOR2X1_101 ( .A(core__abc_21302_new_n3489_), .B(core__abc_21302_new_n1938_), .Y(core__abc_21302_new_n3490_));
XNOR2X1 XNOR2X1_102 ( .A(core_v3_reg_20_), .B(core_mi_20_), .Y(core__abc_21302_new_n3494_));
XNOR2X1 XNOR2X1_103 ( .A(core__abc_21302_new_n3521_), .B(core__abc_21302_new_n3520_), .Y(core__abc_21302_new_n3522_));
XNOR2X1 XNOR2X1_104 ( .A(core_v3_reg_21_), .B(core_mi_21_), .Y(core__abc_21302_new_n3526_));
XNOR2X1 XNOR2X1_105 ( .A(core_v3_reg_22_), .B(core_mi_22_), .Y(core__abc_21302_new_n3568_));
XNOR2X1 XNOR2X1_106 ( .A(core_v3_reg_23_), .B(core_mi_23_), .Y(core__abc_21302_new_n3599_));
XNOR2X1 XNOR2X1_107 ( .A(core__abc_21302_new_n3638_), .B(core_v3_reg_8_), .Y(core__abc_21302_new_n3639_));
XNOR2X1 XNOR2X1_108 ( .A(core__abc_21302_new_n3616_), .B(core__abc_21302_new_n3645_), .Y(core__abc_21302_new_n3646_));
XNOR2X1 XNOR2X1_109 ( .A(core__abc_21302_new_n3704_), .B(core__abc_21302_new_n1502_), .Y(core__abc_21302_new_n3708_));
XNOR2X1 XNOR2X1_11 ( .A(core__abc_21302_new_n1265_), .B(core__abc_21302_new_n1268_), .Y(core__abc_21302_new_n1269_));
XNOR2X1 XNOR2X1_110 ( .A(core__abc_21302_new_n3693_), .B(core__abc_21302_new_n3716_), .Y(core__abc_21302_new_n3717_));
XNOR2X1 XNOR2X1_111 ( .A(core_v3_reg_26_), .B(core_mi_26_), .Y(core__abc_21302_new_n3720_));
XNOR2X1 XNOR2X1_112 ( .A(core__abc_21302_new_n3773_), .B(core__abc_21302_new_n3768_), .Y(core__abc_21302_new_n3774_));
XNOR2X1 XNOR2X1_113 ( .A(core__abc_21302_new_n3776_), .B(core__abc_21302_new_n1526_), .Y(core__abc_21302_new_n3777_));
XNOR2X1 XNOR2X1_114 ( .A(core__abc_21302_new_n3777_), .B(core__abc_21302_new_n1339_), .Y(core__abc_21302_new_n3778_));
XNOR2X1 XNOR2X1_115 ( .A(core_v3_reg_28_), .B(core_mi_28_), .Y(core__abc_21302_new_n3786_));
XNOR2X1 XNOR2X1_116 ( .A(core_v3_reg_30_), .B(core_mi_30_), .Y(core__abc_21302_new_n3872_));
XNOR2X1 XNOR2X1_117 ( .A(core_v3_reg_31_), .B(core_mi_31_), .Y(core__abc_21302_new_n3903_));
XNOR2X1 XNOR2X1_118 ( .A(core__abc_21302_new_n3925_), .B(core_v3_reg_16_), .Y(core__abc_21302_new_n3926_));
XNOR2X1 XNOR2X1_119 ( .A(core_v3_reg_32_), .B(core_mi_32_), .Y(core__abc_21302_new_n3938_));
XNOR2X1 XNOR2X1_12 ( .A(core__abc_21302_new_n1275_), .B(core__abc_21302_new_n1278_), .Y(core__abc_21302_new_n1279_));
XNOR2X1 XNOR2X1_120 ( .A(core__abc_21302_new_n3962_), .B(core__abc_21302_new_n3108_), .Y(core__abc_21302_new_n3963_));
XNOR2X1 XNOR2X1_121 ( .A(core_v3_reg_33_), .B(core_mi_33_), .Y(core__abc_21302_new_n3965_));
XNOR2X1 XNOR2X1_122 ( .A(core__abc_21302_new_n3995_), .B(core__abc_21302_new_n3270_), .Y(core__abc_21302_new_n3996_));
XNOR2X1 XNOR2X1_123 ( .A(core_v3_reg_34_), .B(core_mi_34_), .Y(core__abc_21302_new_n3997_));
XNOR2X1 XNOR2X1_124 ( .A(core__abc_21302_new_n4004_), .B(core__abc_21302_new_n1243_), .Y(core__abc_21302_new_n4005_));
XNOR2X1 XNOR2X1_125 ( .A(core__abc_21302_new_n4045_), .B(core__abc_21302_new_n1620_), .Y(core__abc_21302_new_n4046_));
XNOR2X1 XNOR2X1_126 ( .A(core__abc_21302_new_n4045_), .B(core__abc_21302_new_n4048_), .Y(core__abc_21302_new_n4049_));
XNOR2X1 XNOR2X1_127 ( .A(core__abc_21302_new_n4040_), .B(core__abc_21302_new_n4055_), .Y(core__abc_21302_new_n4056_));
XNOR2X1 XNOR2X1_128 ( .A(core__abc_21302_new_n4056_), .B(core__abc_21302_new_n3240_), .Y(core__abc_21302_new_n4057_));
XNOR2X1 XNOR2X1_129 ( .A(core_v3_reg_36_), .B(core_mi_36_), .Y(core__abc_21302_new_n4058_));
XNOR2X1 XNOR2X1_13 ( .A(core__abc_21302_new_n1285_), .B(core__abc_21302_new_n1288_), .Y(core__abc_21302_new_n1289_));
XNOR2X1 XNOR2X1_130 ( .A(core__abc_21302_new_n4063_), .B(core__abc_21302_new_n1265_), .Y(core__abc_21302_new_n4064_));
XNOR2X1 XNOR2X1_131 ( .A(core_v3_reg_37_), .B(core_mi_37_), .Y(core__abc_21302_new_n4086_));
XNOR2X1 XNOR2X1_132 ( .A(core_v3_reg_38_), .B(core_mi_38_), .Y(core__abc_21302_new_n4121_));
XNOR2X1 XNOR2X1_133 ( .A(core__abc_21302_new_n4125_), .B(core__abc_21302_new_n1285_), .Y(core__abc_21302_new_n4126_));
XNOR2X1 XNOR2X1_134 ( .A(core__abc_21302_new_n4125_), .B(core__abc_21302_new_n2384_), .Y(core__abc_21302_new_n4135_));
XNOR2X1 XNOR2X1_135 ( .A(core_v3_reg_39_), .B(core_mi_39_), .Y(core__abc_21302_new_n4148_));
XNOR2X1 XNOR2X1_136 ( .A(core__abc_21302_new_n4174_), .B(core__abc_21302_new_n1664_), .Y(core__abc_21302_new_n4175_));
XNOR2X1 XNOR2X1_137 ( .A(core__abc_21302_new_n4175_), .B(core_v3_reg_24_), .Y(core__abc_21302_new_n4176_));
XNOR2X1 XNOR2X1_138 ( .A(core__abc_21302_new_n4184_), .B(core__abc_21302_new_n3432_), .Y(core__abc_21302_new_n4185_));
XNOR2X1 XNOR2X1_139 ( .A(core_v3_reg_40_), .B(core_mi_40_), .Y(core__abc_21302_new_n4186_));
XNOR2X1 XNOR2X1_14 ( .A(core__abc_21302_new_n1293_), .B(core__abc_21302_new_n1296_), .Y(core__abc_21302_new_n1297_));
XNOR2X1 XNOR2X1_140 ( .A(core__abc_21302_new_n4193_), .B(core__abc_21302_new_n1303_), .Y(core__abc_21302_new_n4194_));
XNOR2X1 XNOR2X1_141 ( .A(core__abc_21302_new_n4197_), .B(core__abc_21302_new_n1675_), .Y(core__abc_21302_new_n4198_));
XNOR2X1 XNOR2X1_142 ( .A(core__abc_21302_new_n4197_), .B(core__abc_21302_new_n4200_), .Y(core__abc_21302_new_n4201_));
XNOR2X1 XNOR2X1_143 ( .A(core_v3_reg_41_), .B(core_mi_41_), .Y(core__abc_21302_new_n4213_));
XNOR2X1 XNOR2X1_144 ( .A(core__abc_21302_new_n4218_), .B(core__abc_21302_new_n1314_), .Y(core__abc_21302_new_n4219_));
XNOR2X1 XNOR2X1_145 ( .A(core_v3_reg_42_), .B(core_mi_42_), .Y(core__abc_21302_new_n4244_));
XNOR2X1 XNOR2X1_146 ( .A(core__abc_21302_new_n4251_), .B(core__abc_21302_new_n1326_), .Y(core__abc_21302_new_n4257_));
XNOR2X1 XNOR2X1_147 ( .A(core__abc_21302_new_n4284_), .B(core__abc_21302_new_n1336_), .Y(core__abc_21302_new_n4285_));
XNOR2X1 XNOR2X1_148 ( .A(core__abc_21302_new_n4283_), .B(core__abc_21302_new_n4290_), .Y(core__abc_21302_new_n4291_));
XNOR2X1 XNOR2X1_149 ( .A(core__abc_21302_new_n4291_), .B(core__abc_21302_new_n3587_), .Y(core__abc_21302_new_n4292_));
XNOR2X1 XNOR2X1_15 ( .A(core__abc_21302_new_n1307_), .B(core__abc_21302_new_n1303_), .Y(core__abc_21302_new_n1308_));
XNOR2X1 XNOR2X1_150 ( .A(core_v3_reg_44_), .B(core_mi_44_), .Y(core__abc_21302_new_n4295_));
XNOR2X1 XNOR2X1_151 ( .A(core_v3_reg_45_), .B(core_mi_45_), .Y(core__abc_21302_new_n4318_));
XNOR2X1 XNOR2X1_152 ( .A(core__abc_21302_new_n4330_), .B(core__abc_21302_new_n4342_), .Y(core__abc_21302_new_n4343_));
XNOR2X1 XNOR2X1_153 ( .A(core_v3_reg_46_), .B(core_mi_46_), .Y(core__abc_21302_new_n4353_));
XNOR2X1 XNOR2X1_154 ( .A(core__abc_21302_new_n4362_), .B(core__abc_21302_new_n1372_), .Y(core__abc_21302_new_n4365_));
XNOR2X1 XNOR2X1_155 ( .A(core_v3_reg_47_), .B(core_mi_47_), .Y(core__abc_21302_new_n4380_));
XNOR2X1 XNOR2X1_156 ( .A(core__abc_21302_new_n2420_), .B(core__abc_21302_new_n4397_), .Y(core__abc_21302_new_n4398_));
XNOR2X1 XNOR2X1_157 ( .A(core__abc_21302_new_n4396_), .B(core__abc_21302_new_n4403_), .Y(core__abc_21302_new_n4404_));
XNOR2X1 XNOR2X1_158 ( .A(core__abc_21302_new_n4404_), .B(core__abc_21302_new_n3742_), .Y(core__abc_21302_new_n4405_));
XNOR2X1 XNOR2X1_159 ( .A(core_v3_reg_48_), .B(core_mi_48_), .Y(core__abc_21302_new_n4406_));
XNOR2X1 XNOR2X1_16 ( .A(core__abc_21302_new_n1319_), .B(core__abc_21302_new_n1314_), .Y(core__abc_21302_new_n1320_));
XNOR2X1 XNOR2X1_160 ( .A(core__abc_21302_new_n4412_), .B(core__abc_21302_new_n1395_), .Y(core__abc_21302_new_n4413_));
XNOR2X1 XNOR2X1_161 ( .A(core_v3_reg_49_), .B(core_mi_49_), .Y(core__abc_21302_new_n4438_));
XNOR2X1 XNOR2X1_162 ( .A(core_v3_reg_50_), .B(core_mi_50_), .Y(core__abc_21302_new_n4465_));
XNOR2X1 XNOR2X1_163 ( .A(core_v3_reg_51_), .B(core_mi_51_), .Y(core__abc_21302_new_n4487_));
XNOR2X1 XNOR2X1_164 ( .A(core__abc_21302_new_n4499_), .B(core__abc_21302_new_n4507_), .Y(core__abc_21302_new_n4508_));
XNOR2X1 XNOR2X1_165 ( .A(core__abc_21302_new_n4508_), .B(core__abc_21302_new_n3894_), .Y(core__abc_21302_new_n4509_));
XNOR2X1 XNOR2X1_166 ( .A(core_v3_reg_52_), .B(core_mi_52_), .Y(core__abc_21302_new_n4510_));
XNOR2X1 XNOR2X1_167 ( .A(core_v3_reg_53_), .B(core_mi_53_), .Y(core__abc_21302_new_n4534_));
XNOR2X1 XNOR2X1_168 ( .A(core_v3_reg_54_), .B(core_mi_54_), .Y(core__abc_21302_new_n4559_));
XNOR2X1 XNOR2X1_169 ( .A(core_v3_reg_55_), .B(core_mi_55_), .Y(core__abc_21302_new_n4588_));
XNOR2X1 XNOR2X1_17 ( .A(core__abc_21302_new_n1331_), .B(core__abc_21302_new_n1326_), .Y(core__abc_21302_new_n1332_));
XNOR2X1 XNOR2X1_170 ( .A(core__abc_21302_new_n3167_), .B(core__abc_21302_new_n4608_), .Y(core__abc_21302_new_n4609_));
XNOR2X1 XNOR2X1_171 ( .A(core__abc_21302_new_n4603_), .B(core__abc_21302_new_n4609_), .Y(core__abc_21302_new_n4610_));
XNOR2X1 XNOR2X1_172 ( .A(core__abc_21302_new_n4610_), .B(core__abc_21302_new_n4014_), .Y(core__abc_21302_new_n4611_));
XNOR2X1 XNOR2X1_173 ( .A(core_v3_reg_56_), .B(core_mi_56_), .Y(core__abc_21302_new_n4612_));
XNOR2X1 XNOR2X1_174 ( .A(core__abc_21302_new_n4623_), .B(core__abc_21302_new_n1485_), .Y(core__abc_21302_new_n4624_));
XNOR2X1 XNOR2X1_175 ( .A(core_v3_reg_57_), .B(core_mi_57_), .Y(core__abc_21302_new_n4637_));
XNOR2X1 XNOR2X1_176 ( .A(core__abc_21302_new_n4650_), .B(core__abc_21302_new_n1497_), .Y(core__abc_21302_new_n4651_));
XNOR2X1 XNOR2X1_177 ( .A(core_v3_reg_58_), .B(core_mi_58_), .Y(core__abc_21302_new_n4667_));
XNOR2X1 XNOR2X1_178 ( .A(core_v3_reg_60_), .B(core_mi_60_), .Y(core__abc_21302_new_n4726_));
XNOR2X1 XNOR2X1_179 ( .A(core_v3_reg_61_), .B(core_mi_61_), .Y(core__abc_21302_new_n4758_));
XNOR2X1 XNOR2X1_18 ( .A(core__abc_21302_new_n1388_), .B(core__abc_21302_new_n1384_), .Y(core__abc_21302_new_n1389_));
XNOR2X1 XNOR2X1_180 ( .A(core_v3_reg_62_), .B(core_mi_62_), .Y(core__abc_21302_new_n4791_));
XNOR2X1 XNOR2X1_181 ( .A(core__abc_21302_new_n3490_), .B(core_v3_reg_47_), .Y(core__abc_21302_new_n4804_));
XNOR2X1 XNOR2X1_182 ( .A(core__abc_21302_new_n4804_), .B(core__abc_21302_new_n4802_), .Y(core__abc_21302_new_n4808_));
XNOR2X1 XNOR2X1_183 ( .A(core__abc_21302_new_n4836_), .B(core__abc_21302_new_n4832_), .Y(core__abc_21302_new_n4837_));
XNOR2X1 XNOR2X1_184 ( .A(core__abc_21302_new_n4850_), .B(core__abc_21302_new_n3777_), .Y(core__abc_21302_new_n4851_));
XNOR2X1 XNOR2X1_185 ( .A(core__abc_21302_new_n4651_), .B(core_v1_reg_13_), .Y(core__abc_21302_new_n4862_));
XNOR2X1 XNOR2X1_186 ( .A(core__abc_21302_new_n4624_), .B(core__abc_21302_new_n4868_), .Y(core__abc_21302_new_n4869_));
XNOR2X1 XNOR2X1_187 ( .A(core__abc_21302_new_n4608_), .B(core__abc_21302_new_n4871_), .Y(core__abc_21302_new_n4872_));
XNOR2X1 XNOR2X1_188 ( .A(core__abc_21302_new_n4869_), .B(core__abc_21302_new_n3667_), .Y(core__abc_21302_new_n4890_));
XNOR2X1 XNOR2X1_189 ( .A(core__abc_21302_new_n4504_), .B(core__abc_21302_new_n4924_), .Y(core__abc_21302_new_n4925_));
XNOR2X1 XNOR2X1_19 ( .A(core__abc_21302_new_n1412_), .B(core__abc_21302_new_n1407_), .Y(core__abc_21302_new_n1413_));
XNOR2X1 XNOR2X1_190 ( .A(core__abc_21302_new_n4449_), .B(core_v1_reg_5_), .Y(core__abc_21302_new_n4930_));
XNOR2X1 XNOR2X1_191 ( .A(core__abc_21302_new_n4930_), .B(core__abc_21302_new_n4929_), .Y(core__abc_21302_new_n4931_));
XNOR2X1 XNOR2X1_192 ( .A(core__abc_21302_new_n4416_), .B(core_v1_reg_4_), .Y(core__abc_21302_new_n4944_));
XNOR2X1 XNOR2X1_193 ( .A(core__abc_21302_new_n4413_), .B(core_v1_reg_4_), .Y(core__abc_21302_new_n4945_));
XNOR2X1 XNOR2X1_194 ( .A(core__abc_21302_new_n4337_), .B(core__abc_21302_new_n4970_), .Y(core__abc_21302_new_n4971_));
XNOR2X1 XNOR2X1_195 ( .A(core__abc_21302_new_n4305_), .B(core_v1_reg_0_), .Y(core__abc_21302_new_n4977_));
XNOR2X1 XNOR2X1_196 ( .A(core__abc_21302_new_n4285_), .B(core__abc_21302_new_n4978_), .Y(core__abc_21302_new_n4979_));
XNOR2X1 XNOR2X1_197 ( .A(core__abc_21302_new_n4219_), .B(core__abc_21302_new_n1911_), .Y(core__abc_21302_new_n5001_));
XNOR2X1 XNOR2X1_198 ( .A(core__abc_21302_new_n4194_), .B(core_v1_reg_60_), .Y(core__abc_21302_new_n5010_));
XNOR2X1 XNOR2X1_199 ( .A(core__abc_21302_new_n4173_), .B(core_v1_reg_59_), .Y(core__abc_21302_new_n5012_));
XNOR2X1 XNOR2X1_2 ( .A(core_loop_ctr_reg_1_), .B(core_compression_rounds_1_), .Y(core__abc_21302_new_n1139_));
XNOR2X1 XNOR2X1_20 ( .A(core__abc_21302_new_n1424_), .B(core__abc_21302_new_n1419_), .Y(core__abc_21302_new_n1425_));
XNOR2X1 XNOR2X1_200 ( .A(core__abc_21302_new_n5010_), .B(core__abc_21302_new_n2970_), .Y(core__abc_21302_new_n5014_));
XNOR2X1 XNOR2X1_201 ( .A(core__abc_21302_new_n4099_), .B(core__abc_21302_new_n5024_), .Y(core__abc_21302_new_n5025_));
XNOR2X1 XNOR2X1_202 ( .A(core__abc_21302_new_n4064_), .B(core__abc_21302_new_n1845_), .Y(core__abc_21302_new_n5030_));
XNOR2X1 XNOR2X1_203 ( .A(core__abc_21302_new_n4043_), .B(core__abc_21302_new_n5034_), .Y(core__abc_21302_new_n5035_));
XNOR2X1 XNOR2X1_204 ( .A(core__abc_21302_new_n3978_), .B(core__abc_21302_new_n1807_), .Y(core__abc_21302_new_n5041_));
XNOR2X1 XNOR2X1_205 ( .A(core__abc_21302_new_n1211_), .B(core_v1_reg_51_), .Y(core__abc_21302_new_n5047_));
XNOR2X1 XNOR2X1_206 ( .A(core__abc_21302_new_n4944_), .B(core__abc_21302_new_n4943_), .Y(core__abc_21302_new_n5065_));
XNOR2X1 XNOR2X1_207 ( .A(core__abc_21302_new_n2509_), .B(core_v1_reg_19_), .Y(core__abc_21302_new_n5074_));
XNOR2X1 XNOR2X1_208 ( .A(core__abc_21302_new_n5073_), .B(core__abc_21302_new_n5078_), .Y(core__abc_21302_new_n5079_));
XNOR2X1 XNOR2X1_209 ( .A(core__abc_21302_new_n5088_), .B(core_v1_reg_20_), .Y(core__abc_21302_new_n5089_));
XNOR2X1 XNOR2X1_21 ( .A(core__abc_21302_new_n1436_), .B(core__abc_21302_new_n1431_), .Y(core__abc_21302_new_n1437_));
XNOR2X1 XNOR2X1_210 ( .A(core__abc_21302_new_n5096_), .B(core__abc_21302_new_n5090_), .Y(core__abc_21302_new_n5097_));
XNOR2X1 XNOR2X1_211 ( .A(core__abc_21302_new_n5134_), .B(core__abc_21302_new_n5144_), .Y(core__abc_21302_new_n5145_));
XNOR2X1 XNOR2X1_212 ( .A(core__abc_21302_new_n2777_), .B(core_v1_reg_23_), .Y(core__abc_21302_new_n5151_));
XNOR2X1 XNOR2X1_213 ( .A(core_v2_reg_4_), .B(core_long), .Y(core__abc_21302_new_n5169_));
XNOR2X1 XNOR2X1_214 ( .A(core__abc_21302_new_n2809_), .B(core_v1_reg_24_), .Y(core__abc_21302_new_n5176_));
XNOR2X1 XNOR2X1_215 ( .A(core__abc_21302_new_n2809_), .B(core__abc_21302_new_n2453_), .Y(core__abc_21302_new_n5178_));
XNOR2X1 XNOR2X1_216 ( .A(core__abc_21302_new_n2853_), .B(core_v1_reg_25_), .Y(core__abc_21302_new_n5188_));
XNOR2X1 XNOR2X1_217 ( .A(core__abc_21302_new_n2937_), .B(core_v1_reg_27_), .Y(core__abc_21302_new_n5237_));
XNOR2X1 XNOR2X1_218 ( .A(core__abc_21302_new_n5255_), .B(core__abc_21302_new_n5254_), .Y(core__abc_21302_new_n5256_));
XNOR2X1 XNOR2X1_219 ( .A(core__abc_21302_new_n3101_), .B(core__abc_21302_new_n5311_), .Y(core__abc_21302_new_n5312_));
XNOR2X1 XNOR2X1_22 ( .A(core__abc_21302_new_n1448_), .B(core__abc_21302_new_n1443_), .Y(core__abc_21302_new_n1449_));
XNOR2X1 XNOR2X1_220 ( .A(core__abc_21302_new_n5310_), .B(core__abc_21302_new_n5315_), .Y(core__abc_21302_new_n5316_));
XNOR2X1 XNOR2X1_221 ( .A(core__abc_21302_new_n3303_), .B(core_v1_reg_35_), .Y(core__abc_21302_new_n5404_));
XNOR2X1 XNOR2X1_222 ( .A(core__abc_21302_new_n5403_), .B(core__abc_21302_new_n5408_), .Y(core__abc_21302_new_n5409_));
XNOR2X1 XNOR2X1_223 ( .A(core__abc_21302_new_n3337_), .B(core__abc_21302_new_n5422_), .Y(core__abc_21302_new_n5423_));
XNOR2X1 XNOR2X1_224 ( .A(core__abc_21302_new_n5421_), .B(core__abc_21302_new_n5426_), .Y(core__abc_21302_new_n5427_));
XNOR2X1 XNOR2X1_225 ( .A(core__abc_21302_new_n5434_), .B(core__abc_21302_new_n1625_), .Y(core__abc_21302_new_n5435_));
XNOR2X1 XNOR2X1_226 ( .A(core__abc_21302_new_n3476_), .B(core__abc_21302_new_n5478_), .Y(core__abc_21302_new_n5479_));
XNOR2X1 XNOR2X1_227 ( .A(core__abc_21302_new_n5477_), .B(core__abc_21302_new_n5484_), .Y(core__abc_21302_new_n5485_));
XNOR2X1 XNOR2X1_228 ( .A(core__abc_21302_new_n3518_), .B(core_v1_reg_40_), .Y(core__abc_21302_new_n5493_));
XNOR2X1 XNOR2X1_229 ( .A(core__abc_21302_new_n5508_), .B(core__abc_21302_new_n5507_), .Y(core__abc_21302_new_n5509_));
XNOR2X1 XNOR2X1_23 ( .A(core__abc_21302_new_n1460_), .B(core__abc_21302_new_n1455_), .Y(core__abc_21302_new_n1461_));
XNOR2X1 XNOR2X1_230 ( .A(core__abc_21302_new_n5529_), .B(core__abc_21302_new_n5528_), .Y(core__abc_21302_new_n5530_));
XNOR2X1 XNOR2X1_231 ( .A(core__abc_21302_new_n5529_), .B(core_v1_reg_42_), .Y(core__abc_21302_new_n5532_));
XNOR2X1 XNOR2X1_232 ( .A(core__abc_21302_new_n3642_), .B(core_v1_reg_43_), .Y(core__abc_21302_new_n5554_));
XNOR2X1 XNOR2X1_233 ( .A(core__abc_21302_new_n3660_), .B(core_v1_reg_44_), .Y(core__abc_21302_new_n5572_));
XNOR2X1 XNOR2X1_234 ( .A(core__abc_21302_new_n3725_), .B(core_v1_reg_45_), .Y(core__abc_21302_new_n5584_));
XNOR2X1 XNOR2X1_235 ( .A(core__abc_21302_new_n5602_), .B(core__abc_21302_new_n5601_), .Y(core__abc_21302_new_n5603_));
XNOR2X1 XNOR2X1_236 ( .A(core__abc_21302_new_n3774_), .B(core_v1_reg_47_), .Y(core__abc_21302_new_n5625_));
XNOR2X1 XNOR2X1_237 ( .A(core__abc_21302_new_n3859_), .B(core__abc_21302_new_n5646_), .Y(core__abc_21302_new_n5647_));
XNOR2X1 XNOR2X1_238 ( .A(core__abc_21302_new_n5668_), .B(core_v1_reg_49_), .Y(core__abc_21302_new_n5669_));
XNOR2X1 XNOR2X1_239 ( .A(core__abc_21302_new_n5686_), .B(core__abc_21302_new_n5685_), .Y(core__abc_21302_new_n5687_));
XNOR2X1 XNOR2X1_24 ( .A(core_v2_reg_23_), .B(core_v3_reg_23_), .Y(core__abc_21302_new_n1468_));
XNOR2X1 XNOR2X1_240 ( .A(core__abc_21302_new_n3490_), .B(core__abc_21302_new_n5687_), .Y(core__abc_21302_new_n5688_));
XNOR2X1 XNOR2X1_241 ( .A(core__abc_21302_new_n5047_), .B(core__abc_21302_new_n1215_), .Y(core__abc_21302_new_n5700_));
XNOR2X1 XNOR2X1_242 ( .A(core__abc_21302_new_n5709_), .B(core__abc_21302_new_n5048_), .Y(core__abc_21302_new_n5710_));
XNOR2X1 XNOR2X1_243 ( .A(core__abc_21302_new_n5720_), .B(core__abc_21302_new_n5053_), .Y(core__abc_21302_new_n5721_));
XNOR2X1 XNOR2X1_244 ( .A(core__abc_21302_new_n5058_), .B(core__abc_21302_new_n5028_), .Y(core__abc_21302_new_n5745_));
XNOR2X1 XNOR2X1_245 ( .A(core__abc_21302_new_n5755_), .B(core__abc_21302_new_n5752_), .Y(core__abc_21302_new_n5756_));
XNOR2X1 XNOR2X1_246 ( .A(core__abc_21302_new_n5059_), .B(core__abc_21302_new_n5061_), .Y(core__abc_21302_new_n5764_));
XNOR2X1 XNOR2X1_247 ( .A(core__abc_21302_new_n5774_), .B(core__abc_21302_new_n5014_), .Y(core__abc_21302_new_n5775_));
XNOR2X1 XNOR2X1_248 ( .A(core__abc_21302_new_n5790_), .B(core__abc_21302_new_n5005_), .Y(core__abc_21302_new_n5791_));
XNOR2X1 XNOR2X1_249 ( .A(core__abc_21302_new_n5819_), .B(core__abc_21302_new_n4974_), .Y(core__abc_21302_new_n5820_));
XNOR2X1 XNOR2X1_25 ( .A(core__abc_21302_new_n1468_), .B(core__abc_21302_new_n1467_), .Y(core__abc_21302_new_n1469_));
XNOR2X1 XNOR2X1_250 ( .A(core__abc_21302_new_n5831_), .B(core__abc_21302_new_n5829_), .Y(core__abc_21302_new_n5832_));
XNOR2X1 XNOR2X1_251 ( .A(core__abc_21302_new_n5841_), .B(core__abc_21302_new_n5067_), .Y(core__abc_21302_new_n5842_));
XNOR2X1 XNOR2X1_252 ( .A(core__abc_21302_new_n5891_), .B(core__abc_21302_new_n5889_), .Y(core__abc_21302_new_n5892_));
XNOR2X1 XNOR2X1_253 ( .A(core__abc_21302_new_n5930_), .B(core__abc_21302_new_n4890_), .Y(core__abc_21302_new_n5931_));
XNOR2X1 XNOR2X1_254 ( .A(core__abc_21302_new_n5946_), .B(core__abc_21302_new_n4861_), .Y(core__abc_21302_new_n5947_));
XNOR2X1 XNOR2X1_255 ( .A(core_key_66_), .B(core_long), .Y(core__abc_21302_new_n6017_));
XNOR2X1 XNOR2X1_256 ( .A(core_key_69_), .B(core_long), .Y(core__abc_21302_new_n6041_));
XNOR2X1 XNOR2X1_257 ( .A(core__abc_21302_new_n5493_), .B(core__abc_21302_new_n5745_), .Y(core__abc_21302_new_n6049_));
XNOR2X1 XNOR2X1_258 ( .A(core_key_71_), .B(core_long), .Y(core__abc_21302_new_n6057_));
XNOR2X1 XNOR2X1_26 ( .A(core__abc_21302_new_n1502_), .B(core__abc_21302_new_n1497_), .Y(core__abc_21302_new_n1503_));
XNOR2X1 XNOR2X1_27 ( .A(core__abc_21302_new_n1514_), .B(core__abc_21302_new_n1509_), .Y(core__abc_21302_new_n1515_));
XNOR2X1 XNOR2X1_28 ( .A(core__abc_21302_new_n1526_), .B(core__abc_21302_new_n1521_), .Y(core__abc_21302_new_n1527_));
XNOR2X1 XNOR2X1_29 ( .A(core__abc_21302_new_n1534_), .B(core__abc_21302_new_n1539_), .Y(core__abc_21302_new_n1540_));
XNOR2X1 XNOR2X1_3 ( .A(core__abc_21302_new_n1142_), .B(core_loop_ctr_reg_2_), .Y(core__abc_21302_new_n1143_));
XNOR2X1 XNOR2X1_30 ( .A(core__abc_21302_new_n1551_), .B(core__abc_21302_new_n1546_), .Y(core__abc_21302_new_n1552_));
XNOR2X1 XNOR2X1_31 ( .A(core_v2_reg_31_), .B(core_v3_reg_31_), .Y(core__abc_21302_new_n1559_));
XNOR2X1 XNOR2X1_32 ( .A(core__abc_21302_new_n1559_), .B(core__abc_21302_new_n1558_), .Y(core__abc_21302_new_n1560_));
XNOR2X1 XNOR2X1_33 ( .A(core__abc_21302_new_n1571_), .B(core__abc_21302_new_n1567_), .Y(core__abc_21302_new_n1572_));
XNOR2X1 XNOR2X1_34 ( .A(core__abc_21302_new_n1620_), .B(core__abc_21302_new_n1616_), .Y(core__abc_21302_new_n1621_));
XNOR2X1 XNOR2X1_35 ( .A(core_v1_reg_38_), .B(core_v0_reg_38_), .Y(core__abc_21302_new_n1638_));
XNOR2X1 XNOR2X1_36 ( .A(core__abc_21302_new_n1664_), .B(core__abc_21302_new_n1660_), .Y(core__abc_21302_new_n1665_));
XNOR2X1 XNOR2X1_37 ( .A(core__abc_21302_new_n1675_), .B(core__abc_21302_new_n1671_), .Y(core__abc_21302_new_n1676_));
XNOR2X1 XNOR2X1_38 ( .A(core__abc_21302_new_n1720_), .B(core__abc_21302_new_n1716_), .Y(core__abc_21302_new_n1721_));
XNOR2X1 XNOR2X1_39 ( .A(core__abc_21302_new_n1732_), .B(core__abc_21302_new_n1728_), .Y(core__abc_21302_new_n1733_));
XNOR2X1 XNOR2X1_4 ( .A(core__abc_21302_new_n1162_), .B(core_final_rounds_3_), .Y(core__abc_21302_new_n1163_));
XNOR2X1 XNOR2X1_40 ( .A(core__abc_21302_new_n1743_), .B(core__abc_21302_new_n1739_), .Y(core__abc_21302_new_n1744_));
XNOR2X1 XNOR2X1_41 ( .A(core__abc_21302_new_n1766_), .B(core__abc_21302_new_n1761_), .Y(core__abc_21302_new_n1767_));
XNOR2X1 XNOR2X1_42 ( .A(core__abc_21302_new_n1811_), .B(core__abc_21302_new_n1814_), .Y(core__abc_21302_new_n1815_));
XNOR2X1 XNOR2X1_43 ( .A(core_v1_reg_63_), .B(core_v0_reg_63_), .Y(core__abc_21302_new_n1937_));
XNOR2X1 XNOR2X1_44 ( .A(core__abc_21302_new_n1938_), .B(core__abc_21302_new_n1937_), .Y(core__abc_21302_new_n1939_));
XNOR2X1 XNOR2X1_45 ( .A(core__abc_21302_new_n1215_), .B(core_v3_reg_48_), .Y(core__abc_21302_new_n2507_));
XNOR2X1 XNOR2X1_46 ( .A(core_v3_reg_0_), .B(core_mi_0_), .Y(core__abc_21302_new_n2642_));
XNOR2X1 XNOR2X1_47 ( .A(core__abc_21302_new_n1227_), .B(core__abc_21302_new_n1214_), .Y(core__abc_21302_new_n2651_));
XNOR2X1 XNOR2X1_48 ( .A(core__abc_21302_new_n2651_), .B(core__abc_21302_new_n1764_), .Y(core__abc_21302_new_n2652_));
XNOR2X1 XNOR2X1_49 ( .A(core__abc_21302_new_n2657_), .B(core__abc_21302_new_n2511_), .Y(core__abc_21302_new_n2658_));
XNOR2X1 XNOR2X1_5 ( .A(core__abc_21302_new_n1163_), .B(core_loop_ctr_reg_3_), .Y(core__abc_21302_new_n1164_));
XNOR2X1 XNOR2X1_50 ( .A(core_v3_reg_1_), .B(core_mi_1_), .Y(core__abc_21302_new_n2676_));
XNOR2X1 XNOR2X1_51 ( .A(core__abc_21302_new_n2699_), .B(core__abc_21302_new_n2681_), .Y(core__abc_21302_new_n2700_));
XNOR2X1 XNOR2X1_52 ( .A(core__abc_21302_new_n2704_), .B(core__abc_21302_new_n2701_), .Y(core__abc_21302_new_n2705_));
XNOR2X1 XNOR2X1_53 ( .A(core__abc_21302_new_n2704_), .B(core__abc_21302_new_n1720_), .Y(core__abc_21302_new_n2707_));
XNOR2X1 XNOR2X1_54 ( .A(core__abc_21302_new_n2744_), .B(core__abc_21302_new_n2740_), .Y(core__abc_21302_new_n2745_));
XNOR2X1 XNOR2X1_55 ( .A(core__abc_21302_new_n2750_), .B(core__abc_21302_new_n2734_), .Y(core__abc_21302_new_n2751_));
XNOR2X1 XNOR2X1_56 ( .A(core__abc_21302_new_n2773_), .B(core_v3_reg_52_), .Y(core__abc_21302_new_n2774_));
XNOR2X1 XNOR2X1_57 ( .A(core__abc_21302_new_n2805_), .B(core__abc_21302_new_n1268_), .Y(core__abc_21302_new_n2806_));
XNOR2X1 XNOR2X1_58 ( .A(core__abc_21302_new_n2806_), .B(core__abc_21302_new_n2804_), .Y(core__abc_21302_new_n2807_));
XNOR2X1 XNOR2X1_59 ( .A(core__abc_21302_new_n2799_), .B(core__abc_21302_new_n2812_), .Y(core__abc_21302_new_n2813_));
XNOR2X1 XNOR2X1_6 ( .A(core__abc_21302_new_n1167_), .B(core_loop_ctr_reg_2_), .Y(core__abc_21302_new_n1168_));
XNOR2X1 XNOR2X1_60 ( .A(core__abc_21302_new_n2829_), .B(core_v3_reg_32_), .Y(core__abc_21302_new_n2830_));
XNOR2X1 XNOR2X1_61 ( .A(core__abc_21302_new_n2850_), .B(core__abc_21302_new_n1824_), .Y(core__abc_21302_new_n2851_));
XNOR2X1 XNOR2X1_62 ( .A(core__abc_21302_new_n2862_), .B(core__abc_21302_new_n2857_), .Y(core__abc_21302_new_n2863_));
XNOR2X1 XNOR2X1_63 ( .A(core__abc_21302_new_n2880_), .B(core__abc_21302_new_n1649_), .Y(core__abc_21302_new_n2881_));
XNOR2X1 XNOR2X1_64 ( .A(core__abc_21302_new_n2885_), .B(core__abc_21302_new_n1837_), .Y(core__abc_21302_new_n2886_));
XNOR2X1 XNOR2X1_65 ( .A(core__abc_21302_new_n2880_), .B(core__abc_21302_new_n2889_), .Y(core__abc_21302_new_n2890_));
XNOR2X1 XNOR2X1_66 ( .A(core_v3_reg_7_), .B(core_mi_7_), .Y(core__abc_21302_new_n2909_));
XNOR2X1 XNOR2X1_67 ( .A(core__abc_21302_new_n2526_), .B(core__abc_21302_new_n2938_), .Y(core__abc_21302_new_n2939_));
XNOR2X1 XNOR2X1_68 ( .A(core__abc_21302_new_n2939_), .B(core_v3_reg_56_), .Y(core__abc_21302_new_n2940_));
XNOR2X1 XNOR2X1_69 ( .A(core_v3_reg_8_), .B(core_mi_8_), .Y(core__abc_21302_new_n2959_));
XNOR2X1 XNOR2X1_7 ( .A(core_final_rounds_1_), .B(core_loop_ctr_reg_1_), .Y(core__abc_21302_new_n1172_));
XNOR2X1 XNOR2X1_70 ( .A(core__abc_21302_new_n2969_), .B(core__abc_21302_new_n1307_), .Y(core__abc_21302_new_n2970_));
XNOR2X1 XNOR2X1_71 ( .A(core__abc_21302_new_n2978_), .B(core__abc_21302_new_n2976_), .Y(core__abc_21302_new_n2979_));
XNOR2X1 XNOR2X1_72 ( .A(core__abc_21302_new_n2990_), .B(core__abc_21302_new_n2980_), .Y(core__abc_21302_new_n2991_));
XNOR2X1 XNOR2X1_73 ( .A(core_v3_reg_9_), .B(core_mi_9_), .Y(core__abc_21302_new_n2994_));
XNOR2X1 XNOR2X1_74 ( .A(core__abc_21302_new_n3017_), .B(core__abc_21302_new_n2534_), .Y(core__abc_21302_new_n3018_));
XNOR2X1 XNOR2X1_75 ( .A(core__abc_21302_new_n3018_), .B(core__abc_21302_new_n1877_), .Y(core__abc_21302_new_n3019_));
XNOR2X1 XNOR2X1_76 ( .A(core_v3_reg_10_), .B(core_mi_10_), .Y(core__abc_21302_new_n3037_));
XNOR2X1 XNOR2X1_77 ( .A(core__abc_21302_new_n3044_), .B(core__abc_21302_new_n3061_), .Y(core__abc_21302_new_n3062_));
XNOR2X1 XNOR2X1_78 ( .A(core_v3_reg_11_), .B(core_mi_11_), .Y(core__abc_21302_new_n3077_));
XNOR2X1 XNOR2X1_79 ( .A(core__abc_21302_new_n3107_), .B(core_v3_reg_60_), .Y(core__abc_21302_new_n3108_));
XNOR2X1 XNOR2X1_8 ( .A(core__abc_21302_new_n1234_), .B(core__abc_21302_new_n1237_), .Y(core__abc_21302_new_n1238_));
XNOR2X1 XNOR2X1_80 ( .A(core_v3_reg_12_), .B(core_mi_12_), .Y(core__abc_21302_new_n3124_));
XNOR2X1 XNOR2X1_81 ( .A(core_v3_reg_13_), .B(core_mi_13_), .Y(core__abc_21302_new_n3170_));
XNOR2X1 XNOR2X1_82 ( .A(core__abc_21302_new_n3176_), .B(core__abc_21302_new_n3204_), .Y(core__abc_21302_new_n3205_));
XNOR2X1 XNOR2X1_83 ( .A(core__abc_21302_new_n3206_), .B(core__abc_21302_new_n1865_), .Y(core__abc_21302_new_n3213_));
XNOR2X1 XNOR2X1_84 ( .A(core_v3_reg_14_), .B(core_mi_14_), .Y(core__abc_21302_new_n3218_));
XNOR2X1 XNOR2X1_85 ( .A(core_v3_reg_15_), .B(core_mi_15_), .Y(core__abc_21302_new_n3260_));
XNOR2X1 XNOR2X1_86 ( .A(core__abc_21302_new_n2548_), .B(core__abc_21302_new_n1388_), .Y(core__abc_21302_new_n3299_));
XNOR2X1 XNOR2X1_87 ( .A(core__abc_21302_new_n3299_), .B(core_v3_reg_0_), .Y(core__abc_21302_new_n3300_));
XNOR2X1 XNOR2X1_88 ( .A(core__abc_21302_new_n3310_), .B(core__abc_21302_new_n3322_), .Y(core__abc_21302_new_n3323_));
XNOR2X1 XNOR2X1_89 ( .A(core_v3_reg_16_), .B(core_mi_16_), .Y(core__abc_21302_new_n3324_));
XNOR2X1 XNOR2X1_9 ( .A(core__abc_21302_new_n1243_), .B(core__abc_21302_new_n1246_), .Y(core__abc_21302_new_n1247_));
XNOR2X1 XNOR2X1_90 ( .A(core__abc_21302_new_n3339_), .B(core__abc_21302_new_n2563_), .Y(core__abc_21302_new_n3340_));
XNOR2X1 XNOR2X1_91 ( .A(core__abc_21302_new_n3353_), .B(core__abc_21302_new_n3357_), .Y(core__abc_21302_new_n3358_));
XNOR2X1 XNOR2X1_92 ( .A(core_v3_reg_17_), .B(core_mi_17_), .Y(core__abc_21302_new_n3363_));
XNOR2X1 XNOR2X1_93 ( .A(core__abc_21302_new_n3386_), .B(core__abc_21302_new_n2560_), .Y(core__abc_21302_new_n3387_));
XNOR2X1 XNOR2X1_94 ( .A(core__abc_21302_new_n3387_), .B(core__abc_21302_new_n2742_), .Y(core__abc_21302_new_n3388_));
XNOR2X1 XNOR2X1_95 ( .A(core__abc_21302_new_n3387_), .B(core_v3_reg_2_), .Y(core__abc_21302_new_n3392_));
XNOR2X1 XNOR2X1_96 ( .A(core__abc_21302_new_n3376_), .B(core__abc_21302_new_n3394_), .Y(core__abc_21302_new_n3395_));
XNOR2X1 XNOR2X1_97 ( .A(core_v3_reg_18_), .B(core_mi_18_), .Y(core__abc_21302_new_n3410_));
XNOR2X1 XNOR2X1_98 ( .A(core__abc_21302_new_n3475_), .B(core__abc_21302_new_n1797_), .Y(core__abc_21302_new_n3476_));
XNOR2X1 XNOR2X1_99 ( .A(core__abc_21302_new_n3481_), .B(core_v3_reg_4_), .Y(core__abc_21302_new_n3482_));
XOR2X1 XOR2X1_1 ( .A(core__abc_21302_new_n1130_), .B(core_compression_rounds_2_), .Y(core__abc_21302_new_n1142_));
XOR2X1 XOR2X1_10 ( .A(core__abc_21302_new_n1395_), .B(core__abc_21302_new_n1400_), .Y(core__abc_21302_new_n1401_));
XOR2X1 XOR2X1_100 ( .A(core_v0_reg_0_), .B(core_mi_reg_0_), .Y(core__abc_21302_new_n6452_));
XOR2X1 XOR2X1_101 ( .A(core_v0_reg_1_), .B(core_mi_reg_1_), .Y(core__abc_21302_new_n6458_));
XOR2X1 XOR2X1_102 ( .A(core_v0_reg_2_), .B(core_mi_reg_2_), .Y(core__abc_21302_new_n6466_));
XOR2X1 XOR2X1_103 ( .A(core_v0_reg_3_), .B(core_mi_reg_3_), .Y(core__abc_21302_new_n6473_));
XOR2X1 XOR2X1_104 ( .A(core_v0_reg_4_), .B(core_mi_reg_4_), .Y(core__abc_21302_new_n6479_));
XOR2X1 XOR2X1_105 ( .A(core_v0_reg_5_), .B(core_mi_reg_5_), .Y(core__abc_21302_new_n6486_));
XOR2X1 XOR2X1_106 ( .A(core_v0_reg_6_), .B(core_mi_reg_6_), .Y(core__abc_21302_new_n6493_));
XOR2X1 XOR2X1_107 ( .A(core_v0_reg_7_), .B(core_mi_reg_7_), .Y(core__abc_21302_new_n6500_));
XOR2X1 XOR2X1_108 ( .A(core_v0_reg_8_), .B(core_mi_reg_8_), .Y(core__abc_21302_new_n6507_));
XOR2X1 XOR2X1_109 ( .A(core_v0_reg_9_), .B(core_mi_reg_9_), .Y(core__abc_21302_new_n6515_));
XOR2X1 XOR2X1_11 ( .A(core__abc_21302_new_n1480_), .B(core__abc_21302_new_n1475_), .Y(core__abc_21302_new_n1481_));
XOR2X1 XOR2X1_110 ( .A(core_v0_reg_10_), .B(core_mi_reg_10_), .Y(core__abc_21302_new_n6522_));
XOR2X1 XOR2X1_111 ( .A(core_v0_reg_11_), .B(core_mi_reg_11_), .Y(core__abc_21302_new_n6529_));
XOR2X1 XOR2X1_112 ( .A(core_v0_reg_12_), .B(core_mi_reg_12_), .Y(core__abc_21302_new_n6537_));
XOR2X1 XOR2X1_113 ( .A(core_v0_reg_13_), .B(core_mi_reg_13_), .Y(core__abc_21302_new_n6544_));
XOR2X1 XOR2X1_114 ( .A(core_v0_reg_14_), .B(core_mi_reg_14_), .Y(core__abc_21302_new_n6551_));
XOR2X1 XOR2X1_115 ( .A(core_v0_reg_15_), .B(core_mi_reg_15_), .Y(core__abc_21302_new_n6558_));
XOR2X1 XOR2X1_116 ( .A(core_v0_reg_16_), .B(core_mi_reg_16_), .Y(core__abc_21302_new_n6565_));
XOR2X1 XOR2X1_117 ( .A(core_v0_reg_17_), .B(core_mi_reg_17_), .Y(core__abc_21302_new_n6572_));
XOR2X1 XOR2X1_118 ( .A(core_v0_reg_18_), .B(core_mi_reg_18_), .Y(core__abc_21302_new_n6580_));
XOR2X1 XOR2X1_119 ( .A(core_v0_reg_19_), .B(core_mi_reg_19_), .Y(core__abc_21302_new_n6587_));
XOR2X1 XOR2X1_12 ( .A(core_v1_reg_25_), .B(core_v0_reg_25_), .Y(core__abc_21302_new_n1485_));
XOR2X1 XOR2X1_120 ( .A(core_v0_reg_20_), .B(core_mi_reg_20_), .Y(core__abc_21302_new_n6594_));
XOR2X1 XOR2X1_121 ( .A(core_v0_reg_21_), .B(core_mi_reg_21_), .Y(core__abc_21302_new_n6601_));
XOR2X1 XOR2X1_122 ( .A(core_v0_reg_22_), .B(core_mi_reg_22_), .Y(core__abc_21302_new_n6608_));
XOR2X1 XOR2X1_123 ( .A(core_v0_reg_23_), .B(core_mi_reg_23_), .Y(core__abc_21302_new_n6615_));
XOR2X1 XOR2X1_124 ( .A(core_v0_reg_24_), .B(core_mi_reg_24_), .Y(core__abc_21302_new_n6621_));
XOR2X1 XOR2X1_125 ( .A(core_v0_reg_25_), .B(core_mi_reg_25_), .Y(core__abc_21302_new_n6630_));
XOR2X1 XOR2X1_126 ( .A(core_v0_reg_26_), .B(core_mi_reg_26_), .Y(core__abc_21302_new_n6638_));
XOR2X1 XOR2X1_127 ( .A(core_v0_reg_27_), .B(core_mi_reg_27_), .Y(core__abc_21302_new_n6646_));
XOR2X1 XOR2X1_128 ( .A(core_v0_reg_28_), .B(core_mi_reg_28_), .Y(core__abc_21302_new_n6653_));
XOR2X1 XOR2X1_129 ( .A(core_v0_reg_29_), .B(core_mi_reg_29_), .Y(core__abc_21302_new_n6660_));
XOR2X1 XOR2X1_13 ( .A(core__abc_21302_new_n1490_), .B(core__abc_21302_new_n1485_), .Y(core__abc_21302_new_n1491_));
XOR2X1 XOR2X1_130 ( .A(core_v0_reg_30_), .B(core_mi_reg_30_), .Y(core__abc_21302_new_n6667_));
XOR2X1 XOR2X1_131 ( .A(core_v0_reg_31_), .B(core_mi_reg_31_), .Y(core__abc_21302_new_n6674_));
XOR2X1 XOR2X1_132 ( .A(core_v0_reg_32_), .B(core_mi_reg_32_), .Y(core__abc_21302_new_n6680_));
XOR2X1 XOR2X1_133 ( .A(core_v0_reg_33_), .B(core_mi_reg_33_), .Y(core__abc_21302_new_n6686_));
XOR2X1 XOR2X1_134 ( .A(core_v0_reg_34_), .B(core_mi_reg_34_), .Y(core__abc_21302_new_n6693_));
XOR2X1 XOR2X1_135 ( .A(core_v0_reg_35_), .B(core_mi_reg_35_), .Y(core__abc_21302_new_n6700_));
XOR2X1 XOR2X1_136 ( .A(core_v0_reg_36_), .B(core_mi_reg_36_), .Y(core__abc_21302_new_n6707_));
XOR2X1 XOR2X1_137 ( .A(core_v0_reg_37_), .B(core_mi_reg_37_), .Y(core__abc_21302_new_n6713_));
XOR2X1 XOR2X1_138 ( .A(core_v0_reg_38_), .B(core_mi_reg_38_), .Y(core__abc_21302_new_n6720_));
XOR2X1 XOR2X1_139 ( .A(core_v0_reg_39_), .B(core_mi_reg_39_), .Y(core__abc_21302_new_n6727_));
XOR2X1 XOR2X1_14 ( .A(core__abc_21302_new_n1580_), .B(core__abc_21302_new_n1583_), .Y(core__abc_21302_new_n1584_));
XOR2X1 XOR2X1_140 ( .A(core_v0_reg_40_), .B(core_mi_reg_40_), .Y(core__abc_21302_new_n6733_));
XOR2X1 XOR2X1_141 ( .A(core_v0_reg_41_), .B(core_mi_reg_41_), .Y(core__abc_21302_new_n6741_));
XOR2X1 XOR2X1_142 ( .A(core_v0_reg_42_), .B(core_mi_reg_42_), .Y(core__abc_21302_new_n6748_));
XOR2X1 XOR2X1_143 ( .A(core_v0_reg_43_), .B(core_mi_reg_43_), .Y(core__abc_21302_new_n6755_));
XOR2X1 XOR2X1_144 ( .A(core_v0_reg_44_), .B(core_mi_reg_44_), .Y(core__abc_21302_new_n6762_));
XOR2X1 XOR2X1_145 ( .A(core_v0_reg_45_), .B(core_mi_reg_45_), .Y(core__abc_21302_new_n6769_));
XOR2X1 XOR2X1_146 ( .A(core_v0_reg_46_), .B(core_mi_reg_46_), .Y(core__abc_21302_new_n6776_));
XOR2X1 XOR2X1_147 ( .A(core_v0_reg_47_), .B(core_mi_reg_47_), .Y(core__abc_21302_new_n6783_));
XOR2X1 XOR2X1_148 ( .A(core_v0_reg_48_), .B(core_mi_reg_48_), .Y(core__abc_21302_new_n6789_));
XOR2X1 XOR2X1_149 ( .A(core_v0_reg_49_), .B(core_mi_reg_49_), .Y(core__abc_21302_new_n6796_));
XOR2X1 XOR2X1_15 ( .A(core__abc_21302_new_n1592_), .B(core__abc_21302_new_n1597_), .Y(core__abc_21302_new_n1598_));
XOR2X1 XOR2X1_150 ( .A(core_v0_reg_50_), .B(core_mi_reg_50_), .Y(core__abc_21302_new_n6803_));
XOR2X1 XOR2X1_151 ( .A(core_v0_reg_51_), .B(core_mi_reg_51_), .Y(core__abc_21302_new_n6810_));
XOR2X1 XOR2X1_152 ( .A(core_v0_reg_52_), .B(core_mi_reg_52_), .Y(core__abc_21302_new_n6818_));
XOR2X1 XOR2X1_153 ( .A(core_v0_reg_53_), .B(core_mi_reg_53_), .Y(core__abc_21302_new_n6825_));
XOR2X1 XOR2X1_154 ( .A(core_v0_reg_54_), .B(core_mi_reg_54_), .Y(core__abc_21302_new_n6832_));
XOR2X1 XOR2X1_155 ( .A(core_v0_reg_55_), .B(core_mi_reg_55_), .Y(core__abc_21302_new_n6839_));
XOR2X1 XOR2X1_156 ( .A(core_v0_reg_56_), .B(core_mi_reg_56_), .Y(core__abc_21302_new_n6846_));
XOR2X1 XOR2X1_157 ( .A(core_v0_reg_57_), .B(core_mi_reg_57_), .Y(core__abc_21302_new_n6854_));
XOR2X1 XOR2X1_158 ( .A(core_v0_reg_58_), .B(core_mi_reg_58_), .Y(core__abc_21302_new_n6862_));
XOR2X1 XOR2X1_159 ( .A(core_v0_reg_59_), .B(core_mi_reg_59_), .Y(core__abc_21302_new_n6870_));
XOR2X1 XOR2X1_16 ( .A(core__abc_21302_new_n1604_), .B(core__abc_21302_new_n1609_), .Y(core__abc_21302_new_n1610_));
XOR2X1 XOR2X1_160 ( .A(core_v0_reg_60_), .B(core_mi_reg_60_), .Y(core__abc_21302_new_n6877_));
XOR2X1 XOR2X1_161 ( .A(core_v0_reg_61_), .B(core_mi_reg_61_), .Y(core__abc_21302_new_n6884_));
XOR2X1 XOR2X1_162 ( .A(core_v0_reg_62_), .B(core_mi_reg_62_), .Y(core__abc_21302_new_n6892_));
XOR2X1 XOR2X1_163 ( .A(core_v0_reg_63_), .B(core_mi_reg_63_), .Y(core__abc_21302_new_n6899_));
XOR2X1 XOR2X1_17 ( .A(core__abc_21302_new_n1633_), .B(core__abc_21302_new_n1629_), .Y(core__abc_21302_new_n1634_));
XOR2X1 XOR2X1_18 ( .A(core__abc_21302_new_n1642_), .B(core__abc_21302_new_n1638_), .Y(core__abc_21302_new_n1643_));
XOR2X1 XOR2X1_19 ( .A(core__abc_21302_new_n1653_), .B(core__abc_21302_new_n1649_), .Y(core__abc_21302_new_n1654_));
XOR2X1 XOR2X1_2 ( .A(core__abc_21302_new_n1211_), .B(core__abc_21302_new_n1215_), .Y(core__abc_21302_new_n1216_));
XOR2X1 XOR2X1_20 ( .A(core__abc_21302_new_n1686_), .B(core__abc_21302_new_n1682_), .Y(core__abc_21302_new_n1687_));
XOR2X1 XOR2X1_21 ( .A(core__abc_21302_new_n1697_), .B(core__abc_21302_new_n1693_), .Y(core__abc_21302_new_n1698_));
XOR2X1 XOR2X1_22 ( .A(core__abc_21302_new_n1705_), .B(core__abc_21302_new_n1709_), .Y(core__abc_21302_new_n1710_));
XOR2X1 XOR2X1_23 ( .A(core__abc_21302_new_n1756_), .B(core__abc_21302_new_n1751_), .Y(core__abc_21302_new_n1757_));
XOR2X1 XOR2X1_24 ( .A(core_v1_reg_49_), .B(core_v0_reg_49_), .Y(core__abc_21302_new_n1761_));
XOR2X1 XOR2X1_25 ( .A(core__abc_21302_new_n1773_), .B(core__abc_21302_new_n1777_), .Y(core__abc_21302_new_n1778_));
XOR2X1 XOR2X1_26 ( .A(core__abc_21302_new_n1785_), .B(core__abc_21302_new_n1788_), .Y(core__abc_21302_new_n1789_));
XOR2X1 XOR2X1_27 ( .A(core__abc_21302_new_n1797_), .B(core__abc_21302_new_n1802_), .Y(core__abc_21302_new_n1803_));
XOR2X1 XOR2X1_28 ( .A(core__abc_21302_new_n1826_), .B(core__abc_21302_new_n1821_), .Y(core__abc_21302_new_n1827_));
XOR2X1 XOR2X1_29 ( .A(core__abc_21302_new_n1839_), .B(core__abc_21302_new_n1834_), .Y(core__abc_21302_new_n1840_));
XOR2X1 XOR2X1_3 ( .A(core__abc_21302_new_n1223_), .B(core__abc_21302_new_n1227_), .Y(core__abc_21302_new_n1228_));
XOR2X1 XOR2X1_30 ( .A(core__abc_21302_new_n1848_), .B(core__abc_21302_new_n1853_), .Y(core__abc_21302_new_n1854_));
XOR2X1 XOR2X1_31 ( .A(core__abc_21302_new_n1861_), .B(core__abc_21302_new_n1865_), .Y(core__abc_21302_new_n1866_));
XOR2X1 XOR2X1_32 ( .A(core__abc_21302_new_n1874_), .B(core__abc_21302_new_n1879_), .Y(core__abc_21302_new_n1880_));
XOR2X1 XOR2X1_33 ( .A(core__abc_21302_new_n1887_), .B(core__abc_21302_new_n1891_), .Y(core__abc_21302_new_n1892_));
XOR2X1 XOR2X1_34 ( .A(core__abc_21302_new_n1900_), .B(core__abc_21302_new_n1905_), .Y(core__abc_21302_new_n1906_));
XOR2X1 XOR2X1_35 ( .A(core__abc_21302_new_n1914_), .B(core__abc_21302_new_n1919_), .Y(core__abc_21302_new_n1920_));
XOR2X1 XOR2X1_36 ( .A(core__abc_21302_new_n1932_), .B(core__abc_21302_new_n1927_), .Y(core__abc_21302_new_n1933_));
XOR2X1 XOR2X1_37 ( .A(core_v2_reg_63_), .B(core_v3_reg_63_), .Y(core__abc_21302_new_n1938_));
XOR2X1 XOR2X1_38 ( .A(core_v1_reg_4_), .B(core_v0_reg_4_), .Y(core__abc_21302_new_n2386_));
XOR2X1 XOR2X1_39 ( .A(core__abc_21302_new_n2692_), .B(core_v3_reg_50_), .Y(core__abc_21302_new_n2693_));
XOR2X1 XOR2X1_4 ( .A(core_v1_reg_8_), .B(core_v0_reg_8_), .Y(core__abc_21302_new_n1293_));
XOR2X1 XOR2X1_40 ( .A(core_v3_reg_2_), .B(core_mi_2_), .Y(core__abc_21302_new_n2713_));
XOR2X1 XOR2X1_41 ( .A(core__abc_21302_new_n2743_), .B(core__abc_21302_new_n1246_), .Y(core__abc_21302_new_n2744_));
XOR2X1 XOR2X1_42 ( .A(core_v3_reg_3_), .B(core_mi_3_), .Y(core__abc_21302_new_n2756_));
XOR2X1 XOR2X1_43 ( .A(core__abc_21302_new_n2780_), .B(core__abc_21302_new_n2779_), .Y(core__abc_21302_new_n2781_));
XOR2X1 XOR2X1_44 ( .A(core_v3_reg_4_), .B(core_mi_4_), .Y(core__abc_21302_new_n2792_));
XOR2X1 XOR2X1_45 ( .A(core_v3_reg_5_), .B(core_mi_5_), .Y(core__abc_21302_new_n2833_));
XOR2X1 XOR2X1_46 ( .A(core_v3_reg_6_), .B(core_mi_6_), .Y(core__abc_21302_new_n2874_));
XOR2X1 XOR2X1_47 ( .A(core__abc_21302_new_n2884_), .B(core__abc_21302_new_n1288_), .Y(core__abc_21302_new_n2885_));
XOR2X1 XOR2X1_48 ( .A(core__abc_21302_new_n2893_), .B(core__abc_21302_new_n2892_), .Y(core__abc_21302_new_n2894_));
XOR2X1 XOR2X1_49 ( .A(core__abc_21302_new_n2970_), .B(core_v3_reg_57_), .Y(core__abc_21302_new_n2971_));
XOR2X1 XOR2X1_5 ( .A(core_v1_reg_12_), .B(core_v0_reg_12_), .Y(core__abc_21302_new_n1336_));
XOR2X1 XOR2X1_50 ( .A(core__abc_21302_new_n3005_), .B(core__abc_21302_new_n3024_), .Y(core__abc_21302_new_n3025_));
XOR2X1 XOR2X1_51 ( .A(core__abc_21302_new_n3101_), .B(core__abc_21302_new_n3108_), .Y(core__abc_21302_new_n3109_));
XOR2X1 XOR2X1_52 ( .A(core__abc_21302_new_n3090_), .B(core__abc_21302_new_n3109_), .Y(core__abc_21302_new_n3110_));
XOR2X1 XOR2X1_53 ( .A(core__abc_21302_new_n3340_), .B(core_v3_reg_1_), .Y(core__abc_21302_new_n3341_));
XOR2X1 XOR2X1_54 ( .A(core__abc_21302_new_n3438_), .B(core__abc_21302_new_n3449_), .Y(core__abc_21302_new_n3450_));
XOR2X1 XOR2X1_55 ( .A(core_v3_reg_19_), .B(core_mi_19_), .Y(core__abc_21302_new_n3451_));
XOR2X1 XOR2X1_56 ( .A(core__abc_21302_new_n3490_), .B(core_v3_reg_47_), .Y(core__abc_21302_new_n3491_));
XOR2X1 XOR2X1_57 ( .A(core_v3_reg_24_), .B(core_mi_24_), .Y(core__abc_21302_new_n3649_));
XOR2X1 XOR2X1_58 ( .A(core__abc_21302_new_n3677_), .B(core__abc_21302_new_n3676_), .Y(core__abc_21302_new_n3678_));
XOR2X1 XOR2X1_59 ( .A(core_v3_reg_25_), .B(core_mi_25_), .Y(core__abc_21302_new_n3681_));
XOR2X1 XOR2X1_6 ( .A(core__abc_21302_new_n1341_), .B(core__abc_21302_new_n1336_), .Y(core__abc_21302_new_n1342_));
XOR2X1 XOR2X1_60 ( .A(core_v3_reg_27_), .B(core_mi_27_), .Y(core__abc_21302_new_n3754_));
XOR2X1 XOR2X1_61 ( .A(core__abc_21302_new_n3774_), .B(core__abc_21302_new_n3778_), .Y(core__abc_21302_new_n3779_));
XOR2X1 XOR2X1_62 ( .A(core__abc_21302_new_n3790_), .B(core__abc_21302_new_n3820_), .Y(core__abc_21302_new_n3821_));
XOR2X1 XOR2X1_63 ( .A(core_v3_reg_29_), .B(core_mi_29_), .Y(core__abc_21302_new_n3824_));
XOR2X1 XOR2X1_64 ( .A(core__abc_21302_new_n3944_), .B(core__abc_21302_new_n3961_), .Y(core__abc_21302_new_n3962_));
XOR2X1 XOR2X1_65 ( .A(core__abc_21302_new_n3975_), .B(core__abc_21302_new_n3994_), .Y(core__abc_21302_new_n3995_));
XOR2X1 XOR2X1_66 ( .A(core_v3_reg_35_), .B(core_mi_35_), .Y(core__abc_21302_new_n4024_));
XOR2X1 XOR2X1_67 ( .A(core__abc_21302_new_n4100_), .B(core__abc_21302_new_n1642_), .Y(core__abc_21302_new_n4105_));
XOR2X1 XOR2X1_68 ( .A(core__abc_21302_new_n2397_), .B(core__abc_21302_new_n1293_), .Y(core__abc_21302_new_n4173_));
XOR2X1 XOR2X1_69 ( .A(core__abc_21302_new_n4191_), .B(core__abc_21302_new_n4207_), .Y(core__abc_21302_new_n4208_));
XOR2X1 XOR2X1_7 ( .A(core__abc_21302_new_n1353_), .B(core__abc_21302_new_n1348_), .Y(core__abc_21302_new_n1354_));
XOR2X1 XOR2X1_70 ( .A(core__abc_21302_new_n4251_), .B(core__abc_21302_new_n1326_), .Y(core__abc_21302_new_n4252_));
XOR2X1 XOR2X1_71 ( .A(core_v3_reg_43_), .B(core_mi_43_), .Y(core__abc_21302_new_n4267_));
XOR2X1 XOR2X1_72 ( .A(core__abc_21302_new_n4304_), .B(core__abc_21302_new_n1348_), .Y(core__abc_21302_new_n4305_));
XOR2X1 XOR2X1_73 ( .A(core__abc_21302_new_n4362_), .B(core__abc_21302_new_n1372_), .Y(core__abc_21302_new_n4363_));
XOR2X1 XOR2X1_74 ( .A(core__abc_21302_new_n4412_), .B(core__abc_21302_new_n1395_), .Y(core__abc_21302_new_n4416_));
XOR2X1 XOR2X1_75 ( .A(core_v3_reg_59_), .B(core_mi_59_), .Y(core__abc_21302_new_n4691_));
XOR2X1 XOR2X1_76 ( .A(core_v3_reg_63_), .B(core_mi_63_), .Y(core__abc_21302_new_n4816_));
XOR2X1 XOR2X1_77 ( .A(core__abc_21302_new_n4925_), .B(core__abc_21302_new_n3481_), .Y(core__abc_21302_new_n4926_));
XOR2X1 XOR2X1_78 ( .A(core__abc_21302_new_n4398_), .B(core_v1_reg_3_), .Y(core__abc_21302_new_n4946_));
XOR2X1 XOR2X1_79 ( .A(core__abc_21302_new_n4305_), .B(core_v1_reg_0_), .Y(core__abc_21302_new_n4976_));
XOR2X1 XOR2X1_8 ( .A(core__abc_21302_new_n1365_), .B(core__abc_21302_new_n1360_), .Y(core__abc_21302_new_n1366_));
XOR2X1 XOR2X1_80 ( .A(core__abc_21302_new_n5025_), .B(core__abc_21302_new_n2850_), .Y(core__abc_21302_new_n5028_));
XOR2X1 XOR2X1_81 ( .A(core__abc_21302_new_n4005_), .B(core_v1_reg_54_), .Y(core__abc_21302_new_n5037_));
XOR2X1 XOR2X1_82 ( .A(core_v2_reg_0_), .B(core_long), .Y(core__abc_21302_new_n5081_));
XOR2X1 XOR2X1_83 ( .A(core__abc_21302_new_n5089_), .B(core__abc_21302_new_n3954_), .Y(core__abc_21302_new_n5090_));
XOR2X1 XOR2X1_84 ( .A(core__abc_21302_new_n5175_), .B(core__abc_21302_new_n5180_), .Y(core__abc_21302_new_n5181_));
XOR2X1 XOR2X1_85 ( .A(core__abc_21302_new_n5235_), .B(core__abc_21302_new_n5241_), .Y(core__abc_21302_new_n5242_));
XOR2X1 XOR2X1_86 ( .A(core__abc_21302_new_n3458_), .B(core_v1_reg_38_), .Y(core__abc_21302_new_n5455_));
XOR2X1 XOR2X1_87 ( .A(core__abc_21302_new_n5455_), .B(core__abc_21302_new_n2952_), .Y(core__abc_21302_new_n5456_));
XOR2X1 XOR2X1_88 ( .A(core__abc_21302_new_n5052_), .B(core__abc_21302_new_n5050_), .Y(core__abc_21302_new_n5714_));
XOR2X1 XOR2X1_89 ( .A(core__abc_21302_new_n5054_), .B(core__abc_21302_new_n5056_), .Y(core__abc_21302_new_n5729_));
XOR2X1 XOR2X1_9 ( .A(core__abc_21302_new_n1377_), .B(core__abc_21302_new_n1372_), .Y(core__abc_21302_new_n1378_));
XOR2X1 XOR2X1_90 ( .A(core__abc_21302_new_n5057_), .B(core__abc_21302_new_n5738_), .Y(core__abc_21302_new_n5739_));
XOR2X1 XOR2X1_91 ( .A(core__abc_21302_new_n5782_), .B(core__abc_21302_new_n5008_), .Y(core__abc_21302_new_n5783_));
XOR2X1 XOR2X1_92 ( .A(core__abc_21302_new_n5812_), .B(core__abc_21302_new_n4990_), .Y(core__abc_21302_new_n5813_));
XOR2X1 XOR2X1_93 ( .A(core__abc_21302_new_n5850_), .B(core__abc_21302_new_n5065_), .Y(core__abc_21302_new_n5851_));
XOR2X1 XOR2X1_94 ( .A(core__abc_21302_new_n5871_), .B(core__abc_21302_new_n4941_), .Y(core__abc_21302_new_n5872_));
XOR2X1 XOR2X1_95 ( .A(core__abc_21302_new_n5937_), .B(core__abc_21302_new_n4866_), .Y(core__abc_21302_new_n5938_));
XOR2X1 XOR2X1_96 ( .A(core__abc_21302_new_n5988_), .B(core__abc_21302_new_n5987_), .Y(core__abc_21302_new_n5989_));
XOR2X1 XOR2X1_97 ( .A(core_key_65_), .B(core_long), .Y(core__abc_21302_new_n6008_));
XOR2X1 XOR2X1_98 ( .A(core_key_67_), .B(core_long), .Y(core__abc_21302_new_n6026_));
XOR2X1 XOR2X1_99 ( .A(core_key_70_), .B(core_long), .Y(core__abc_21302_new_n6047_));


endmodule