module spi_axi_master(CEB, SCLK, DATA, RST, CLK, axi_awready, axi_wready, axi_bvalid, axi_arready, axi_rvalid, \axi_rdata[0] , \axi_rdata[1] , \axi_rdata[2] , \axi_rdata[3] , \axi_rdata[4] , \axi_rdata[5] , \axi_rdata[6] , \axi_rdata[7] , \axi_rdata[8] , \axi_rdata[9] , \axi_rdata[10] , \axi_rdata[11] , \axi_rdata[12] , \axi_rdata[13] , \axi_rdata[14] , \axi_rdata[15] , \axi_rdata[16] , \axi_rdata[17] , \axi_rdata[18] , \axi_rdata[19] , \axi_rdata[20] , \axi_rdata[21] , \axi_rdata[22] , \axi_rdata[23] , \axi_rdata[24] , \axi_rdata[25] , \axi_rdata[26] , \axi_rdata[27] , \axi_rdata[28] , \axi_rdata[29] , \axi_rdata[30] , \axi_rdata[31] , DOUT, PICORV_RST, axi_awvalid, \axi_awaddr[0] , \axi_awaddr[1] , \axi_awaddr[2] , \axi_awaddr[3] , \axi_awaddr[4] , \axi_awaddr[5] , \axi_awaddr[6] , \axi_awaddr[7] , \axi_awaddr[8] , \axi_awaddr[9] , \axi_awaddr[10] , \axi_awaddr[11] , \axi_awaddr[12] , \axi_awaddr[13] , \axi_awaddr[14] , \axi_awaddr[15] , \axi_awaddr[16] , \axi_awaddr[17] , \axi_awaddr[18] , \axi_awaddr[19] , \axi_awaddr[20] , \axi_awaddr[21] , \axi_awaddr[22] , \axi_awaddr[23] , \axi_awaddr[24] , \axi_awaddr[25] , \axi_awaddr[26] , \axi_awaddr[27] , \axi_awaddr[28] , \axi_awaddr[29] , \axi_awaddr[30] , \axi_awaddr[31] , \axi_awprot[0] , \axi_awprot[1] , \axi_awprot[2] , axi_wvalid, \axi_wdata[0] , \axi_wdata[1] , \axi_wdata[2] , \axi_wdata[3] , \axi_wdata[4] , \axi_wdata[5] , \axi_wdata[6] , \axi_wdata[7] , \axi_wdata[8] , \axi_wdata[9] , \axi_wdata[10] , \axi_wdata[11] , \axi_wdata[12] , \axi_wdata[13] , \axi_wdata[14] , \axi_wdata[15] , \axi_wdata[16] , \axi_wdata[17] , \axi_wdata[18] , \axi_wdata[19] , \axi_wdata[20] , \axi_wdata[21] , \axi_wdata[22] , \axi_wdata[23] , \axi_wdata[24] , \axi_wdata[25] , \axi_wdata[26] , \axi_wdata[27] , \axi_wdata[28] , \axi_wdata[29] , \axi_wdata[30] , \axi_wdata[31] , \axi_wstrb[0] , \axi_wstrb[1] , \axi_wstrb[2] , \axi_wstrb[3] , axi_bready, axi_arvalid, \axi_araddr[0] , \axi_araddr[1] , \axi_araddr[2] , \axi_araddr[3] , \axi_araddr[4] , \axi_araddr[5] , \axi_araddr[6] , \axi_araddr[7] , \axi_araddr[8] , \axi_araddr[9] , \axi_araddr[10] , \axi_araddr[11] , \axi_araddr[12] , \axi_araddr[13] , \axi_araddr[14] , \axi_araddr[15] , \axi_araddr[16] , \axi_araddr[17] , \axi_araddr[18] , \axi_araddr[19] , \axi_araddr[20] , \axi_araddr[21] , \axi_araddr[22] , \axi_araddr[23] , \axi_araddr[24] , \axi_araddr[25] , \axi_araddr[26] , \axi_araddr[27] , \axi_araddr[28] , \axi_araddr[29] , \axi_araddr[30] , \axi_araddr[31] , \axi_arprot[0] , \axi_arprot[1] , \axi_arprot[2] , axi_rready);

wire A_ADDR_0_; 
wire A_ADDR_10_; 
wire A_ADDR_11_; 
wire A_ADDR_12_; 
wire A_ADDR_13_; 
wire A_ADDR_14_; 
wire A_ADDR_15_; 
wire A_ADDR_16_; 
wire A_ADDR_17_; 
wire A_ADDR_18_; 
wire A_ADDR_19_; 
wire A_ADDR_1_; 
wire A_ADDR_20_; 
wire A_ADDR_21_; 
wire A_ADDR_22_; 
wire A_ADDR_23_; 
wire A_ADDR_24_; 
wire A_ADDR_25_; 
wire A_ADDR_26_; 
wire A_ADDR_27_; 
wire A_ADDR_28_; 
wire A_ADDR_29_; 
wire A_ADDR_2_; 
wire A_ADDR_30_; 
wire A_ADDR_31_; 
wire A_ADDR_3_; 
wire A_ADDR_4_; 
wire A_ADDR_5_; 
wire A_ADDR_6_; 
wire A_ADDR_7_; 
wire A_ADDR_8_; 
wire A_ADDR_9_; 
input CEB;
input CLK;
input DATA;
output DOUT;
output PICORV_RST;
wire PICORV_RST_SPI; 
input RST;
input SCLK;
wire WDATA_0_; 
wire WDATA_10_; 
wire WDATA_11_; 
wire WDATA_12_; 
wire WDATA_13_; 
wire WDATA_14_; 
wire WDATA_15_; 
wire WDATA_16_; 
wire WDATA_17_; 
wire WDATA_18_; 
wire WDATA_19_; 
wire WDATA_1_; 
wire WDATA_20_; 
wire WDATA_21_; 
wire WDATA_22_; 
wire WDATA_23_; 
wire WDATA_24_; 
wire WDATA_25_; 
wire WDATA_26_; 
wire WDATA_27_; 
wire WDATA_28_; 
wire WDATA_29_; 
wire WDATA_2_; 
wire WDATA_30_; 
wire WDATA_31_; 
wire WDATA_3_; 
wire WDATA_4_; 
wire WDATA_5_; 
wire WDATA_6_; 
wire WDATA_7_; 
wire WDATA_8_; 
wire WDATA_9_; 
wire _0A_ADDR_31_0__0_; 
wire _0A_ADDR_31_0__10_; 
wire _0A_ADDR_31_0__11_; 
wire _0A_ADDR_31_0__12_; 
wire _0A_ADDR_31_0__13_; 
wire _0A_ADDR_31_0__14_; 
wire _0A_ADDR_31_0__15_; 
wire _0A_ADDR_31_0__16_; 
wire _0A_ADDR_31_0__17_; 
wire _0A_ADDR_31_0__18_; 
wire _0A_ADDR_31_0__19_; 
wire _0A_ADDR_31_0__1_; 
wire _0A_ADDR_31_0__20_; 
wire _0A_ADDR_31_0__21_; 
wire _0A_ADDR_31_0__22_; 
wire _0A_ADDR_31_0__23_; 
wire _0A_ADDR_31_0__24_; 
wire _0A_ADDR_31_0__25_; 
wire _0A_ADDR_31_0__26_; 
wire _0A_ADDR_31_0__27_; 
wire _0A_ADDR_31_0__28_; 
wire _0A_ADDR_31_0__29_; 
wire _0A_ADDR_31_0__2_; 
wire _0A_ADDR_31_0__30_; 
wire _0A_ADDR_31_0__31_; 
wire _0A_ADDR_31_0__3_; 
wire _0A_ADDR_31_0__4_; 
wire _0A_ADDR_31_0__5_; 
wire _0A_ADDR_31_0__6_; 
wire _0A_ADDR_31_0__7_; 
wire _0A_ADDR_31_0__8_; 
wire _0A_ADDR_31_0__9_; 
wire _0PICORV_RST_SPI_0_0_; 
wire _0WDATA_31_0__0_; 
wire _0WDATA_31_0__10_; 
wire _0WDATA_31_0__11_; 
wire _0WDATA_31_0__12_; 
wire _0WDATA_31_0__13_; 
wire _0WDATA_31_0__14_; 
wire _0WDATA_31_0__15_; 
wire _0WDATA_31_0__16_; 
wire _0WDATA_31_0__17_; 
wire _0WDATA_31_0__18_; 
wire _0WDATA_31_0__19_; 
wire _0WDATA_31_0__1_; 
wire _0WDATA_31_0__20_; 
wire _0WDATA_31_0__21_; 
wire _0WDATA_31_0__22_; 
wire _0WDATA_31_0__23_; 
wire _0WDATA_31_0__24_; 
wire _0WDATA_31_0__25_; 
wire _0WDATA_31_0__26_; 
wire _0WDATA_31_0__27_; 
wire _0WDATA_31_0__28_; 
wire _0WDATA_31_0__29_; 
wire _0WDATA_31_0__2_; 
wire _0WDATA_31_0__30_; 
wire _0WDATA_31_0__31_; 
wire _0WDATA_31_0__3_; 
wire _0WDATA_31_0__4_; 
wire _0WDATA_31_0__5_; 
wire _0WDATA_31_0__6_; 
wire _0WDATA_31_0__7_; 
wire _0WDATA_31_0__8_; 
wire _0WDATA_31_0__9_; 
wire _0bus_cap_31_0__0_; 
wire _0bus_cap_31_0__10_; 
wire _0bus_cap_31_0__11_; 
wire _0bus_cap_31_0__12_; 
wire _0bus_cap_31_0__13_; 
wire _0bus_cap_31_0__14_; 
wire _0bus_cap_31_0__15_; 
wire _0bus_cap_31_0__16_; 
wire _0bus_cap_31_0__17_; 
wire _0bus_cap_31_0__18_; 
wire _0bus_cap_31_0__19_; 
wire _0bus_cap_31_0__1_; 
wire _0bus_cap_31_0__20_; 
wire _0bus_cap_31_0__21_; 
wire _0bus_cap_31_0__22_; 
wire _0bus_cap_31_0__23_; 
wire _0bus_cap_31_0__24_; 
wire _0bus_cap_31_0__25_; 
wire _0bus_cap_31_0__26_; 
wire _0bus_cap_31_0__27_; 
wire _0bus_cap_31_0__28_; 
wire _0bus_cap_31_0__29_; 
wire _0bus_cap_31_0__2_; 
wire _0bus_cap_31_0__30_; 
wire _0bus_cap_31_0__31_; 
wire _0bus_cap_31_0__3_; 
wire _0bus_cap_31_0__4_; 
wire _0bus_cap_31_0__5_; 
wire _0bus_cap_31_0__6_; 
wire _0bus_cap_31_0__7_; 
wire _0bus_cap_31_0__8_; 
wire _0bus_cap_31_0__9_; 
wire _0counter_65_0__0_; 
wire _0counter_65_0__10_; 
wire _0counter_65_0__11_; 
wire _0counter_65_0__12_; 
wire _0counter_65_0__13_; 
wire _0counter_65_0__14_; 
wire _0counter_65_0__15_; 
wire _0counter_65_0__16_; 
wire _0counter_65_0__17_; 
wire _0counter_65_0__18_; 
wire _0counter_65_0__19_; 
wire _0counter_65_0__1_; 
wire _0counter_65_0__20_; 
wire _0counter_65_0__21_; 
wire _0counter_65_0__22_; 
wire _0counter_65_0__23_; 
wire _0counter_65_0__24_; 
wire _0counter_65_0__25_; 
wire _0counter_65_0__26_; 
wire _0counter_65_0__27_; 
wire _0counter_65_0__28_; 
wire _0counter_65_0__29_; 
wire _0counter_65_0__2_; 
wire _0counter_65_0__30_; 
wire _0counter_65_0__31_; 
wire _0counter_65_0__32_; 
wire _0counter_65_0__33_; 
wire _0counter_65_0__34_; 
wire _0counter_65_0__35_; 
wire _0counter_65_0__36_; 
wire _0counter_65_0__37_; 
wire _0counter_65_0__38_; 
wire _0counter_65_0__39_; 
wire _0counter_65_0__3_; 
wire _0counter_65_0__40_; 
wire _0counter_65_0__41_; 
wire _0counter_65_0__42_; 
wire _0counter_65_0__43_; 
wire _0counter_65_0__44_; 
wire _0counter_65_0__45_; 
wire _0counter_65_0__46_; 
wire _0counter_65_0__47_; 
wire _0counter_65_0__48_; 
wire _0counter_65_0__49_; 
wire _0counter_65_0__4_; 
wire _0counter_65_0__50_; 
wire _0counter_65_0__51_; 
wire _0counter_65_0__52_; 
wire _0counter_65_0__53_; 
wire _0counter_65_0__54_; 
wire _0counter_65_0__55_; 
wire _0counter_65_0__56_; 
wire _0counter_65_0__57_; 
wire _0counter_65_0__58_; 
wire _0counter_65_0__59_; 
wire _0counter_65_0__5_; 
wire _0counter_65_0__60_; 
wire _0counter_65_0__61_; 
wire _0counter_65_0__62_; 
wire _0counter_65_0__63_; 
wire _0counter_65_0__64_; 
wire _0counter_65_0__65_; 
wire _0counter_65_0__6_; 
wire _0counter_65_0__7_; 
wire _0counter_65_0__8_; 
wire _0counter_65_0__9_; 
wire _0fini_spi_0_0_; 
wire _0rdata_31_0__0_; 
wire _0rdata_31_0__10_; 
wire _0rdata_31_0__11_; 
wire _0rdata_31_0__12_; 
wire _0rdata_31_0__13_; 
wire _0rdata_31_0__14_; 
wire _0rdata_31_0__15_; 
wire _0rdata_31_0__16_; 
wire _0rdata_31_0__17_; 
wire _0rdata_31_0__18_; 
wire _0rdata_31_0__19_; 
wire _0rdata_31_0__1_; 
wire _0rdata_31_0__20_; 
wire _0rdata_31_0__21_; 
wire _0rdata_31_0__22_; 
wire _0rdata_31_0__23_; 
wire _0rdata_31_0__24_; 
wire _0rdata_31_0__25_; 
wire _0rdata_31_0__26_; 
wire _0rdata_31_0__27_; 
wire _0rdata_31_0__28_; 
wire _0rdata_31_0__29_; 
wire _0rdata_31_0__2_; 
wire _0rdata_31_0__30_; 
wire _0rdata_31_0__31_; 
wire _0rdata_31_0__3_; 
wire _0rdata_31_0__4_; 
wire _0rdata_31_0__5_; 
wire _0rdata_31_0__6_; 
wire _0rdata_31_0__7_; 
wire _0rdata_31_0__8_; 
wire _0rdata_31_0__9_; 
wire _0re_0_0_; 
wire _0sft_reg_65_0__0_; 
wire _0sft_reg_65_0__10_; 
wire _0sft_reg_65_0__11_; 
wire _0sft_reg_65_0__12_; 
wire _0sft_reg_65_0__13_; 
wire _0sft_reg_65_0__14_; 
wire _0sft_reg_65_0__15_; 
wire _0sft_reg_65_0__16_; 
wire _0sft_reg_65_0__17_; 
wire _0sft_reg_65_0__18_; 
wire _0sft_reg_65_0__19_; 
wire _0sft_reg_65_0__1_; 
wire _0sft_reg_65_0__20_; 
wire _0sft_reg_65_0__21_; 
wire _0sft_reg_65_0__22_; 
wire _0sft_reg_65_0__23_; 
wire _0sft_reg_65_0__24_; 
wire _0sft_reg_65_0__25_; 
wire _0sft_reg_65_0__26_; 
wire _0sft_reg_65_0__27_; 
wire _0sft_reg_65_0__28_; 
wire _0sft_reg_65_0__29_; 
wire _0sft_reg_65_0__2_; 
wire _0sft_reg_65_0__30_; 
wire _0sft_reg_65_0__3_; 
wire _0sft_reg_65_0__4_; 
wire _0sft_reg_65_0__5_; 
wire _0sft_reg_65_0__6_; 
wire _0sft_reg_65_0__7_; 
wire _0sft_reg_65_0__8_; 
wire _0sft_reg_65_0__9_; 
wire _0we_0_0_; 
wire _abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_430; 
wire _abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_479; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_0_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_1_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_3_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_4_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_5_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_6_; 
wire _abc_2903_auto_fsm_map_cc_170_map_fsm_402_7_; 
wire _abc_4268_new_n1000_; 
wire _abc_4268_new_n1001_; 
wire _abc_4268_new_n1003_; 
wire _abc_4268_new_n1004_; 
wire _abc_4268_new_n1005_; 
wire _abc_4268_new_n1007_; 
wire _abc_4268_new_n1008_; 
wire _abc_4268_new_n1009_; 
wire _abc_4268_new_n1011_; 
wire _abc_4268_new_n1012_; 
wire _abc_4268_new_n1013_; 
wire _abc_4268_new_n1015_; 
wire _abc_4268_new_n1016_; 
wire _abc_4268_new_n1017_; 
wire _abc_4268_new_n1019_; 
wire _abc_4268_new_n1020_; 
wire _abc_4268_new_n1021_; 
wire _abc_4268_new_n1023_; 
wire _abc_4268_new_n1024_; 
wire _abc_4268_new_n1025_; 
wire _abc_4268_new_n1027_; 
wire _abc_4268_new_n1028_; 
wire _abc_4268_new_n1029_; 
wire _abc_4268_new_n1031_; 
wire _abc_4268_new_n1032_; 
wire _abc_4268_new_n1033_; 
wire _abc_4268_new_n1035_; 
wire _abc_4268_new_n1036_; 
wire _abc_4268_new_n1037_; 
wire _abc_4268_new_n1039_; 
wire _abc_4268_new_n1040_; 
wire _abc_4268_new_n1041_; 
wire _abc_4268_new_n1043_; 
wire _abc_4268_new_n1044_; 
wire _abc_4268_new_n1045_; 
wire _abc_4268_new_n1047_; 
wire _abc_4268_new_n1048_; 
wire _abc_4268_new_n1049_; 
wire _abc_4268_new_n1051_; 
wire _abc_4268_new_n1052_; 
wire _abc_4268_new_n1053_; 
wire _abc_4268_new_n1055_; 
wire _abc_4268_new_n1056_; 
wire _abc_4268_new_n1057_; 
wire _abc_4268_new_n1059_; 
wire _abc_4268_new_n1060_; 
wire _abc_4268_new_n1061_; 
wire _abc_4268_new_n1063_; 
wire _abc_4268_new_n1064_; 
wire _abc_4268_new_n1065_; 
wire _abc_4268_new_n1067_; 
wire _abc_4268_new_n1068_; 
wire _abc_4268_new_n1069_; 
wire _abc_4268_new_n1071_; 
wire _abc_4268_new_n1072_; 
wire _abc_4268_new_n1073_; 
wire _abc_4268_new_n1075_; 
wire _abc_4268_new_n1076_; 
wire _abc_4268_new_n1077_; 
wire _abc_4268_new_n1079_; 
wire _abc_4268_new_n1080_; 
wire _abc_4268_new_n1081_; 
wire _abc_4268_new_n1083_; 
wire _abc_4268_new_n1084_; 
wire _abc_4268_new_n1085_; 
wire _abc_4268_new_n1086_; 
wire _abc_4268_new_n1087_; 
wire _abc_4268_new_n1088_; 
wire _abc_4268_new_n1089_; 
wire _abc_4268_new_n1091_; 
wire _abc_4268_new_n1092_; 
wire _abc_4268_new_n1093_; 
wire _abc_4268_new_n1095_; 
wire _abc_4268_new_n1096_; 
wire _abc_4268_new_n1097_; 
wire _abc_4268_new_n1099_; 
wire _abc_4268_new_n1100_; 
wire _abc_4268_new_n1101_; 
wire _abc_4268_new_n1103_; 
wire _abc_4268_new_n1104_; 
wire _abc_4268_new_n1105_; 
wire _abc_4268_new_n1107_; 
wire _abc_4268_new_n1108_; 
wire _abc_4268_new_n1109_; 
wire _abc_4268_new_n1111_; 
wire _abc_4268_new_n1112_; 
wire _abc_4268_new_n1113_; 
wire _abc_4268_new_n1115_; 
wire _abc_4268_new_n1116_; 
wire _abc_4268_new_n1117_; 
wire _abc_4268_new_n1119_; 
wire _abc_4268_new_n1120_; 
wire _abc_4268_new_n1121_; 
wire _abc_4268_new_n1123_; 
wire _abc_4268_new_n1124_; 
wire _abc_4268_new_n1125_; 
wire _abc_4268_new_n1127_; 
wire _abc_4268_new_n1128_; 
wire _abc_4268_new_n1129_; 
wire _abc_4268_new_n1131_; 
wire _abc_4268_new_n1132_; 
wire _abc_4268_new_n1133_; 
wire _abc_4268_new_n1135_; 
wire _abc_4268_new_n1136_; 
wire _abc_4268_new_n1137_; 
wire _abc_4268_new_n1139_; 
wire _abc_4268_new_n1140_; 
wire _abc_4268_new_n1141_; 
wire _abc_4268_new_n1143_; 
wire _abc_4268_new_n1144_; 
wire _abc_4268_new_n1145_; 
wire _abc_4268_new_n1147_; 
wire _abc_4268_new_n1148_; 
wire _abc_4268_new_n1149_; 
wire _abc_4268_new_n1151_; 
wire _abc_4268_new_n1152_; 
wire _abc_4268_new_n1153_; 
wire _abc_4268_new_n1155_; 
wire _abc_4268_new_n1156_; 
wire _abc_4268_new_n1157_; 
wire _abc_4268_new_n1159_; 
wire _abc_4268_new_n1160_; 
wire _abc_4268_new_n1161_; 
wire _abc_4268_new_n1163_; 
wire _abc_4268_new_n1164_; 
wire _abc_4268_new_n1165_; 
wire _abc_4268_new_n1167_; 
wire _abc_4268_new_n1168_; 
wire _abc_4268_new_n1169_; 
wire _abc_4268_new_n1171_; 
wire _abc_4268_new_n1172_; 
wire _abc_4268_new_n1173_; 
wire _abc_4268_new_n1175_; 
wire _abc_4268_new_n1176_; 
wire _abc_4268_new_n1177_; 
wire _abc_4268_new_n1179_; 
wire _abc_4268_new_n1180_; 
wire _abc_4268_new_n1181_; 
wire _abc_4268_new_n1183_; 
wire _abc_4268_new_n1184_; 
wire _abc_4268_new_n1185_; 
wire _abc_4268_new_n1187_; 
wire _abc_4268_new_n1188_; 
wire _abc_4268_new_n1189_; 
wire _abc_4268_new_n1191_; 
wire _abc_4268_new_n1192_; 
wire _abc_4268_new_n1193_; 
wire _abc_4268_new_n1195_; 
wire _abc_4268_new_n1196_; 
wire _abc_4268_new_n1197_; 
wire _abc_4268_new_n1199_; 
wire _abc_4268_new_n1200_; 
wire _abc_4268_new_n1201_; 
wire _abc_4268_new_n1203_; 
wire _abc_4268_new_n1204_; 
wire _abc_4268_new_n1205_; 
wire _abc_4268_new_n1207_; 
wire _abc_4268_new_n1208_; 
wire _abc_4268_new_n1209_; 
wire _abc_4268_new_n1211_; 
wire _abc_4268_new_n1212_; 
wire _abc_4268_new_n1213_; 
wire _abc_4268_new_n1215_; 
wire _abc_4268_new_n1216_; 
wire _abc_4268_new_n1217_; 
wire _abc_4268_new_n1218_; 
wire _abc_4268_new_n1219_; 
wire _abc_4268_new_n1220_; 
wire _abc_4268_new_n1222_; 
wire _abc_4268_new_n1223_; 
wire _abc_4268_new_n1224_; 
wire _abc_4268_new_n1226_; 
wire _abc_4268_new_n1227_; 
wire _abc_4268_new_n1228_; 
wire _abc_4268_new_n1230_; 
wire _abc_4268_new_n1231_; 
wire _abc_4268_new_n1232_; 
wire _abc_4268_new_n1234_; 
wire _abc_4268_new_n1235_; 
wire _abc_4268_new_n1236_; 
wire _abc_4268_new_n1238_; 
wire _abc_4268_new_n1239_; 
wire _abc_4268_new_n1240_; 
wire _abc_4268_new_n1242_; 
wire _abc_4268_new_n1243_; 
wire _abc_4268_new_n1244_; 
wire _abc_4268_new_n1246_; 
wire _abc_4268_new_n1247_; 
wire _abc_4268_new_n1248_; 
wire _abc_4268_new_n1250_; 
wire _abc_4268_new_n1251_; 
wire _abc_4268_new_n1252_; 
wire _abc_4268_new_n1254_; 
wire _abc_4268_new_n1255_; 
wire _abc_4268_new_n1256_; 
wire _abc_4268_new_n1258_; 
wire _abc_4268_new_n1259_; 
wire _abc_4268_new_n1260_; 
wire _abc_4268_new_n1262_; 
wire _abc_4268_new_n1263_; 
wire _abc_4268_new_n1264_; 
wire _abc_4268_new_n1266_; 
wire _abc_4268_new_n1267_; 
wire _abc_4268_new_n1268_; 
wire _abc_4268_new_n1270_; 
wire _abc_4268_new_n1271_; 
wire _abc_4268_new_n1272_; 
wire _abc_4268_new_n1274_; 
wire _abc_4268_new_n1275_; 
wire _abc_4268_new_n1276_; 
wire _abc_4268_new_n1278_; 
wire _abc_4268_new_n1279_; 
wire _abc_4268_new_n1280_; 
wire _abc_4268_new_n1282_; 
wire _abc_4268_new_n1283_; 
wire _abc_4268_new_n1284_; 
wire _abc_4268_new_n1286_; 
wire _abc_4268_new_n1287_; 
wire _abc_4268_new_n1288_; 
wire _abc_4268_new_n1290_; 
wire _abc_4268_new_n1291_; 
wire _abc_4268_new_n1292_; 
wire _abc_4268_new_n1294_; 
wire _abc_4268_new_n1295_; 
wire _abc_4268_new_n1296_; 
wire _abc_4268_new_n1298_; 
wire _abc_4268_new_n1299_; 
wire _abc_4268_new_n1300_; 
wire _abc_4268_new_n1302_; 
wire _abc_4268_new_n1303_; 
wire _abc_4268_new_n1304_; 
wire _abc_4268_new_n1306_; 
wire _abc_4268_new_n1307_; 
wire _abc_4268_new_n1308_; 
wire _abc_4268_new_n1310_; 
wire _abc_4268_new_n1311_; 
wire _abc_4268_new_n1312_; 
wire _abc_4268_new_n1314_; 
wire _abc_4268_new_n1315_; 
wire _abc_4268_new_n1316_; 
wire _abc_4268_new_n1318_; 
wire _abc_4268_new_n1319_; 
wire _abc_4268_new_n1320_; 
wire _abc_4268_new_n1322_; 
wire _abc_4268_new_n1323_; 
wire _abc_4268_new_n1324_; 
wire _abc_4268_new_n1326_; 
wire _abc_4268_new_n1327_; 
wire _abc_4268_new_n1328_; 
wire _abc_4268_new_n1330_; 
wire _abc_4268_new_n1331_; 
wire _abc_4268_new_n1332_; 
wire _abc_4268_new_n1334_; 
wire _abc_4268_new_n1335_; 
wire _abc_4268_new_n1336_; 
wire _abc_4268_new_n1338_; 
wire _abc_4268_new_n1339_; 
wire _abc_4268_new_n1340_; 
wire _abc_4268_new_n1342_; 
wire _abc_4268_new_n1343_; 
wire _abc_4268_new_n1344_; 
wire _abc_4268_new_n1346_; 
wire _abc_4268_new_n1347_; 
wire _abc_4268_new_n1348_; 
wire _abc_4268_new_n1350_; 
wire _abc_4268_new_n1351_; 
wire _abc_4268_new_n1352_; 
wire _abc_4268_new_n1354_; 
wire _abc_4268_new_n1355_; 
wire _abc_4268_new_n1356_; 
wire _abc_4268_new_n1358_; 
wire _abc_4268_new_n1359_; 
wire _abc_4268_new_n1360_; 
wire _abc_4268_new_n1362_; 
wire _abc_4268_new_n1363_; 
wire _abc_4268_new_n1364_; 
wire _abc_4268_new_n1366_; 
wire _abc_4268_new_n1367_; 
wire _abc_4268_new_n1368_; 
wire _abc_4268_new_n1370_; 
wire _abc_4268_new_n1371_; 
wire _abc_4268_new_n1372_; 
wire _abc_4268_new_n1374_; 
wire _abc_4268_new_n1375_; 
wire _abc_4268_new_n1376_; 
wire _abc_4268_new_n1378_; 
wire _abc_4268_new_n1379_; 
wire _abc_4268_new_n1380_; 
wire _abc_4268_new_n1382_; 
wire _abc_4268_new_n1383_; 
wire _abc_4268_new_n1384_; 
wire _abc_4268_new_n1386_; 
wire _abc_4268_new_n1387_; 
wire _abc_4268_new_n1388_; 
wire _abc_4268_new_n1390_; 
wire _abc_4268_new_n1391_; 
wire _abc_4268_new_n1392_; 
wire _abc_4268_new_n1394_; 
wire _abc_4268_new_n1395_; 
wire _abc_4268_new_n1396_; 
wire _abc_4268_new_n1398_; 
wire _abc_4268_new_n1399_; 
wire _abc_4268_new_n1400_; 
wire _abc_4268_new_n1402_; 
wire _abc_4268_new_n1403_; 
wire _abc_4268_new_n1404_; 
wire _abc_4268_new_n1406_; 
wire _abc_4268_new_n1407_; 
wire _abc_4268_new_n1408_; 
wire _abc_4268_new_n1410_; 
wire _abc_4268_new_n1411_; 
wire _abc_4268_new_n1412_; 
wire _abc_4268_new_n1414_; 
wire _abc_4268_new_n1415_; 
wire _abc_4268_new_n1416_; 
wire _abc_4268_new_n1418_; 
wire _abc_4268_new_n1419_; 
wire _abc_4268_new_n1420_; 
wire _abc_4268_new_n1422_; 
wire _abc_4268_new_n1423_; 
wire _abc_4268_new_n1424_; 
wire _abc_4268_new_n1426_; 
wire _abc_4268_new_n1427_; 
wire _abc_4268_new_n1428_; 
wire _abc_4268_new_n1430_; 
wire _abc_4268_new_n1431_; 
wire _abc_4268_new_n1432_; 
wire _abc_4268_new_n1434_; 
wire _abc_4268_new_n1435_; 
wire _abc_4268_new_n1436_; 
wire _abc_4268_new_n1438_; 
wire _abc_4268_new_n1439_; 
wire _abc_4268_new_n1440_; 
wire _abc_4268_new_n1442_; 
wire _abc_4268_new_n1443_; 
wire _abc_4268_new_n1444_; 
wire _abc_4268_new_n1446_; 
wire _abc_4268_new_n1447_; 
wire _abc_4268_new_n1448_; 
wire _abc_4268_new_n1450_; 
wire _abc_4268_new_n1451_; 
wire _abc_4268_new_n1452_; 
wire _abc_4268_new_n1454_; 
wire _abc_4268_new_n1455_; 
wire _abc_4268_new_n1456_; 
wire _abc_4268_new_n1458_; 
wire _abc_4268_new_n1459_; 
wire _abc_4268_new_n1460_; 
wire _abc_4268_new_n1462_; 
wire _abc_4268_new_n1463_; 
wire _abc_4268_new_n1464_; 
wire _abc_4268_new_n1466_; 
wire _abc_4268_new_n1467_; 
wire _abc_4268_new_n1468_; 
wire _abc_4268_new_n1470_; 
wire _abc_4268_new_n1537_; 
wire _abc_4268_new_n1538_; 
wire _abc_4268_new_n1539_; 
wire _abc_4268_new_n1540_; 
wire _abc_4268_new_n1541_; 
wire _abc_4268_new_n1543_; 
wire _abc_4268_new_n1544_; 
wire _abc_4268_new_n1545_; 
wire _abc_4268_new_n1547_; 
wire _abc_4268_new_n1548_; 
wire _abc_4268_new_n1549_; 
wire _abc_4268_new_n1550_; 
wire _abc_4268_new_n558_; 
wire _abc_4268_new_n559_; 
wire _abc_4268_new_n560_; 
wire _abc_4268_new_n561_; 
wire _abc_4268_new_n562_; 
wire _abc_4268_new_n564_; 
wire _abc_4268_new_n566_; 
wire _abc_4268_new_n567_; 
wire _abc_4268_new_n568_; 
wire _abc_4268_new_n569_; 
wire _abc_4268_new_n571_; 
wire _abc_4268_new_n572_; 
wire _abc_4268_new_n573_; 
wire _abc_4268_new_n575_; 
wire _abc_4268_new_n576_; 
wire _abc_4268_new_n577_; 
wire _abc_4268_new_n578_; 
wire _abc_4268_new_n579_; 
wire _abc_4268_new_n580_; 
wire _abc_4268_new_n581_; 
wire _abc_4268_new_n582_; 
wire _abc_4268_new_n583_; 
wire _abc_4268_new_n584_; 
wire _abc_4268_new_n585_; 
wire _abc_4268_new_n586_; 
wire _abc_4268_new_n587_; 
wire _abc_4268_new_n589_; 
wire _abc_4268_new_n590_; 
wire _abc_4268_new_n591_; 
wire _abc_4268_new_n592_; 
wire _abc_4268_new_n594_; 
wire _abc_4268_new_n596_; 
wire _abc_4268_new_n598_; 
wire _abc_4268_new_n599_; 
wire _abc_4268_new_n600_; 
wire _abc_4268_new_n602_; 
wire _abc_4268_new_n603_; 
wire _abc_4268_new_n604_; 
wire _abc_4268_new_n605_; 
wire _abc_4268_new_n606_; 
wire _abc_4268_new_n607_; 
wire _abc_4268_new_n608_; 
wire _abc_4268_new_n610_; 
wire _abc_4268_new_n611_; 
wire _abc_4268_new_n612_; 
wire _abc_4268_new_n613_; 
wire _abc_4268_new_n615_; 
wire _abc_4268_new_n616_; 
wire _abc_4268_new_n617_; 
wire _abc_4268_new_n618_; 
wire _abc_4268_new_n619_; 
wire _abc_4268_new_n620_; 
wire _abc_4268_new_n621_; 
wire _abc_4268_new_n622_; 
wire _abc_4268_new_n623_; 
wire _abc_4268_new_n624_; 
wire _abc_4268_new_n625_; 
wire _abc_4268_new_n626_; 
wire _abc_4268_new_n627_; 
wire _abc_4268_new_n628_; 
wire _abc_4268_new_n629_; 
wire _abc_4268_new_n630_; 
wire _abc_4268_new_n631_; 
wire _abc_4268_new_n632_; 
wire _abc_4268_new_n633_; 
wire _abc_4268_new_n634_; 
wire _abc_4268_new_n635_; 
wire _abc_4268_new_n636_; 
wire _abc_4268_new_n637_; 
wire _abc_4268_new_n638_; 
wire _abc_4268_new_n639_; 
wire _abc_4268_new_n640_; 
wire _abc_4268_new_n641_; 
wire _abc_4268_new_n642_; 
wire _abc_4268_new_n643_; 
wire _abc_4268_new_n644_; 
wire _abc_4268_new_n645_; 
wire _abc_4268_new_n646_; 
wire _abc_4268_new_n647_; 
wire _abc_4268_new_n648_; 
wire _abc_4268_new_n649_; 
wire _abc_4268_new_n650_; 
wire _abc_4268_new_n651_; 
wire _abc_4268_new_n652_; 
wire _abc_4268_new_n653_; 
wire _abc_4268_new_n654_; 
wire _abc_4268_new_n655_; 
wire _abc_4268_new_n656_; 
wire _abc_4268_new_n657_; 
wire _abc_4268_new_n658_; 
wire _abc_4268_new_n659_; 
wire _abc_4268_new_n660_; 
wire _abc_4268_new_n661_; 
wire _abc_4268_new_n662_; 
wire _abc_4268_new_n663_; 
wire _abc_4268_new_n664_; 
wire _abc_4268_new_n665_; 
wire _abc_4268_new_n666_; 
wire _abc_4268_new_n667_; 
wire _abc_4268_new_n668_; 
wire _abc_4268_new_n669_; 
wire _abc_4268_new_n670_; 
wire _abc_4268_new_n671_; 
wire _abc_4268_new_n672_; 
wire _abc_4268_new_n673_; 
wire _abc_4268_new_n674_; 
wire _abc_4268_new_n675_; 
wire _abc_4268_new_n676_; 
wire _abc_4268_new_n677_; 
wire _abc_4268_new_n678_; 
wire _abc_4268_new_n679_; 
wire _abc_4268_new_n680_; 
wire _abc_4268_new_n681_; 
wire _abc_4268_new_n682_; 
wire _abc_4268_new_n683_; 
wire _abc_4268_new_n685_; 
wire _abc_4268_new_n686_; 
wire _abc_4268_new_n687_; 
wire _abc_4268_new_n688_; 
wire _abc_4268_new_n689_; 
wire _abc_4268_new_n690_; 
wire _abc_4268_new_n691_; 
wire _abc_4268_new_n692_; 
wire _abc_4268_new_n693_; 
wire _abc_4268_new_n694_; 
wire _abc_4268_new_n695_; 
wire _abc_4268_new_n696_; 
wire _abc_4268_new_n697_; 
wire _abc_4268_new_n698_; 
wire _abc_4268_new_n699_; 
wire _abc_4268_new_n700_; 
wire _abc_4268_new_n701_; 
wire _abc_4268_new_n702_; 
wire _abc_4268_new_n703_; 
wire _abc_4268_new_n704_; 
wire _abc_4268_new_n705_; 
wire _abc_4268_new_n706_; 
wire _abc_4268_new_n707_; 
wire _abc_4268_new_n708_; 
wire _abc_4268_new_n709_; 
wire _abc_4268_new_n710_; 
wire _abc_4268_new_n712_; 
wire _abc_4268_new_n713_; 
wire _abc_4268_new_n714_; 
wire _abc_4268_new_n715_; 
wire _abc_4268_new_n716_; 
wire _abc_4268_new_n717_; 
wire _abc_4268_new_n718_; 
wire _abc_4268_new_n719_; 
wire _abc_4268_new_n720_; 
wire _abc_4268_new_n722_; 
wire _abc_4268_new_n723_; 
wire _abc_4268_new_n724_; 
wire _abc_4268_new_n725_; 
wire _abc_4268_new_n726_; 
wire _abc_4268_new_n727_; 
wire _abc_4268_new_n728_; 
wire _abc_4268_new_n730_; 
wire _abc_4268_new_n731_; 
wire _abc_4268_new_n732_; 
wire _abc_4268_new_n733_; 
wire _abc_4268_new_n734_; 
wire _abc_4268_new_n735_; 
wire _abc_4268_new_n736_; 
wire _abc_4268_new_n738_; 
wire _abc_4268_new_n739_; 
wire _abc_4268_new_n740_; 
wire _abc_4268_new_n741_; 
wire _abc_4268_new_n742_; 
wire _abc_4268_new_n743_; 
wire _abc_4268_new_n744_; 
wire _abc_4268_new_n746_; 
wire _abc_4268_new_n747_; 
wire _abc_4268_new_n748_; 
wire _abc_4268_new_n749_; 
wire _abc_4268_new_n750_; 
wire _abc_4268_new_n751_; 
wire _abc_4268_new_n752_; 
wire _abc_4268_new_n754_; 
wire _abc_4268_new_n755_; 
wire _abc_4268_new_n756_; 
wire _abc_4268_new_n757_; 
wire _abc_4268_new_n758_; 
wire _abc_4268_new_n759_; 
wire _abc_4268_new_n760_; 
wire _abc_4268_new_n762_; 
wire _abc_4268_new_n763_; 
wire _abc_4268_new_n764_; 
wire _abc_4268_new_n765_; 
wire _abc_4268_new_n766_; 
wire _abc_4268_new_n767_; 
wire _abc_4268_new_n768_; 
wire _abc_4268_new_n770_; 
wire _abc_4268_new_n771_; 
wire _abc_4268_new_n772_; 
wire _abc_4268_new_n773_; 
wire _abc_4268_new_n774_; 
wire _abc_4268_new_n775_; 
wire _abc_4268_new_n776_; 
wire _abc_4268_new_n778_; 
wire _abc_4268_new_n779_; 
wire _abc_4268_new_n780_; 
wire _abc_4268_new_n781_; 
wire _abc_4268_new_n782_; 
wire _abc_4268_new_n783_; 
wire _abc_4268_new_n784_; 
wire _abc_4268_new_n786_; 
wire _abc_4268_new_n787_; 
wire _abc_4268_new_n788_; 
wire _abc_4268_new_n789_; 
wire _abc_4268_new_n790_; 
wire _abc_4268_new_n791_; 
wire _abc_4268_new_n792_; 
wire _abc_4268_new_n794_; 
wire _abc_4268_new_n795_; 
wire _abc_4268_new_n796_; 
wire _abc_4268_new_n797_; 
wire _abc_4268_new_n798_; 
wire _abc_4268_new_n799_; 
wire _abc_4268_new_n800_; 
wire _abc_4268_new_n802_; 
wire _abc_4268_new_n803_; 
wire _abc_4268_new_n804_; 
wire _abc_4268_new_n805_; 
wire _abc_4268_new_n806_; 
wire _abc_4268_new_n807_; 
wire _abc_4268_new_n808_; 
wire _abc_4268_new_n810_; 
wire _abc_4268_new_n811_; 
wire _abc_4268_new_n812_; 
wire _abc_4268_new_n813_; 
wire _abc_4268_new_n814_; 
wire _abc_4268_new_n815_; 
wire _abc_4268_new_n816_; 
wire _abc_4268_new_n818_; 
wire _abc_4268_new_n819_; 
wire _abc_4268_new_n820_; 
wire _abc_4268_new_n821_; 
wire _abc_4268_new_n822_; 
wire _abc_4268_new_n823_; 
wire _abc_4268_new_n824_; 
wire _abc_4268_new_n826_; 
wire _abc_4268_new_n827_; 
wire _abc_4268_new_n828_; 
wire _abc_4268_new_n829_; 
wire _abc_4268_new_n830_; 
wire _abc_4268_new_n831_; 
wire _abc_4268_new_n832_; 
wire _abc_4268_new_n834_; 
wire _abc_4268_new_n835_; 
wire _abc_4268_new_n836_; 
wire _abc_4268_new_n837_; 
wire _abc_4268_new_n838_; 
wire _abc_4268_new_n839_; 
wire _abc_4268_new_n840_; 
wire _abc_4268_new_n842_; 
wire _abc_4268_new_n843_; 
wire _abc_4268_new_n844_; 
wire _abc_4268_new_n845_; 
wire _abc_4268_new_n846_; 
wire _abc_4268_new_n847_; 
wire _abc_4268_new_n848_; 
wire _abc_4268_new_n850_; 
wire _abc_4268_new_n851_; 
wire _abc_4268_new_n852_; 
wire _abc_4268_new_n853_; 
wire _abc_4268_new_n854_; 
wire _abc_4268_new_n855_; 
wire _abc_4268_new_n856_; 
wire _abc_4268_new_n858_; 
wire _abc_4268_new_n859_; 
wire _abc_4268_new_n860_; 
wire _abc_4268_new_n861_; 
wire _abc_4268_new_n862_; 
wire _abc_4268_new_n863_; 
wire _abc_4268_new_n864_; 
wire _abc_4268_new_n866_; 
wire _abc_4268_new_n867_; 
wire _abc_4268_new_n868_; 
wire _abc_4268_new_n869_; 
wire _abc_4268_new_n870_; 
wire _abc_4268_new_n871_; 
wire _abc_4268_new_n872_; 
wire _abc_4268_new_n874_; 
wire _abc_4268_new_n875_; 
wire _abc_4268_new_n876_; 
wire _abc_4268_new_n877_; 
wire _abc_4268_new_n878_; 
wire _abc_4268_new_n879_; 
wire _abc_4268_new_n880_; 
wire _abc_4268_new_n882_; 
wire _abc_4268_new_n883_; 
wire _abc_4268_new_n884_; 
wire _abc_4268_new_n885_; 
wire _abc_4268_new_n886_; 
wire _abc_4268_new_n887_; 
wire _abc_4268_new_n888_; 
wire _abc_4268_new_n890_; 
wire _abc_4268_new_n891_; 
wire _abc_4268_new_n892_; 
wire _abc_4268_new_n893_; 
wire _abc_4268_new_n894_; 
wire _abc_4268_new_n895_; 
wire _abc_4268_new_n896_; 
wire _abc_4268_new_n898_; 
wire _abc_4268_new_n899_; 
wire _abc_4268_new_n900_; 
wire _abc_4268_new_n901_; 
wire _abc_4268_new_n902_; 
wire _abc_4268_new_n903_; 
wire _abc_4268_new_n904_; 
wire _abc_4268_new_n906_; 
wire _abc_4268_new_n907_; 
wire _abc_4268_new_n908_; 
wire _abc_4268_new_n909_; 
wire _abc_4268_new_n910_; 
wire _abc_4268_new_n911_; 
wire _abc_4268_new_n912_; 
wire _abc_4268_new_n914_; 
wire _abc_4268_new_n915_; 
wire _abc_4268_new_n916_; 
wire _abc_4268_new_n917_; 
wire _abc_4268_new_n918_; 
wire _abc_4268_new_n919_; 
wire _abc_4268_new_n920_; 
wire _abc_4268_new_n922_; 
wire _abc_4268_new_n923_; 
wire _abc_4268_new_n924_; 
wire _abc_4268_new_n925_; 
wire _abc_4268_new_n926_; 
wire _abc_4268_new_n927_; 
wire _abc_4268_new_n928_; 
wire _abc_4268_new_n930_; 
wire _abc_4268_new_n931_; 
wire _abc_4268_new_n932_; 
wire _abc_4268_new_n933_; 
wire _abc_4268_new_n934_; 
wire _abc_4268_new_n935_; 
wire _abc_4268_new_n936_; 
wire _abc_4268_new_n938_; 
wire _abc_4268_new_n939_; 
wire _abc_4268_new_n940_; 
wire _abc_4268_new_n941_; 
wire _abc_4268_new_n942_; 
wire _abc_4268_new_n943_; 
wire _abc_4268_new_n944_; 
wire _abc_4268_new_n946_; 
wire _abc_4268_new_n947_; 
wire _abc_4268_new_n948_; 
wire _abc_4268_new_n949_; 
wire _abc_4268_new_n950_; 
wire _abc_4268_new_n951_; 
wire _abc_4268_new_n952_; 
wire _abc_4268_new_n954_; 
wire _abc_4268_new_n955_; 
wire _abc_4268_new_n956_; 
wire _abc_4268_new_n957_; 
wire _abc_4268_new_n959_; 
wire _abc_4268_new_n960_; 
wire _abc_4268_new_n961_; 
wire _abc_4268_new_n963_; 
wire _abc_4268_new_n964_; 
wire _abc_4268_new_n965_; 
wire _abc_4268_new_n967_; 
wire _abc_4268_new_n968_; 
wire _abc_4268_new_n969_; 
wire _abc_4268_new_n971_; 
wire _abc_4268_new_n972_; 
wire _abc_4268_new_n973_; 
wire _abc_4268_new_n975_; 
wire _abc_4268_new_n976_; 
wire _abc_4268_new_n977_; 
wire _abc_4268_new_n979_; 
wire _abc_4268_new_n980_; 
wire _abc_4268_new_n981_; 
wire _abc_4268_new_n983_; 
wire _abc_4268_new_n984_; 
wire _abc_4268_new_n985_; 
wire _abc_4268_new_n987_; 
wire _abc_4268_new_n988_; 
wire _abc_4268_new_n989_; 
wire _abc_4268_new_n991_; 
wire _abc_4268_new_n992_; 
wire _abc_4268_new_n993_; 
wire _abc_4268_new_n995_; 
wire _abc_4268_new_n996_; 
wire _abc_4268_new_n997_; 
wire _abc_4268_new_n999_; 
output \axi_araddr[0] ;
output \axi_araddr[10] ;
output \axi_araddr[11] ;
output \axi_araddr[12] ;
output \axi_araddr[13] ;
output \axi_araddr[14] ;
output \axi_araddr[15] ;
output \axi_araddr[16] ;
output \axi_araddr[17] ;
output \axi_araddr[18] ;
output \axi_araddr[19] ;
output \axi_araddr[1] ;
output \axi_araddr[20] ;
output \axi_araddr[21] ;
output \axi_araddr[22] ;
output \axi_araddr[23] ;
output \axi_araddr[24] ;
output \axi_araddr[25] ;
output \axi_araddr[26] ;
output \axi_araddr[27] ;
output \axi_araddr[28] ;
output \axi_araddr[29] ;
output \axi_araddr[2] ;
output \axi_araddr[30] ;
output \axi_araddr[31] ;
output \axi_araddr[3] ;
output \axi_araddr[4] ;
output \axi_araddr[5] ;
output \axi_araddr[6] ;
output \axi_araddr[7] ;
output \axi_araddr[8] ;
output \axi_araddr[9] ;
output \axi_arprot[0] ;
output \axi_arprot[1] ;
output \axi_arprot[2] ;
input axi_arready;
output axi_arvalid;
output \axi_awaddr[0] ;
output \axi_awaddr[10] ;
output \axi_awaddr[11] ;
output \axi_awaddr[12] ;
output \axi_awaddr[13] ;
output \axi_awaddr[14] ;
output \axi_awaddr[15] ;
output \axi_awaddr[16] ;
output \axi_awaddr[17] ;
output \axi_awaddr[18] ;
output \axi_awaddr[19] ;
output \axi_awaddr[1] ;
output \axi_awaddr[20] ;
output \axi_awaddr[21] ;
output \axi_awaddr[22] ;
output \axi_awaddr[23] ;
output \axi_awaddr[24] ;
output \axi_awaddr[25] ;
output \axi_awaddr[26] ;
output \axi_awaddr[27] ;
output \axi_awaddr[28] ;
output \axi_awaddr[29] ;
output \axi_awaddr[2] ;
output \axi_awaddr[30] ;
output \axi_awaddr[31] ;
output \axi_awaddr[3] ;
output \axi_awaddr[4] ;
output \axi_awaddr[5] ;
output \axi_awaddr[6] ;
output \axi_awaddr[7] ;
output \axi_awaddr[8] ;
output \axi_awaddr[9] ;
output \axi_awprot[0] ;
output \axi_awprot[1] ;
output \axi_awprot[2] ;
input axi_awready;
output axi_awvalid;
output axi_bready;
input axi_bvalid;
input \axi_rdata[0] ;
input \axi_rdata[10] ;
input \axi_rdata[11] ;
input \axi_rdata[12] ;
input \axi_rdata[13] ;
input \axi_rdata[14] ;
input \axi_rdata[15] ;
input \axi_rdata[16] ;
input \axi_rdata[17] ;
input \axi_rdata[18] ;
input \axi_rdata[19] ;
input \axi_rdata[1] ;
input \axi_rdata[20] ;
input \axi_rdata[21] ;
input \axi_rdata[22] ;
input \axi_rdata[23] ;
input \axi_rdata[24] ;
input \axi_rdata[25] ;
input \axi_rdata[26] ;
input \axi_rdata[27] ;
input \axi_rdata[28] ;
input \axi_rdata[29] ;
input \axi_rdata[2] ;
input \axi_rdata[30] ;
input \axi_rdata[31] ;
input \axi_rdata[3] ;
input \axi_rdata[4] ;
input \axi_rdata[5] ;
input \axi_rdata[6] ;
input \axi_rdata[7] ;
input \axi_rdata[8] ;
input \axi_rdata[9] ;
output axi_rready;
input axi_rvalid;
output \axi_wdata[0] ;
output \axi_wdata[10] ;
output \axi_wdata[11] ;
output \axi_wdata[12] ;
output \axi_wdata[13] ;
output \axi_wdata[14] ;
output \axi_wdata[15] ;
output \axi_wdata[16] ;
output \axi_wdata[17] ;
output \axi_wdata[18] ;
output \axi_wdata[19] ;
output \axi_wdata[1] ;
output \axi_wdata[20] ;
output \axi_wdata[21] ;
output \axi_wdata[22] ;
output \axi_wdata[23] ;
output \axi_wdata[24] ;
output \axi_wdata[25] ;
output \axi_wdata[26] ;
output \axi_wdata[27] ;
output \axi_wdata[28] ;
output \axi_wdata[29] ;
output \axi_wdata[2] ;
output \axi_wdata[30] ;
output \axi_wdata[31] ;
output \axi_wdata[3] ;
output \axi_wdata[4] ;
output \axi_wdata[5] ;
output \axi_wdata[6] ;
output \axi_wdata[7] ;
output \axi_wdata[8] ;
output \axi_wdata[9] ;
input axi_wready;
output \axi_wstrb[0] ;
output \axi_wstrb[1] ;
output \axi_wstrb[2] ;
output \axi_wstrb[3] ;
output axi_wvalid;
wire bus_cap_0_; 
wire bus_cap_10_; 
wire bus_cap_11_; 
wire bus_cap_12_; 
wire bus_cap_13_; 
wire bus_cap_14_; 
wire bus_cap_15_; 
wire bus_cap_16_; 
wire bus_cap_17_; 
wire bus_cap_18_; 
wire bus_cap_19_; 
wire bus_cap_1_; 
wire bus_cap_20_; 
wire bus_cap_21_; 
wire bus_cap_22_; 
wire bus_cap_23_; 
wire bus_cap_24_; 
wire bus_cap_25_; 
wire bus_cap_26_; 
wire bus_cap_27_; 
wire bus_cap_28_; 
wire bus_cap_29_; 
wire bus_cap_2_; 
wire bus_cap_30_; 
wire bus_cap_3_; 
wire bus_cap_4_; 
wire bus_cap_5_; 
wire bus_cap_6_; 
wire bus_cap_7_; 
wire bus_cap_8_; 
wire bus_cap_9_; 
wire bus_sync_axi_bus_ECLK1; 
wire bus_sync_axi_bus_EECLK1; 
wire bus_sync_axi_bus_NCLK2; 
wire bus_sync_axi_bus__0ECLK1_0_0_; 
wire bus_sync_axi_bus__0EECLK1_0_0_; 
wire bus_sync_axi_bus__0reg_data1_63_0__0_; 
wire bus_sync_axi_bus__0reg_data1_63_0__10_; 
wire bus_sync_axi_bus__0reg_data1_63_0__11_; 
wire bus_sync_axi_bus__0reg_data1_63_0__12_; 
wire bus_sync_axi_bus__0reg_data1_63_0__13_; 
wire bus_sync_axi_bus__0reg_data1_63_0__14_; 
wire bus_sync_axi_bus__0reg_data1_63_0__15_; 
wire bus_sync_axi_bus__0reg_data1_63_0__16_; 
wire bus_sync_axi_bus__0reg_data1_63_0__17_; 
wire bus_sync_axi_bus__0reg_data1_63_0__18_; 
wire bus_sync_axi_bus__0reg_data1_63_0__19_; 
wire bus_sync_axi_bus__0reg_data1_63_0__1_; 
wire bus_sync_axi_bus__0reg_data1_63_0__20_; 
wire bus_sync_axi_bus__0reg_data1_63_0__21_; 
wire bus_sync_axi_bus__0reg_data1_63_0__22_; 
wire bus_sync_axi_bus__0reg_data1_63_0__23_; 
wire bus_sync_axi_bus__0reg_data1_63_0__24_; 
wire bus_sync_axi_bus__0reg_data1_63_0__25_; 
wire bus_sync_axi_bus__0reg_data1_63_0__26_; 
wire bus_sync_axi_bus__0reg_data1_63_0__27_; 
wire bus_sync_axi_bus__0reg_data1_63_0__28_; 
wire bus_sync_axi_bus__0reg_data1_63_0__29_; 
wire bus_sync_axi_bus__0reg_data1_63_0__2_; 
wire bus_sync_axi_bus__0reg_data1_63_0__30_; 
wire bus_sync_axi_bus__0reg_data1_63_0__31_; 
wire bus_sync_axi_bus__0reg_data1_63_0__32_; 
wire bus_sync_axi_bus__0reg_data1_63_0__33_; 
wire bus_sync_axi_bus__0reg_data1_63_0__34_; 
wire bus_sync_axi_bus__0reg_data1_63_0__35_; 
wire bus_sync_axi_bus__0reg_data1_63_0__36_; 
wire bus_sync_axi_bus__0reg_data1_63_0__37_; 
wire bus_sync_axi_bus__0reg_data1_63_0__38_; 
wire bus_sync_axi_bus__0reg_data1_63_0__39_; 
wire bus_sync_axi_bus__0reg_data1_63_0__3_; 
wire bus_sync_axi_bus__0reg_data1_63_0__40_; 
wire bus_sync_axi_bus__0reg_data1_63_0__41_; 
wire bus_sync_axi_bus__0reg_data1_63_0__42_; 
wire bus_sync_axi_bus__0reg_data1_63_0__43_; 
wire bus_sync_axi_bus__0reg_data1_63_0__44_; 
wire bus_sync_axi_bus__0reg_data1_63_0__45_; 
wire bus_sync_axi_bus__0reg_data1_63_0__46_; 
wire bus_sync_axi_bus__0reg_data1_63_0__47_; 
wire bus_sync_axi_bus__0reg_data1_63_0__48_; 
wire bus_sync_axi_bus__0reg_data1_63_0__49_; 
wire bus_sync_axi_bus__0reg_data1_63_0__4_; 
wire bus_sync_axi_bus__0reg_data1_63_0__50_; 
wire bus_sync_axi_bus__0reg_data1_63_0__51_; 
wire bus_sync_axi_bus__0reg_data1_63_0__52_; 
wire bus_sync_axi_bus__0reg_data1_63_0__53_; 
wire bus_sync_axi_bus__0reg_data1_63_0__54_; 
wire bus_sync_axi_bus__0reg_data1_63_0__55_; 
wire bus_sync_axi_bus__0reg_data1_63_0__56_; 
wire bus_sync_axi_bus__0reg_data1_63_0__57_; 
wire bus_sync_axi_bus__0reg_data1_63_0__58_; 
wire bus_sync_axi_bus__0reg_data1_63_0__59_; 
wire bus_sync_axi_bus__0reg_data1_63_0__5_; 
wire bus_sync_axi_bus__0reg_data1_63_0__60_; 
wire bus_sync_axi_bus__0reg_data1_63_0__61_; 
wire bus_sync_axi_bus__0reg_data1_63_0__62_; 
wire bus_sync_axi_bus__0reg_data1_63_0__63_; 
wire bus_sync_axi_bus__0reg_data1_63_0__6_; 
wire bus_sync_axi_bus__0reg_data1_63_0__7_; 
wire bus_sync_axi_bus__0reg_data1_63_0__8_; 
wire bus_sync_axi_bus__0reg_data1_63_0__9_; 
wire bus_sync_axi_bus__0reg_data2_63_0__0_; 
wire bus_sync_axi_bus__0reg_data2_63_0__10_; 
wire bus_sync_axi_bus__0reg_data2_63_0__11_; 
wire bus_sync_axi_bus__0reg_data2_63_0__12_; 
wire bus_sync_axi_bus__0reg_data2_63_0__13_; 
wire bus_sync_axi_bus__0reg_data2_63_0__14_; 
wire bus_sync_axi_bus__0reg_data2_63_0__15_; 
wire bus_sync_axi_bus__0reg_data2_63_0__16_; 
wire bus_sync_axi_bus__0reg_data2_63_0__17_; 
wire bus_sync_axi_bus__0reg_data2_63_0__18_; 
wire bus_sync_axi_bus__0reg_data2_63_0__19_; 
wire bus_sync_axi_bus__0reg_data2_63_0__1_; 
wire bus_sync_axi_bus__0reg_data2_63_0__20_; 
wire bus_sync_axi_bus__0reg_data2_63_0__21_; 
wire bus_sync_axi_bus__0reg_data2_63_0__22_; 
wire bus_sync_axi_bus__0reg_data2_63_0__23_; 
wire bus_sync_axi_bus__0reg_data2_63_0__24_; 
wire bus_sync_axi_bus__0reg_data2_63_0__25_; 
wire bus_sync_axi_bus__0reg_data2_63_0__26_; 
wire bus_sync_axi_bus__0reg_data2_63_0__27_; 
wire bus_sync_axi_bus__0reg_data2_63_0__28_; 
wire bus_sync_axi_bus__0reg_data2_63_0__29_; 
wire bus_sync_axi_bus__0reg_data2_63_0__2_; 
wire bus_sync_axi_bus__0reg_data2_63_0__30_; 
wire bus_sync_axi_bus__0reg_data2_63_0__31_; 
wire bus_sync_axi_bus__0reg_data2_63_0__32_; 
wire bus_sync_axi_bus__0reg_data2_63_0__33_; 
wire bus_sync_axi_bus__0reg_data2_63_0__34_; 
wire bus_sync_axi_bus__0reg_data2_63_0__35_; 
wire bus_sync_axi_bus__0reg_data2_63_0__36_; 
wire bus_sync_axi_bus__0reg_data2_63_0__37_; 
wire bus_sync_axi_bus__0reg_data2_63_0__38_; 
wire bus_sync_axi_bus__0reg_data2_63_0__39_; 
wire bus_sync_axi_bus__0reg_data2_63_0__3_; 
wire bus_sync_axi_bus__0reg_data2_63_0__40_; 
wire bus_sync_axi_bus__0reg_data2_63_0__41_; 
wire bus_sync_axi_bus__0reg_data2_63_0__42_; 
wire bus_sync_axi_bus__0reg_data2_63_0__43_; 
wire bus_sync_axi_bus__0reg_data2_63_0__44_; 
wire bus_sync_axi_bus__0reg_data2_63_0__45_; 
wire bus_sync_axi_bus__0reg_data2_63_0__46_; 
wire bus_sync_axi_bus__0reg_data2_63_0__47_; 
wire bus_sync_axi_bus__0reg_data2_63_0__48_; 
wire bus_sync_axi_bus__0reg_data2_63_0__49_; 
wire bus_sync_axi_bus__0reg_data2_63_0__4_; 
wire bus_sync_axi_bus__0reg_data2_63_0__50_; 
wire bus_sync_axi_bus__0reg_data2_63_0__51_; 
wire bus_sync_axi_bus__0reg_data2_63_0__52_; 
wire bus_sync_axi_bus__0reg_data2_63_0__53_; 
wire bus_sync_axi_bus__0reg_data2_63_0__54_; 
wire bus_sync_axi_bus__0reg_data2_63_0__55_; 
wire bus_sync_axi_bus__0reg_data2_63_0__56_; 
wire bus_sync_axi_bus__0reg_data2_63_0__57_; 
wire bus_sync_axi_bus__0reg_data2_63_0__58_; 
wire bus_sync_axi_bus__0reg_data2_63_0__59_; 
wire bus_sync_axi_bus__0reg_data2_63_0__5_; 
wire bus_sync_axi_bus__0reg_data2_63_0__60_; 
wire bus_sync_axi_bus__0reg_data2_63_0__61_; 
wire bus_sync_axi_bus__0reg_data2_63_0__62_; 
wire bus_sync_axi_bus__0reg_data2_63_0__63_; 
wire bus_sync_axi_bus__0reg_data2_63_0__6_; 
wire bus_sync_axi_bus__0reg_data2_63_0__7_; 
wire bus_sync_axi_bus__0reg_data2_63_0__8_; 
wire bus_sync_axi_bus__0reg_data2_63_0__9_; 
wire bus_sync_axi_bus__0reg_data3_63_0__0_; 
wire bus_sync_axi_bus__0reg_data3_63_0__10_; 
wire bus_sync_axi_bus__0reg_data3_63_0__11_; 
wire bus_sync_axi_bus__0reg_data3_63_0__12_; 
wire bus_sync_axi_bus__0reg_data3_63_0__13_; 
wire bus_sync_axi_bus__0reg_data3_63_0__14_; 
wire bus_sync_axi_bus__0reg_data3_63_0__15_; 
wire bus_sync_axi_bus__0reg_data3_63_0__16_; 
wire bus_sync_axi_bus__0reg_data3_63_0__17_; 
wire bus_sync_axi_bus__0reg_data3_63_0__18_; 
wire bus_sync_axi_bus__0reg_data3_63_0__19_; 
wire bus_sync_axi_bus__0reg_data3_63_0__1_; 
wire bus_sync_axi_bus__0reg_data3_63_0__20_; 
wire bus_sync_axi_bus__0reg_data3_63_0__21_; 
wire bus_sync_axi_bus__0reg_data3_63_0__22_; 
wire bus_sync_axi_bus__0reg_data3_63_0__23_; 
wire bus_sync_axi_bus__0reg_data3_63_0__24_; 
wire bus_sync_axi_bus__0reg_data3_63_0__25_; 
wire bus_sync_axi_bus__0reg_data3_63_0__26_; 
wire bus_sync_axi_bus__0reg_data3_63_0__27_; 
wire bus_sync_axi_bus__0reg_data3_63_0__28_; 
wire bus_sync_axi_bus__0reg_data3_63_0__29_; 
wire bus_sync_axi_bus__0reg_data3_63_0__2_; 
wire bus_sync_axi_bus__0reg_data3_63_0__30_; 
wire bus_sync_axi_bus__0reg_data3_63_0__31_; 
wire bus_sync_axi_bus__0reg_data3_63_0__32_; 
wire bus_sync_axi_bus__0reg_data3_63_0__33_; 
wire bus_sync_axi_bus__0reg_data3_63_0__34_; 
wire bus_sync_axi_bus__0reg_data3_63_0__35_; 
wire bus_sync_axi_bus__0reg_data3_63_0__36_; 
wire bus_sync_axi_bus__0reg_data3_63_0__37_; 
wire bus_sync_axi_bus__0reg_data3_63_0__38_; 
wire bus_sync_axi_bus__0reg_data3_63_0__39_; 
wire bus_sync_axi_bus__0reg_data3_63_0__3_; 
wire bus_sync_axi_bus__0reg_data3_63_0__40_; 
wire bus_sync_axi_bus__0reg_data3_63_0__41_; 
wire bus_sync_axi_bus__0reg_data3_63_0__42_; 
wire bus_sync_axi_bus__0reg_data3_63_0__43_; 
wire bus_sync_axi_bus__0reg_data3_63_0__44_; 
wire bus_sync_axi_bus__0reg_data3_63_0__45_; 
wire bus_sync_axi_bus__0reg_data3_63_0__46_; 
wire bus_sync_axi_bus__0reg_data3_63_0__47_; 
wire bus_sync_axi_bus__0reg_data3_63_0__48_; 
wire bus_sync_axi_bus__0reg_data3_63_0__49_; 
wire bus_sync_axi_bus__0reg_data3_63_0__4_; 
wire bus_sync_axi_bus__0reg_data3_63_0__50_; 
wire bus_sync_axi_bus__0reg_data3_63_0__51_; 
wire bus_sync_axi_bus__0reg_data3_63_0__52_; 
wire bus_sync_axi_bus__0reg_data3_63_0__53_; 
wire bus_sync_axi_bus__0reg_data3_63_0__54_; 
wire bus_sync_axi_bus__0reg_data3_63_0__55_; 
wire bus_sync_axi_bus__0reg_data3_63_0__56_; 
wire bus_sync_axi_bus__0reg_data3_63_0__57_; 
wire bus_sync_axi_bus__0reg_data3_63_0__58_; 
wire bus_sync_axi_bus__0reg_data3_63_0__59_; 
wire bus_sync_axi_bus__0reg_data3_63_0__5_; 
wire bus_sync_axi_bus__0reg_data3_63_0__60_; 
wire bus_sync_axi_bus__0reg_data3_63_0__61_; 
wire bus_sync_axi_bus__0reg_data3_63_0__62_; 
wire bus_sync_axi_bus__0reg_data3_63_0__63_; 
wire bus_sync_axi_bus__0reg_data3_63_0__6_; 
wire bus_sync_axi_bus__0reg_data3_63_0__7_; 
wire bus_sync_axi_bus__0reg_data3_63_0__8_; 
wire bus_sync_axi_bus__0reg_data3_63_0__9_; 
wire bus_sync_axi_bus__abc_3879_new_n393_; 
wire bus_sync_axi_bus__abc_3879_new_n394_; 
wire bus_sync_axi_bus__abc_3879_new_n395_; 
wire bus_sync_axi_bus__abc_3879_new_n396_; 
wire bus_sync_axi_bus__abc_3879_new_n398_; 
wire bus_sync_axi_bus__abc_3879_new_n399_; 
wire bus_sync_axi_bus__abc_3879_new_n400_; 
wire bus_sync_axi_bus__abc_3879_new_n402_; 
wire bus_sync_axi_bus__abc_3879_new_n403_; 
wire bus_sync_axi_bus__abc_3879_new_n404_; 
wire bus_sync_axi_bus__abc_3879_new_n406_; 
wire bus_sync_axi_bus__abc_3879_new_n407_; 
wire bus_sync_axi_bus__abc_3879_new_n408_; 
wire bus_sync_axi_bus__abc_3879_new_n410_; 
wire bus_sync_axi_bus__abc_3879_new_n411_; 
wire bus_sync_axi_bus__abc_3879_new_n412_; 
wire bus_sync_axi_bus__abc_3879_new_n414_; 
wire bus_sync_axi_bus__abc_3879_new_n415_; 
wire bus_sync_axi_bus__abc_3879_new_n416_; 
wire bus_sync_axi_bus__abc_3879_new_n418_; 
wire bus_sync_axi_bus__abc_3879_new_n419_; 
wire bus_sync_axi_bus__abc_3879_new_n420_; 
wire bus_sync_axi_bus__abc_3879_new_n422_; 
wire bus_sync_axi_bus__abc_3879_new_n423_; 
wire bus_sync_axi_bus__abc_3879_new_n424_; 
wire bus_sync_axi_bus__abc_3879_new_n426_; 
wire bus_sync_axi_bus__abc_3879_new_n427_; 
wire bus_sync_axi_bus__abc_3879_new_n428_; 
wire bus_sync_axi_bus__abc_3879_new_n430_; 
wire bus_sync_axi_bus__abc_3879_new_n431_; 
wire bus_sync_axi_bus__abc_3879_new_n432_; 
wire bus_sync_axi_bus__abc_3879_new_n434_; 
wire bus_sync_axi_bus__abc_3879_new_n435_; 
wire bus_sync_axi_bus__abc_3879_new_n436_; 
wire bus_sync_axi_bus__abc_3879_new_n438_; 
wire bus_sync_axi_bus__abc_3879_new_n439_; 
wire bus_sync_axi_bus__abc_3879_new_n440_; 
wire bus_sync_axi_bus__abc_3879_new_n442_; 
wire bus_sync_axi_bus__abc_3879_new_n443_; 
wire bus_sync_axi_bus__abc_3879_new_n444_; 
wire bus_sync_axi_bus__abc_3879_new_n446_; 
wire bus_sync_axi_bus__abc_3879_new_n447_; 
wire bus_sync_axi_bus__abc_3879_new_n448_; 
wire bus_sync_axi_bus__abc_3879_new_n450_; 
wire bus_sync_axi_bus__abc_3879_new_n451_; 
wire bus_sync_axi_bus__abc_3879_new_n452_; 
wire bus_sync_axi_bus__abc_3879_new_n454_; 
wire bus_sync_axi_bus__abc_3879_new_n455_; 
wire bus_sync_axi_bus__abc_3879_new_n456_; 
wire bus_sync_axi_bus__abc_3879_new_n458_; 
wire bus_sync_axi_bus__abc_3879_new_n459_; 
wire bus_sync_axi_bus__abc_3879_new_n460_; 
wire bus_sync_axi_bus__abc_3879_new_n462_; 
wire bus_sync_axi_bus__abc_3879_new_n463_; 
wire bus_sync_axi_bus__abc_3879_new_n464_; 
wire bus_sync_axi_bus__abc_3879_new_n466_; 
wire bus_sync_axi_bus__abc_3879_new_n467_; 
wire bus_sync_axi_bus__abc_3879_new_n468_; 
wire bus_sync_axi_bus__abc_3879_new_n470_; 
wire bus_sync_axi_bus__abc_3879_new_n471_; 
wire bus_sync_axi_bus__abc_3879_new_n472_; 
wire bus_sync_axi_bus__abc_3879_new_n474_; 
wire bus_sync_axi_bus__abc_3879_new_n475_; 
wire bus_sync_axi_bus__abc_3879_new_n476_; 
wire bus_sync_axi_bus__abc_3879_new_n478_; 
wire bus_sync_axi_bus__abc_3879_new_n479_; 
wire bus_sync_axi_bus__abc_3879_new_n480_; 
wire bus_sync_axi_bus__abc_3879_new_n482_; 
wire bus_sync_axi_bus__abc_3879_new_n483_; 
wire bus_sync_axi_bus__abc_3879_new_n484_; 
wire bus_sync_axi_bus__abc_3879_new_n486_; 
wire bus_sync_axi_bus__abc_3879_new_n487_; 
wire bus_sync_axi_bus__abc_3879_new_n488_; 
wire bus_sync_axi_bus__abc_3879_new_n490_; 
wire bus_sync_axi_bus__abc_3879_new_n491_; 
wire bus_sync_axi_bus__abc_3879_new_n492_; 
wire bus_sync_axi_bus__abc_3879_new_n494_; 
wire bus_sync_axi_bus__abc_3879_new_n495_; 
wire bus_sync_axi_bus__abc_3879_new_n496_; 
wire bus_sync_axi_bus__abc_3879_new_n498_; 
wire bus_sync_axi_bus__abc_3879_new_n499_; 
wire bus_sync_axi_bus__abc_3879_new_n500_; 
wire bus_sync_axi_bus__abc_3879_new_n502_; 
wire bus_sync_axi_bus__abc_3879_new_n503_; 
wire bus_sync_axi_bus__abc_3879_new_n504_; 
wire bus_sync_axi_bus__abc_3879_new_n506_; 
wire bus_sync_axi_bus__abc_3879_new_n507_; 
wire bus_sync_axi_bus__abc_3879_new_n508_; 
wire bus_sync_axi_bus__abc_3879_new_n510_; 
wire bus_sync_axi_bus__abc_3879_new_n511_; 
wire bus_sync_axi_bus__abc_3879_new_n512_; 
wire bus_sync_axi_bus__abc_3879_new_n514_; 
wire bus_sync_axi_bus__abc_3879_new_n515_; 
wire bus_sync_axi_bus__abc_3879_new_n516_; 
wire bus_sync_axi_bus__abc_3879_new_n518_; 
wire bus_sync_axi_bus__abc_3879_new_n519_; 
wire bus_sync_axi_bus__abc_3879_new_n520_; 
wire bus_sync_axi_bus__abc_3879_new_n522_; 
wire bus_sync_axi_bus__abc_3879_new_n523_; 
wire bus_sync_axi_bus__abc_3879_new_n524_; 
wire bus_sync_axi_bus__abc_3879_new_n526_; 
wire bus_sync_axi_bus__abc_3879_new_n527_; 
wire bus_sync_axi_bus__abc_3879_new_n528_; 
wire bus_sync_axi_bus__abc_3879_new_n530_; 
wire bus_sync_axi_bus__abc_3879_new_n531_; 
wire bus_sync_axi_bus__abc_3879_new_n532_; 
wire bus_sync_axi_bus__abc_3879_new_n534_; 
wire bus_sync_axi_bus__abc_3879_new_n535_; 
wire bus_sync_axi_bus__abc_3879_new_n536_; 
wire bus_sync_axi_bus__abc_3879_new_n538_; 
wire bus_sync_axi_bus__abc_3879_new_n539_; 
wire bus_sync_axi_bus__abc_3879_new_n540_; 
wire bus_sync_axi_bus__abc_3879_new_n542_; 
wire bus_sync_axi_bus__abc_3879_new_n543_; 
wire bus_sync_axi_bus__abc_3879_new_n544_; 
wire bus_sync_axi_bus__abc_3879_new_n546_; 
wire bus_sync_axi_bus__abc_3879_new_n547_; 
wire bus_sync_axi_bus__abc_3879_new_n548_; 
wire bus_sync_axi_bus__abc_3879_new_n550_; 
wire bus_sync_axi_bus__abc_3879_new_n551_; 
wire bus_sync_axi_bus__abc_3879_new_n552_; 
wire bus_sync_axi_bus__abc_3879_new_n554_; 
wire bus_sync_axi_bus__abc_3879_new_n555_; 
wire bus_sync_axi_bus__abc_3879_new_n556_; 
wire bus_sync_axi_bus__abc_3879_new_n558_; 
wire bus_sync_axi_bus__abc_3879_new_n559_; 
wire bus_sync_axi_bus__abc_3879_new_n560_; 
wire bus_sync_axi_bus__abc_3879_new_n562_; 
wire bus_sync_axi_bus__abc_3879_new_n563_; 
wire bus_sync_axi_bus__abc_3879_new_n564_; 
wire bus_sync_axi_bus__abc_3879_new_n566_; 
wire bus_sync_axi_bus__abc_3879_new_n567_; 
wire bus_sync_axi_bus__abc_3879_new_n568_; 
wire bus_sync_axi_bus__abc_3879_new_n570_; 
wire bus_sync_axi_bus__abc_3879_new_n571_; 
wire bus_sync_axi_bus__abc_3879_new_n572_; 
wire bus_sync_axi_bus__abc_3879_new_n574_; 
wire bus_sync_axi_bus__abc_3879_new_n575_; 
wire bus_sync_axi_bus__abc_3879_new_n576_; 
wire bus_sync_axi_bus__abc_3879_new_n578_; 
wire bus_sync_axi_bus__abc_3879_new_n579_; 
wire bus_sync_axi_bus__abc_3879_new_n580_; 
wire bus_sync_axi_bus__abc_3879_new_n582_; 
wire bus_sync_axi_bus__abc_3879_new_n583_; 
wire bus_sync_axi_bus__abc_3879_new_n584_; 
wire bus_sync_axi_bus__abc_3879_new_n586_; 
wire bus_sync_axi_bus__abc_3879_new_n587_; 
wire bus_sync_axi_bus__abc_3879_new_n588_; 
wire bus_sync_axi_bus__abc_3879_new_n590_; 
wire bus_sync_axi_bus__abc_3879_new_n591_; 
wire bus_sync_axi_bus__abc_3879_new_n592_; 
wire bus_sync_axi_bus__abc_3879_new_n594_; 
wire bus_sync_axi_bus__abc_3879_new_n595_; 
wire bus_sync_axi_bus__abc_3879_new_n596_; 
wire bus_sync_axi_bus__abc_3879_new_n598_; 
wire bus_sync_axi_bus__abc_3879_new_n599_; 
wire bus_sync_axi_bus__abc_3879_new_n600_; 
wire bus_sync_axi_bus__abc_3879_new_n602_; 
wire bus_sync_axi_bus__abc_3879_new_n603_; 
wire bus_sync_axi_bus__abc_3879_new_n604_; 
wire bus_sync_axi_bus__abc_3879_new_n606_; 
wire bus_sync_axi_bus__abc_3879_new_n607_; 
wire bus_sync_axi_bus__abc_3879_new_n608_; 
wire bus_sync_axi_bus__abc_3879_new_n610_; 
wire bus_sync_axi_bus__abc_3879_new_n611_; 
wire bus_sync_axi_bus__abc_3879_new_n612_; 
wire bus_sync_axi_bus__abc_3879_new_n614_; 
wire bus_sync_axi_bus__abc_3879_new_n615_; 
wire bus_sync_axi_bus__abc_3879_new_n616_; 
wire bus_sync_axi_bus__abc_3879_new_n618_; 
wire bus_sync_axi_bus__abc_3879_new_n619_; 
wire bus_sync_axi_bus__abc_3879_new_n620_; 
wire bus_sync_axi_bus__abc_3879_new_n622_; 
wire bus_sync_axi_bus__abc_3879_new_n623_; 
wire bus_sync_axi_bus__abc_3879_new_n624_; 
wire bus_sync_axi_bus__abc_3879_new_n626_; 
wire bus_sync_axi_bus__abc_3879_new_n627_; 
wire bus_sync_axi_bus__abc_3879_new_n628_; 
wire bus_sync_axi_bus__abc_3879_new_n630_; 
wire bus_sync_axi_bus__abc_3879_new_n631_; 
wire bus_sync_axi_bus__abc_3879_new_n632_; 
wire bus_sync_axi_bus__abc_3879_new_n634_; 
wire bus_sync_axi_bus__abc_3879_new_n635_; 
wire bus_sync_axi_bus__abc_3879_new_n636_; 
wire bus_sync_axi_bus__abc_3879_new_n638_; 
wire bus_sync_axi_bus__abc_3879_new_n639_; 
wire bus_sync_axi_bus__abc_3879_new_n640_; 
wire bus_sync_axi_bus__abc_3879_new_n642_; 
wire bus_sync_axi_bus__abc_3879_new_n643_; 
wire bus_sync_axi_bus__abc_3879_new_n644_; 
wire bus_sync_axi_bus__abc_3879_new_n646_; 
wire bus_sync_axi_bus__abc_3879_new_n647_; 
wire bus_sync_axi_bus__abc_3879_new_n648_; 
wire bus_sync_axi_bus_reg_data1_0_; 
wire bus_sync_axi_bus_reg_data1_10_; 
wire bus_sync_axi_bus_reg_data1_11_; 
wire bus_sync_axi_bus_reg_data1_12_; 
wire bus_sync_axi_bus_reg_data1_13_; 
wire bus_sync_axi_bus_reg_data1_14_; 
wire bus_sync_axi_bus_reg_data1_15_; 
wire bus_sync_axi_bus_reg_data1_16_; 
wire bus_sync_axi_bus_reg_data1_17_; 
wire bus_sync_axi_bus_reg_data1_18_; 
wire bus_sync_axi_bus_reg_data1_19_; 
wire bus_sync_axi_bus_reg_data1_1_; 
wire bus_sync_axi_bus_reg_data1_20_; 
wire bus_sync_axi_bus_reg_data1_21_; 
wire bus_sync_axi_bus_reg_data1_22_; 
wire bus_sync_axi_bus_reg_data1_23_; 
wire bus_sync_axi_bus_reg_data1_24_; 
wire bus_sync_axi_bus_reg_data1_25_; 
wire bus_sync_axi_bus_reg_data1_26_; 
wire bus_sync_axi_bus_reg_data1_27_; 
wire bus_sync_axi_bus_reg_data1_28_; 
wire bus_sync_axi_bus_reg_data1_29_; 
wire bus_sync_axi_bus_reg_data1_2_; 
wire bus_sync_axi_bus_reg_data1_30_; 
wire bus_sync_axi_bus_reg_data1_31_; 
wire bus_sync_axi_bus_reg_data1_32_; 
wire bus_sync_axi_bus_reg_data1_33_; 
wire bus_sync_axi_bus_reg_data1_34_; 
wire bus_sync_axi_bus_reg_data1_35_; 
wire bus_sync_axi_bus_reg_data1_36_; 
wire bus_sync_axi_bus_reg_data1_37_; 
wire bus_sync_axi_bus_reg_data1_38_; 
wire bus_sync_axi_bus_reg_data1_39_; 
wire bus_sync_axi_bus_reg_data1_3_; 
wire bus_sync_axi_bus_reg_data1_40_; 
wire bus_sync_axi_bus_reg_data1_41_; 
wire bus_sync_axi_bus_reg_data1_42_; 
wire bus_sync_axi_bus_reg_data1_43_; 
wire bus_sync_axi_bus_reg_data1_44_; 
wire bus_sync_axi_bus_reg_data1_45_; 
wire bus_sync_axi_bus_reg_data1_46_; 
wire bus_sync_axi_bus_reg_data1_47_; 
wire bus_sync_axi_bus_reg_data1_48_; 
wire bus_sync_axi_bus_reg_data1_49_; 
wire bus_sync_axi_bus_reg_data1_4_; 
wire bus_sync_axi_bus_reg_data1_50_; 
wire bus_sync_axi_bus_reg_data1_51_; 
wire bus_sync_axi_bus_reg_data1_52_; 
wire bus_sync_axi_bus_reg_data1_53_; 
wire bus_sync_axi_bus_reg_data1_54_; 
wire bus_sync_axi_bus_reg_data1_55_; 
wire bus_sync_axi_bus_reg_data1_56_; 
wire bus_sync_axi_bus_reg_data1_57_; 
wire bus_sync_axi_bus_reg_data1_58_; 
wire bus_sync_axi_bus_reg_data1_59_; 
wire bus_sync_axi_bus_reg_data1_5_; 
wire bus_sync_axi_bus_reg_data1_60_; 
wire bus_sync_axi_bus_reg_data1_61_; 
wire bus_sync_axi_bus_reg_data1_62_; 
wire bus_sync_axi_bus_reg_data1_63_; 
wire bus_sync_axi_bus_reg_data1_6_; 
wire bus_sync_axi_bus_reg_data1_7_; 
wire bus_sync_axi_bus_reg_data1_8_; 
wire bus_sync_axi_bus_reg_data1_9_; 
wire bus_sync_axi_bus_reg_data2_0_; 
wire bus_sync_axi_bus_reg_data2_10_; 
wire bus_sync_axi_bus_reg_data2_11_; 
wire bus_sync_axi_bus_reg_data2_12_; 
wire bus_sync_axi_bus_reg_data2_13_; 
wire bus_sync_axi_bus_reg_data2_14_; 
wire bus_sync_axi_bus_reg_data2_15_; 
wire bus_sync_axi_bus_reg_data2_16_; 
wire bus_sync_axi_bus_reg_data2_17_; 
wire bus_sync_axi_bus_reg_data2_18_; 
wire bus_sync_axi_bus_reg_data2_19_; 
wire bus_sync_axi_bus_reg_data2_1_; 
wire bus_sync_axi_bus_reg_data2_20_; 
wire bus_sync_axi_bus_reg_data2_21_; 
wire bus_sync_axi_bus_reg_data2_22_; 
wire bus_sync_axi_bus_reg_data2_23_; 
wire bus_sync_axi_bus_reg_data2_24_; 
wire bus_sync_axi_bus_reg_data2_25_; 
wire bus_sync_axi_bus_reg_data2_26_; 
wire bus_sync_axi_bus_reg_data2_27_; 
wire bus_sync_axi_bus_reg_data2_28_; 
wire bus_sync_axi_bus_reg_data2_29_; 
wire bus_sync_axi_bus_reg_data2_2_; 
wire bus_sync_axi_bus_reg_data2_30_; 
wire bus_sync_axi_bus_reg_data2_31_; 
wire bus_sync_axi_bus_reg_data2_32_; 
wire bus_sync_axi_bus_reg_data2_33_; 
wire bus_sync_axi_bus_reg_data2_34_; 
wire bus_sync_axi_bus_reg_data2_35_; 
wire bus_sync_axi_bus_reg_data2_36_; 
wire bus_sync_axi_bus_reg_data2_37_; 
wire bus_sync_axi_bus_reg_data2_38_; 
wire bus_sync_axi_bus_reg_data2_39_; 
wire bus_sync_axi_bus_reg_data2_3_; 
wire bus_sync_axi_bus_reg_data2_40_; 
wire bus_sync_axi_bus_reg_data2_41_; 
wire bus_sync_axi_bus_reg_data2_42_; 
wire bus_sync_axi_bus_reg_data2_43_; 
wire bus_sync_axi_bus_reg_data2_44_; 
wire bus_sync_axi_bus_reg_data2_45_; 
wire bus_sync_axi_bus_reg_data2_46_; 
wire bus_sync_axi_bus_reg_data2_47_; 
wire bus_sync_axi_bus_reg_data2_48_; 
wire bus_sync_axi_bus_reg_data2_49_; 
wire bus_sync_axi_bus_reg_data2_4_; 
wire bus_sync_axi_bus_reg_data2_50_; 
wire bus_sync_axi_bus_reg_data2_51_; 
wire bus_sync_axi_bus_reg_data2_52_; 
wire bus_sync_axi_bus_reg_data2_53_; 
wire bus_sync_axi_bus_reg_data2_54_; 
wire bus_sync_axi_bus_reg_data2_55_; 
wire bus_sync_axi_bus_reg_data2_56_; 
wire bus_sync_axi_bus_reg_data2_57_; 
wire bus_sync_axi_bus_reg_data2_58_; 
wire bus_sync_axi_bus_reg_data2_59_; 
wire bus_sync_axi_bus_reg_data2_5_; 
wire bus_sync_axi_bus_reg_data2_60_; 
wire bus_sync_axi_bus_reg_data2_61_; 
wire bus_sync_axi_bus_reg_data2_62_; 
wire bus_sync_axi_bus_reg_data2_63_; 
wire bus_sync_axi_bus_reg_data2_6_; 
wire bus_sync_axi_bus_reg_data2_7_; 
wire bus_sync_axi_bus_reg_data2_8_; 
wire bus_sync_axi_bus_reg_data2_9_; 
wire bus_sync_rdata_ECLK2; 
wire bus_sync_rdata_EECLK2; 
wire bus_sync_rdata_NCLK1; 
wire bus_sync_rdata__0ECLK2_0_0_; 
wire bus_sync_rdata__0EECLK2_0_0_; 
wire bus_sync_rdata__0reg_data1_31_0__0_; 
wire bus_sync_rdata__0reg_data1_31_0__10_; 
wire bus_sync_rdata__0reg_data1_31_0__11_; 
wire bus_sync_rdata__0reg_data1_31_0__12_; 
wire bus_sync_rdata__0reg_data1_31_0__13_; 
wire bus_sync_rdata__0reg_data1_31_0__14_; 
wire bus_sync_rdata__0reg_data1_31_0__15_; 
wire bus_sync_rdata__0reg_data1_31_0__16_; 
wire bus_sync_rdata__0reg_data1_31_0__17_; 
wire bus_sync_rdata__0reg_data1_31_0__18_; 
wire bus_sync_rdata__0reg_data1_31_0__19_; 
wire bus_sync_rdata__0reg_data1_31_0__1_; 
wire bus_sync_rdata__0reg_data1_31_0__20_; 
wire bus_sync_rdata__0reg_data1_31_0__21_; 
wire bus_sync_rdata__0reg_data1_31_0__22_; 
wire bus_sync_rdata__0reg_data1_31_0__23_; 
wire bus_sync_rdata__0reg_data1_31_0__24_; 
wire bus_sync_rdata__0reg_data1_31_0__25_; 
wire bus_sync_rdata__0reg_data1_31_0__26_; 
wire bus_sync_rdata__0reg_data1_31_0__27_; 
wire bus_sync_rdata__0reg_data1_31_0__28_; 
wire bus_sync_rdata__0reg_data1_31_0__29_; 
wire bus_sync_rdata__0reg_data1_31_0__2_; 
wire bus_sync_rdata__0reg_data1_31_0__30_; 
wire bus_sync_rdata__0reg_data1_31_0__31_; 
wire bus_sync_rdata__0reg_data1_31_0__3_; 
wire bus_sync_rdata__0reg_data1_31_0__4_; 
wire bus_sync_rdata__0reg_data1_31_0__5_; 
wire bus_sync_rdata__0reg_data1_31_0__6_; 
wire bus_sync_rdata__0reg_data1_31_0__7_; 
wire bus_sync_rdata__0reg_data1_31_0__8_; 
wire bus_sync_rdata__0reg_data1_31_0__9_; 
wire bus_sync_rdata__0reg_data2_31_0__0_; 
wire bus_sync_rdata__0reg_data2_31_0__10_; 
wire bus_sync_rdata__0reg_data2_31_0__11_; 
wire bus_sync_rdata__0reg_data2_31_0__12_; 
wire bus_sync_rdata__0reg_data2_31_0__13_; 
wire bus_sync_rdata__0reg_data2_31_0__14_; 
wire bus_sync_rdata__0reg_data2_31_0__15_; 
wire bus_sync_rdata__0reg_data2_31_0__16_; 
wire bus_sync_rdata__0reg_data2_31_0__17_; 
wire bus_sync_rdata__0reg_data2_31_0__18_; 
wire bus_sync_rdata__0reg_data2_31_0__19_; 
wire bus_sync_rdata__0reg_data2_31_0__1_; 
wire bus_sync_rdata__0reg_data2_31_0__20_; 
wire bus_sync_rdata__0reg_data2_31_0__21_; 
wire bus_sync_rdata__0reg_data2_31_0__22_; 
wire bus_sync_rdata__0reg_data2_31_0__23_; 
wire bus_sync_rdata__0reg_data2_31_0__24_; 
wire bus_sync_rdata__0reg_data2_31_0__25_; 
wire bus_sync_rdata__0reg_data2_31_0__26_; 
wire bus_sync_rdata__0reg_data2_31_0__27_; 
wire bus_sync_rdata__0reg_data2_31_0__28_; 
wire bus_sync_rdata__0reg_data2_31_0__29_; 
wire bus_sync_rdata__0reg_data2_31_0__2_; 
wire bus_sync_rdata__0reg_data2_31_0__30_; 
wire bus_sync_rdata__0reg_data2_31_0__31_; 
wire bus_sync_rdata__0reg_data2_31_0__3_; 
wire bus_sync_rdata__0reg_data2_31_0__4_; 
wire bus_sync_rdata__0reg_data2_31_0__5_; 
wire bus_sync_rdata__0reg_data2_31_0__6_; 
wire bus_sync_rdata__0reg_data2_31_0__7_; 
wire bus_sync_rdata__0reg_data2_31_0__8_; 
wire bus_sync_rdata__0reg_data2_31_0__9_; 
wire bus_sync_rdata__0reg_data3_31_0__0_; 
wire bus_sync_rdata__0reg_data3_31_0__10_; 
wire bus_sync_rdata__0reg_data3_31_0__11_; 
wire bus_sync_rdata__0reg_data3_31_0__12_; 
wire bus_sync_rdata__0reg_data3_31_0__13_; 
wire bus_sync_rdata__0reg_data3_31_0__14_; 
wire bus_sync_rdata__0reg_data3_31_0__15_; 
wire bus_sync_rdata__0reg_data3_31_0__16_; 
wire bus_sync_rdata__0reg_data3_31_0__17_; 
wire bus_sync_rdata__0reg_data3_31_0__18_; 
wire bus_sync_rdata__0reg_data3_31_0__19_; 
wire bus_sync_rdata__0reg_data3_31_0__1_; 
wire bus_sync_rdata__0reg_data3_31_0__20_; 
wire bus_sync_rdata__0reg_data3_31_0__21_; 
wire bus_sync_rdata__0reg_data3_31_0__22_; 
wire bus_sync_rdata__0reg_data3_31_0__23_; 
wire bus_sync_rdata__0reg_data3_31_0__24_; 
wire bus_sync_rdata__0reg_data3_31_0__25_; 
wire bus_sync_rdata__0reg_data3_31_0__26_; 
wire bus_sync_rdata__0reg_data3_31_0__27_; 
wire bus_sync_rdata__0reg_data3_31_0__28_; 
wire bus_sync_rdata__0reg_data3_31_0__29_; 
wire bus_sync_rdata__0reg_data3_31_0__2_; 
wire bus_sync_rdata__0reg_data3_31_0__30_; 
wire bus_sync_rdata__0reg_data3_31_0__31_; 
wire bus_sync_rdata__0reg_data3_31_0__3_; 
wire bus_sync_rdata__0reg_data3_31_0__4_; 
wire bus_sync_rdata__0reg_data3_31_0__5_; 
wire bus_sync_rdata__0reg_data3_31_0__6_; 
wire bus_sync_rdata__0reg_data3_31_0__7_; 
wire bus_sync_rdata__0reg_data3_31_0__8_; 
wire bus_sync_rdata__0reg_data3_31_0__9_; 
wire bus_sync_rdata__abc_3653_new_n265_; 
wire bus_sync_rdata__abc_3653_new_n266_; 
wire bus_sync_rdata__abc_3653_new_n267_; 
wire bus_sync_rdata__abc_3653_new_n268_; 
wire bus_sync_rdata__abc_3653_new_n270_; 
wire bus_sync_rdata__abc_3653_new_n271_; 
wire bus_sync_rdata__abc_3653_new_n272_; 
wire bus_sync_rdata__abc_3653_new_n274_; 
wire bus_sync_rdata__abc_3653_new_n275_; 
wire bus_sync_rdata__abc_3653_new_n276_; 
wire bus_sync_rdata__abc_3653_new_n278_; 
wire bus_sync_rdata__abc_3653_new_n279_; 
wire bus_sync_rdata__abc_3653_new_n280_; 
wire bus_sync_rdata__abc_3653_new_n282_; 
wire bus_sync_rdata__abc_3653_new_n283_; 
wire bus_sync_rdata__abc_3653_new_n284_; 
wire bus_sync_rdata__abc_3653_new_n286_; 
wire bus_sync_rdata__abc_3653_new_n287_; 
wire bus_sync_rdata__abc_3653_new_n288_; 
wire bus_sync_rdata__abc_3653_new_n290_; 
wire bus_sync_rdata__abc_3653_new_n291_; 
wire bus_sync_rdata__abc_3653_new_n292_; 
wire bus_sync_rdata__abc_3653_new_n294_; 
wire bus_sync_rdata__abc_3653_new_n295_; 
wire bus_sync_rdata__abc_3653_new_n296_; 
wire bus_sync_rdata__abc_3653_new_n298_; 
wire bus_sync_rdata__abc_3653_new_n299_; 
wire bus_sync_rdata__abc_3653_new_n300_; 
wire bus_sync_rdata__abc_3653_new_n302_; 
wire bus_sync_rdata__abc_3653_new_n303_; 
wire bus_sync_rdata__abc_3653_new_n304_; 
wire bus_sync_rdata__abc_3653_new_n306_; 
wire bus_sync_rdata__abc_3653_new_n307_; 
wire bus_sync_rdata__abc_3653_new_n308_; 
wire bus_sync_rdata__abc_3653_new_n310_; 
wire bus_sync_rdata__abc_3653_new_n311_; 
wire bus_sync_rdata__abc_3653_new_n312_; 
wire bus_sync_rdata__abc_3653_new_n314_; 
wire bus_sync_rdata__abc_3653_new_n315_; 
wire bus_sync_rdata__abc_3653_new_n316_; 
wire bus_sync_rdata__abc_3653_new_n318_; 
wire bus_sync_rdata__abc_3653_new_n319_; 
wire bus_sync_rdata__abc_3653_new_n320_; 
wire bus_sync_rdata__abc_3653_new_n322_; 
wire bus_sync_rdata__abc_3653_new_n323_; 
wire bus_sync_rdata__abc_3653_new_n324_; 
wire bus_sync_rdata__abc_3653_new_n326_; 
wire bus_sync_rdata__abc_3653_new_n327_; 
wire bus_sync_rdata__abc_3653_new_n328_; 
wire bus_sync_rdata__abc_3653_new_n330_; 
wire bus_sync_rdata__abc_3653_new_n331_; 
wire bus_sync_rdata__abc_3653_new_n332_; 
wire bus_sync_rdata__abc_3653_new_n334_; 
wire bus_sync_rdata__abc_3653_new_n335_; 
wire bus_sync_rdata__abc_3653_new_n336_; 
wire bus_sync_rdata__abc_3653_new_n338_; 
wire bus_sync_rdata__abc_3653_new_n339_; 
wire bus_sync_rdata__abc_3653_new_n340_; 
wire bus_sync_rdata__abc_3653_new_n342_; 
wire bus_sync_rdata__abc_3653_new_n343_; 
wire bus_sync_rdata__abc_3653_new_n344_; 
wire bus_sync_rdata__abc_3653_new_n346_; 
wire bus_sync_rdata__abc_3653_new_n347_; 
wire bus_sync_rdata__abc_3653_new_n348_; 
wire bus_sync_rdata__abc_3653_new_n350_; 
wire bus_sync_rdata__abc_3653_new_n351_; 
wire bus_sync_rdata__abc_3653_new_n352_; 
wire bus_sync_rdata__abc_3653_new_n354_; 
wire bus_sync_rdata__abc_3653_new_n355_; 
wire bus_sync_rdata__abc_3653_new_n356_; 
wire bus_sync_rdata__abc_3653_new_n358_; 
wire bus_sync_rdata__abc_3653_new_n359_; 
wire bus_sync_rdata__abc_3653_new_n360_; 
wire bus_sync_rdata__abc_3653_new_n362_; 
wire bus_sync_rdata__abc_3653_new_n363_; 
wire bus_sync_rdata__abc_3653_new_n364_; 
wire bus_sync_rdata__abc_3653_new_n366_; 
wire bus_sync_rdata__abc_3653_new_n367_; 
wire bus_sync_rdata__abc_3653_new_n368_; 
wire bus_sync_rdata__abc_3653_new_n370_; 
wire bus_sync_rdata__abc_3653_new_n371_; 
wire bus_sync_rdata__abc_3653_new_n372_; 
wire bus_sync_rdata__abc_3653_new_n374_; 
wire bus_sync_rdata__abc_3653_new_n375_; 
wire bus_sync_rdata__abc_3653_new_n376_; 
wire bus_sync_rdata__abc_3653_new_n378_; 
wire bus_sync_rdata__abc_3653_new_n379_; 
wire bus_sync_rdata__abc_3653_new_n380_; 
wire bus_sync_rdata__abc_3653_new_n382_; 
wire bus_sync_rdata__abc_3653_new_n383_; 
wire bus_sync_rdata__abc_3653_new_n384_; 
wire bus_sync_rdata__abc_3653_new_n386_; 
wire bus_sync_rdata__abc_3653_new_n387_; 
wire bus_sync_rdata__abc_3653_new_n388_; 
wire bus_sync_rdata__abc_3653_new_n390_; 
wire bus_sync_rdata__abc_3653_new_n391_; 
wire bus_sync_rdata__abc_3653_new_n392_; 
wire bus_sync_rdata_data_in_0_; 
wire bus_sync_rdata_data_in_10_; 
wire bus_sync_rdata_data_in_11_; 
wire bus_sync_rdata_data_in_12_; 
wire bus_sync_rdata_data_in_13_; 
wire bus_sync_rdata_data_in_14_; 
wire bus_sync_rdata_data_in_15_; 
wire bus_sync_rdata_data_in_16_; 
wire bus_sync_rdata_data_in_17_; 
wire bus_sync_rdata_data_in_18_; 
wire bus_sync_rdata_data_in_19_; 
wire bus_sync_rdata_data_in_1_; 
wire bus_sync_rdata_data_in_20_; 
wire bus_sync_rdata_data_in_21_; 
wire bus_sync_rdata_data_in_22_; 
wire bus_sync_rdata_data_in_23_; 
wire bus_sync_rdata_data_in_24_; 
wire bus_sync_rdata_data_in_25_; 
wire bus_sync_rdata_data_in_26_; 
wire bus_sync_rdata_data_in_27_; 
wire bus_sync_rdata_data_in_28_; 
wire bus_sync_rdata_data_in_29_; 
wire bus_sync_rdata_data_in_2_; 
wire bus_sync_rdata_data_in_30_; 
wire bus_sync_rdata_data_in_31_; 
wire bus_sync_rdata_data_in_3_; 
wire bus_sync_rdata_data_in_4_; 
wire bus_sync_rdata_data_in_5_; 
wire bus_sync_rdata_data_in_6_; 
wire bus_sync_rdata_data_in_7_; 
wire bus_sync_rdata_data_in_8_; 
wire bus_sync_rdata_data_in_9_; 
wire bus_sync_rdata_data_out_0_; 
wire bus_sync_rdata_data_out_10_; 
wire bus_sync_rdata_data_out_11_; 
wire bus_sync_rdata_data_out_12_; 
wire bus_sync_rdata_data_out_13_; 
wire bus_sync_rdata_data_out_14_; 
wire bus_sync_rdata_data_out_15_; 
wire bus_sync_rdata_data_out_16_; 
wire bus_sync_rdata_data_out_17_; 
wire bus_sync_rdata_data_out_18_; 
wire bus_sync_rdata_data_out_19_; 
wire bus_sync_rdata_data_out_1_; 
wire bus_sync_rdata_data_out_20_; 
wire bus_sync_rdata_data_out_21_; 
wire bus_sync_rdata_data_out_22_; 
wire bus_sync_rdata_data_out_23_; 
wire bus_sync_rdata_data_out_24_; 
wire bus_sync_rdata_data_out_25_; 
wire bus_sync_rdata_data_out_26_; 
wire bus_sync_rdata_data_out_27_; 
wire bus_sync_rdata_data_out_28_; 
wire bus_sync_rdata_data_out_29_; 
wire bus_sync_rdata_data_out_2_; 
wire bus_sync_rdata_data_out_30_; 
wire bus_sync_rdata_data_out_31_; 
wire bus_sync_rdata_data_out_3_; 
wire bus_sync_rdata_data_out_4_; 
wire bus_sync_rdata_data_out_5_; 
wire bus_sync_rdata_data_out_6_; 
wire bus_sync_rdata_data_out_7_; 
wire bus_sync_rdata_data_out_8_; 
wire bus_sync_rdata_data_out_9_; 
wire bus_sync_rdata_reg_data1_0_; 
wire bus_sync_rdata_reg_data1_10_; 
wire bus_sync_rdata_reg_data1_11_; 
wire bus_sync_rdata_reg_data1_12_; 
wire bus_sync_rdata_reg_data1_13_; 
wire bus_sync_rdata_reg_data1_14_; 
wire bus_sync_rdata_reg_data1_15_; 
wire bus_sync_rdata_reg_data1_16_; 
wire bus_sync_rdata_reg_data1_17_; 
wire bus_sync_rdata_reg_data1_18_; 
wire bus_sync_rdata_reg_data1_19_; 
wire bus_sync_rdata_reg_data1_1_; 
wire bus_sync_rdata_reg_data1_20_; 
wire bus_sync_rdata_reg_data1_21_; 
wire bus_sync_rdata_reg_data1_22_; 
wire bus_sync_rdata_reg_data1_23_; 
wire bus_sync_rdata_reg_data1_24_; 
wire bus_sync_rdata_reg_data1_25_; 
wire bus_sync_rdata_reg_data1_26_; 
wire bus_sync_rdata_reg_data1_27_; 
wire bus_sync_rdata_reg_data1_28_; 
wire bus_sync_rdata_reg_data1_29_; 
wire bus_sync_rdata_reg_data1_2_; 
wire bus_sync_rdata_reg_data1_30_; 
wire bus_sync_rdata_reg_data1_31_; 
wire bus_sync_rdata_reg_data1_3_; 
wire bus_sync_rdata_reg_data1_4_; 
wire bus_sync_rdata_reg_data1_5_; 
wire bus_sync_rdata_reg_data1_6_; 
wire bus_sync_rdata_reg_data1_7_; 
wire bus_sync_rdata_reg_data1_8_; 
wire bus_sync_rdata_reg_data1_9_; 
wire bus_sync_rdata_reg_data2_0_; 
wire bus_sync_rdata_reg_data2_10_; 
wire bus_sync_rdata_reg_data2_11_; 
wire bus_sync_rdata_reg_data2_12_; 
wire bus_sync_rdata_reg_data2_13_; 
wire bus_sync_rdata_reg_data2_14_; 
wire bus_sync_rdata_reg_data2_15_; 
wire bus_sync_rdata_reg_data2_16_; 
wire bus_sync_rdata_reg_data2_17_; 
wire bus_sync_rdata_reg_data2_18_; 
wire bus_sync_rdata_reg_data2_19_; 
wire bus_sync_rdata_reg_data2_1_; 
wire bus_sync_rdata_reg_data2_20_; 
wire bus_sync_rdata_reg_data2_21_; 
wire bus_sync_rdata_reg_data2_22_; 
wire bus_sync_rdata_reg_data2_23_; 
wire bus_sync_rdata_reg_data2_24_; 
wire bus_sync_rdata_reg_data2_25_; 
wire bus_sync_rdata_reg_data2_26_; 
wire bus_sync_rdata_reg_data2_27_; 
wire bus_sync_rdata_reg_data2_28_; 
wire bus_sync_rdata_reg_data2_29_; 
wire bus_sync_rdata_reg_data2_2_; 
wire bus_sync_rdata_reg_data2_30_; 
wire bus_sync_rdata_reg_data2_31_; 
wire bus_sync_rdata_reg_data2_3_; 
wire bus_sync_rdata_reg_data2_4_; 
wire bus_sync_rdata_reg_data2_5_; 
wire bus_sync_rdata_reg_data2_6_; 
wire bus_sync_rdata_reg_data2_7_; 
wire bus_sync_rdata_reg_data2_8_; 
wire bus_sync_rdata_reg_data2_9_; 
wire bus_sync_state_machine_ECLK1; 
wire bus_sync_state_machine_EECLK1; 
wire bus_sync_state_machine_NCLK2; 
wire bus_sync_state_machine__0ECLK1_0_0_; 
wire bus_sync_state_machine__0EECLK1_0_0_; 
wire bus_sync_state_machine__0reg_data1_3_0__0_; 
wire bus_sync_state_machine__0reg_data1_3_0__1_; 
wire bus_sync_state_machine__0reg_data1_3_0__2_; 
wire bus_sync_state_machine__0reg_data1_3_0__3_; 
wire bus_sync_state_machine__0reg_data2_3_0__0_; 
wire bus_sync_state_machine__0reg_data2_3_0__1_; 
wire bus_sync_state_machine__0reg_data2_3_0__2_; 
wire bus_sync_state_machine__0reg_data2_3_0__3_; 
wire bus_sync_state_machine__0reg_data3_3_0__0_; 
wire bus_sync_state_machine__0reg_data3_3_0__1_; 
wire bus_sync_state_machine__0reg_data3_3_0__2_; 
wire bus_sync_state_machine__0reg_data3_3_0__3_; 
wire bus_sync_state_machine__abc_3850_new_n33_; 
wire bus_sync_state_machine__abc_3850_new_n34_; 
wire bus_sync_state_machine__abc_3850_new_n35_; 
wire bus_sync_state_machine__abc_3850_new_n36_; 
wire bus_sync_state_machine__abc_3850_new_n38_; 
wire bus_sync_state_machine__abc_3850_new_n39_; 
wire bus_sync_state_machine__abc_3850_new_n40_; 
wire bus_sync_state_machine__abc_3850_new_n42_; 
wire bus_sync_state_machine__abc_3850_new_n43_; 
wire bus_sync_state_machine__abc_3850_new_n44_; 
wire bus_sync_state_machine__abc_3850_new_n46_; 
wire bus_sync_state_machine__abc_3850_new_n47_; 
wire bus_sync_state_machine__abc_3850_new_n48_; 
wire bus_sync_state_machine_reg_data1_0_; 
wire bus_sync_state_machine_reg_data1_1_; 
wire bus_sync_state_machine_reg_data1_2_; 
wire bus_sync_state_machine_reg_data1_3_; 
wire bus_sync_state_machine_reg_data2_0_; 
wire bus_sync_state_machine_reg_data2_1_; 
wire bus_sync_state_machine_reg_data2_2_; 
wire bus_sync_state_machine_reg_data2_3_; 
wire bus_sync_status_ECLK2; 
wire bus_sync_status_EECLK2; 
wire bus_sync_status_NCLK1; 
wire bus_sync_status__0ECLK2_0_0_; 
wire bus_sync_status__0EECLK2_0_0_; 
wire bus_sync_status__0reg_data1_2_0__0_; 
wire bus_sync_status__0reg_data1_2_0__1_; 
wire bus_sync_status__0reg_data1_2_0__2_; 
wire bus_sync_status__0reg_data2_2_0__0_; 
wire bus_sync_status__0reg_data2_2_0__1_; 
wire bus_sync_status__0reg_data2_2_0__2_; 
wire bus_sync_status__0reg_data3_2_0__0_; 
wire bus_sync_status__0reg_data3_2_0__1_; 
wire bus_sync_status__0reg_data3_2_0__2_; 
wire bus_sync_status__abc_3630_new_n27_; 
wire bus_sync_status__abc_3630_new_n28_; 
wire bus_sync_status__abc_3630_new_n29_; 
wire bus_sync_status__abc_3630_new_n30_; 
wire bus_sync_status__abc_3630_new_n32_; 
wire bus_sync_status__abc_3630_new_n33_; 
wire bus_sync_status__abc_3630_new_n34_; 
wire bus_sync_status__abc_3630_new_n36_; 
wire bus_sync_status__abc_3630_new_n37_; 
wire bus_sync_status__abc_3630_new_n38_; 
wire bus_sync_status_data_out_0_; 
wire bus_sync_status_data_out_1_; 
wire bus_sync_status_data_out_2_; 
wire bus_sync_status_reg_data1_0_; 
wire bus_sync_status_reg_data1_1_; 
wire bus_sync_status_reg_data1_2_; 
wire bus_sync_status_reg_data2_0_; 
wire bus_sync_status_reg_data2_1_; 
wire bus_sync_status_reg_data2_2_; 
wire busy; 
wire counter_0_; 
wire counter_10_; 
wire counter_11_; 
wire counter_12_; 
wire counter_13_; 
wire counter_14_; 
wire counter_15_; 
wire counter_16_; 
wire counter_17_; 
wire counter_18_; 
wire counter_19_; 
wire counter_1_; 
wire counter_20_; 
wire counter_21_; 
wire counter_22_; 
wire counter_23_; 
wire counter_24_; 
wire counter_25_; 
wire counter_26_; 
wire counter_27_; 
wire counter_28_; 
wire counter_29_; 
wire counter_2_; 
wire counter_30_; 
wire counter_31_; 
wire counter_32_; 
wire counter_33_; 
wire counter_34_; 
wire counter_35_; 
wire counter_36_; 
wire counter_37_; 
wire counter_38_; 
wire counter_39_; 
wire counter_3_; 
wire counter_40_; 
wire counter_41_; 
wire counter_42_; 
wire counter_43_; 
wire counter_44_; 
wire counter_45_; 
wire counter_46_; 
wire counter_47_; 
wire counter_48_; 
wire counter_49_; 
wire counter_4_; 
wire counter_50_; 
wire counter_51_; 
wire counter_52_; 
wire counter_53_; 
wire counter_54_; 
wire counter_55_; 
wire counter_56_; 
wire counter_57_; 
wire counter_58_; 
wire counter_59_; 
wire counter_5_; 
wire counter_60_; 
wire counter_61_; 
wire counter_62_; 
wire counter_63_; 
wire counter_64_; 
wire counter_65_; 
wire counter_6_; 
wire counter_7_; 
wire counter_8_; 
wire counter_9_; 
wire fini_spi; 
wire fini_spi_clk; 
wire re; 
wire re_clk; 
wire sft_reg_0_; 
wire sft_reg_10_; 
wire sft_reg_11_; 
wire sft_reg_12_; 
wire sft_reg_13_; 
wire sft_reg_14_; 
wire sft_reg_15_; 
wire sft_reg_16_; 
wire sft_reg_17_; 
wire sft_reg_18_; 
wire sft_reg_19_; 
wire sft_reg_1_; 
wire sft_reg_20_; 
wire sft_reg_21_; 
wire sft_reg_22_; 
wire sft_reg_23_; 
wire sft_reg_24_; 
wire sft_reg_25_; 
wire sft_reg_26_; 
wire sft_reg_27_; 
wire sft_reg_28_; 
wire sft_reg_29_; 
wire sft_reg_2_; 
wire sft_reg_30_; 
wire sft_reg_3_; 
wire sft_reg_4_; 
wire sft_reg_5_; 
wire sft_reg_6_; 
wire sft_reg_7_; 
wire sft_reg_8_; 
wire sft_reg_9_; 
wire state_0_; 
wire state_1_; 
wire state_3_; 
wire state_4_; 
wire state_5_; 
wire state_6_; 
wire state_7_; 
wire we; 
wire we_clk; 
AND2X2 AND2X2_1 ( .A(state_3_), .B(RST), .Y(_abc_4268_new_n558_));
AND2X2 AND2X2_10 ( .A(RST), .B(state_6_), .Y(_abc_4268_new_n576_));
AND2X2 AND2X2_100 ( .A(_abc_4268_new_n794_), .B(_abc_4268_new_n795_), .Y(_abc_4268_new_n796_));
AND2X2 AND2X2_1000 ( .A(bus_sync_rdata__abc_3653_new_n312_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__11_));
AND2X2 AND2X2_1001 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_12_), .Y(bus_sync_rdata__abc_3653_new_n314_));
AND2X2 AND2X2_1002 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_12_), .Y(bus_sync_rdata__abc_3653_new_n315_));
AND2X2 AND2X2_1003 ( .A(bus_sync_rdata__abc_3653_new_n316_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__12_));
AND2X2 AND2X2_1004 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_13_), .Y(bus_sync_rdata__abc_3653_new_n318_));
AND2X2 AND2X2_1005 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_13_), .Y(bus_sync_rdata__abc_3653_new_n319_));
AND2X2 AND2X2_1006 ( .A(bus_sync_rdata__abc_3653_new_n320_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__13_));
AND2X2 AND2X2_1007 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_14_), .Y(bus_sync_rdata__abc_3653_new_n322_));
AND2X2 AND2X2_1008 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_14_), .Y(bus_sync_rdata__abc_3653_new_n323_));
AND2X2 AND2X2_1009 ( .A(bus_sync_rdata__abc_3653_new_n324_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__14_));
AND2X2 AND2X2_101 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_12_), .Y(_abc_4268_new_n798_));
AND2X2 AND2X2_1010 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_15_), .Y(bus_sync_rdata__abc_3653_new_n326_));
AND2X2 AND2X2_1011 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_15_), .Y(bus_sync_rdata__abc_3653_new_n327_));
AND2X2 AND2X2_1012 ( .A(bus_sync_rdata__abc_3653_new_n328_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__15_));
AND2X2 AND2X2_1013 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_16_), .Y(bus_sync_rdata__abc_3653_new_n330_));
AND2X2 AND2X2_1014 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_16_), .Y(bus_sync_rdata__abc_3653_new_n331_));
AND2X2 AND2X2_1015 ( .A(bus_sync_rdata__abc_3653_new_n332_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__16_));
AND2X2 AND2X2_1016 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_17_), .Y(bus_sync_rdata__abc_3653_new_n334_));
AND2X2 AND2X2_1017 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_17_), .Y(bus_sync_rdata__abc_3653_new_n335_));
AND2X2 AND2X2_1018 ( .A(bus_sync_rdata__abc_3653_new_n336_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__17_));
AND2X2 AND2X2_1019 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_18_), .Y(bus_sync_rdata__abc_3653_new_n338_));
AND2X2 AND2X2_102 ( .A(_abc_4268_new_n799_), .B(RST), .Y(_abc_4268_new_n800_));
AND2X2 AND2X2_1020 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_18_), .Y(bus_sync_rdata__abc_3653_new_n339_));
AND2X2 AND2X2_1021 ( .A(bus_sync_rdata__abc_3653_new_n340_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__18_));
AND2X2 AND2X2_1022 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_19_), .Y(bus_sync_rdata__abc_3653_new_n342_));
AND2X2 AND2X2_1023 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_19_), .Y(bus_sync_rdata__abc_3653_new_n343_));
AND2X2 AND2X2_1024 ( .A(bus_sync_rdata__abc_3653_new_n344_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__19_));
AND2X2 AND2X2_1025 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_20_), .Y(bus_sync_rdata__abc_3653_new_n346_));
AND2X2 AND2X2_1026 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_20_), .Y(bus_sync_rdata__abc_3653_new_n347_));
AND2X2 AND2X2_1027 ( .A(bus_sync_rdata__abc_3653_new_n348_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__20_));
AND2X2 AND2X2_1028 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_21_), .Y(bus_sync_rdata__abc_3653_new_n350_));
AND2X2 AND2X2_1029 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_21_), .Y(bus_sync_rdata__abc_3653_new_n351_));
AND2X2 AND2X2_103 ( .A(_abc_4268_new_n797_), .B(_abc_4268_new_n800_), .Y(_0bus_cap_31_0__12_));
AND2X2 AND2X2_1030 ( .A(bus_sync_rdata__abc_3653_new_n352_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__21_));
AND2X2 AND2X2_1031 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_22_), .Y(bus_sync_rdata__abc_3653_new_n354_));
AND2X2 AND2X2_1032 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_22_), .Y(bus_sync_rdata__abc_3653_new_n355_));
AND2X2 AND2X2_1033 ( .A(bus_sync_rdata__abc_3653_new_n356_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__22_));
AND2X2 AND2X2_1034 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_23_), .Y(bus_sync_rdata__abc_3653_new_n358_));
AND2X2 AND2X2_1035 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_23_), .Y(bus_sync_rdata__abc_3653_new_n359_));
AND2X2 AND2X2_1036 ( .A(bus_sync_rdata__abc_3653_new_n360_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__23_));
AND2X2 AND2X2_1037 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_24_), .Y(bus_sync_rdata__abc_3653_new_n362_));
AND2X2 AND2X2_1038 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_24_), .Y(bus_sync_rdata__abc_3653_new_n363_));
AND2X2 AND2X2_1039 ( .A(bus_sync_rdata__abc_3653_new_n364_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__24_));
AND2X2 AND2X2_104 ( .A(_abc_4268_new_n802_), .B(_abc_4268_new_n803_), .Y(_abc_4268_new_n804_));
AND2X2 AND2X2_1040 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_25_), .Y(bus_sync_rdata__abc_3653_new_n366_));
AND2X2 AND2X2_1041 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_25_), .Y(bus_sync_rdata__abc_3653_new_n367_));
AND2X2 AND2X2_1042 ( .A(bus_sync_rdata__abc_3653_new_n368_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__25_));
AND2X2 AND2X2_1043 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_26_), .Y(bus_sync_rdata__abc_3653_new_n370_));
AND2X2 AND2X2_1044 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_26_), .Y(bus_sync_rdata__abc_3653_new_n371_));
AND2X2 AND2X2_1045 ( .A(bus_sync_rdata__abc_3653_new_n372_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__26_));
AND2X2 AND2X2_1046 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_27_), .Y(bus_sync_rdata__abc_3653_new_n374_));
AND2X2 AND2X2_1047 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_27_), .Y(bus_sync_rdata__abc_3653_new_n375_));
AND2X2 AND2X2_1048 ( .A(bus_sync_rdata__abc_3653_new_n376_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__27_));
AND2X2 AND2X2_1049 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_28_), .Y(bus_sync_rdata__abc_3653_new_n378_));
AND2X2 AND2X2_105 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_13_), .Y(_abc_4268_new_n806_));
AND2X2 AND2X2_1050 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_28_), .Y(bus_sync_rdata__abc_3653_new_n379_));
AND2X2 AND2X2_1051 ( .A(bus_sync_rdata__abc_3653_new_n380_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__28_));
AND2X2 AND2X2_1052 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_29_), .Y(bus_sync_rdata__abc_3653_new_n382_));
AND2X2 AND2X2_1053 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_29_), .Y(bus_sync_rdata__abc_3653_new_n383_));
AND2X2 AND2X2_1054 ( .A(bus_sync_rdata__abc_3653_new_n384_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__29_));
AND2X2 AND2X2_1055 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_30_), .Y(bus_sync_rdata__abc_3653_new_n386_));
AND2X2 AND2X2_1056 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_30_), .Y(bus_sync_rdata__abc_3653_new_n387_));
AND2X2 AND2X2_1057 ( .A(bus_sync_rdata__abc_3653_new_n388_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__30_));
AND2X2 AND2X2_1058 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_31_), .Y(bus_sync_rdata__abc_3653_new_n390_));
AND2X2 AND2X2_1059 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_31_), .Y(bus_sync_rdata__abc_3653_new_n391_));
AND2X2 AND2X2_106 ( .A(_abc_4268_new_n807_), .B(RST), .Y(_abc_4268_new_n808_));
AND2X2 AND2X2_1060 ( .A(bus_sync_rdata__abc_3653_new_n392_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__31_));
AND2X2 AND2X2_1061 ( .A(RST), .B(SCLK), .Y(bus_sync_rdata__0ECLK2_0_0_));
AND2X2 AND2X2_1062 ( .A(RST), .B(bus_sync_rdata_ECLK2), .Y(bus_sync_rdata__0EECLK2_0_0_));
AND2X2 AND2X2_1063 ( .A(bus_sync_state_machine__abc_3850_new_n33_), .B(bus_sync_state_machine_reg_data2_0_), .Y(bus_sync_state_machine__abc_3850_new_n34_));
AND2X2 AND2X2_1064 ( .A(bus_sync_state_machine_reg_data1_0_), .B(bus_sync_state_machine_EECLK1), .Y(bus_sync_state_machine__abc_3850_new_n35_));
AND2X2 AND2X2_1065 ( .A(bus_sync_state_machine__abc_3850_new_n36_), .B(RST), .Y(bus_sync_state_machine__0reg_data2_3_0__0_));
AND2X2 AND2X2_1066 ( .A(bus_sync_state_machine__abc_3850_new_n33_), .B(bus_sync_state_machine_reg_data2_1_), .Y(bus_sync_state_machine__abc_3850_new_n38_));
AND2X2 AND2X2_1067 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_1_), .Y(bus_sync_state_machine__abc_3850_new_n39_));
AND2X2 AND2X2_1068 ( .A(bus_sync_state_machine__abc_3850_new_n40_), .B(RST), .Y(bus_sync_state_machine__0reg_data2_3_0__1_));
AND2X2 AND2X2_1069 ( .A(bus_sync_state_machine__abc_3850_new_n33_), .B(bus_sync_state_machine_reg_data2_2_), .Y(bus_sync_state_machine__abc_3850_new_n42_));
AND2X2 AND2X2_107 ( .A(_abc_4268_new_n805_), .B(_abc_4268_new_n808_), .Y(_0bus_cap_31_0__13_));
AND2X2 AND2X2_1070 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_2_), .Y(bus_sync_state_machine__abc_3850_new_n43_));
AND2X2 AND2X2_1071 ( .A(bus_sync_state_machine__abc_3850_new_n44_), .B(RST), .Y(bus_sync_state_machine__0reg_data2_3_0__2_));
AND2X2 AND2X2_1072 ( .A(bus_sync_state_machine__abc_3850_new_n33_), .B(bus_sync_state_machine_reg_data2_3_), .Y(bus_sync_state_machine__abc_3850_new_n46_));
AND2X2 AND2X2_1073 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_3_), .Y(bus_sync_state_machine__abc_3850_new_n47_));
AND2X2 AND2X2_1074 ( .A(bus_sync_state_machine__abc_3850_new_n48_), .B(RST), .Y(bus_sync_state_machine__0reg_data2_3_0__3_));
AND2X2 AND2X2_1075 ( .A(RST), .B(bus_sync_state_machine_reg_data2_0_), .Y(bus_sync_state_machine__0reg_data3_3_0__0_));
AND2X2 AND2X2_1076 ( .A(RST), .B(bus_sync_state_machine_reg_data2_1_), .Y(bus_sync_state_machine__0reg_data3_3_0__1_));
AND2X2 AND2X2_1077 ( .A(RST), .B(bus_sync_state_machine_reg_data2_2_), .Y(bus_sync_state_machine__0reg_data3_3_0__2_));
AND2X2 AND2X2_1078 ( .A(RST), .B(bus_sync_state_machine_reg_data2_3_), .Y(bus_sync_state_machine__0reg_data3_3_0__3_));
AND2X2 AND2X2_1079 ( .A(RST), .B(fini_spi), .Y(bus_sync_state_machine__0reg_data1_3_0__0_));
AND2X2 AND2X2_108 ( .A(_abc_4268_new_n810_), .B(_abc_4268_new_n811_), .Y(_abc_4268_new_n812_));
AND2X2 AND2X2_1080 ( .A(RST), .B(re), .Y(bus_sync_state_machine__0reg_data1_3_0__1_));
AND2X2 AND2X2_1081 ( .A(RST), .B(we), .Y(bus_sync_state_machine__0reg_data1_3_0__2_));
AND2X2 AND2X2_1082 ( .A(RST), .B(PICORV_RST_SPI), .Y(bus_sync_state_machine__0reg_data1_3_0__3_));
AND2X2 AND2X2_1083 ( .A(RST), .B(SCLK), .Y(bus_sync_state_machine__0ECLK1_0_0_));
AND2X2 AND2X2_1084 ( .A(RST), .B(bus_sync_state_machine_ECLK1), .Y(bus_sync_state_machine__0EECLK1_0_0_));
AND2X2 AND2X2_1085 ( .A(bus_sync_status__abc_3630_new_n27_), .B(bus_sync_status_reg_data2_0_), .Y(bus_sync_status__abc_3630_new_n28_));
AND2X2 AND2X2_1086 ( .A(bus_sync_status_reg_data1_0_), .B(bus_sync_status_EECLK2), .Y(bus_sync_status__abc_3630_new_n29_));
AND2X2 AND2X2_1087 ( .A(bus_sync_status__abc_3630_new_n30_), .B(RST), .Y(bus_sync_status__0reg_data2_2_0__0_));
AND2X2 AND2X2_1088 ( .A(bus_sync_status__abc_3630_new_n27_), .B(bus_sync_status_reg_data2_1_), .Y(bus_sync_status__abc_3630_new_n32_));
AND2X2 AND2X2_1089 ( .A(bus_sync_status_EECLK2), .B(bus_sync_status_reg_data1_1_), .Y(bus_sync_status__abc_3630_new_n33_));
AND2X2 AND2X2_109 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_14_), .Y(_abc_4268_new_n814_));
AND2X2 AND2X2_1090 ( .A(bus_sync_status__abc_3630_new_n34_), .B(RST), .Y(bus_sync_status__0reg_data2_2_0__1_));
AND2X2 AND2X2_1091 ( .A(bus_sync_status__abc_3630_new_n27_), .B(bus_sync_status_reg_data2_2_), .Y(bus_sync_status__abc_3630_new_n36_));
AND2X2 AND2X2_1092 ( .A(bus_sync_status_EECLK2), .B(bus_sync_status_reg_data1_2_), .Y(bus_sync_status__abc_3630_new_n37_));
AND2X2 AND2X2_1093 ( .A(bus_sync_status__abc_3630_new_n38_), .B(RST), .Y(bus_sync_status__0reg_data2_2_0__2_));
AND2X2 AND2X2_1094 ( .A(RST), .B(bus_sync_status_reg_data2_0_), .Y(bus_sync_status__0reg_data3_2_0__0_));
AND2X2 AND2X2_1095 ( .A(RST), .B(bus_sync_status_reg_data2_1_), .Y(bus_sync_status__0reg_data3_2_0__1_));
AND2X2 AND2X2_1096 ( .A(RST), .B(bus_sync_status_reg_data2_2_), .Y(bus_sync_status__0reg_data3_2_0__2_));
AND2X2 AND2X2_1097 ( .A(RST), .B(busy), .Y(bus_sync_status__0reg_data1_2_0__0_));
AND2X2 AND2X2_1098 ( .A(RST), .B(axi_awvalid), .Y(bus_sync_status__0reg_data1_2_0__1_));
AND2X2 AND2X2_1099 ( .A(RST), .B(axi_arvalid), .Y(bus_sync_status__0reg_data1_2_0__2_));
AND2X2 AND2X2_11 ( .A(_abc_4268_new_n576_), .B(_abc_4268_new_n575_), .Y(_abc_4268_new_n577_));
AND2X2 AND2X2_110 ( .A(_abc_4268_new_n815_), .B(RST), .Y(_abc_4268_new_n816_));
AND2X2 AND2X2_1100 ( .A(RST), .B(bus_sync_status_ECLK2), .Y(bus_sync_status__0EECLK2_0_0_));
AND2X2 AND2X2_1101 ( .A(RST), .B(SCLK), .Y(bus_sync_status__0ECLK2_0_0_));
AND2X2 AND2X2_111 ( .A(_abc_4268_new_n813_), .B(_abc_4268_new_n816_), .Y(_0bus_cap_31_0__14_));
AND2X2 AND2X2_112 ( .A(_abc_4268_new_n818_), .B(_abc_4268_new_n819_), .Y(_abc_4268_new_n820_));
AND2X2 AND2X2_113 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_15_), .Y(_abc_4268_new_n822_));
AND2X2 AND2X2_114 ( .A(_abc_4268_new_n823_), .B(RST), .Y(_abc_4268_new_n824_));
AND2X2 AND2X2_115 ( .A(_abc_4268_new_n821_), .B(_abc_4268_new_n824_), .Y(_0bus_cap_31_0__15_));
AND2X2 AND2X2_116 ( .A(_abc_4268_new_n826_), .B(_abc_4268_new_n827_), .Y(_abc_4268_new_n828_));
AND2X2 AND2X2_117 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_16_), .Y(_abc_4268_new_n830_));
AND2X2 AND2X2_118 ( .A(_abc_4268_new_n831_), .B(RST), .Y(_abc_4268_new_n832_));
AND2X2 AND2X2_119 ( .A(_abc_4268_new_n829_), .B(_abc_4268_new_n832_), .Y(_0bus_cap_31_0__16_));
AND2X2 AND2X2_12 ( .A(fini_spi_clk), .B(we_clk), .Y(_abc_4268_new_n579_));
AND2X2 AND2X2_120 ( .A(_abc_4268_new_n834_), .B(_abc_4268_new_n835_), .Y(_abc_4268_new_n836_));
AND2X2 AND2X2_121 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_17_), .Y(_abc_4268_new_n838_));
AND2X2 AND2X2_122 ( .A(_abc_4268_new_n839_), .B(RST), .Y(_abc_4268_new_n840_));
AND2X2 AND2X2_123 ( .A(_abc_4268_new_n837_), .B(_abc_4268_new_n840_), .Y(_0bus_cap_31_0__17_));
AND2X2 AND2X2_124 ( .A(_abc_4268_new_n842_), .B(_abc_4268_new_n843_), .Y(_abc_4268_new_n844_));
AND2X2 AND2X2_125 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_18_), .Y(_abc_4268_new_n846_));
AND2X2 AND2X2_126 ( .A(_abc_4268_new_n847_), .B(RST), .Y(_abc_4268_new_n848_));
AND2X2 AND2X2_127 ( .A(_abc_4268_new_n845_), .B(_abc_4268_new_n848_), .Y(_0bus_cap_31_0__18_));
AND2X2 AND2X2_128 ( .A(_abc_4268_new_n850_), .B(_abc_4268_new_n851_), .Y(_abc_4268_new_n852_));
AND2X2 AND2X2_129 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_19_), .Y(_abc_4268_new_n854_));
AND2X2 AND2X2_13 ( .A(_abc_4268_new_n579_), .B(_abc_4268_new_n578_), .Y(_abc_4268_new_n580_));
AND2X2 AND2X2_130 ( .A(_abc_4268_new_n855_), .B(RST), .Y(_abc_4268_new_n856_));
AND2X2 AND2X2_131 ( .A(_abc_4268_new_n853_), .B(_abc_4268_new_n856_), .Y(_0bus_cap_31_0__19_));
AND2X2 AND2X2_132 ( .A(_abc_4268_new_n858_), .B(_abc_4268_new_n859_), .Y(_abc_4268_new_n860_));
AND2X2 AND2X2_133 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_20_), .Y(_abc_4268_new_n862_));
AND2X2 AND2X2_134 ( .A(_abc_4268_new_n863_), .B(RST), .Y(_abc_4268_new_n864_));
AND2X2 AND2X2_135 ( .A(_abc_4268_new_n861_), .B(_abc_4268_new_n864_), .Y(_0bus_cap_31_0__20_));
AND2X2 AND2X2_136 ( .A(_abc_4268_new_n866_), .B(_abc_4268_new_n867_), .Y(_abc_4268_new_n868_));
AND2X2 AND2X2_137 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_21_), .Y(_abc_4268_new_n870_));
AND2X2 AND2X2_138 ( .A(_abc_4268_new_n871_), .B(RST), .Y(_abc_4268_new_n872_));
AND2X2 AND2X2_139 ( .A(_abc_4268_new_n869_), .B(_abc_4268_new_n872_), .Y(_0bus_cap_31_0__21_));
AND2X2 AND2X2_14 ( .A(_abc_4268_new_n581_), .B(RST), .Y(_abc_4268_new_n582_));
AND2X2 AND2X2_140 ( .A(_abc_4268_new_n874_), .B(_abc_4268_new_n875_), .Y(_abc_4268_new_n876_));
AND2X2 AND2X2_141 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_22_), .Y(_abc_4268_new_n878_));
AND2X2 AND2X2_142 ( .A(_abc_4268_new_n879_), .B(RST), .Y(_abc_4268_new_n880_));
AND2X2 AND2X2_143 ( .A(_abc_4268_new_n877_), .B(_abc_4268_new_n880_), .Y(_0bus_cap_31_0__22_));
AND2X2 AND2X2_144 ( .A(_abc_4268_new_n882_), .B(_abc_4268_new_n883_), .Y(_abc_4268_new_n884_));
AND2X2 AND2X2_145 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_23_), .Y(_abc_4268_new_n886_));
AND2X2 AND2X2_146 ( .A(_abc_4268_new_n887_), .B(RST), .Y(_abc_4268_new_n888_));
AND2X2 AND2X2_147 ( .A(_abc_4268_new_n885_), .B(_abc_4268_new_n888_), .Y(_0bus_cap_31_0__23_));
AND2X2 AND2X2_148 ( .A(_abc_4268_new_n890_), .B(_abc_4268_new_n891_), .Y(_abc_4268_new_n892_));
AND2X2 AND2X2_149 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_24_), .Y(_abc_4268_new_n894_));
AND2X2 AND2X2_15 ( .A(fini_spi_clk), .B(re_clk), .Y(_abc_4268_new_n584_));
AND2X2 AND2X2_150 ( .A(_abc_4268_new_n895_), .B(RST), .Y(_abc_4268_new_n896_));
AND2X2 AND2X2_151 ( .A(_abc_4268_new_n893_), .B(_abc_4268_new_n896_), .Y(_0bus_cap_31_0__24_));
AND2X2 AND2X2_152 ( .A(_abc_4268_new_n898_), .B(_abc_4268_new_n899_), .Y(_abc_4268_new_n900_));
AND2X2 AND2X2_153 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_25_), .Y(_abc_4268_new_n902_));
AND2X2 AND2X2_154 ( .A(_abc_4268_new_n903_), .B(RST), .Y(_abc_4268_new_n904_));
AND2X2 AND2X2_155 ( .A(_abc_4268_new_n901_), .B(_abc_4268_new_n904_), .Y(_0bus_cap_31_0__25_));
AND2X2 AND2X2_156 ( .A(_abc_4268_new_n906_), .B(_abc_4268_new_n907_), .Y(_abc_4268_new_n908_));
AND2X2 AND2X2_157 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_26_), .Y(_abc_4268_new_n910_));
AND2X2 AND2X2_158 ( .A(_abc_4268_new_n911_), .B(RST), .Y(_abc_4268_new_n912_));
AND2X2 AND2X2_159 ( .A(_abc_4268_new_n909_), .B(_abc_4268_new_n912_), .Y(_0bus_cap_31_0__26_));
AND2X2 AND2X2_16 ( .A(_abc_4268_new_n584_), .B(_abc_4268_new_n583_), .Y(_abc_4268_new_n585_));
AND2X2 AND2X2_160 ( .A(_abc_4268_new_n914_), .B(_abc_4268_new_n915_), .Y(_abc_4268_new_n916_));
AND2X2 AND2X2_161 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_27_), .Y(_abc_4268_new_n918_));
AND2X2 AND2X2_162 ( .A(_abc_4268_new_n919_), .B(RST), .Y(_abc_4268_new_n920_));
AND2X2 AND2X2_163 ( .A(_abc_4268_new_n917_), .B(_abc_4268_new_n920_), .Y(_0bus_cap_31_0__27_));
AND2X2 AND2X2_164 ( .A(_abc_4268_new_n922_), .B(_abc_4268_new_n923_), .Y(_abc_4268_new_n924_));
AND2X2 AND2X2_165 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_28_), .Y(_abc_4268_new_n926_));
AND2X2 AND2X2_166 ( .A(_abc_4268_new_n927_), .B(RST), .Y(_abc_4268_new_n928_));
AND2X2 AND2X2_167 ( .A(_abc_4268_new_n925_), .B(_abc_4268_new_n928_), .Y(_0bus_cap_31_0__28_));
AND2X2 AND2X2_168 ( .A(_abc_4268_new_n930_), .B(_abc_4268_new_n931_), .Y(_abc_4268_new_n932_));
AND2X2 AND2X2_169 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_29_), .Y(_abc_4268_new_n934_));
AND2X2 AND2X2_17 ( .A(_abc_4268_new_n585_), .B(state_0_), .Y(_abc_4268_new_n586_));
AND2X2 AND2X2_170 ( .A(_abc_4268_new_n935_), .B(RST), .Y(_abc_4268_new_n936_));
AND2X2 AND2X2_171 ( .A(_abc_4268_new_n933_), .B(_abc_4268_new_n936_), .Y(_0bus_cap_31_0__29_));
AND2X2 AND2X2_172 ( .A(_abc_4268_new_n938_), .B(_abc_4268_new_n939_), .Y(_abc_4268_new_n940_));
AND2X2 AND2X2_173 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_30_), .Y(_abc_4268_new_n942_));
AND2X2 AND2X2_174 ( .A(_abc_4268_new_n943_), .B(RST), .Y(_abc_4268_new_n944_));
AND2X2 AND2X2_175 ( .A(_abc_4268_new_n941_), .B(_abc_4268_new_n944_), .Y(_0bus_cap_31_0__30_));
AND2X2 AND2X2_176 ( .A(_abc_4268_new_n946_), .B(_abc_4268_new_n947_), .Y(_abc_4268_new_n948_));
AND2X2 AND2X2_177 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_31_), .Y(_abc_4268_new_n950_));
AND2X2 AND2X2_178 ( .A(_abc_4268_new_n951_), .B(RST), .Y(_abc_4268_new_n952_));
AND2X2 AND2X2_179 ( .A(_abc_4268_new_n949_), .B(_abc_4268_new_n952_), .Y(_0bus_cap_31_0__31_));
AND2X2 AND2X2_18 ( .A(_abc_4268_new_n582_), .B(_abc_4268_new_n586_), .Y(_abc_4268_new_n587_));
AND2X2 AND2X2_180 ( .A(axi_rready), .B(\axi_rdata[0] ), .Y(_abc_4268_new_n954_));
AND2X2 AND2X2_181 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_0_), .Y(_abc_4268_new_n956_));
AND2X2 AND2X2_182 ( .A(_abc_4268_new_n957_), .B(RST), .Y(_0rdata_31_0__0_));
AND2X2 AND2X2_183 ( .A(axi_rready), .B(\axi_rdata[1] ), .Y(_abc_4268_new_n959_));
AND2X2 AND2X2_184 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_1_), .Y(_abc_4268_new_n960_));
AND2X2 AND2X2_185 ( .A(_abc_4268_new_n961_), .B(RST), .Y(_0rdata_31_0__1_));
AND2X2 AND2X2_186 ( .A(axi_rready), .B(\axi_rdata[2] ), .Y(_abc_4268_new_n963_));
AND2X2 AND2X2_187 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_2_), .Y(_abc_4268_new_n964_));
AND2X2 AND2X2_188 ( .A(_abc_4268_new_n965_), .B(RST), .Y(_0rdata_31_0__2_));
AND2X2 AND2X2_189 ( .A(axi_rready), .B(\axi_rdata[3] ), .Y(_abc_4268_new_n967_));
AND2X2 AND2X2_19 ( .A(_abc_4268_new_n576_), .B(axi_arready), .Y(_abc_4268_new_n589_));
AND2X2 AND2X2_190 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_3_), .Y(_abc_4268_new_n968_));
AND2X2 AND2X2_191 ( .A(_abc_4268_new_n969_), .B(RST), .Y(_0rdata_31_0__3_));
AND2X2 AND2X2_192 ( .A(axi_rready), .B(\axi_rdata[4] ), .Y(_abc_4268_new_n971_));
AND2X2 AND2X2_193 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_4_), .Y(_abc_4268_new_n972_));
AND2X2 AND2X2_194 ( .A(_abc_4268_new_n973_), .B(RST), .Y(_0rdata_31_0__4_));
AND2X2 AND2X2_195 ( .A(axi_rready), .B(\axi_rdata[5] ), .Y(_abc_4268_new_n975_));
AND2X2 AND2X2_196 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_5_), .Y(_abc_4268_new_n976_));
AND2X2 AND2X2_197 ( .A(_abc_4268_new_n977_), .B(RST), .Y(_0rdata_31_0__5_));
AND2X2 AND2X2_198 ( .A(axi_rready), .B(\axi_rdata[6] ), .Y(_abc_4268_new_n979_));
AND2X2 AND2X2_199 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_6_), .Y(_abc_4268_new_n980_));
AND2X2 AND2X2_2 ( .A(_abc_4268_new_n558_), .B(axi_wready), .Y(_abc_4268_new_n559_));
AND2X2 AND2X2_20 ( .A(RST), .B(state_4_), .Y(_abc_4268_new_n591_));
AND2X2 AND2X2_200 ( .A(_abc_4268_new_n981_), .B(RST), .Y(_0rdata_31_0__6_));
AND2X2 AND2X2_201 ( .A(axi_rready), .B(\axi_rdata[7] ), .Y(_abc_4268_new_n983_));
AND2X2 AND2X2_202 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_7_), .Y(_abc_4268_new_n984_));
AND2X2 AND2X2_203 ( .A(_abc_4268_new_n985_), .B(RST), .Y(_0rdata_31_0__7_));
AND2X2 AND2X2_204 ( .A(axi_rready), .B(\axi_rdata[8] ), .Y(_abc_4268_new_n987_));
AND2X2 AND2X2_205 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_8_), .Y(_abc_4268_new_n988_));
AND2X2 AND2X2_206 ( .A(_abc_4268_new_n989_), .B(RST), .Y(_0rdata_31_0__8_));
AND2X2 AND2X2_207 ( .A(axi_rready), .B(\axi_rdata[9] ), .Y(_abc_4268_new_n991_));
AND2X2 AND2X2_208 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_9_), .Y(_abc_4268_new_n992_));
AND2X2 AND2X2_209 ( .A(_abc_4268_new_n993_), .B(RST), .Y(_0rdata_31_0__9_));
AND2X2 AND2X2_21 ( .A(_abc_4268_new_n591_), .B(_abc_4268_new_n590_), .Y(_abc_4268_new_n592_));
AND2X2 AND2X2_210 ( .A(axi_rready), .B(\axi_rdata[10] ), .Y(_abc_4268_new_n995_));
AND2X2 AND2X2_211 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_10_), .Y(_abc_4268_new_n996_));
AND2X2 AND2X2_212 ( .A(_abc_4268_new_n997_), .B(RST), .Y(_0rdata_31_0__10_));
AND2X2 AND2X2_213 ( .A(axi_rready), .B(\axi_rdata[11] ), .Y(_abc_4268_new_n999_));
AND2X2 AND2X2_214 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_11_), .Y(_abc_4268_new_n1000_));
AND2X2 AND2X2_215 ( .A(_abc_4268_new_n1001_), .B(RST), .Y(_0rdata_31_0__11_));
AND2X2 AND2X2_216 ( .A(axi_rready), .B(\axi_rdata[12] ), .Y(_abc_4268_new_n1003_));
AND2X2 AND2X2_217 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_12_), .Y(_abc_4268_new_n1004_));
AND2X2 AND2X2_218 ( .A(_abc_4268_new_n1005_), .B(RST), .Y(_0rdata_31_0__12_));
AND2X2 AND2X2_219 ( .A(axi_rready), .B(\axi_rdata[13] ), .Y(_abc_4268_new_n1007_));
AND2X2 AND2X2_22 ( .A(_abc_4268_new_n602_), .B(state_0_), .Y(_abc_4268_new_n603_));
AND2X2 AND2X2_220 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_13_), .Y(_abc_4268_new_n1008_));
AND2X2 AND2X2_221 ( .A(_abc_4268_new_n1009_), .B(RST), .Y(_0rdata_31_0__13_));
AND2X2 AND2X2_222 ( .A(axi_rready), .B(\axi_rdata[14] ), .Y(_abc_4268_new_n1011_));
AND2X2 AND2X2_223 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_14_), .Y(_abc_4268_new_n1012_));
AND2X2 AND2X2_224 ( .A(_abc_4268_new_n1013_), .B(RST), .Y(_0rdata_31_0__14_));
AND2X2 AND2X2_225 ( .A(axi_rready), .B(\axi_rdata[15] ), .Y(_abc_4268_new_n1015_));
AND2X2 AND2X2_226 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_15_), .Y(_abc_4268_new_n1016_));
AND2X2 AND2X2_227 ( .A(_abc_4268_new_n1017_), .B(RST), .Y(_0rdata_31_0__15_));
AND2X2 AND2X2_228 ( .A(axi_rready), .B(\axi_rdata[16] ), .Y(_abc_4268_new_n1019_));
AND2X2 AND2X2_229 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_16_), .Y(_abc_4268_new_n1020_));
AND2X2 AND2X2_23 ( .A(_abc_4268_new_n582_), .B(_abc_4268_new_n603_), .Y(_abc_4268_new_n604_));
AND2X2 AND2X2_230 ( .A(_abc_4268_new_n1021_), .B(RST), .Y(_0rdata_31_0__16_));
AND2X2 AND2X2_231 ( .A(axi_rready), .B(\axi_rdata[17] ), .Y(_abc_4268_new_n1023_));
AND2X2 AND2X2_232 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_17_), .Y(_abc_4268_new_n1024_));
AND2X2 AND2X2_233 ( .A(_abc_4268_new_n1025_), .B(RST), .Y(_0rdata_31_0__17_));
AND2X2 AND2X2_234 ( .A(axi_rready), .B(\axi_rdata[18] ), .Y(_abc_4268_new_n1027_));
AND2X2 AND2X2_235 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_18_), .Y(_abc_4268_new_n1028_));
AND2X2 AND2X2_236 ( .A(_abc_4268_new_n1029_), .B(RST), .Y(_0rdata_31_0__18_));
AND2X2 AND2X2_237 ( .A(axi_rready), .B(\axi_rdata[19] ), .Y(_abc_4268_new_n1031_));
AND2X2 AND2X2_238 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_19_), .Y(_abc_4268_new_n1032_));
AND2X2 AND2X2_239 ( .A(_abc_4268_new_n1033_), .B(RST), .Y(_0rdata_31_0__19_));
AND2X2 AND2X2_24 ( .A(_abc_4268_new_n606_), .B(state_1_), .Y(_abc_4268_new_n607_));
AND2X2 AND2X2_240 ( .A(axi_rready), .B(\axi_rdata[20] ), .Y(_abc_4268_new_n1035_));
AND2X2 AND2X2_241 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_20_), .Y(_abc_4268_new_n1036_));
AND2X2 AND2X2_242 ( .A(_abc_4268_new_n1037_), .B(RST), .Y(_0rdata_31_0__20_));
AND2X2 AND2X2_243 ( .A(axi_rready), .B(\axi_rdata[21] ), .Y(_abc_4268_new_n1039_));
AND2X2 AND2X2_244 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_21_), .Y(_abc_4268_new_n1040_));
AND2X2 AND2X2_245 ( .A(_abc_4268_new_n1041_), .B(RST), .Y(_0rdata_31_0__21_));
AND2X2 AND2X2_246 ( .A(axi_rready), .B(\axi_rdata[22] ), .Y(_abc_4268_new_n1043_));
AND2X2 AND2X2_247 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_22_), .Y(_abc_4268_new_n1044_));
AND2X2 AND2X2_248 ( .A(_abc_4268_new_n1045_), .B(RST), .Y(_0rdata_31_0__22_));
AND2X2 AND2X2_249 ( .A(axi_rready), .B(\axi_rdata[23] ), .Y(_abc_4268_new_n1047_));
AND2X2 AND2X2_25 ( .A(_abc_4268_new_n610_), .B(state_5_), .Y(_abc_4268_new_n611_));
AND2X2 AND2X2_250 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_23_), .Y(_abc_4268_new_n1048_));
AND2X2 AND2X2_251 ( .A(_abc_4268_new_n1049_), .B(RST), .Y(_0rdata_31_0__23_));
AND2X2 AND2X2_252 ( .A(axi_rready), .B(\axi_rdata[24] ), .Y(_abc_4268_new_n1051_));
AND2X2 AND2X2_253 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_24_), .Y(_abc_4268_new_n1052_));
AND2X2 AND2X2_254 ( .A(_abc_4268_new_n1053_), .B(RST), .Y(_0rdata_31_0__24_));
AND2X2 AND2X2_255 ( .A(axi_rready), .B(\axi_rdata[25] ), .Y(_abc_4268_new_n1055_));
AND2X2 AND2X2_256 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_25_), .Y(_abc_4268_new_n1056_));
AND2X2 AND2X2_257 ( .A(_abc_4268_new_n1057_), .B(RST), .Y(_0rdata_31_0__25_));
AND2X2 AND2X2_258 ( .A(axi_rready), .B(\axi_rdata[26] ), .Y(_abc_4268_new_n1059_));
AND2X2 AND2X2_259 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_26_), .Y(_abc_4268_new_n1060_));
AND2X2 AND2X2_26 ( .A(_abc_4268_new_n580_), .B(state_0_), .Y(_abc_4268_new_n612_));
AND2X2 AND2X2_260 ( .A(_abc_4268_new_n1061_), .B(RST), .Y(_0rdata_31_0__26_));
AND2X2 AND2X2_261 ( .A(axi_rready), .B(\axi_rdata[27] ), .Y(_abc_4268_new_n1063_));
AND2X2 AND2X2_262 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_27_), .Y(_abc_4268_new_n1064_));
AND2X2 AND2X2_263 ( .A(_abc_4268_new_n1065_), .B(RST), .Y(_0rdata_31_0__27_));
AND2X2 AND2X2_264 ( .A(axi_rready), .B(\axi_rdata[28] ), .Y(_abc_4268_new_n1067_));
AND2X2 AND2X2_265 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_28_), .Y(_abc_4268_new_n1068_));
AND2X2 AND2X2_266 ( .A(_abc_4268_new_n1069_), .B(RST), .Y(_0rdata_31_0__28_));
AND2X2 AND2X2_267 ( .A(axi_rready), .B(\axi_rdata[29] ), .Y(_abc_4268_new_n1071_));
AND2X2 AND2X2_268 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_29_), .Y(_abc_4268_new_n1072_));
AND2X2 AND2X2_269 ( .A(_abc_4268_new_n1073_), .B(RST), .Y(_0rdata_31_0__29_));
AND2X2 AND2X2_27 ( .A(_abc_4268_new_n613_), .B(RST), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_5_));
AND2X2 AND2X2_270 ( .A(axi_rready), .B(\axi_rdata[30] ), .Y(_abc_4268_new_n1075_));
AND2X2 AND2X2_271 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_30_), .Y(_abc_4268_new_n1076_));
AND2X2 AND2X2_272 ( .A(_abc_4268_new_n1077_), .B(RST), .Y(_0rdata_31_0__30_));
AND2X2 AND2X2_273 ( .A(axi_rready), .B(\axi_rdata[31] ), .Y(_abc_4268_new_n1079_));
AND2X2 AND2X2_274 ( .A(_abc_4268_new_n955_), .B(bus_sync_rdata_data_in_31_), .Y(_abc_4268_new_n1080_));
AND2X2 AND2X2_275 ( .A(_abc_4268_new_n1081_), .B(RST), .Y(_0rdata_31_0__31_));
AND2X2 AND2X2_276 ( .A(_abc_4268_new_n1083_), .B(counter_65_), .Y(_abc_4268_new_n1084_));
AND2X2 AND2X2_277 ( .A(_abc_4268_new_n1084_), .B(we), .Y(_abc_4268_new_n1085_));
AND2X2 AND2X2_278 ( .A(_abc_4268_new_n1085_), .B(DATA), .Y(_abc_4268_new_n1086_));
AND2X2 AND2X2_279 ( .A(_abc_4268_new_n1087_), .B(WDATA_0_), .Y(_abc_4268_new_n1088_));
AND2X2 AND2X2_28 ( .A(we), .B(DATA), .Y(_abc_4268_new_n615_));
AND2X2 AND2X2_280 ( .A(_abc_4268_new_n1089_), .B(RST), .Y(_0WDATA_31_0__0_));
AND2X2 AND2X2_281 ( .A(_abc_4268_new_n1085_), .B(sft_reg_0_), .Y(_abc_4268_new_n1091_));
AND2X2 AND2X2_282 ( .A(_abc_4268_new_n1087_), .B(WDATA_1_), .Y(_abc_4268_new_n1092_));
AND2X2 AND2X2_283 ( .A(_abc_4268_new_n1093_), .B(RST), .Y(_0WDATA_31_0__1_));
AND2X2 AND2X2_284 ( .A(_abc_4268_new_n1085_), .B(sft_reg_1_), .Y(_abc_4268_new_n1095_));
AND2X2 AND2X2_285 ( .A(_abc_4268_new_n1087_), .B(WDATA_2_), .Y(_abc_4268_new_n1096_));
AND2X2 AND2X2_286 ( .A(_abc_4268_new_n1097_), .B(RST), .Y(_0WDATA_31_0__2_));
AND2X2 AND2X2_287 ( .A(_abc_4268_new_n1085_), .B(sft_reg_2_), .Y(_abc_4268_new_n1099_));
AND2X2 AND2X2_288 ( .A(_abc_4268_new_n1087_), .B(WDATA_3_), .Y(_abc_4268_new_n1100_));
AND2X2 AND2X2_289 ( .A(_abc_4268_new_n1101_), .B(RST), .Y(_0WDATA_31_0__3_));
AND2X2 AND2X2_29 ( .A(_abc_4268_new_n615_), .B(counter_1_), .Y(_abc_4268_new_n616_));
AND2X2 AND2X2_290 ( .A(_abc_4268_new_n1085_), .B(sft_reg_3_), .Y(_abc_4268_new_n1103_));
AND2X2 AND2X2_291 ( .A(_abc_4268_new_n1087_), .B(WDATA_4_), .Y(_abc_4268_new_n1104_));
AND2X2 AND2X2_292 ( .A(_abc_4268_new_n1105_), .B(RST), .Y(_0WDATA_31_0__4_));
AND2X2 AND2X2_293 ( .A(_abc_4268_new_n1085_), .B(sft_reg_4_), .Y(_abc_4268_new_n1107_));
AND2X2 AND2X2_294 ( .A(_abc_4268_new_n1087_), .B(WDATA_5_), .Y(_abc_4268_new_n1108_));
AND2X2 AND2X2_295 ( .A(_abc_4268_new_n1109_), .B(RST), .Y(_0WDATA_31_0__5_));
AND2X2 AND2X2_296 ( .A(_abc_4268_new_n1085_), .B(sft_reg_5_), .Y(_abc_4268_new_n1111_));
AND2X2 AND2X2_297 ( .A(_abc_4268_new_n1087_), .B(WDATA_6_), .Y(_abc_4268_new_n1112_));
AND2X2 AND2X2_298 ( .A(_abc_4268_new_n1113_), .B(RST), .Y(_0WDATA_31_0__6_));
AND2X2 AND2X2_299 ( .A(_abc_4268_new_n1085_), .B(sft_reg_6_), .Y(_abc_4268_new_n1115_));
AND2X2 AND2X2_3 ( .A(state_7_), .B(RST), .Y(_abc_4268_new_n561_));
AND2X2 AND2X2_30 ( .A(_abc_4268_new_n617_), .B(_abc_4268_new_n620_), .Y(_abc_4268_new_n621_));
AND2X2 AND2X2_300 ( .A(_abc_4268_new_n1087_), .B(WDATA_7_), .Y(_abc_4268_new_n1116_));
AND2X2 AND2X2_301 ( .A(_abc_4268_new_n1117_), .B(RST), .Y(_0WDATA_31_0__7_));
AND2X2 AND2X2_302 ( .A(_abc_4268_new_n1085_), .B(sft_reg_7_), .Y(_abc_4268_new_n1119_));
AND2X2 AND2X2_303 ( .A(_abc_4268_new_n1087_), .B(WDATA_8_), .Y(_abc_4268_new_n1120_));
AND2X2 AND2X2_304 ( .A(_abc_4268_new_n1121_), .B(RST), .Y(_0WDATA_31_0__8_));
AND2X2 AND2X2_305 ( .A(_abc_4268_new_n1085_), .B(sft_reg_8_), .Y(_abc_4268_new_n1123_));
AND2X2 AND2X2_306 ( .A(_abc_4268_new_n1087_), .B(WDATA_9_), .Y(_abc_4268_new_n1124_));
AND2X2 AND2X2_307 ( .A(_abc_4268_new_n1125_), .B(RST), .Y(_0WDATA_31_0__9_));
AND2X2 AND2X2_308 ( .A(_abc_4268_new_n1085_), .B(sft_reg_9_), .Y(_abc_4268_new_n1127_));
AND2X2 AND2X2_309 ( .A(_abc_4268_new_n1087_), .B(WDATA_10_), .Y(_abc_4268_new_n1128_));
AND2X2 AND2X2_31 ( .A(re), .B(we), .Y(_abc_4268_new_n623_));
AND2X2 AND2X2_310 ( .A(_abc_4268_new_n1129_), .B(RST), .Y(_0WDATA_31_0__10_));
AND2X2 AND2X2_311 ( .A(_abc_4268_new_n1085_), .B(sft_reg_10_), .Y(_abc_4268_new_n1131_));
AND2X2 AND2X2_312 ( .A(_abc_4268_new_n1087_), .B(WDATA_11_), .Y(_abc_4268_new_n1132_));
AND2X2 AND2X2_313 ( .A(_abc_4268_new_n1133_), .B(RST), .Y(_0WDATA_31_0__11_));
AND2X2 AND2X2_314 ( .A(_abc_4268_new_n1085_), .B(sft_reg_11_), .Y(_abc_4268_new_n1135_));
AND2X2 AND2X2_315 ( .A(_abc_4268_new_n1087_), .B(WDATA_12_), .Y(_abc_4268_new_n1136_));
AND2X2 AND2X2_316 ( .A(_abc_4268_new_n1137_), .B(RST), .Y(_0WDATA_31_0__12_));
AND2X2 AND2X2_317 ( .A(_abc_4268_new_n1085_), .B(sft_reg_12_), .Y(_abc_4268_new_n1139_));
AND2X2 AND2X2_318 ( .A(_abc_4268_new_n1087_), .B(WDATA_13_), .Y(_abc_4268_new_n1140_));
AND2X2 AND2X2_319 ( .A(_abc_4268_new_n1141_), .B(RST), .Y(_0WDATA_31_0__13_));
AND2X2 AND2X2_32 ( .A(_abc_4268_new_n629_), .B(_abc_4268_new_n631_), .Y(_abc_4268_new_n632_));
AND2X2 AND2X2_320 ( .A(_abc_4268_new_n1085_), .B(sft_reg_13_), .Y(_abc_4268_new_n1143_));
AND2X2 AND2X2_321 ( .A(_abc_4268_new_n1087_), .B(WDATA_14_), .Y(_abc_4268_new_n1144_));
AND2X2 AND2X2_322 ( .A(_abc_4268_new_n1145_), .B(RST), .Y(_0WDATA_31_0__14_));
AND2X2 AND2X2_323 ( .A(_abc_4268_new_n1085_), .B(sft_reg_14_), .Y(_abc_4268_new_n1147_));
AND2X2 AND2X2_324 ( .A(_abc_4268_new_n1087_), .B(WDATA_15_), .Y(_abc_4268_new_n1148_));
AND2X2 AND2X2_325 ( .A(_abc_4268_new_n1149_), .B(RST), .Y(_0WDATA_31_0__15_));
AND2X2 AND2X2_326 ( .A(_abc_4268_new_n1085_), .B(sft_reg_15_), .Y(_abc_4268_new_n1151_));
AND2X2 AND2X2_327 ( .A(_abc_4268_new_n1087_), .B(WDATA_16_), .Y(_abc_4268_new_n1152_));
AND2X2 AND2X2_328 ( .A(_abc_4268_new_n1153_), .B(RST), .Y(_0WDATA_31_0__16_));
AND2X2 AND2X2_329 ( .A(_abc_4268_new_n1085_), .B(sft_reg_16_), .Y(_abc_4268_new_n1155_));
AND2X2 AND2X2_33 ( .A(_abc_4268_new_n634_), .B(_abc_4268_new_n636_), .Y(_abc_4268_new_n637_));
AND2X2 AND2X2_330 ( .A(_abc_4268_new_n1087_), .B(WDATA_17_), .Y(_abc_4268_new_n1156_));
AND2X2 AND2X2_331 ( .A(_abc_4268_new_n1157_), .B(RST), .Y(_0WDATA_31_0__17_));
AND2X2 AND2X2_332 ( .A(_abc_4268_new_n1085_), .B(sft_reg_17_), .Y(_abc_4268_new_n1159_));
AND2X2 AND2X2_333 ( .A(_abc_4268_new_n1087_), .B(WDATA_18_), .Y(_abc_4268_new_n1160_));
AND2X2 AND2X2_334 ( .A(_abc_4268_new_n1161_), .B(RST), .Y(_0WDATA_31_0__18_));
AND2X2 AND2X2_335 ( .A(_abc_4268_new_n1085_), .B(sft_reg_18_), .Y(_abc_4268_new_n1163_));
AND2X2 AND2X2_336 ( .A(_abc_4268_new_n1087_), .B(WDATA_19_), .Y(_abc_4268_new_n1164_));
AND2X2 AND2X2_337 ( .A(_abc_4268_new_n1165_), .B(RST), .Y(_0WDATA_31_0__19_));
AND2X2 AND2X2_338 ( .A(_abc_4268_new_n1085_), .B(sft_reg_19_), .Y(_abc_4268_new_n1167_));
AND2X2 AND2X2_339 ( .A(_abc_4268_new_n1087_), .B(WDATA_20_), .Y(_abc_4268_new_n1168_));
AND2X2 AND2X2_34 ( .A(_abc_4268_new_n632_), .B(_abc_4268_new_n637_), .Y(_abc_4268_new_n638_));
AND2X2 AND2X2_340 ( .A(_abc_4268_new_n1169_), .B(RST), .Y(_0WDATA_31_0__20_));
AND2X2 AND2X2_341 ( .A(_abc_4268_new_n1085_), .B(sft_reg_20_), .Y(_abc_4268_new_n1171_));
AND2X2 AND2X2_342 ( .A(_abc_4268_new_n1087_), .B(WDATA_21_), .Y(_abc_4268_new_n1172_));
AND2X2 AND2X2_343 ( .A(_abc_4268_new_n1173_), .B(RST), .Y(_0WDATA_31_0__21_));
AND2X2 AND2X2_344 ( .A(_abc_4268_new_n1085_), .B(sft_reg_21_), .Y(_abc_4268_new_n1175_));
AND2X2 AND2X2_345 ( .A(_abc_4268_new_n1087_), .B(WDATA_22_), .Y(_abc_4268_new_n1176_));
AND2X2 AND2X2_346 ( .A(_abc_4268_new_n1177_), .B(RST), .Y(_0WDATA_31_0__22_));
AND2X2 AND2X2_347 ( .A(_abc_4268_new_n1085_), .B(sft_reg_22_), .Y(_abc_4268_new_n1179_));
AND2X2 AND2X2_348 ( .A(_abc_4268_new_n1087_), .B(WDATA_23_), .Y(_abc_4268_new_n1180_));
AND2X2 AND2X2_349 ( .A(_abc_4268_new_n1181_), .B(RST), .Y(_0WDATA_31_0__23_));
AND2X2 AND2X2_35 ( .A(_abc_4268_new_n640_), .B(_abc_4268_new_n642_), .Y(_abc_4268_new_n643_));
AND2X2 AND2X2_350 ( .A(_abc_4268_new_n1085_), .B(sft_reg_23_), .Y(_abc_4268_new_n1183_));
AND2X2 AND2X2_351 ( .A(_abc_4268_new_n1087_), .B(WDATA_24_), .Y(_abc_4268_new_n1184_));
AND2X2 AND2X2_352 ( .A(_abc_4268_new_n1185_), .B(RST), .Y(_0WDATA_31_0__24_));
AND2X2 AND2X2_353 ( .A(_abc_4268_new_n1085_), .B(sft_reg_24_), .Y(_abc_4268_new_n1187_));
AND2X2 AND2X2_354 ( .A(_abc_4268_new_n1087_), .B(WDATA_25_), .Y(_abc_4268_new_n1188_));
AND2X2 AND2X2_355 ( .A(_abc_4268_new_n1189_), .B(RST), .Y(_0WDATA_31_0__25_));
AND2X2 AND2X2_356 ( .A(_abc_4268_new_n1085_), .B(sft_reg_25_), .Y(_abc_4268_new_n1191_));
AND2X2 AND2X2_357 ( .A(_abc_4268_new_n1087_), .B(WDATA_26_), .Y(_abc_4268_new_n1192_));
AND2X2 AND2X2_358 ( .A(_abc_4268_new_n1193_), .B(RST), .Y(_0WDATA_31_0__26_));
AND2X2 AND2X2_359 ( .A(_abc_4268_new_n1085_), .B(sft_reg_26_), .Y(_abc_4268_new_n1195_));
AND2X2 AND2X2_36 ( .A(_abc_4268_new_n645_), .B(_abc_4268_new_n647_), .Y(_abc_4268_new_n648_));
AND2X2 AND2X2_360 ( .A(_abc_4268_new_n1087_), .B(WDATA_27_), .Y(_abc_4268_new_n1196_));
AND2X2 AND2X2_361 ( .A(_abc_4268_new_n1197_), .B(RST), .Y(_0WDATA_31_0__27_));
AND2X2 AND2X2_362 ( .A(_abc_4268_new_n1085_), .B(sft_reg_27_), .Y(_abc_4268_new_n1199_));
AND2X2 AND2X2_363 ( .A(_abc_4268_new_n1087_), .B(WDATA_28_), .Y(_abc_4268_new_n1200_));
AND2X2 AND2X2_364 ( .A(_abc_4268_new_n1201_), .B(RST), .Y(_0WDATA_31_0__28_));
AND2X2 AND2X2_365 ( .A(_abc_4268_new_n1085_), .B(sft_reg_28_), .Y(_abc_4268_new_n1203_));
AND2X2 AND2X2_366 ( .A(_abc_4268_new_n1087_), .B(WDATA_29_), .Y(_abc_4268_new_n1204_));
AND2X2 AND2X2_367 ( .A(_abc_4268_new_n1205_), .B(RST), .Y(_0WDATA_31_0__29_));
AND2X2 AND2X2_368 ( .A(_abc_4268_new_n1085_), .B(sft_reg_29_), .Y(_abc_4268_new_n1207_));
AND2X2 AND2X2_369 ( .A(_abc_4268_new_n1087_), .B(WDATA_30_), .Y(_abc_4268_new_n1208_));
AND2X2 AND2X2_37 ( .A(_abc_4268_new_n643_), .B(_abc_4268_new_n648_), .Y(_abc_4268_new_n649_));
AND2X2 AND2X2_370 ( .A(_abc_4268_new_n1209_), .B(RST), .Y(_0WDATA_31_0__30_));
AND2X2 AND2X2_371 ( .A(_abc_4268_new_n1085_), .B(sft_reg_30_), .Y(_abc_4268_new_n1211_));
AND2X2 AND2X2_372 ( .A(_abc_4268_new_n1087_), .B(WDATA_31_), .Y(_abc_4268_new_n1212_));
AND2X2 AND2X2_373 ( .A(_abc_4268_new_n1213_), .B(RST), .Y(_0WDATA_31_0__31_));
AND2X2 AND2X2_374 ( .A(_abc_4268_new_n627_), .B(counter_33_), .Y(_abc_4268_new_n1215_));
AND2X2 AND2X2_375 ( .A(_abc_4268_new_n1215_), .B(_abc_4268_new_n1083_), .Y(_abc_4268_new_n1216_));
AND2X2 AND2X2_376 ( .A(_abc_4268_new_n1219_), .B(RST), .Y(_abc_4268_new_n1220_));
AND2X2 AND2X2_377 ( .A(_abc_4268_new_n1220_), .B(_abc_4268_new_n1217_), .Y(_0A_ADDR_31_0__0_));
AND2X2 AND2X2_378 ( .A(_abc_4268_new_n1223_), .B(RST), .Y(_abc_4268_new_n1224_));
AND2X2 AND2X2_379 ( .A(_abc_4268_new_n1224_), .B(_abc_4268_new_n1222_), .Y(_0A_ADDR_31_0__1_));
AND2X2 AND2X2_38 ( .A(_abc_4268_new_n638_), .B(_abc_4268_new_n649_), .Y(_abc_4268_new_n650_));
AND2X2 AND2X2_380 ( .A(_abc_4268_new_n1227_), .B(RST), .Y(_abc_4268_new_n1228_));
AND2X2 AND2X2_381 ( .A(_abc_4268_new_n1228_), .B(_abc_4268_new_n1226_), .Y(_0A_ADDR_31_0__2_));
AND2X2 AND2X2_382 ( .A(_abc_4268_new_n1231_), .B(RST), .Y(_abc_4268_new_n1232_));
AND2X2 AND2X2_383 ( .A(_abc_4268_new_n1232_), .B(_abc_4268_new_n1230_), .Y(_0A_ADDR_31_0__3_));
AND2X2 AND2X2_384 ( .A(_abc_4268_new_n1235_), .B(RST), .Y(_abc_4268_new_n1236_));
AND2X2 AND2X2_385 ( .A(_abc_4268_new_n1236_), .B(_abc_4268_new_n1234_), .Y(_0A_ADDR_31_0__4_));
AND2X2 AND2X2_386 ( .A(_abc_4268_new_n1239_), .B(RST), .Y(_abc_4268_new_n1240_));
AND2X2 AND2X2_387 ( .A(_abc_4268_new_n1240_), .B(_abc_4268_new_n1238_), .Y(_0A_ADDR_31_0__5_));
AND2X2 AND2X2_388 ( .A(_abc_4268_new_n1243_), .B(RST), .Y(_abc_4268_new_n1244_));
AND2X2 AND2X2_389 ( .A(_abc_4268_new_n1244_), .B(_abc_4268_new_n1242_), .Y(_0A_ADDR_31_0__6_));
AND2X2 AND2X2_39 ( .A(_abc_4268_new_n652_), .B(_abc_4268_new_n654_), .Y(_abc_4268_new_n655_));
AND2X2 AND2X2_390 ( .A(_abc_4268_new_n1247_), .B(RST), .Y(_abc_4268_new_n1248_));
AND2X2 AND2X2_391 ( .A(_abc_4268_new_n1248_), .B(_abc_4268_new_n1246_), .Y(_0A_ADDR_31_0__7_));
AND2X2 AND2X2_392 ( .A(_abc_4268_new_n1251_), .B(RST), .Y(_abc_4268_new_n1252_));
AND2X2 AND2X2_393 ( .A(_abc_4268_new_n1252_), .B(_abc_4268_new_n1250_), .Y(_0A_ADDR_31_0__8_));
AND2X2 AND2X2_394 ( .A(_abc_4268_new_n1255_), .B(RST), .Y(_abc_4268_new_n1256_));
AND2X2 AND2X2_395 ( .A(_abc_4268_new_n1256_), .B(_abc_4268_new_n1254_), .Y(_0A_ADDR_31_0__9_));
AND2X2 AND2X2_396 ( .A(_abc_4268_new_n1259_), .B(RST), .Y(_abc_4268_new_n1260_));
AND2X2 AND2X2_397 ( .A(_abc_4268_new_n1260_), .B(_abc_4268_new_n1258_), .Y(_0A_ADDR_31_0__10_));
AND2X2 AND2X2_398 ( .A(_abc_4268_new_n1263_), .B(RST), .Y(_abc_4268_new_n1264_));
AND2X2 AND2X2_399 ( .A(_abc_4268_new_n1264_), .B(_abc_4268_new_n1262_), .Y(_0A_ADDR_31_0__11_));
AND2X2 AND2X2_4 ( .A(_abc_4268_new_n561_), .B(_abc_4268_new_n560_), .Y(_abc_4268_new_n562_));
AND2X2 AND2X2_40 ( .A(_abc_4268_new_n657_), .B(_abc_4268_new_n659_), .Y(_abc_4268_new_n660_));
AND2X2 AND2X2_400 ( .A(_abc_4268_new_n1267_), .B(RST), .Y(_abc_4268_new_n1268_));
AND2X2 AND2X2_401 ( .A(_abc_4268_new_n1268_), .B(_abc_4268_new_n1266_), .Y(_0A_ADDR_31_0__12_));
AND2X2 AND2X2_402 ( .A(_abc_4268_new_n1271_), .B(RST), .Y(_abc_4268_new_n1272_));
AND2X2 AND2X2_403 ( .A(_abc_4268_new_n1272_), .B(_abc_4268_new_n1270_), .Y(_0A_ADDR_31_0__13_));
AND2X2 AND2X2_404 ( .A(_abc_4268_new_n1275_), .B(RST), .Y(_abc_4268_new_n1276_));
AND2X2 AND2X2_405 ( .A(_abc_4268_new_n1276_), .B(_abc_4268_new_n1274_), .Y(_0A_ADDR_31_0__14_));
AND2X2 AND2X2_406 ( .A(_abc_4268_new_n1279_), .B(RST), .Y(_abc_4268_new_n1280_));
AND2X2 AND2X2_407 ( .A(_abc_4268_new_n1280_), .B(_abc_4268_new_n1278_), .Y(_0A_ADDR_31_0__15_));
AND2X2 AND2X2_408 ( .A(_abc_4268_new_n1283_), .B(RST), .Y(_abc_4268_new_n1284_));
AND2X2 AND2X2_409 ( .A(_abc_4268_new_n1284_), .B(_abc_4268_new_n1282_), .Y(_0A_ADDR_31_0__16_));
AND2X2 AND2X2_41 ( .A(_abc_4268_new_n655_), .B(_abc_4268_new_n660_), .Y(_abc_4268_new_n661_));
AND2X2 AND2X2_410 ( .A(_abc_4268_new_n1287_), .B(RST), .Y(_abc_4268_new_n1288_));
AND2X2 AND2X2_411 ( .A(_abc_4268_new_n1288_), .B(_abc_4268_new_n1286_), .Y(_0A_ADDR_31_0__17_));
AND2X2 AND2X2_412 ( .A(_abc_4268_new_n1291_), .B(RST), .Y(_abc_4268_new_n1292_));
AND2X2 AND2X2_413 ( .A(_abc_4268_new_n1292_), .B(_abc_4268_new_n1290_), .Y(_0A_ADDR_31_0__18_));
AND2X2 AND2X2_414 ( .A(_abc_4268_new_n1295_), .B(RST), .Y(_abc_4268_new_n1296_));
AND2X2 AND2X2_415 ( .A(_abc_4268_new_n1296_), .B(_abc_4268_new_n1294_), .Y(_0A_ADDR_31_0__19_));
AND2X2 AND2X2_416 ( .A(_abc_4268_new_n1299_), .B(RST), .Y(_abc_4268_new_n1300_));
AND2X2 AND2X2_417 ( .A(_abc_4268_new_n1300_), .B(_abc_4268_new_n1298_), .Y(_0A_ADDR_31_0__20_));
AND2X2 AND2X2_418 ( .A(_abc_4268_new_n1303_), .B(RST), .Y(_abc_4268_new_n1304_));
AND2X2 AND2X2_419 ( .A(_abc_4268_new_n1304_), .B(_abc_4268_new_n1302_), .Y(_0A_ADDR_31_0__21_));
AND2X2 AND2X2_42 ( .A(_abc_4268_new_n663_), .B(_abc_4268_new_n665_), .Y(_abc_4268_new_n666_));
AND2X2 AND2X2_420 ( .A(_abc_4268_new_n1307_), .B(RST), .Y(_abc_4268_new_n1308_));
AND2X2 AND2X2_421 ( .A(_abc_4268_new_n1308_), .B(_abc_4268_new_n1306_), .Y(_0A_ADDR_31_0__22_));
AND2X2 AND2X2_422 ( .A(_abc_4268_new_n1311_), .B(RST), .Y(_abc_4268_new_n1312_));
AND2X2 AND2X2_423 ( .A(_abc_4268_new_n1312_), .B(_abc_4268_new_n1310_), .Y(_0A_ADDR_31_0__23_));
AND2X2 AND2X2_424 ( .A(_abc_4268_new_n1315_), .B(RST), .Y(_abc_4268_new_n1316_));
AND2X2 AND2X2_425 ( .A(_abc_4268_new_n1316_), .B(_abc_4268_new_n1314_), .Y(_0A_ADDR_31_0__24_));
AND2X2 AND2X2_426 ( .A(_abc_4268_new_n1319_), .B(RST), .Y(_abc_4268_new_n1320_));
AND2X2 AND2X2_427 ( .A(_abc_4268_new_n1320_), .B(_abc_4268_new_n1318_), .Y(_0A_ADDR_31_0__25_));
AND2X2 AND2X2_428 ( .A(_abc_4268_new_n1323_), .B(RST), .Y(_abc_4268_new_n1324_));
AND2X2 AND2X2_429 ( .A(_abc_4268_new_n1324_), .B(_abc_4268_new_n1322_), .Y(_0A_ADDR_31_0__26_));
AND2X2 AND2X2_43 ( .A(_abc_4268_new_n669_), .B(_abc_4268_new_n670_), .Y(_abc_4268_new_n671_));
AND2X2 AND2X2_430 ( .A(_abc_4268_new_n1327_), .B(RST), .Y(_abc_4268_new_n1328_));
AND2X2 AND2X2_431 ( .A(_abc_4268_new_n1328_), .B(_abc_4268_new_n1326_), .Y(_0A_ADDR_31_0__27_));
AND2X2 AND2X2_432 ( .A(_abc_4268_new_n1331_), .B(RST), .Y(_abc_4268_new_n1332_));
AND2X2 AND2X2_433 ( .A(_abc_4268_new_n1332_), .B(_abc_4268_new_n1330_), .Y(_0A_ADDR_31_0__28_));
AND2X2 AND2X2_434 ( .A(_abc_4268_new_n1335_), .B(RST), .Y(_abc_4268_new_n1336_));
AND2X2 AND2X2_435 ( .A(_abc_4268_new_n1336_), .B(_abc_4268_new_n1334_), .Y(_0A_ADDR_31_0__29_));
AND2X2 AND2X2_436 ( .A(_abc_4268_new_n1339_), .B(RST), .Y(_abc_4268_new_n1340_));
AND2X2 AND2X2_437 ( .A(_abc_4268_new_n1340_), .B(_abc_4268_new_n1338_), .Y(_0A_ADDR_31_0__30_));
AND2X2 AND2X2_438 ( .A(_abc_4268_new_n1216_), .B(sft_reg_30_), .Y(_abc_4268_new_n1342_));
AND2X2 AND2X2_439 ( .A(_abc_4268_new_n1218_), .B(A_ADDR_31_), .Y(_abc_4268_new_n1343_));
AND2X2 AND2X2_44 ( .A(_abc_4268_new_n668_), .B(_abc_4268_new_n671_), .Y(_abc_4268_new_n672_));
AND2X2 AND2X2_440 ( .A(_abc_4268_new_n1344_), .B(RST), .Y(_0A_ADDR_31_0__31_));
AND2X2 AND2X2_441 ( .A(_abc_4268_new_n1347_), .B(RST), .Y(_abc_4268_new_n1348_));
AND2X2 AND2X2_442 ( .A(_abc_4268_new_n1348_), .B(_abc_4268_new_n1346_), .Y(_0sft_reg_65_0__0_));
AND2X2 AND2X2_443 ( .A(_abc_4268_new_n1351_), .B(RST), .Y(_abc_4268_new_n1352_));
AND2X2 AND2X2_444 ( .A(_abc_4268_new_n1352_), .B(_abc_4268_new_n1350_), .Y(_0sft_reg_65_0__1_));
AND2X2 AND2X2_445 ( .A(_abc_4268_new_n1355_), .B(RST), .Y(_abc_4268_new_n1356_));
AND2X2 AND2X2_446 ( .A(_abc_4268_new_n1356_), .B(_abc_4268_new_n1354_), .Y(_0sft_reg_65_0__2_));
AND2X2 AND2X2_447 ( .A(_abc_4268_new_n1359_), .B(RST), .Y(_abc_4268_new_n1360_));
AND2X2 AND2X2_448 ( .A(_abc_4268_new_n1360_), .B(_abc_4268_new_n1358_), .Y(_0sft_reg_65_0__3_));
AND2X2 AND2X2_449 ( .A(_abc_4268_new_n1363_), .B(RST), .Y(_abc_4268_new_n1364_));
AND2X2 AND2X2_45 ( .A(_abc_4268_new_n666_), .B(_abc_4268_new_n672_), .Y(_abc_4268_new_n673_));
AND2X2 AND2X2_450 ( .A(_abc_4268_new_n1364_), .B(_abc_4268_new_n1362_), .Y(_0sft_reg_65_0__4_));
AND2X2 AND2X2_451 ( .A(_abc_4268_new_n1367_), .B(RST), .Y(_abc_4268_new_n1368_));
AND2X2 AND2X2_452 ( .A(_abc_4268_new_n1368_), .B(_abc_4268_new_n1366_), .Y(_0sft_reg_65_0__5_));
AND2X2 AND2X2_453 ( .A(_abc_4268_new_n1371_), .B(RST), .Y(_abc_4268_new_n1372_));
AND2X2 AND2X2_454 ( .A(_abc_4268_new_n1372_), .B(_abc_4268_new_n1370_), .Y(_0sft_reg_65_0__6_));
AND2X2 AND2X2_455 ( .A(_abc_4268_new_n1375_), .B(RST), .Y(_abc_4268_new_n1376_));
AND2X2 AND2X2_456 ( .A(_abc_4268_new_n1376_), .B(_abc_4268_new_n1374_), .Y(_0sft_reg_65_0__7_));
AND2X2 AND2X2_457 ( .A(_abc_4268_new_n1379_), .B(RST), .Y(_abc_4268_new_n1380_));
AND2X2 AND2X2_458 ( .A(_abc_4268_new_n1380_), .B(_abc_4268_new_n1378_), .Y(_0sft_reg_65_0__8_));
AND2X2 AND2X2_459 ( .A(_abc_4268_new_n1383_), .B(RST), .Y(_abc_4268_new_n1384_));
AND2X2 AND2X2_46 ( .A(_abc_4268_new_n661_), .B(_abc_4268_new_n673_), .Y(_abc_4268_new_n674_));
AND2X2 AND2X2_460 ( .A(_abc_4268_new_n1384_), .B(_abc_4268_new_n1382_), .Y(_0sft_reg_65_0__9_));
AND2X2 AND2X2_461 ( .A(_abc_4268_new_n1387_), .B(RST), .Y(_abc_4268_new_n1388_));
AND2X2 AND2X2_462 ( .A(_abc_4268_new_n1388_), .B(_abc_4268_new_n1386_), .Y(_0sft_reg_65_0__10_));
AND2X2 AND2X2_463 ( .A(_abc_4268_new_n1391_), .B(RST), .Y(_abc_4268_new_n1392_));
AND2X2 AND2X2_464 ( .A(_abc_4268_new_n1392_), .B(_abc_4268_new_n1390_), .Y(_0sft_reg_65_0__11_));
AND2X2 AND2X2_465 ( .A(_abc_4268_new_n1395_), .B(RST), .Y(_abc_4268_new_n1396_));
AND2X2 AND2X2_466 ( .A(_abc_4268_new_n1396_), .B(_abc_4268_new_n1394_), .Y(_0sft_reg_65_0__12_));
AND2X2 AND2X2_467 ( .A(_abc_4268_new_n1399_), .B(RST), .Y(_abc_4268_new_n1400_));
AND2X2 AND2X2_468 ( .A(_abc_4268_new_n1400_), .B(_abc_4268_new_n1398_), .Y(_0sft_reg_65_0__13_));
AND2X2 AND2X2_469 ( .A(_abc_4268_new_n1403_), .B(RST), .Y(_abc_4268_new_n1404_));
AND2X2 AND2X2_47 ( .A(_abc_4268_new_n650_), .B(_abc_4268_new_n674_), .Y(_abc_4268_new_n675_));
AND2X2 AND2X2_470 ( .A(_abc_4268_new_n1404_), .B(_abc_4268_new_n1402_), .Y(_0sft_reg_65_0__14_));
AND2X2 AND2X2_471 ( .A(_abc_4268_new_n1407_), .B(RST), .Y(_abc_4268_new_n1408_));
AND2X2 AND2X2_472 ( .A(_abc_4268_new_n1408_), .B(_abc_4268_new_n1406_), .Y(_0sft_reg_65_0__15_));
AND2X2 AND2X2_473 ( .A(_abc_4268_new_n1411_), .B(RST), .Y(_abc_4268_new_n1412_));
AND2X2 AND2X2_474 ( .A(_abc_4268_new_n1412_), .B(_abc_4268_new_n1410_), .Y(_0sft_reg_65_0__16_));
AND2X2 AND2X2_475 ( .A(_abc_4268_new_n1415_), .B(RST), .Y(_abc_4268_new_n1416_));
AND2X2 AND2X2_476 ( .A(_abc_4268_new_n1416_), .B(_abc_4268_new_n1414_), .Y(_0sft_reg_65_0__17_));
AND2X2 AND2X2_477 ( .A(_abc_4268_new_n1419_), .B(RST), .Y(_abc_4268_new_n1420_));
AND2X2 AND2X2_478 ( .A(_abc_4268_new_n1420_), .B(_abc_4268_new_n1418_), .Y(_0sft_reg_65_0__18_));
AND2X2 AND2X2_479 ( .A(_abc_4268_new_n1423_), .B(RST), .Y(_abc_4268_new_n1424_));
AND2X2 AND2X2_48 ( .A(_abc_4268_new_n676_), .B(bus_cap_0_), .Y(_abc_4268_new_n677_));
AND2X2 AND2X2_480 ( .A(_abc_4268_new_n1424_), .B(_abc_4268_new_n1422_), .Y(_0sft_reg_65_0__19_));
AND2X2 AND2X2_481 ( .A(_abc_4268_new_n1427_), .B(RST), .Y(_abc_4268_new_n1428_));
AND2X2 AND2X2_482 ( .A(_abc_4268_new_n1428_), .B(_abc_4268_new_n1426_), .Y(_0sft_reg_65_0__20_));
AND2X2 AND2X2_483 ( .A(_abc_4268_new_n1431_), .B(RST), .Y(_abc_4268_new_n1432_));
AND2X2 AND2X2_484 ( .A(_abc_4268_new_n1432_), .B(_abc_4268_new_n1430_), .Y(_0sft_reg_65_0__21_));
AND2X2 AND2X2_485 ( .A(_abc_4268_new_n1435_), .B(RST), .Y(_abc_4268_new_n1436_));
AND2X2 AND2X2_486 ( .A(_abc_4268_new_n1436_), .B(_abc_4268_new_n1434_), .Y(_0sft_reg_65_0__22_));
AND2X2 AND2X2_487 ( .A(_abc_4268_new_n1439_), .B(RST), .Y(_abc_4268_new_n1440_));
AND2X2 AND2X2_488 ( .A(_abc_4268_new_n1440_), .B(_abc_4268_new_n1438_), .Y(_0sft_reg_65_0__23_));
AND2X2 AND2X2_489 ( .A(_abc_4268_new_n1443_), .B(RST), .Y(_abc_4268_new_n1444_));
AND2X2 AND2X2_49 ( .A(_abc_4268_new_n617_), .B(bus_sync_status_data_out_0_), .Y(_abc_4268_new_n679_));
AND2X2 AND2X2_490 ( .A(_abc_4268_new_n1444_), .B(_abc_4268_new_n1442_), .Y(_0sft_reg_65_0__24_));
AND2X2 AND2X2_491 ( .A(_abc_4268_new_n1447_), .B(RST), .Y(_abc_4268_new_n1448_));
AND2X2 AND2X2_492 ( .A(_abc_4268_new_n1448_), .B(_abc_4268_new_n1446_), .Y(_0sft_reg_65_0__25_));
AND2X2 AND2X2_493 ( .A(_abc_4268_new_n1451_), .B(RST), .Y(_abc_4268_new_n1452_));
AND2X2 AND2X2_494 ( .A(_abc_4268_new_n1452_), .B(_abc_4268_new_n1450_), .Y(_0sft_reg_65_0__26_));
AND2X2 AND2X2_495 ( .A(_abc_4268_new_n1455_), .B(RST), .Y(_abc_4268_new_n1456_));
AND2X2 AND2X2_496 ( .A(_abc_4268_new_n1456_), .B(_abc_4268_new_n1454_), .Y(_0sft_reg_65_0__27_));
AND2X2 AND2X2_497 ( .A(_abc_4268_new_n1459_), .B(RST), .Y(_abc_4268_new_n1460_));
AND2X2 AND2X2_498 ( .A(_abc_4268_new_n1460_), .B(_abc_4268_new_n1458_), .Y(_0sft_reg_65_0__28_));
AND2X2 AND2X2_499 ( .A(_abc_4268_new_n1463_), .B(RST), .Y(_abc_4268_new_n1464_));
AND2X2 AND2X2_5 ( .A(_abc_4268_new_n566_), .B(state_3_), .Y(_abc_4268_new_n567_));
AND2X2 AND2X2_50 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_0_), .Y(_abc_4268_new_n680_));
AND2X2 AND2X2_500 ( .A(_abc_4268_new_n1464_), .B(_abc_4268_new_n1462_), .Y(_0sft_reg_65_0__29_));
AND2X2 AND2X2_501 ( .A(_abc_4268_new_n1467_), .B(RST), .Y(_abc_4268_new_n1468_));
AND2X2 AND2X2_502 ( .A(_abc_4268_new_n1468_), .B(_abc_4268_new_n1466_), .Y(_0sft_reg_65_0__30_));
AND2X2 AND2X2_503 ( .A(_abc_4268_new_n1083_), .B(RST), .Y(_abc_4268_new_n1470_));
AND2X2 AND2X2_504 ( .A(_abc_4268_new_n1470_), .B(counter_0_), .Y(_0counter_65_0__1_));
AND2X2 AND2X2_505 ( .A(_abc_4268_new_n1470_), .B(counter_1_), .Y(_0counter_65_0__2_));
AND2X2 AND2X2_506 ( .A(_abc_4268_new_n1470_), .B(counter_2_), .Y(_0counter_65_0__3_));
AND2X2 AND2X2_507 ( .A(_abc_4268_new_n1470_), .B(counter_3_), .Y(_0counter_65_0__4_));
AND2X2 AND2X2_508 ( .A(_abc_4268_new_n1470_), .B(counter_4_), .Y(_0counter_65_0__5_));
AND2X2 AND2X2_509 ( .A(_abc_4268_new_n1470_), .B(counter_5_), .Y(_0counter_65_0__6_));
AND2X2 AND2X2_51 ( .A(_abc_4268_new_n682_), .B(RST), .Y(_abc_4268_new_n683_));
AND2X2 AND2X2_510 ( .A(_abc_4268_new_n1470_), .B(counter_6_), .Y(_0counter_65_0__7_));
AND2X2 AND2X2_511 ( .A(_abc_4268_new_n1470_), .B(counter_7_), .Y(_0counter_65_0__8_));
AND2X2 AND2X2_512 ( .A(_abc_4268_new_n1470_), .B(counter_8_), .Y(_0counter_65_0__9_));
AND2X2 AND2X2_513 ( .A(_abc_4268_new_n1470_), .B(counter_9_), .Y(_0counter_65_0__10_));
AND2X2 AND2X2_514 ( .A(_abc_4268_new_n1470_), .B(counter_10_), .Y(_0counter_65_0__11_));
AND2X2 AND2X2_515 ( .A(_abc_4268_new_n1470_), .B(counter_11_), .Y(_0counter_65_0__12_));
AND2X2 AND2X2_516 ( .A(_abc_4268_new_n1470_), .B(counter_12_), .Y(_0counter_65_0__13_));
AND2X2 AND2X2_517 ( .A(_abc_4268_new_n1470_), .B(counter_13_), .Y(_0counter_65_0__14_));
AND2X2 AND2X2_518 ( .A(_abc_4268_new_n1470_), .B(counter_14_), .Y(_0counter_65_0__15_));
AND2X2 AND2X2_519 ( .A(_abc_4268_new_n1470_), .B(counter_15_), .Y(_0counter_65_0__16_));
AND2X2 AND2X2_52 ( .A(_abc_4268_new_n678_), .B(_abc_4268_new_n683_), .Y(_0bus_cap_31_0__0_));
AND2X2 AND2X2_520 ( .A(_abc_4268_new_n1470_), .B(counter_16_), .Y(_0counter_65_0__17_));
AND2X2 AND2X2_521 ( .A(_abc_4268_new_n1470_), .B(counter_17_), .Y(_0counter_65_0__18_));
AND2X2 AND2X2_522 ( .A(_abc_4268_new_n1470_), .B(counter_18_), .Y(_0counter_65_0__19_));
AND2X2 AND2X2_523 ( .A(_abc_4268_new_n1470_), .B(counter_19_), .Y(_0counter_65_0__20_));
AND2X2 AND2X2_524 ( .A(_abc_4268_new_n1470_), .B(counter_20_), .Y(_0counter_65_0__21_));
AND2X2 AND2X2_525 ( .A(_abc_4268_new_n1470_), .B(counter_21_), .Y(_0counter_65_0__22_));
AND2X2 AND2X2_526 ( .A(_abc_4268_new_n1470_), .B(counter_22_), .Y(_0counter_65_0__23_));
AND2X2 AND2X2_527 ( .A(_abc_4268_new_n1470_), .B(counter_23_), .Y(_0counter_65_0__24_));
AND2X2 AND2X2_528 ( .A(_abc_4268_new_n1470_), .B(counter_24_), .Y(_0counter_65_0__25_));
AND2X2 AND2X2_529 ( .A(_abc_4268_new_n1470_), .B(counter_25_), .Y(_0counter_65_0__26_));
AND2X2 AND2X2_53 ( .A(_abc_4268_new_n700_), .B(_abc_4268_new_n626_), .Y(_abc_4268_new_n701_));
AND2X2 AND2X2_530 ( .A(_abc_4268_new_n1470_), .B(counter_26_), .Y(_0counter_65_0__27_));
AND2X2 AND2X2_531 ( .A(_abc_4268_new_n1470_), .B(counter_27_), .Y(_0counter_65_0__28_));
AND2X2 AND2X2_532 ( .A(_abc_4268_new_n1470_), .B(counter_28_), .Y(_0counter_65_0__29_));
AND2X2 AND2X2_533 ( .A(_abc_4268_new_n1470_), .B(counter_29_), .Y(_0counter_65_0__30_));
AND2X2 AND2X2_534 ( .A(_abc_4268_new_n1470_), .B(counter_30_), .Y(_0counter_65_0__31_));
AND2X2 AND2X2_535 ( .A(_abc_4268_new_n1470_), .B(counter_31_), .Y(_0counter_65_0__32_));
AND2X2 AND2X2_536 ( .A(_abc_4268_new_n1470_), .B(counter_32_), .Y(_0counter_65_0__33_));
AND2X2 AND2X2_537 ( .A(_abc_4268_new_n1470_), .B(counter_33_), .Y(_0counter_65_0__34_));
AND2X2 AND2X2_538 ( .A(_abc_4268_new_n1470_), .B(counter_34_), .Y(_0counter_65_0__35_));
AND2X2 AND2X2_539 ( .A(_abc_4268_new_n1470_), .B(counter_35_), .Y(_0counter_65_0__36_));
AND2X2 AND2X2_54 ( .A(_abc_4268_new_n702_), .B(_abc_4268_new_n703_), .Y(_abc_4268_new_n704_));
AND2X2 AND2X2_540 ( .A(_abc_4268_new_n1470_), .B(counter_36_), .Y(_0counter_65_0__37_));
AND2X2 AND2X2_541 ( .A(_abc_4268_new_n1470_), .B(counter_37_), .Y(_0counter_65_0__38_));
AND2X2 AND2X2_542 ( .A(_abc_4268_new_n1470_), .B(counter_38_), .Y(_0counter_65_0__39_));
AND2X2 AND2X2_543 ( .A(_abc_4268_new_n1470_), .B(counter_39_), .Y(_0counter_65_0__40_));
AND2X2 AND2X2_544 ( .A(_abc_4268_new_n1470_), .B(counter_40_), .Y(_0counter_65_0__41_));
AND2X2 AND2X2_545 ( .A(_abc_4268_new_n1470_), .B(counter_41_), .Y(_0counter_65_0__42_));
AND2X2 AND2X2_546 ( .A(_abc_4268_new_n1470_), .B(counter_42_), .Y(_0counter_65_0__43_));
AND2X2 AND2X2_547 ( .A(_abc_4268_new_n1470_), .B(counter_43_), .Y(_0counter_65_0__44_));
AND2X2 AND2X2_548 ( .A(_abc_4268_new_n1470_), .B(counter_44_), .Y(_0counter_65_0__45_));
AND2X2 AND2X2_549 ( .A(_abc_4268_new_n1470_), .B(counter_45_), .Y(_0counter_65_0__46_));
AND2X2 AND2X2_55 ( .A(_abc_4268_new_n617_), .B(bus_sync_status_data_out_1_), .Y(_abc_4268_new_n706_));
AND2X2 AND2X2_550 ( .A(_abc_4268_new_n1470_), .B(counter_46_), .Y(_0counter_65_0__47_));
AND2X2 AND2X2_551 ( .A(_abc_4268_new_n1470_), .B(counter_47_), .Y(_0counter_65_0__48_));
AND2X2 AND2X2_552 ( .A(_abc_4268_new_n1470_), .B(counter_48_), .Y(_0counter_65_0__49_));
AND2X2 AND2X2_553 ( .A(_abc_4268_new_n1470_), .B(counter_49_), .Y(_0counter_65_0__50_));
AND2X2 AND2X2_554 ( .A(_abc_4268_new_n1470_), .B(counter_50_), .Y(_0counter_65_0__51_));
AND2X2 AND2X2_555 ( .A(_abc_4268_new_n1470_), .B(counter_51_), .Y(_0counter_65_0__52_));
AND2X2 AND2X2_556 ( .A(_abc_4268_new_n1470_), .B(counter_52_), .Y(_0counter_65_0__53_));
AND2X2 AND2X2_557 ( .A(_abc_4268_new_n1470_), .B(counter_53_), .Y(_0counter_65_0__54_));
AND2X2 AND2X2_558 ( .A(_abc_4268_new_n1470_), .B(counter_54_), .Y(_0counter_65_0__55_));
AND2X2 AND2X2_559 ( .A(_abc_4268_new_n1470_), .B(counter_55_), .Y(_0counter_65_0__56_));
AND2X2 AND2X2_56 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_1_), .Y(_abc_4268_new_n707_));
AND2X2 AND2X2_560 ( .A(_abc_4268_new_n1470_), .B(counter_56_), .Y(_0counter_65_0__57_));
AND2X2 AND2X2_561 ( .A(_abc_4268_new_n1470_), .B(counter_57_), .Y(_0counter_65_0__58_));
AND2X2 AND2X2_562 ( .A(_abc_4268_new_n1470_), .B(counter_58_), .Y(_0counter_65_0__59_));
AND2X2 AND2X2_563 ( .A(_abc_4268_new_n1470_), .B(counter_59_), .Y(_0counter_65_0__60_));
AND2X2 AND2X2_564 ( .A(_abc_4268_new_n1470_), .B(counter_60_), .Y(_0counter_65_0__61_));
AND2X2 AND2X2_565 ( .A(_abc_4268_new_n1470_), .B(counter_61_), .Y(_0counter_65_0__62_));
AND2X2 AND2X2_566 ( .A(_abc_4268_new_n1470_), .B(counter_62_), .Y(_0counter_65_0__63_));
AND2X2 AND2X2_567 ( .A(_abc_4268_new_n1470_), .B(counter_63_), .Y(_0counter_65_0__64_));
AND2X2 AND2X2_568 ( .A(_abc_4268_new_n1470_), .B(counter_64_), .Y(_0counter_65_0__65_));
AND2X2 AND2X2_569 ( .A(_abc_4268_new_n625_), .B(_abc_4268_new_n1084_), .Y(_abc_4268_new_n1537_));
AND2X2 AND2X2_57 ( .A(_abc_4268_new_n709_), .B(RST), .Y(_abc_4268_new_n710_));
AND2X2 AND2X2_570 ( .A(_abc_4268_new_n1540_), .B(RST), .Y(_abc_4268_new_n1541_));
AND2X2 AND2X2_571 ( .A(_abc_4268_new_n1541_), .B(_abc_4268_new_n1539_), .Y(_0PICORV_RST_SPI_0_0_));
AND2X2 AND2X2_572 ( .A(RST), .B(re), .Y(_abc_4268_new_n1544_));
AND2X2 AND2X2_573 ( .A(_abc_4268_new_n1545_), .B(_abc_4268_new_n1543_), .Y(_0re_0_0_));
AND2X2 AND2X2_574 ( .A(RST), .B(we), .Y(_abc_4268_new_n1549_));
AND2X2 AND2X2_575 ( .A(_abc_4268_new_n1550_), .B(_abc_4268_new_n1548_), .Y(_0we_0_0_));
AND2X2 AND2X2_576 ( .A(_abc_4268_new_n591_), .B(axi_rvalid), .Y(_abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_479));
AND2X2 AND2X2_577 ( .A(_abc_4268_new_n561_), .B(axi_bvalid), .Y(_abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_430));
AND2X2 AND2X2_578 ( .A(RST), .B(counter_65_), .Y(_0fini_spi_0_0_));
AND2X2 AND2X2_579 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_0_), .Y(bus_sync_axi_bus__abc_3879_new_n394_));
AND2X2 AND2X2_58 ( .A(_abc_4268_new_n705_), .B(_abc_4268_new_n710_), .Y(_0bus_cap_31_0__1_));
AND2X2 AND2X2_580 ( .A(bus_sync_axi_bus_reg_data1_0_), .B(bus_sync_axi_bus_EECLK1), .Y(bus_sync_axi_bus__abc_3879_new_n395_));
AND2X2 AND2X2_581 ( .A(bus_sync_axi_bus__abc_3879_new_n396_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__0_));
AND2X2 AND2X2_582 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_1_), .Y(bus_sync_axi_bus__abc_3879_new_n398_));
AND2X2 AND2X2_583 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_1_), .Y(bus_sync_axi_bus__abc_3879_new_n399_));
AND2X2 AND2X2_584 ( .A(bus_sync_axi_bus__abc_3879_new_n400_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__1_));
AND2X2 AND2X2_585 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_2_), .Y(bus_sync_axi_bus__abc_3879_new_n402_));
AND2X2 AND2X2_586 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_2_), .Y(bus_sync_axi_bus__abc_3879_new_n403_));
AND2X2 AND2X2_587 ( .A(bus_sync_axi_bus__abc_3879_new_n404_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__2_));
AND2X2 AND2X2_588 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_3_), .Y(bus_sync_axi_bus__abc_3879_new_n406_));
AND2X2 AND2X2_589 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_3_), .Y(bus_sync_axi_bus__abc_3879_new_n407_));
AND2X2 AND2X2_59 ( .A(_abc_4268_new_n712_), .B(_abc_4268_new_n713_), .Y(_abc_4268_new_n714_));
AND2X2 AND2X2_590 ( .A(bus_sync_axi_bus__abc_3879_new_n408_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__3_));
AND2X2 AND2X2_591 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_4_), .Y(bus_sync_axi_bus__abc_3879_new_n410_));
AND2X2 AND2X2_592 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_4_), .Y(bus_sync_axi_bus__abc_3879_new_n411_));
AND2X2 AND2X2_593 ( .A(bus_sync_axi_bus__abc_3879_new_n412_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__4_));
AND2X2 AND2X2_594 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_5_), .Y(bus_sync_axi_bus__abc_3879_new_n414_));
AND2X2 AND2X2_595 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_5_), .Y(bus_sync_axi_bus__abc_3879_new_n415_));
AND2X2 AND2X2_596 ( .A(bus_sync_axi_bus__abc_3879_new_n416_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__5_));
AND2X2 AND2X2_597 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_6_), .Y(bus_sync_axi_bus__abc_3879_new_n418_));
AND2X2 AND2X2_598 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_6_), .Y(bus_sync_axi_bus__abc_3879_new_n419_));
AND2X2 AND2X2_599 ( .A(bus_sync_axi_bus__abc_3879_new_n420_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__6_));
AND2X2 AND2X2_6 ( .A(state_5_), .B(axi_awready), .Y(_abc_4268_new_n568_));
AND2X2 AND2X2_60 ( .A(_abc_4268_new_n617_), .B(bus_sync_status_data_out_2_), .Y(_abc_4268_new_n716_));
AND2X2 AND2X2_600 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_7_), .Y(bus_sync_axi_bus__abc_3879_new_n422_));
AND2X2 AND2X2_601 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_7_), .Y(bus_sync_axi_bus__abc_3879_new_n423_));
AND2X2 AND2X2_602 ( .A(bus_sync_axi_bus__abc_3879_new_n424_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__7_));
AND2X2 AND2X2_603 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_8_), .Y(bus_sync_axi_bus__abc_3879_new_n426_));
AND2X2 AND2X2_604 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_8_), .Y(bus_sync_axi_bus__abc_3879_new_n427_));
AND2X2 AND2X2_605 ( .A(bus_sync_axi_bus__abc_3879_new_n428_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__8_));
AND2X2 AND2X2_606 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_9_), .Y(bus_sync_axi_bus__abc_3879_new_n430_));
AND2X2 AND2X2_607 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_9_), .Y(bus_sync_axi_bus__abc_3879_new_n431_));
AND2X2 AND2X2_608 ( .A(bus_sync_axi_bus__abc_3879_new_n432_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__9_));
AND2X2 AND2X2_609 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_10_), .Y(bus_sync_axi_bus__abc_3879_new_n434_));
AND2X2 AND2X2_61 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_2_), .Y(_abc_4268_new_n717_));
AND2X2 AND2X2_610 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_10_), .Y(bus_sync_axi_bus__abc_3879_new_n435_));
AND2X2 AND2X2_611 ( .A(bus_sync_axi_bus__abc_3879_new_n436_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__10_));
AND2X2 AND2X2_612 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_11_), .Y(bus_sync_axi_bus__abc_3879_new_n438_));
AND2X2 AND2X2_613 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_11_), .Y(bus_sync_axi_bus__abc_3879_new_n439_));
AND2X2 AND2X2_614 ( .A(bus_sync_axi_bus__abc_3879_new_n440_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__11_));
AND2X2 AND2X2_615 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_12_), .Y(bus_sync_axi_bus__abc_3879_new_n442_));
AND2X2 AND2X2_616 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_12_), .Y(bus_sync_axi_bus__abc_3879_new_n443_));
AND2X2 AND2X2_617 ( .A(bus_sync_axi_bus__abc_3879_new_n444_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__12_));
AND2X2 AND2X2_618 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_13_), .Y(bus_sync_axi_bus__abc_3879_new_n446_));
AND2X2 AND2X2_619 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_13_), .Y(bus_sync_axi_bus__abc_3879_new_n447_));
AND2X2 AND2X2_62 ( .A(_abc_4268_new_n719_), .B(RST), .Y(_abc_4268_new_n720_));
AND2X2 AND2X2_620 ( .A(bus_sync_axi_bus__abc_3879_new_n448_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__13_));
AND2X2 AND2X2_621 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_14_), .Y(bus_sync_axi_bus__abc_3879_new_n450_));
AND2X2 AND2X2_622 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_14_), .Y(bus_sync_axi_bus__abc_3879_new_n451_));
AND2X2 AND2X2_623 ( .A(bus_sync_axi_bus__abc_3879_new_n452_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__14_));
AND2X2 AND2X2_624 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_15_), .Y(bus_sync_axi_bus__abc_3879_new_n454_));
AND2X2 AND2X2_625 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_15_), .Y(bus_sync_axi_bus__abc_3879_new_n455_));
AND2X2 AND2X2_626 ( .A(bus_sync_axi_bus__abc_3879_new_n456_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__15_));
AND2X2 AND2X2_627 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_16_), .Y(bus_sync_axi_bus__abc_3879_new_n458_));
AND2X2 AND2X2_628 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_16_), .Y(bus_sync_axi_bus__abc_3879_new_n459_));
AND2X2 AND2X2_629 ( .A(bus_sync_axi_bus__abc_3879_new_n460_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__16_));
AND2X2 AND2X2_63 ( .A(_abc_4268_new_n715_), .B(_abc_4268_new_n720_), .Y(_0bus_cap_31_0__2_));
AND2X2 AND2X2_630 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_17_), .Y(bus_sync_axi_bus__abc_3879_new_n462_));
AND2X2 AND2X2_631 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_17_), .Y(bus_sync_axi_bus__abc_3879_new_n463_));
AND2X2 AND2X2_632 ( .A(bus_sync_axi_bus__abc_3879_new_n464_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__17_));
AND2X2 AND2X2_633 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_18_), .Y(bus_sync_axi_bus__abc_3879_new_n466_));
AND2X2 AND2X2_634 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_18_), .Y(bus_sync_axi_bus__abc_3879_new_n467_));
AND2X2 AND2X2_635 ( .A(bus_sync_axi_bus__abc_3879_new_n468_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__18_));
AND2X2 AND2X2_636 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_19_), .Y(bus_sync_axi_bus__abc_3879_new_n470_));
AND2X2 AND2X2_637 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_19_), .Y(bus_sync_axi_bus__abc_3879_new_n471_));
AND2X2 AND2X2_638 ( .A(bus_sync_axi_bus__abc_3879_new_n472_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__19_));
AND2X2 AND2X2_639 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_20_), .Y(bus_sync_axi_bus__abc_3879_new_n474_));
AND2X2 AND2X2_64 ( .A(_abc_4268_new_n722_), .B(_abc_4268_new_n723_), .Y(_abc_4268_new_n724_));
AND2X2 AND2X2_640 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_20_), .Y(bus_sync_axi_bus__abc_3879_new_n475_));
AND2X2 AND2X2_641 ( .A(bus_sync_axi_bus__abc_3879_new_n476_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__20_));
AND2X2 AND2X2_642 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_21_), .Y(bus_sync_axi_bus__abc_3879_new_n478_));
AND2X2 AND2X2_643 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_21_), .Y(bus_sync_axi_bus__abc_3879_new_n479_));
AND2X2 AND2X2_644 ( .A(bus_sync_axi_bus__abc_3879_new_n480_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__21_));
AND2X2 AND2X2_645 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_22_), .Y(bus_sync_axi_bus__abc_3879_new_n482_));
AND2X2 AND2X2_646 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_22_), .Y(bus_sync_axi_bus__abc_3879_new_n483_));
AND2X2 AND2X2_647 ( .A(bus_sync_axi_bus__abc_3879_new_n484_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__22_));
AND2X2 AND2X2_648 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_23_), .Y(bus_sync_axi_bus__abc_3879_new_n486_));
AND2X2 AND2X2_649 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_23_), .Y(bus_sync_axi_bus__abc_3879_new_n487_));
AND2X2 AND2X2_65 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_3_), .Y(_abc_4268_new_n726_));
AND2X2 AND2X2_650 ( .A(bus_sync_axi_bus__abc_3879_new_n488_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__23_));
AND2X2 AND2X2_651 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_24_), .Y(bus_sync_axi_bus__abc_3879_new_n490_));
AND2X2 AND2X2_652 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_24_), .Y(bus_sync_axi_bus__abc_3879_new_n491_));
AND2X2 AND2X2_653 ( .A(bus_sync_axi_bus__abc_3879_new_n492_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__24_));
AND2X2 AND2X2_654 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_25_), .Y(bus_sync_axi_bus__abc_3879_new_n494_));
AND2X2 AND2X2_655 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_25_), .Y(bus_sync_axi_bus__abc_3879_new_n495_));
AND2X2 AND2X2_656 ( .A(bus_sync_axi_bus__abc_3879_new_n496_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__25_));
AND2X2 AND2X2_657 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_26_), .Y(bus_sync_axi_bus__abc_3879_new_n498_));
AND2X2 AND2X2_658 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_26_), .Y(bus_sync_axi_bus__abc_3879_new_n499_));
AND2X2 AND2X2_659 ( .A(bus_sync_axi_bus__abc_3879_new_n500_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__26_));
AND2X2 AND2X2_66 ( .A(_abc_4268_new_n727_), .B(RST), .Y(_abc_4268_new_n728_));
AND2X2 AND2X2_660 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_27_), .Y(bus_sync_axi_bus__abc_3879_new_n502_));
AND2X2 AND2X2_661 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_27_), .Y(bus_sync_axi_bus__abc_3879_new_n503_));
AND2X2 AND2X2_662 ( .A(bus_sync_axi_bus__abc_3879_new_n504_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__27_));
AND2X2 AND2X2_663 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_28_), .Y(bus_sync_axi_bus__abc_3879_new_n506_));
AND2X2 AND2X2_664 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_28_), .Y(bus_sync_axi_bus__abc_3879_new_n507_));
AND2X2 AND2X2_665 ( .A(bus_sync_axi_bus__abc_3879_new_n508_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__28_));
AND2X2 AND2X2_666 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_29_), .Y(bus_sync_axi_bus__abc_3879_new_n510_));
AND2X2 AND2X2_667 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_29_), .Y(bus_sync_axi_bus__abc_3879_new_n511_));
AND2X2 AND2X2_668 ( .A(bus_sync_axi_bus__abc_3879_new_n512_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__29_));
AND2X2 AND2X2_669 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_30_), .Y(bus_sync_axi_bus__abc_3879_new_n514_));
AND2X2 AND2X2_67 ( .A(_abc_4268_new_n725_), .B(_abc_4268_new_n728_), .Y(_0bus_cap_31_0__3_));
AND2X2 AND2X2_670 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_30_), .Y(bus_sync_axi_bus__abc_3879_new_n515_));
AND2X2 AND2X2_671 ( .A(bus_sync_axi_bus__abc_3879_new_n516_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__30_));
AND2X2 AND2X2_672 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_31_), .Y(bus_sync_axi_bus__abc_3879_new_n518_));
AND2X2 AND2X2_673 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_31_), .Y(bus_sync_axi_bus__abc_3879_new_n519_));
AND2X2 AND2X2_674 ( .A(bus_sync_axi_bus__abc_3879_new_n520_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__31_));
AND2X2 AND2X2_675 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_32_), .Y(bus_sync_axi_bus__abc_3879_new_n522_));
AND2X2 AND2X2_676 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_32_), .Y(bus_sync_axi_bus__abc_3879_new_n523_));
AND2X2 AND2X2_677 ( .A(bus_sync_axi_bus__abc_3879_new_n524_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__32_));
AND2X2 AND2X2_678 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_33_), .Y(bus_sync_axi_bus__abc_3879_new_n526_));
AND2X2 AND2X2_679 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_33_), .Y(bus_sync_axi_bus__abc_3879_new_n527_));
AND2X2 AND2X2_68 ( .A(_abc_4268_new_n730_), .B(_abc_4268_new_n731_), .Y(_abc_4268_new_n732_));
AND2X2 AND2X2_680 ( .A(bus_sync_axi_bus__abc_3879_new_n528_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__33_));
AND2X2 AND2X2_681 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_34_), .Y(bus_sync_axi_bus__abc_3879_new_n530_));
AND2X2 AND2X2_682 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_34_), .Y(bus_sync_axi_bus__abc_3879_new_n531_));
AND2X2 AND2X2_683 ( .A(bus_sync_axi_bus__abc_3879_new_n532_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__34_));
AND2X2 AND2X2_684 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_35_), .Y(bus_sync_axi_bus__abc_3879_new_n534_));
AND2X2 AND2X2_685 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_35_), .Y(bus_sync_axi_bus__abc_3879_new_n535_));
AND2X2 AND2X2_686 ( .A(bus_sync_axi_bus__abc_3879_new_n536_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__35_));
AND2X2 AND2X2_687 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_36_), .Y(bus_sync_axi_bus__abc_3879_new_n538_));
AND2X2 AND2X2_688 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_36_), .Y(bus_sync_axi_bus__abc_3879_new_n539_));
AND2X2 AND2X2_689 ( .A(bus_sync_axi_bus__abc_3879_new_n540_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__36_));
AND2X2 AND2X2_69 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_4_), .Y(_abc_4268_new_n734_));
AND2X2 AND2X2_690 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_37_), .Y(bus_sync_axi_bus__abc_3879_new_n542_));
AND2X2 AND2X2_691 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_37_), .Y(bus_sync_axi_bus__abc_3879_new_n543_));
AND2X2 AND2X2_692 ( .A(bus_sync_axi_bus__abc_3879_new_n544_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__37_));
AND2X2 AND2X2_693 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_38_), .Y(bus_sync_axi_bus__abc_3879_new_n546_));
AND2X2 AND2X2_694 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_38_), .Y(bus_sync_axi_bus__abc_3879_new_n547_));
AND2X2 AND2X2_695 ( .A(bus_sync_axi_bus__abc_3879_new_n548_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__38_));
AND2X2 AND2X2_696 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_39_), .Y(bus_sync_axi_bus__abc_3879_new_n550_));
AND2X2 AND2X2_697 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_39_), .Y(bus_sync_axi_bus__abc_3879_new_n551_));
AND2X2 AND2X2_698 ( .A(bus_sync_axi_bus__abc_3879_new_n552_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__39_));
AND2X2 AND2X2_699 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_40_), .Y(bus_sync_axi_bus__abc_3879_new_n554_));
AND2X2 AND2X2_7 ( .A(_abc_4268_new_n569_), .B(RST), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_3_));
AND2X2 AND2X2_70 ( .A(_abc_4268_new_n735_), .B(RST), .Y(_abc_4268_new_n736_));
AND2X2 AND2X2_700 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_40_), .Y(bus_sync_axi_bus__abc_3879_new_n555_));
AND2X2 AND2X2_701 ( .A(bus_sync_axi_bus__abc_3879_new_n556_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__40_));
AND2X2 AND2X2_702 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_41_), .Y(bus_sync_axi_bus__abc_3879_new_n558_));
AND2X2 AND2X2_703 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_41_), .Y(bus_sync_axi_bus__abc_3879_new_n559_));
AND2X2 AND2X2_704 ( .A(bus_sync_axi_bus__abc_3879_new_n560_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__41_));
AND2X2 AND2X2_705 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_42_), .Y(bus_sync_axi_bus__abc_3879_new_n562_));
AND2X2 AND2X2_706 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_42_), .Y(bus_sync_axi_bus__abc_3879_new_n563_));
AND2X2 AND2X2_707 ( .A(bus_sync_axi_bus__abc_3879_new_n564_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__42_));
AND2X2 AND2X2_708 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_43_), .Y(bus_sync_axi_bus__abc_3879_new_n566_));
AND2X2 AND2X2_709 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_43_), .Y(bus_sync_axi_bus__abc_3879_new_n567_));
AND2X2 AND2X2_71 ( .A(_abc_4268_new_n733_), .B(_abc_4268_new_n736_), .Y(_0bus_cap_31_0__4_));
AND2X2 AND2X2_710 ( .A(bus_sync_axi_bus__abc_3879_new_n568_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__43_));
AND2X2 AND2X2_711 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_44_), .Y(bus_sync_axi_bus__abc_3879_new_n570_));
AND2X2 AND2X2_712 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_44_), .Y(bus_sync_axi_bus__abc_3879_new_n571_));
AND2X2 AND2X2_713 ( .A(bus_sync_axi_bus__abc_3879_new_n572_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__44_));
AND2X2 AND2X2_714 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_45_), .Y(bus_sync_axi_bus__abc_3879_new_n574_));
AND2X2 AND2X2_715 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_45_), .Y(bus_sync_axi_bus__abc_3879_new_n575_));
AND2X2 AND2X2_716 ( .A(bus_sync_axi_bus__abc_3879_new_n576_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__45_));
AND2X2 AND2X2_717 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_46_), .Y(bus_sync_axi_bus__abc_3879_new_n578_));
AND2X2 AND2X2_718 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_46_), .Y(bus_sync_axi_bus__abc_3879_new_n579_));
AND2X2 AND2X2_719 ( .A(bus_sync_axi_bus__abc_3879_new_n580_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__46_));
AND2X2 AND2X2_72 ( .A(_abc_4268_new_n738_), .B(_abc_4268_new_n739_), .Y(_abc_4268_new_n740_));
AND2X2 AND2X2_720 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_47_), .Y(bus_sync_axi_bus__abc_3879_new_n582_));
AND2X2 AND2X2_721 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_47_), .Y(bus_sync_axi_bus__abc_3879_new_n583_));
AND2X2 AND2X2_722 ( .A(bus_sync_axi_bus__abc_3879_new_n584_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__47_));
AND2X2 AND2X2_723 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_48_), .Y(bus_sync_axi_bus__abc_3879_new_n586_));
AND2X2 AND2X2_724 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_48_), .Y(bus_sync_axi_bus__abc_3879_new_n587_));
AND2X2 AND2X2_725 ( .A(bus_sync_axi_bus__abc_3879_new_n588_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__48_));
AND2X2 AND2X2_726 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_49_), .Y(bus_sync_axi_bus__abc_3879_new_n590_));
AND2X2 AND2X2_727 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_49_), .Y(bus_sync_axi_bus__abc_3879_new_n591_));
AND2X2 AND2X2_728 ( .A(bus_sync_axi_bus__abc_3879_new_n592_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__49_));
AND2X2 AND2X2_729 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_50_), .Y(bus_sync_axi_bus__abc_3879_new_n594_));
AND2X2 AND2X2_73 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_5_), .Y(_abc_4268_new_n742_));
AND2X2 AND2X2_730 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_50_), .Y(bus_sync_axi_bus__abc_3879_new_n595_));
AND2X2 AND2X2_731 ( .A(bus_sync_axi_bus__abc_3879_new_n596_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__50_));
AND2X2 AND2X2_732 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_51_), .Y(bus_sync_axi_bus__abc_3879_new_n598_));
AND2X2 AND2X2_733 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_51_), .Y(bus_sync_axi_bus__abc_3879_new_n599_));
AND2X2 AND2X2_734 ( .A(bus_sync_axi_bus__abc_3879_new_n600_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__51_));
AND2X2 AND2X2_735 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_52_), .Y(bus_sync_axi_bus__abc_3879_new_n602_));
AND2X2 AND2X2_736 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_52_), .Y(bus_sync_axi_bus__abc_3879_new_n603_));
AND2X2 AND2X2_737 ( .A(bus_sync_axi_bus__abc_3879_new_n604_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__52_));
AND2X2 AND2X2_738 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_53_), .Y(bus_sync_axi_bus__abc_3879_new_n606_));
AND2X2 AND2X2_739 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_53_), .Y(bus_sync_axi_bus__abc_3879_new_n607_));
AND2X2 AND2X2_74 ( .A(_abc_4268_new_n743_), .B(RST), .Y(_abc_4268_new_n744_));
AND2X2 AND2X2_740 ( .A(bus_sync_axi_bus__abc_3879_new_n608_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__53_));
AND2X2 AND2X2_741 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_54_), .Y(bus_sync_axi_bus__abc_3879_new_n610_));
AND2X2 AND2X2_742 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_54_), .Y(bus_sync_axi_bus__abc_3879_new_n611_));
AND2X2 AND2X2_743 ( .A(bus_sync_axi_bus__abc_3879_new_n612_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__54_));
AND2X2 AND2X2_744 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_55_), .Y(bus_sync_axi_bus__abc_3879_new_n614_));
AND2X2 AND2X2_745 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_55_), .Y(bus_sync_axi_bus__abc_3879_new_n615_));
AND2X2 AND2X2_746 ( .A(bus_sync_axi_bus__abc_3879_new_n616_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__55_));
AND2X2 AND2X2_747 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_56_), .Y(bus_sync_axi_bus__abc_3879_new_n618_));
AND2X2 AND2X2_748 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_56_), .Y(bus_sync_axi_bus__abc_3879_new_n619_));
AND2X2 AND2X2_749 ( .A(bus_sync_axi_bus__abc_3879_new_n620_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__56_));
AND2X2 AND2X2_75 ( .A(_abc_4268_new_n741_), .B(_abc_4268_new_n744_), .Y(_0bus_cap_31_0__5_));
AND2X2 AND2X2_750 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_57_), .Y(bus_sync_axi_bus__abc_3879_new_n622_));
AND2X2 AND2X2_751 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_57_), .Y(bus_sync_axi_bus__abc_3879_new_n623_));
AND2X2 AND2X2_752 ( .A(bus_sync_axi_bus__abc_3879_new_n624_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__57_));
AND2X2 AND2X2_753 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_58_), .Y(bus_sync_axi_bus__abc_3879_new_n626_));
AND2X2 AND2X2_754 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_58_), .Y(bus_sync_axi_bus__abc_3879_new_n627_));
AND2X2 AND2X2_755 ( .A(bus_sync_axi_bus__abc_3879_new_n628_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__58_));
AND2X2 AND2X2_756 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_59_), .Y(bus_sync_axi_bus__abc_3879_new_n630_));
AND2X2 AND2X2_757 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_59_), .Y(bus_sync_axi_bus__abc_3879_new_n631_));
AND2X2 AND2X2_758 ( .A(bus_sync_axi_bus__abc_3879_new_n632_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__59_));
AND2X2 AND2X2_759 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_60_), .Y(bus_sync_axi_bus__abc_3879_new_n634_));
AND2X2 AND2X2_76 ( .A(_abc_4268_new_n746_), .B(_abc_4268_new_n747_), .Y(_abc_4268_new_n748_));
AND2X2 AND2X2_760 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_60_), .Y(bus_sync_axi_bus__abc_3879_new_n635_));
AND2X2 AND2X2_761 ( .A(bus_sync_axi_bus__abc_3879_new_n636_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__60_));
AND2X2 AND2X2_762 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_61_), .Y(bus_sync_axi_bus__abc_3879_new_n638_));
AND2X2 AND2X2_763 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_61_), .Y(bus_sync_axi_bus__abc_3879_new_n639_));
AND2X2 AND2X2_764 ( .A(bus_sync_axi_bus__abc_3879_new_n640_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__61_));
AND2X2 AND2X2_765 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_62_), .Y(bus_sync_axi_bus__abc_3879_new_n642_));
AND2X2 AND2X2_766 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_62_), .Y(bus_sync_axi_bus__abc_3879_new_n643_));
AND2X2 AND2X2_767 ( .A(bus_sync_axi_bus__abc_3879_new_n644_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__62_));
AND2X2 AND2X2_768 ( .A(bus_sync_axi_bus__abc_3879_new_n393_), .B(bus_sync_axi_bus_reg_data2_63_), .Y(bus_sync_axi_bus__abc_3879_new_n646_));
AND2X2 AND2X2_769 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_63_), .Y(bus_sync_axi_bus__abc_3879_new_n647_));
AND2X2 AND2X2_77 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_6_), .Y(_abc_4268_new_n750_));
AND2X2 AND2X2_770 ( .A(bus_sync_axi_bus__abc_3879_new_n648_), .B(RST), .Y(bus_sync_axi_bus__0reg_data2_63_0__63_));
AND2X2 AND2X2_771 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_0_), .Y(bus_sync_axi_bus__0reg_data3_63_0__0_));
AND2X2 AND2X2_772 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_1_), .Y(bus_sync_axi_bus__0reg_data3_63_0__1_));
AND2X2 AND2X2_773 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_2_), .Y(bus_sync_axi_bus__0reg_data3_63_0__2_));
AND2X2 AND2X2_774 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_3_), .Y(bus_sync_axi_bus__0reg_data3_63_0__3_));
AND2X2 AND2X2_775 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_4_), .Y(bus_sync_axi_bus__0reg_data3_63_0__4_));
AND2X2 AND2X2_776 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_5_), .Y(bus_sync_axi_bus__0reg_data3_63_0__5_));
AND2X2 AND2X2_777 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_6_), .Y(bus_sync_axi_bus__0reg_data3_63_0__6_));
AND2X2 AND2X2_778 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_7_), .Y(bus_sync_axi_bus__0reg_data3_63_0__7_));
AND2X2 AND2X2_779 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_8_), .Y(bus_sync_axi_bus__0reg_data3_63_0__8_));
AND2X2 AND2X2_78 ( .A(_abc_4268_new_n751_), .B(RST), .Y(_abc_4268_new_n752_));
AND2X2 AND2X2_780 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_9_), .Y(bus_sync_axi_bus__0reg_data3_63_0__9_));
AND2X2 AND2X2_781 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_10_), .Y(bus_sync_axi_bus__0reg_data3_63_0__10_));
AND2X2 AND2X2_782 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_11_), .Y(bus_sync_axi_bus__0reg_data3_63_0__11_));
AND2X2 AND2X2_783 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_12_), .Y(bus_sync_axi_bus__0reg_data3_63_0__12_));
AND2X2 AND2X2_784 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_13_), .Y(bus_sync_axi_bus__0reg_data3_63_0__13_));
AND2X2 AND2X2_785 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_14_), .Y(bus_sync_axi_bus__0reg_data3_63_0__14_));
AND2X2 AND2X2_786 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_15_), .Y(bus_sync_axi_bus__0reg_data3_63_0__15_));
AND2X2 AND2X2_787 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_16_), .Y(bus_sync_axi_bus__0reg_data3_63_0__16_));
AND2X2 AND2X2_788 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_17_), .Y(bus_sync_axi_bus__0reg_data3_63_0__17_));
AND2X2 AND2X2_789 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_18_), .Y(bus_sync_axi_bus__0reg_data3_63_0__18_));
AND2X2 AND2X2_79 ( .A(_abc_4268_new_n749_), .B(_abc_4268_new_n752_), .Y(_0bus_cap_31_0__6_));
AND2X2 AND2X2_790 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_19_), .Y(bus_sync_axi_bus__0reg_data3_63_0__19_));
AND2X2 AND2X2_791 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_20_), .Y(bus_sync_axi_bus__0reg_data3_63_0__20_));
AND2X2 AND2X2_792 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_21_), .Y(bus_sync_axi_bus__0reg_data3_63_0__21_));
AND2X2 AND2X2_793 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_22_), .Y(bus_sync_axi_bus__0reg_data3_63_0__22_));
AND2X2 AND2X2_794 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_23_), .Y(bus_sync_axi_bus__0reg_data3_63_0__23_));
AND2X2 AND2X2_795 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_24_), .Y(bus_sync_axi_bus__0reg_data3_63_0__24_));
AND2X2 AND2X2_796 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_25_), .Y(bus_sync_axi_bus__0reg_data3_63_0__25_));
AND2X2 AND2X2_797 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_26_), .Y(bus_sync_axi_bus__0reg_data3_63_0__26_));
AND2X2 AND2X2_798 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_27_), .Y(bus_sync_axi_bus__0reg_data3_63_0__27_));
AND2X2 AND2X2_799 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_28_), .Y(bus_sync_axi_bus__0reg_data3_63_0__28_));
AND2X2 AND2X2_8 ( .A(state_1_), .B(fini_spi_clk), .Y(_abc_4268_new_n572_));
AND2X2 AND2X2_80 ( .A(_abc_4268_new_n754_), .B(_abc_4268_new_n755_), .Y(_abc_4268_new_n756_));
AND2X2 AND2X2_800 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_29_), .Y(bus_sync_axi_bus__0reg_data3_63_0__29_));
AND2X2 AND2X2_801 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_30_), .Y(bus_sync_axi_bus__0reg_data3_63_0__30_));
AND2X2 AND2X2_802 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_31_), .Y(bus_sync_axi_bus__0reg_data3_63_0__31_));
AND2X2 AND2X2_803 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_32_), .Y(bus_sync_axi_bus__0reg_data3_63_0__32_));
AND2X2 AND2X2_804 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_33_), .Y(bus_sync_axi_bus__0reg_data3_63_0__33_));
AND2X2 AND2X2_805 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_34_), .Y(bus_sync_axi_bus__0reg_data3_63_0__34_));
AND2X2 AND2X2_806 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_35_), .Y(bus_sync_axi_bus__0reg_data3_63_0__35_));
AND2X2 AND2X2_807 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_36_), .Y(bus_sync_axi_bus__0reg_data3_63_0__36_));
AND2X2 AND2X2_808 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_37_), .Y(bus_sync_axi_bus__0reg_data3_63_0__37_));
AND2X2 AND2X2_809 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_38_), .Y(bus_sync_axi_bus__0reg_data3_63_0__38_));
AND2X2 AND2X2_81 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_7_), .Y(_abc_4268_new_n758_));
AND2X2 AND2X2_810 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_39_), .Y(bus_sync_axi_bus__0reg_data3_63_0__39_));
AND2X2 AND2X2_811 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_40_), .Y(bus_sync_axi_bus__0reg_data3_63_0__40_));
AND2X2 AND2X2_812 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_41_), .Y(bus_sync_axi_bus__0reg_data3_63_0__41_));
AND2X2 AND2X2_813 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_42_), .Y(bus_sync_axi_bus__0reg_data3_63_0__42_));
AND2X2 AND2X2_814 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_43_), .Y(bus_sync_axi_bus__0reg_data3_63_0__43_));
AND2X2 AND2X2_815 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_44_), .Y(bus_sync_axi_bus__0reg_data3_63_0__44_));
AND2X2 AND2X2_816 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_45_), .Y(bus_sync_axi_bus__0reg_data3_63_0__45_));
AND2X2 AND2X2_817 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_46_), .Y(bus_sync_axi_bus__0reg_data3_63_0__46_));
AND2X2 AND2X2_818 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_47_), .Y(bus_sync_axi_bus__0reg_data3_63_0__47_));
AND2X2 AND2X2_819 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_48_), .Y(bus_sync_axi_bus__0reg_data3_63_0__48_));
AND2X2 AND2X2_82 ( .A(_abc_4268_new_n759_), .B(RST), .Y(_abc_4268_new_n760_));
AND2X2 AND2X2_820 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_49_), .Y(bus_sync_axi_bus__0reg_data3_63_0__49_));
AND2X2 AND2X2_821 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_50_), .Y(bus_sync_axi_bus__0reg_data3_63_0__50_));
AND2X2 AND2X2_822 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_51_), .Y(bus_sync_axi_bus__0reg_data3_63_0__51_));
AND2X2 AND2X2_823 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_52_), .Y(bus_sync_axi_bus__0reg_data3_63_0__52_));
AND2X2 AND2X2_824 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_53_), .Y(bus_sync_axi_bus__0reg_data3_63_0__53_));
AND2X2 AND2X2_825 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_54_), .Y(bus_sync_axi_bus__0reg_data3_63_0__54_));
AND2X2 AND2X2_826 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_55_), .Y(bus_sync_axi_bus__0reg_data3_63_0__55_));
AND2X2 AND2X2_827 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_56_), .Y(bus_sync_axi_bus__0reg_data3_63_0__56_));
AND2X2 AND2X2_828 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_57_), .Y(bus_sync_axi_bus__0reg_data3_63_0__57_));
AND2X2 AND2X2_829 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_58_), .Y(bus_sync_axi_bus__0reg_data3_63_0__58_));
AND2X2 AND2X2_83 ( .A(_abc_4268_new_n757_), .B(_abc_4268_new_n760_), .Y(_0bus_cap_31_0__7_));
AND2X2 AND2X2_830 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_59_), .Y(bus_sync_axi_bus__0reg_data3_63_0__59_));
AND2X2 AND2X2_831 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_60_), .Y(bus_sync_axi_bus__0reg_data3_63_0__60_));
AND2X2 AND2X2_832 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_61_), .Y(bus_sync_axi_bus__0reg_data3_63_0__61_));
AND2X2 AND2X2_833 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_62_), .Y(bus_sync_axi_bus__0reg_data3_63_0__62_));
AND2X2 AND2X2_834 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_63_), .Y(bus_sync_axi_bus__0reg_data3_63_0__63_));
AND2X2 AND2X2_835 ( .A(RST), .B(WDATA_0_), .Y(bus_sync_axi_bus__0reg_data1_63_0__0_));
AND2X2 AND2X2_836 ( .A(RST), .B(WDATA_1_), .Y(bus_sync_axi_bus__0reg_data1_63_0__1_));
AND2X2 AND2X2_837 ( .A(RST), .B(WDATA_2_), .Y(bus_sync_axi_bus__0reg_data1_63_0__2_));
AND2X2 AND2X2_838 ( .A(RST), .B(WDATA_3_), .Y(bus_sync_axi_bus__0reg_data1_63_0__3_));
AND2X2 AND2X2_839 ( .A(RST), .B(WDATA_4_), .Y(bus_sync_axi_bus__0reg_data1_63_0__4_));
AND2X2 AND2X2_84 ( .A(_abc_4268_new_n762_), .B(_abc_4268_new_n763_), .Y(_abc_4268_new_n764_));
AND2X2 AND2X2_840 ( .A(RST), .B(WDATA_5_), .Y(bus_sync_axi_bus__0reg_data1_63_0__5_));
AND2X2 AND2X2_841 ( .A(RST), .B(WDATA_6_), .Y(bus_sync_axi_bus__0reg_data1_63_0__6_));
AND2X2 AND2X2_842 ( .A(RST), .B(WDATA_7_), .Y(bus_sync_axi_bus__0reg_data1_63_0__7_));
AND2X2 AND2X2_843 ( .A(RST), .B(WDATA_8_), .Y(bus_sync_axi_bus__0reg_data1_63_0__8_));
AND2X2 AND2X2_844 ( .A(RST), .B(WDATA_9_), .Y(bus_sync_axi_bus__0reg_data1_63_0__9_));
AND2X2 AND2X2_845 ( .A(RST), .B(WDATA_10_), .Y(bus_sync_axi_bus__0reg_data1_63_0__10_));
AND2X2 AND2X2_846 ( .A(RST), .B(WDATA_11_), .Y(bus_sync_axi_bus__0reg_data1_63_0__11_));
AND2X2 AND2X2_847 ( .A(RST), .B(WDATA_12_), .Y(bus_sync_axi_bus__0reg_data1_63_0__12_));
AND2X2 AND2X2_848 ( .A(RST), .B(WDATA_13_), .Y(bus_sync_axi_bus__0reg_data1_63_0__13_));
AND2X2 AND2X2_849 ( .A(RST), .B(WDATA_14_), .Y(bus_sync_axi_bus__0reg_data1_63_0__14_));
AND2X2 AND2X2_85 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_8_), .Y(_abc_4268_new_n766_));
AND2X2 AND2X2_850 ( .A(RST), .B(WDATA_15_), .Y(bus_sync_axi_bus__0reg_data1_63_0__15_));
AND2X2 AND2X2_851 ( .A(RST), .B(WDATA_16_), .Y(bus_sync_axi_bus__0reg_data1_63_0__16_));
AND2X2 AND2X2_852 ( .A(RST), .B(WDATA_17_), .Y(bus_sync_axi_bus__0reg_data1_63_0__17_));
AND2X2 AND2X2_853 ( .A(RST), .B(WDATA_18_), .Y(bus_sync_axi_bus__0reg_data1_63_0__18_));
AND2X2 AND2X2_854 ( .A(RST), .B(WDATA_19_), .Y(bus_sync_axi_bus__0reg_data1_63_0__19_));
AND2X2 AND2X2_855 ( .A(RST), .B(WDATA_20_), .Y(bus_sync_axi_bus__0reg_data1_63_0__20_));
AND2X2 AND2X2_856 ( .A(RST), .B(WDATA_21_), .Y(bus_sync_axi_bus__0reg_data1_63_0__21_));
AND2X2 AND2X2_857 ( .A(RST), .B(WDATA_22_), .Y(bus_sync_axi_bus__0reg_data1_63_0__22_));
AND2X2 AND2X2_858 ( .A(RST), .B(WDATA_23_), .Y(bus_sync_axi_bus__0reg_data1_63_0__23_));
AND2X2 AND2X2_859 ( .A(RST), .B(WDATA_24_), .Y(bus_sync_axi_bus__0reg_data1_63_0__24_));
AND2X2 AND2X2_86 ( .A(_abc_4268_new_n767_), .B(RST), .Y(_abc_4268_new_n768_));
AND2X2 AND2X2_860 ( .A(RST), .B(WDATA_25_), .Y(bus_sync_axi_bus__0reg_data1_63_0__25_));
AND2X2 AND2X2_861 ( .A(RST), .B(WDATA_26_), .Y(bus_sync_axi_bus__0reg_data1_63_0__26_));
AND2X2 AND2X2_862 ( .A(RST), .B(WDATA_27_), .Y(bus_sync_axi_bus__0reg_data1_63_0__27_));
AND2X2 AND2X2_863 ( .A(RST), .B(WDATA_28_), .Y(bus_sync_axi_bus__0reg_data1_63_0__28_));
AND2X2 AND2X2_864 ( .A(RST), .B(WDATA_29_), .Y(bus_sync_axi_bus__0reg_data1_63_0__29_));
AND2X2 AND2X2_865 ( .A(RST), .B(WDATA_30_), .Y(bus_sync_axi_bus__0reg_data1_63_0__30_));
AND2X2 AND2X2_866 ( .A(RST), .B(WDATA_31_), .Y(bus_sync_axi_bus__0reg_data1_63_0__31_));
AND2X2 AND2X2_867 ( .A(RST), .B(A_ADDR_0_), .Y(bus_sync_axi_bus__0reg_data1_63_0__32_));
AND2X2 AND2X2_868 ( .A(RST), .B(A_ADDR_1_), .Y(bus_sync_axi_bus__0reg_data1_63_0__33_));
AND2X2 AND2X2_869 ( .A(RST), .B(A_ADDR_2_), .Y(bus_sync_axi_bus__0reg_data1_63_0__34_));
AND2X2 AND2X2_87 ( .A(_abc_4268_new_n765_), .B(_abc_4268_new_n768_), .Y(_0bus_cap_31_0__8_));
AND2X2 AND2X2_870 ( .A(RST), .B(A_ADDR_3_), .Y(bus_sync_axi_bus__0reg_data1_63_0__35_));
AND2X2 AND2X2_871 ( .A(RST), .B(A_ADDR_4_), .Y(bus_sync_axi_bus__0reg_data1_63_0__36_));
AND2X2 AND2X2_872 ( .A(RST), .B(A_ADDR_5_), .Y(bus_sync_axi_bus__0reg_data1_63_0__37_));
AND2X2 AND2X2_873 ( .A(RST), .B(A_ADDR_6_), .Y(bus_sync_axi_bus__0reg_data1_63_0__38_));
AND2X2 AND2X2_874 ( .A(RST), .B(A_ADDR_7_), .Y(bus_sync_axi_bus__0reg_data1_63_0__39_));
AND2X2 AND2X2_875 ( .A(RST), .B(A_ADDR_8_), .Y(bus_sync_axi_bus__0reg_data1_63_0__40_));
AND2X2 AND2X2_876 ( .A(RST), .B(A_ADDR_9_), .Y(bus_sync_axi_bus__0reg_data1_63_0__41_));
AND2X2 AND2X2_877 ( .A(RST), .B(A_ADDR_10_), .Y(bus_sync_axi_bus__0reg_data1_63_0__42_));
AND2X2 AND2X2_878 ( .A(RST), .B(A_ADDR_11_), .Y(bus_sync_axi_bus__0reg_data1_63_0__43_));
AND2X2 AND2X2_879 ( .A(RST), .B(A_ADDR_12_), .Y(bus_sync_axi_bus__0reg_data1_63_0__44_));
AND2X2 AND2X2_88 ( .A(_abc_4268_new_n770_), .B(_abc_4268_new_n771_), .Y(_abc_4268_new_n772_));
AND2X2 AND2X2_880 ( .A(RST), .B(A_ADDR_13_), .Y(bus_sync_axi_bus__0reg_data1_63_0__45_));
AND2X2 AND2X2_881 ( .A(RST), .B(A_ADDR_14_), .Y(bus_sync_axi_bus__0reg_data1_63_0__46_));
AND2X2 AND2X2_882 ( .A(RST), .B(A_ADDR_15_), .Y(bus_sync_axi_bus__0reg_data1_63_0__47_));
AND2X2 AND2X2_883 ( .A(RST), .B(A_ADDR_16_), .Y(bus_sync_axi_bus__0reg_data1_63_0__48_));
AND2X2 AND2X2_884 ( .A(RST), .B(A_ADDR_17_), .Y(bus_sync_axi_bus__0reg_data1_63_0__49_));
AND2X2 AND2X2_885 ( .A(RST), .B(A_ADDR_18_), .Y(bus_sync_axi_bus__0reg_data1_63_0__50_));
AND2X2 AND2X2_886 ( .A(RST), .B(A_ADDR_19_), .Y(bus_sync_axi_bus__0reg_data1_63_0__51_));
AND2X2 AND2X2_887 ( .A(RST), .B(A_ADDR_20_), .Y(bus_sync_axi_bus__0reg_data1_63_0__52_));
AND2X2 AND2X2_888 ( .A(RST), .B(A_ADDR_21_), .Y(bus_sync_axi_bus__0reg_data1_63_0__53_));
AND2X2 AND2X2_889 ( .A(RST), .B(A_ADDR_22_), .Y(bus_sync_axi_bus__0reg_data1_63_0__54_));
AND2X2 AND2X2_89 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_9_), .Y(_abc_4268_new_n774_));
AND2X2 AND2X2_890 ( .A(RST), .B(A_ADDR_23_), .Y(bus_sync_axi_bus__0reg_data1_63_0__55_));
AND2X2 AND2X2_891 ( .A(RST), .B(A_ADDR_24_), .Y(bus_sync_axi_bus__0reg_data1_63_0__56_));
AND2X2 AND2X2_892 ( .A(RST), .B(A_ADDR_25_), .Y(bus_sync_axi_bus__0reg_data1_63_0__57_));
AND2X2 AND2X2_893 ( .A(RST), .B(A_ADDR_26_), .Y(bus_sync_axi_bus__0reg_data1_63_0__58_));
AND2X2 AND2X2_894 ( .A(RST), .B(A_ADDR_27_), .Y(bus_sync_axi_bus__0reg_data1_63_0__59_));
AND2X2 AND2X2_895 ( .A(RST), .B(A_ADDR_28_), .Y(bus_sync_axi_bus__0reg_data1_63_0__60_));
AND2X2 AND2X2_896 ( .A(RST), .B(A_ADDR_29_), .Y(bus_sync_axi_bus__0reg_data1_63_0__61_));
AND2X2 AND2X2_897 ( .A(RST), .B(A_ADDR_30_), .Y(bus_sync_axi_bus__0reg_data1_63_0__62_));
AND2X2 AND2X2_898 ( .A(RST), .B(A_ADDR_31_), .Y(bus_sync_axi_bus__0reg_data1_63_0__63_));
AND2X2 AND2X2_899 ( .A(RST), .B(SCLK), .Y(bus_sync_axi_bus__0ECLK1_0_0_));
AND2X2 AND2X2_9 ( .A(_abc_4268_new_n573_), .B(RST), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_1_));
AND2X2 AND2X2_90 ( .A(_abc_4268_new_n775_), .B(RST), .Y(_abc_4268_new_n776_));
AND2X2 AND2X2_900 ( .A(RST), .B(bus_sync_axi_bus_ECLK1), .Y(bus_sync_axi_bus__0EECLK1_0_0_));
AND2X2 AND2X2_901 ( .A(RST), .B(bus_sync_rdata_data_in_0_), .Y(bus_sync_rdata__0reg_data1_31_0__0_));
AND2X2 AND2X2_902 ( .A(RST), .B(bus_sync_rdata_data_in_1_), .Y(bus_sync_rdata__0reg_data1_31_0__1_));
AND2X2 AND2X2_903 ( .A(RST), .B(bus_sync_rdata_data_in_2_), .Y(bus_sync_rdata__0reg_data1_31_0__2_));
AND2X2 AND2X2_904 ( .A(RST), .B(bus_sync_rdata_data_in_3_), .Y(bus_sync_rdata__0reg_data1_31_0__3_));
AND2X2 AND2X2_905 ( .A(RST), .B(bus_sync_rdata_data_in_4_), .Y(bus_sync_rdata__0reg_data1_31_0__4_));
AND2X2 AND2X2_906 ( .A(RST), .B(bus_sync_rdata_data_in_5_), .Y(bus_sync_rdata__0reg_data1_31_0__5_));
AND2X2 AND2X2_907 ( .A(RST), .B(bus_sync_rdata_data_in_6_), .Y(bus_sync_rdata__0reg_data1_31_0__6_));
AND2X2 AND2X2_908 ( .A(RST), .B(bus_sync_rdata_data_in_7_), .Y(bus_sync_rdata__0reg_data1_31_0__7_));
AND2X2 AND2X2_909 ( .A(RST), .B(bus_sync_rdata_data_in_8_), .Y(bus_sync_rdata__0reg_data1_31_0__8_));
AND2X2 AND2X2_91 ( .A(_abc_4268_new_n773_), .B(_abc_4268_new_n776_), .Y(_0bus_cap_31_0__9_));
AND2X2 AND2X2_910 ( .A(RST), .B(bus_sync_rdata_data_in_9_), .Y(bus_sync_rdata__0reg_data1_31_0__9_));
AND2X2 AND2X2_911 ( .A(RST), .B(bus_sync_rdata_data_in_10_), .Y(bus_sync_rdata__0reg_data1_31_0__10_));
AND2X2 AND2X2_912 ( .A(RST), .B(bus_sync_rdata_data_in_11_), .Y(bus_sync_rdata__0reg_data1_31_0__11_));
AND2X2 AND2X2_913 ( .A(RST), .B(bus_sync_rdata_data_in_12_), .Y(bus_sync_rdata__0reg_data1_31_0__12_));
AND2X2 AND2X2_914 ( .A(RST), .B(bus_sync_rdata_data_in_13_), .Y(bus_sync_rdata__0reg_data1_31_0__13_));
AND2X2 AND2X2_915 ( .A(RST), .B(bus_sync_rdata_data_in_14_), .Y(bus_sync_rdata__0reg_data1_31_0__14_));
AND2X2 AND2X2_916 ( .A(RST), .B(bus_sync_rdata_data_in_15_), .Y(bus_sync_rdata__0reg_data1_31_0__15_));
AND2X2 AND2X2_917 ( .A(RST), .B(bus_sync_rdata_data_in_16_), .Y(bus_sync_rdata__0reg_data1_31_0__16_));
AND2X2 AND2X2_918 ( .A(RST), .B(bus_sync_rdata_data_in_17_), .Y(bus_sync_rdata__0reg_data1_31_0__17_));
AND2X2 AND2X2_919 ( .A(RST), .B(bus_sync_rdata_data_in_18_), .Y(bus_sync_rdata__0reg_data1_31_0__18_));
AND2X2 AND2X2_92 ( .A(_abc_4268_new_n778_), .B(_abc_4268_new_n779_), .Y(_abc_4268_new_n780_));
AND2X2 AND2X2_920 ( .A(RST), .B(bus_sync_rdata_data_in_19_), .Y(bus_sync_rdata__0reg_data1_31_0__19_));
AND2X2 AND2X2_921 ( .A(RST), .B(bus_sync_rdata_data_in_20_), .Y(bus_sync_rdata__0reg_data1_31_0__20_));
AND2X2 AND2X2_922 ( .A(RST), .B(bus_sync_rdata_data_in_21_), .Y(bus_sync_rdata__0reg_data1_31_0__21_));
AND2X2 AND2X2_923 ( .A(RST), .B(bus_sync_rdata_data_in_22_), .Y(bus_sync_rdata__0reg_data1_31_0__22_));
AND2X2 AND2X2_924 ( .A(RST), .B(bus_sync_rdata_data_in_23_), .Y(bus_sync_rdata__0reg_data1_31_0__23_));
AND2X2 AND2X2_925 ( .A(RST), .B(bus_sync_rdata_data_in_24_), .Y(bus_sync_rdata__0reg_data1_31_0__24_));
AND2X2 AND2X2_926 ( .A(RST), .B(bus_sync_rdata_data_in_25_), .Y(bus_sync_rdata__0reg_data1_31_0__25_));
AND2X2 AND2X2_927 ( .A(RST), .B(bus_sync_rdata_data_in_26_), .Y(bus_sync_rdata__0reg_data1_31_0__26_));
AND2X2 AND2X2_928 ( .A(RST), .B(bus_sync_rdata_data_in_27_), .Y(bus_sync_rdata__0reg_data1_31_0__27_));
AND2X2 AND2X2_929 ( .A(RST), .B(bus_sync_rdata_data_in_28_), .Y(bus_sync_rdata__0reg_data1_31_0__28_));
AND2X2 AND2X2_93 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_10_), .Y(_abc_4268_new_n782_));
AND2X2 AND2X2_930 ( .A(RST), .B(bus_sync_rdata_data_in_29_), .Y(bus_sync_rdata__0reg_data1_31_0__29_));
AND2X2 AND2X2_931 ( .A(RST), .B(bus_sync_rdata_data_in_30_), .Y(bus_sync_rdata__0reg_data1_31_0__30_));
AND2X2 AND2X2_932 ( .A(RST), .B(bus_sync_rdata_data_in_31_), .Y(bus_sync_rdata__0reg_data1_31_0__31_));
AND2X2 AND2X2_933 ( .A(RST), .B(bus_sync_rdata_reg_data2_0_), .Y(bus_sync_rdata__0reg_data3_31_0__0_));
AND2X2 AND2X2_934 ( .A(RST), .B(bus_sync_rdata_reg_data2_1_), .Y(bus_sync_rdata__0reg_data3_31_0__1_));
AND2X2 AND2X2_935 ( .A(RST), .B(bus_sync_rdata_reg_data2_2_), .Y(bus_sync_rdata__0reg_data3_31_0__2_));
AND2X2 AND2X2_936 ( .A(RST), .B(bus_sync_rdata_reg_data2_3_), .Y(bus_sync_rdata__0reg_data3_31_0__3_));
AND2X2 AND2X2_937 ( .A(RST), .B(bus_sync_rdata_reg_data2_4_), .Y(bus_sync_rdata__0reg_data3_31_0__4_));
AND2X2 AND2X2_938 ( .A(RST), .B(bus_sync_rdata_reg_data2_5_), .Y(bus_sync_rdata__0reg_data3_31_0__5_));
AND2X2 AND2X2_939 ( .A(RST), .B(bus_sync_rdata_reg_data2_6_), .Y(bus_sync_rdata__0reg_data3_31_0__6_));
AND2X2 AND2X2_94 ( .A(_abc_4268_new_n783_), .B(RST), .Y(_abc_4268_new_n784_));
AND2X2 AND2X2_940 ( .A(RST), .B(bus_sync_rdata_reg_data2_7_), .Y(bus_sync_rdata__0reg_data3_31_0__7_));
AND2X2 AND2X2_941 ( .A(RST), .B(bus_sync_rdata_reg_data2_8_), .Y(bus_sync_rdata__0reg_data3_31_0__8_));
AND2X2 AND2X2_942 ( .A(RST), .B(bus_sync_rdata_reg_data2_9_), .Y(bus_sync_rdata__0reg_data3_31_0__9_));
AND2X2 AND2X2_943 ( .A(RST), .B(bus_sync_rdata_reg_data2_10_), .Y(bus_sync_rdata__0reg_data3_31_0__10_));
AND2X2 AND2X2_944 ( .A(RST), .B(bus_sync_rdata_reg_data2_11_), .Y(bus_sync_rdata__0reg_data3_31_0__11_));
AND2X2 AND2X2_945 ( .A(RST), .B(bus_sync_rdata_reg_data2_12_), .Y(bus_sync_rdata__0reg_data3_31_0__12_));
AND2X2 AND2X2_946 ( .A(RST), .B(bus_sync_rdata_reg_data2_13_), .Y(bus_sync_rdata__0reg_data3_31_0__13_));
AND2X2 AND2X2_947 ( .A(RST), .B(bus_sync_rdata_reg_data2_14_), .Y(bus_sync_rdata__0reg_data3_31_0__14_));
AND2X2 AND2X2_948 ( .A(RST), .B(bus_sync_rdata_reg_data2_15_), .Y(bus_sync_rdata__0reg_data3_31_0__15_));
AND2X2 AND2X2_949 ( .A(RST), .B(bus_sync_rdata_reg_data2_16_), .Y(bus_sync_rdata__0reg_data3_31_0__16_));
AND2X2 AND2X2_95 ( .A(_abc_4268_new_n781_), .B(_abc_4268_new_n784_), .Y(_0bus_cap_31_0__10_));
AND2X2 AND2X2_950 ( .A(RST), .B(bus_sync_rdata_reg_data2_17_), .Y(bus_sync_rdata__0reg_data3_31_0__17_));
AND2X2 AND2X2_951 ( .A(RST), .B(bus_sync_rdata_reg_data2_18_), .Y(bus_sync_rdata__0reg_data3_31_0__18_));
AND2X2 AND2X2_952 ( .A(RST), .B(bus_sync_rdata_reg_data2_19_), .Y(bus_sync_rdata__0reg_data3_31_0__19_));
AND2X2 AND2X2_953 ( .A(RST), .B(bus_sync_rdata_reg_data2_20_), .Y(bus_sync_rdata__0reg_data3_31_0__20_));
AND2X2 AND2X2_954 ( .A(RST), .B(bus_sync_rdata_reg_data2_21_), .Y(bus_sync_rdata__0reg_data3_31_0__21_));
AND2X2 AND2X2_955 ( .A(RST), .B(bus_sync_rdata_reg_data2_22_), .Y(bus_sync_rdata__0reg_data3_31_0__22_));
AND2X2 AND2X2_956 ( .A(RST), .B(bus_sync_rdata_reg_data2_23_), .Y(bus_sync_rdata__0reg_data3_31_0__23_));
AND2X2 AND2X2_957 ( .A(RST), .B(bus_sync_rdata_reg_data2_24_), .Y(bus_sync_rdata__0reg_data3_31_0__24_));
AND2X2 AND2X2_958 ( .A(RST), .B(bus_sync_rdata_reg_data2_25_), .Y(bus_sync_rdata__0reg_data3_31_0__25_));
AND2X2 AND2X2_959 ( .A(RST), .B(bus_sync_rdata_reg_data2_26_), .Y(bus_sync_rdata__0reg_data3_31_0__26_));
AND2X2 AND2X2_96 ( .A(_abc_4268_new_n786_), .B(_abc_4268_new_n787_), .Y(_abc_4268_new_n788_));
AND2X2 AND2X2_960 ( .A(RST), .B(bus_sync_rdata_reg_data2_27_), .Y(bus_sync_rdata__0reg_data3_31_0__27_));
AND2X2 AND2X2_961 ( .A(RST), .B(bus_sync_rdata_reg_data2_28_), .Y(bus_sync_rdata__0reg_data3_31_0__28_));
AND2X2 AND2X2_962 ( .A(RST), .B(bus_sync_rdata_reg_data2_29_), .Y(bus_sync_rdata__0reg_data3_31_0__29_));
AND2X2 AND2X2_963 ( .A(RST), .B(bus_sync_rdata_reg_data2_30_), .Y(bus_sync_rdata__0reg_data3_31_0__30_));
AND2X2 AND2X2_964 ( .A(RST), .B(bus_sync_rdata_reg_data2_31_), .Y(bus_sync_rdata__0reg_data3_31_0__31_));
AND2X2 AND2X2_965 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_0_), .Y(bus_sync_rdata__abc_3653_new_n266_));
AND2X2 AND2X2_966 ( .A(bus_sync_rdata_reg_data1_0_), .B(bus_sync_rdata_EECLK2), .Y(bus_sync_rdata__abc_3653_new_n267_));
AND2X2 AND2X2_967 ( .A(bus_sync_rdata__abc_3653_new_n268_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__0_));
AND2X2 AND2X2_968 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_1_), .Y(bus_sync_rdata__abc_3653_new_n270_));
AND2X2 AND2X2_969 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_1_), .Y(bus_sync_rdata__abc_3653_new_n271_));
AND2X2 AND2X2_97 ( .A(_abc_4268_new_n616_), .B(bus_sync_rdata_data_out_11_), .Y(_abc_4268_new_n790_));
AND2X2 AND2X2_970 ( .A(bus_sync_rdata__abc_3653_new_n272_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__1_));
AND2X2 AND2X2_971 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_2_), .Y(bus_sync_rdata__abc_3653_new_n274_));
AND2X2 AND2X2_972 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_2_), .Y(bus_sync_rdata__abc_3653_new_n275_));
AND2X2 AND2X2_973 ( .A(bus_sync_rdata__abc_3653_new_n276_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__2_));
AND2X2 AND2X2_974 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_3_), .Y(bus_sync_rdata__abc_3653_new_n278_));
AND2X2 AND2X2_975 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_3_), .Y(bus_sync_rdata__abc_3653_new_n279_));
AND2X2 AND2X2_976 ( .A(bus_sync_rdata__abc_3653_new_n280_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__3_));
AND2X2 AND2X2_977 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_4_), .Y(bus_sync_rdata__abc_3653_new_n282_));
AND2X2 AND2X2_978 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_4_), .Y(bus_sync_rdata__abc_3653_new_n283_));
AND2X2 AND2X2_979 ( .A(bus_sync_rdata__abc_3653_new_n284_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__4_));
AND2X2 AND2X2_98 ( .A(_abc_4268_new_n791_), .B(RST), .Y(_abc_4268_new_n792_));
AND2X2 AND2X2_980 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_5_), .Y(bus_sync_rdata__abc_3653_new_n286_));
AND2X2 AND2X2_981 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_5_), .Y(bus_sync_rdata__abc_3653_new_n287_));
AND2X2 AND2X2_982 ( .A(bus_sync_rdata__abc_3653_new_n288_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__5_));
AND2X2 AND2X2_983 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_6_), .Y(bus_sync_rdata__abc_3653_new_n290_));
AND2X2 AND2X2_984 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_6_), .Y(bus_sync_rdata__abc_3653_new_n291_));
AND2X2 AND2X2_985 ( .A(bus_sync_rdata__abc_3653_new_n292_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__6_));
AND2X2 AND2X2_986 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_7_), .Y(bus_sync_rdata__abc_3653_new_n294_));
AND2X2 AND2X2_987 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_7_), .Y(bus_sync_rdata__abc_3653_new_n295_));
AND2X2 AND2X2_988 ( .A(bus_sync_rdata__abc_3653_new_n296_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__7_));
AND2X2 AND2X2_989 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_8_), .Y(bus_sync_rdata__abc_3653_new_n298_));
AND2X2 AND2X2_99 ( .A(_abc_4268_new_n789_), .B(_abc_4268_new_n792_), .Y(_0bus_cap_31_0__11_));
AND2X2 AND2X2_990 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_8_), .Y(bus_sync_rdata__abc_3653_new_n299_));
AND2X2 AND2X2_991 ( .A(bus_sync_rdata__abc_3653_new_n300_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__8_));
AND2X2 AND2X2_992 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_9_), .Y(bus_sync_rdata__abc_3653_new_n302_));
AND2X2 AND2X2_993 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_9_), .Y(bus_sync_rdata__abc_3653_new_n303_));
AND2X2 AND2X2_994 ( .A(bus_sync_rdata__abc_3653_new_n304_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__9_));
AND2X2 AND2X2_995 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_10_), .Y(bus_sync_rdata__abc_3653_new_n306_));
AND2X2 AND2X2_996 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_10_), .Y(bus_sync_rdata__abc_3653_new_n307_));
AND2X2 AND2X2_997 ( .A(bus_sync_rdata__abc_3653_new_n308_), .B(RST), .Y(bus_sync_rdata__0reg_data2_31_0__10_));
AND2X2 AND2X2_998 ( .A(bus_sync_rdata__abc_3653_new_n265_), .B(bus_sync_rdata_reg_data2_11_), .Y(bus_sync_rdata__abc_3653_new_n310_));
AND2X2 AND2X2_999 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_11_), .Y(bus_sync_rdata__abc_3653_new_n311_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(SCLK), .D(_0counter_65_0__0_), .Q(counter_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(SCLK), .D(_0counter_65_0__9_), .Q(counter_9_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(CLK), .D(_0rdata_31_0__0_), .Q(bus_sync_rdata_data_in_0_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(CLK), .D(_0rdata_31_0__1_), .Q(bus_sync_rdata_data_in_1_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(CLK), .D(_0rdata_31_0__2_), .Q(bus_sync_rdata_data_in_2_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(CLK), .D(_0rdata_31_0__3_), .Q(bus_sync_rdata_data_in_3_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(CLK), .D(_0rdata_31_0__4_), .Q(bus_sync_rdata_data_in_4_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(CLK), .D(_0rdata_31_0__5_), .Q(bus_sync_rdata_data_in_5_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(CLK), .D(_0rdata_31_0__6_), .Q(bus_sync_rdata_data_in_6_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(CLK), .D(_0rdata_31_0__7_), .Q(bus_sync_rdata_data_in_7_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(CLK), .D(_0rdata_31_0__8_), .Q(bus_sync_rdata_data_in_8_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(CLK), .D(_0rdata_31_0__9_), .Q(bus_sync_rdata_data_in_9_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(SCLK), .D(_0counter_65_0__10_), .Q(counter_10_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(CLK), .D(_0rdata_31_0__10_), .Q(bus_sync_rdata_data_in_10_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(CLK), .D(_0rdata_31_0__11_), .Q(bus_sync_rdata_data_in_11_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(CLK), .D(_0rdata_31_0__12_), .Q(bus_sync_rdata_data_in_12_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(CLK), .D(_0rdata_31_0__13_), .Q(bus_sync_rdata_data_in_13_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(CLK), .D(_0rdata_31_0__14_), .Q(bus_sync_rdata_data_in_14_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(CLK), .D(_0rdata_31_0__15_), .Q(bus_sync_rdata_data_in_15_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(CLK), .D(_0rdata_31_0__16_), .Q(bus_sync_rdata_data_in_16_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(CLK), .D(_0rdata_31_0__17_), .Q(bus_sync_rdata_data_in_17_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(CLK), .D(_0rdata_31_0__18_), .Q(bus_sync_rdata_data_in_18_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(CLK), .D(_0rdata_31_0__19_), .Q(bus_sync_rdata_data_in_19_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(SCLK), .D(_0counter_65_0__11_), .Q(counter_11_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(CLK), .D(_0rdata_31_0__20_), .Q(bus_sync_rdata_data_in_20_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(CLK), .D(_0rdata_31_0__21_), .Q(bus_sync_rdata_data_in_21_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(CLK), .D(_0rdata_31_0__22_), .Q(bus_sync_rdata_data_in_22_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(CLK), .D(_0rdata_31_0__23_), .Q(bus_sync_rdata_data_in_23_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(CLK), .D(_0rdata_31_0__24_), .Q(bus_sync_rdata_data_in_24_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(CLK), .D(_0rdata_31_0__25_), .Q(bus_sync_rdata_data_in_25_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(CLK), .D(_0rdata_31_0__26_), .Q(bus_sync_rdata_data_in_26_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(CLK), .D(_0rdata_31_0__27_), .Q(bus_sync_rdata_data_in_27_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(CLK), .D(_0rdata_31_0__28_), .Q(bus_sync_rdata_data_in_28_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(CLK), .D(_0rdata_31_0__29_), .Q(bus_sync_rdata_data_in_29_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(SCLK), .D(_0counter_65_0__12_), .Q(counter_12_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(CLK), .D(_0rdata_31_0__30_), .Q(bus_sync_rdata_data_in_30_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(CLK), .D(_0rdata_31_0__31_), .Q(bus_sync_rdata_data_in_31_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(SCLK), .D(_0A_ADDR_31_0__0_), .Q(A_ADDR_0_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(SCLK), .D(_0A_ADDR_31_0__1_), .Q(A_ADDR_1_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(SCLK), .D(_0A_ADDR_31_0__2_), .Q(A_ADDR_2_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(SCLK), .D(_0A_ADDR_31_0__3_), .Q(A_ADDR_3_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(SCLK), .D(_0A_ADDR_31_0__4_), .Q(A_ADDR_4_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(SCLK), .D(_0A_ADDR_31_0__5_), .Q(A_ADDR_5_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(SCLK), .D(_0A_ADDR_31_0__6_), .Q(A_ADDR_6_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(SCLK), .D(_0A_ADDR_31_0__7_), .Q(A_ADDR_7_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(SCLK), .D(_0counter_65_0__13_), .Q(counter_13_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(SCLK), .D(_0A_ADDR_31_0__8_), .Q(A_ADDR_8_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(SCLK), .D(_0A_ADDR_31_0__9_), .Q(A_ADDR_9_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(SCLK), .D(_0A_ADDR_31_0__10_), .Q(A_ADDR_10_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(SCLK), .D(_0A_ADDR_31_0__11_), .Q(A_ADDR_11_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(SCLK), .D(_0A_ADDR_31_0__12_), .Q(A_ADDR_12_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(SCLK), .D(_0A_ADDR_31_0__13_), .Q(A_ADDR_13_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(SCLK), .D(_0A_ADDR_31_0__14_), .Q(A_ADDR_14_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(SCLK), .D(_0A_ADDR_31_0__15_), .Q(A_ADDR_15_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(SCLK), .D(_0A_ADDR_31_0__16_), .Q(A_ADDR_16_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(SCLK), .D(_0A_ADDR_31_0__17_), .Q(A_ADDR_17_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(SCLK), .D(_0counter_65_0__14_), .Q(counter_14_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(SCLK), .D(_0A_ADDR_31_0__18_), .Q(A_ADDR_18_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(SCLK), .D(_0A_ADDR_31_0__19_), .Q(A_ADDR_19_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(SCLK), .D(_0A_ADDR_31_0__20_), .Q(A_ADDR_20_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(SCLK), .D(_0A_ADDR_31_0__21_), .Q(A_ADDR_21_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(SCLK), .D(_0A_ADDR_31_0__22_), .Q(A_ADDR_22_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(SCLK), .D(_0A_ADDR_31_0__23_), .Q(A_ADDR_23_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(SCLK), .D(_0A_ADDR_31_0__24_), .Q(A_ADDR_24_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(SCLK), .D(_0A_ADDR_31_0__25_), .Q(A_ADDR_25_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(SCLK), .D(_0A_ADDR_31_0__26_), .Q(A_ADDR_26_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(SCLK), .D(_0A_ADDR_31_0__27_), .Q(A_ADDR_27_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(SCLK), .D(_0counter_65_0__15_), .Q(counter_15_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(SCLK), .D(_0A_ADDR_31_0__28_), .Q(A_ADDR_28_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(SCLK), .D(_0A_ADDR_31_0__29_), .Q(A_ADDR_29_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(SCLK), .D(_0A_ADDR_31_0__30_), .Q(A_ADDR_30_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(SCLK), .D(_0A_ADDR_31_0__31_), .Q(A_ADDR_31_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(SCLK), .D(_0WDATA_31_0__0_), .Q(WDATA_0_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(SCLK), .D(_0WDATA_31_0__1_), .Q(WDATA_1_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(SCLK), .D(_0WDATA_31_0__2_), .Q(WDATA_2_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(SCLK), .D(_0WDATA_31_0__3_), .Q(WDATA_3_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(SCLK), .D(_0WDATA_31_0__4_), .Q(WDATA_4_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(SCLK), .D(_0WDATA_31_0__5_), .Q(WDATA_5_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(SCLK), .D(_0counter_65_0__16_), .Q(counter_16_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(SCLK), .D(_0WDATA_31_0__6_), .Q(WDATA_6_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(SCLK), .D(_0WDATA_31_0__7_), .Q(WDATA_7_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(SCLK), .D(_0WDATA_31_0__8_), .Q(WDATA_8_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(SCLK), .D(_0WDATA_31_0__9_), .Q(WDATA_9_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(SCLK), .D(_0WDATA_31_0__10_), .Q(WDATA_10_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(SCLK), .D(_0WDATA_31_0__11_), .Q(WDATA_11_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(SCLK), .D(_0WDATA_31_0__12_), .Q(WDATA_12_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(SCLK), .D(_0WDATA_31_0__13_), .Q(WDATA_13_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(SCLK), .D(_0WDATA_31_0__14_), .Q(WDATA_14_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(SCLK), .D(_0WDATA_31_0__15_), .Q(WDATA_15_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(SCLK), .D(_0counter_65_0__17_), .Q(counter_17_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(SCLK), .D(_0WDATA_31_0__16_), .Q(WDATA_16_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(SCLK), .D(_0WDATA_31_0__17_), .Q(WDATA_17_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(SCLK), .D(_0WDATA_31_0__18_), .Q(WDATA_18_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(SCLK), .D(_0WDATA_31_0__19_), .Q(WDATA_19_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(SCLK), .D(_0WDATA_31_0__20_), .Q(WDATA_20_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(SCLK), .D(_0WDATA_31_0__21_), .Q(WDATA_21_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(SCLK), .D(_0WDATA_31_0__22_), .Q(WDATA_22_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(SCLK), .D(_0WDATA_31_0__23_), .Q(WDATA_23_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(SCLK), .D(_0WDATA_31_0__24_), .Q(WDATA_24_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(SCLK), .D(_0WDATA_31_0__25_), .Q(WDATA_25_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(SCLK), .D(_0counter_65_0__18_), .Q(counter_18_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(SCLK), .D(_0WDATA_31_0__26_), .Q(WDATA_26_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(SCLK), .D(_0WDATA_31_0__27_), .Q(WDATA_27_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(SCLK), .D(_0WDATA_31_0__28_), .Q(WDATA_28_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(SCLK), .D(_0WDATA_31_0__29_), .Q(WDATA_29_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(SCLK), .D(_0WDATA_31_0__30_), .Q(WDATA_30_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(SCLK), .D(_0WDATA_31_0__31_), .Q(WDATA_31_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(SCLK), .D(_0PICORV_RST_SPI_0_0_), .Q(PICORV_RST_SPI));
DFFPOSX1 DFFPOSX1_197 ( .CLK(SCLK), .D(_0we_0_0_), .Q(we));
DFFPOSX1 DFFPOSX1_198 ( .CLK(SCLK), .D(_0re_0_0_), .Q(re));
DFFPOSX1 DFFPOSX1_199 ( .CLK(SCLK), .D(_0sft_reg_65_0__0_), .Q(sft_reg_0_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(SCLK), .D(_0counter_65_0__1_), .Q(counter_1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(SCLK), .D(_0counter_65_0__19_), .Q(counter_19_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(SCLK), .D(_0sft_reg_65_0__1_), .Q(sft_reg_1_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(SCLK), .D(_0sft_reg_65_0__2_), .Q(sft_reg_2_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(SCLK), .D(_0sft_reg_65_0__3_), .Q(sft_reg_3_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(SCLK), .D(_0sft_reg_65_0__4_), .Q(sft_reg_4_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(SCLK), .D(_0sft_reg_65_0__5_), .Q(sft_reg_5_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(SCLK), .D(_0sft_reg_65_0__6_), .Q(sft_reg_6_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(SCLK), .D(_0sft_reg_65_0__7_), .Q(sft_reg_7_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(SCLK), .D(_0sft_reg_65_0__8_), .Q(sft_reg_8_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(SCLK), .D(_0sft_reg_65_0__9_), .Q(sft_reg_9_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(SCLK), .D(_0sft_reg_65_0__10_), .Q(sft_reg_10_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(SCLK), .D(_0counter_65_0__20_), .Q(counter_20_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(SCLK), .D(_0sft_reg_65_0__11_), .Q(sft_reg_11_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(SCLK), .D(_0sft_reg_65_0__12_), .Q(sft_reg_12_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(SCLK), .D(_0sft_reg_65_0__13_), .Q(sft_reg_13_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(SCLK), .D(_0sft_reg_65_0__14_), .Q(sft_reg_14_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(SCLK), .D(_0sft_reg_65_0__15_), .Q(sft_reg_15_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(SCLK), .D(_0sft_reg_65_0__16_), .Q(sft_reg_16_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(SCLK), .D(_0sft_reg_65_0__17_), .Q(sft_reg_17_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(SCLK), .D(_0sft_reg_65_0__18_), .Q(sft_reg_18_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(SCLK), .D(_0sft_reg_65_0__19_), .Q(sft_reg_19_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(SCLK), .D(_0sft_reg_65_0__20_), .Q(sft_reg_20_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(SCLK), .D(_0counter_65_0__21_), .Q(counter_21_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(SCLK), .D(_0sft_reg_65_0__21_), .Q(sft_reg_21_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(SCLK), .D(_0sft_reg_65_0__22_), .Q(sft_reg_22_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(SCLK), .D(_0sft_reg_65_0__23_), .Q(sft_reg_23_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(SCLK), .D(_0sft_reg_65_0__24_), .Q(sft_reg_24_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(SCLK), .D(_0sft_reg_65_0__25_), .Q(sft_reg_25_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(SCLK), .D(_0sft_reg_65_0__26_), .Q(sft_reg_26_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(SCLK), .D(_0sft_reg_65_0__27_), .Q(sft_reg_27_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(SCLK), .D(_0sft_reg_65_0__28_), .Q(sft_reg_28_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(SCLK), .D(_0sft_reg_65_0__29_), .Q(sft_reg_29_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(SCLK), .D(_0sft_reg_65_0__30_), .Q(sft_reg_30_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(SCLK), .D(_0counter_65_0__22_), .Q(counter_22_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_0_), .Q(state_0_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_1_), .Q(state_1_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_430), .Q(axi_bready));
DFFPOSX1 DFFPOSX1_233 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_3_), .Q(state_3_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_4_), .Q(state_4_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_5_), .Q(state_5_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_6_), .Q(state_6_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_7_), .Q(state_7_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(CLK), .D(_abc_2903_auto_fsm_map_cc_118_implement_pattern_cache_479), .Q(axi_rready));
DFFPOSX1 DFFPOSX1_239 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__0_), .Q(bus_sync_axi_bus_reg_data2_0_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(SCLK), .D(_0counter_65_0__23_), .Q(counter_23_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__1_), .Q(bus_sync_axi_bus_reg_data2_1_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__2_), .Q(bus_sync_axi_bus_reg_data2_2_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__3_), .Q(bus_sync_axi_bus_reg_data2_3_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__4_), .Q(bus_sync_axi_bus_reg_data2_4_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__5_), .Q(bus_sync_axi_bus_reg_data2_5_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__6_), .Q(bus_sync_axi_bus_reg_data2_6_));
DFFPOSX1 DFFPOSX1_246 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__7_), .Q(bus_sync_axi_bus_reg_data2_7_));
DFFPOSX1 DFFPOSX1_247 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__8_), .Q(bus_sync_axi_bus_reg_data2_8_));
DFFPOSX1 DFFPOSX1_248 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__9_), .Q(bus_sync_axi_bus_reg_data2_9_));
DFFPOSX1 DFFPOSX1_249 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__10_), .Q(bus_sync_axi_bus_reg_data2_10_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(SCLK), .D(_0counter_65_0__24_), .Q(counter_24_));
DFFPOSX1 DFFPOSX1_250 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__11_), .Q(bus_sync_axi_bus_reg_data2_11_));
DFFPOSX1 DFFPOSX1_251 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__12_), .Q(bus_sync_axi_bus_reg_data2_12_));
DFFPOSX1 DFFPOSX1_252 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__13_), .Q(bus_sync_axi_bus_reg_data2_13_));
DFFPOSX1 DFFPOSX1_253 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__14_), .Q(bus_sync_axi_bus_reg_data2_14_));
DFFPOSX1 DFFPOSX1_254 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__15_), .Q(bus_sync_axi_bus_reg_data2_15_));
DFFPOSX1 DFFPOSX1_255 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__16_), .Q(bus_sync_axi_bus_reg_data2_16_));
DFFPOSX1 DFFPOSX1_256 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__17_), .Q(bus_sync_axi_bus_reg_data2_17_));
DFFPOSX1 DFFPOSX1_257 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__18_), .Q(bus_sync_axi_bus_reg_data2_18_));
DFFPOSX1 DFFPOSX1_258 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__19_), .Q(bus_sync_axi_bus_reg_data2_19_));
DFFPOSX1 DFFPOSX1_259 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__20_), .Q(bus_sync_axi_bus_reg_data2_20_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(SCLK), .D(_0counter_65_0__25_), .Q(counter_25_));
DFFPOSX1 DFFPOSX1_260 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__21_), .Q(bus_sync_axi_bus_reg_data2_21_));
DFFPOSX1 DFFPOSX1_261 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__22_), .Q(bus_sync_axi_bus_reg_data2_22_));
DFFPOSX1 DFFPOSX1_262 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__23_), .Q(bus_sync_axi_bus_reg_data2_23_));
DFFPOSX1 DFFPOSX1_263 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__24_), .Q(bus_sync_axi_bus_reg_data2_24_));
DFFPOSX1 DFFPOSX1_264 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__25_), .Q(bus_sync_axi_bus_reg_data2_25_));
DFFPOSX1 DFFPOSX1_265 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__26_), .Q(bus_sync_axi_bus_reg_data2_26_));
DFFPOSX1 DFFPOSX1_266 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__27_), .Q(bus_sync_axi_bus_reg_data2_27_));
DFFPOSX1 DFFPOSX1_267 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__28_), .Q(bus_sync_axi_bus_reg_data2_28_));
DFFPOSX1 DFFPOSX1_268 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__29_), .Q(bus_sync_axi_bus_reg_data2_29_));
DFFPOSX1 DFFPOSX1_269 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__30_), .Q(bus_sync_axi_bus_reg_data2_30_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(SCLK), .D(_0counter_65_0__26_), .Q(counter_26_));
DFFPOSX1 DFFPOSX1_270 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__31_), .Q(bus_sync_axi_bus_reg_data2_31_));
DFFPOSX1 DFFPOSX1_271 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__32_), .Q(bus_sync_axi_bus_reg_data2_32_));
DFFPOSX1 DFFPOSX1_272 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__33_), .Q(bus_sync_axi_bus_reg_data2_33_));
DFFPOSX1 DFFPOSX1_273 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__34_), .Q(bus_sync_axi_bus_reg_data2_34_));
DFFPOSX1 DFFPOSX1_274 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__35_), .Q(bus_sync_axi_bus_reg_data2_35_));
DFFPOSX1 DFFPOSX1_275 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__36_), .Q(bus_sync_axi_bus_reg_data2_36_));
DFFPOSX1 DFFPOSX1_276 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__37_), .Q(bus_sync_axi_bus_reg_data2_37_));
DFFPOSX1 DFFPOSX1_277 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__38_), .Q(bus_sync_axi_bus_reg_data2_38_));
DFFPOSX1 DFFPOSX1_278 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__39_), .Q(bus_sync_axi_bus_reg_data2_39_));
DFFPOSX1 DFFPOSX1_279 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__40_), .Q(bus_sync_axi_bus_reg_data2_40_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(SCLK), .D(_0counter_65_0__27_), .Q(counter_27_));
DFFPOSX1 DFFPOSX1_280 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__41_), .Q(bus_sync_axi_bus_reg_data2_41_));
DFFPOSX1 DFFPOSX1_281 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__42_), .Q(bus_sync_axi_bus_reg_data2_42_));
DFFPOSX1 DFFPOSX1_282 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__43_), .Q(bus_sync_axi_bus_reg_data2_43_));
DFFPOSX1 DFFPOSX1_283 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__44_), .Q(bus_sync_axi_bus_reg_data2_44_));
DFFPOSX1 DFFPOSX1_284 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__45_), .Q(bus_sync_axi_bus_reg_data2_45_));
DFFPOSX1 DFFPOSX1_285 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__46_), .Q(bus_sync_axi_bus_reg_data2_46_));
DFFPOSX1 DFFPOSX1_286 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__47_), .Q(bus_sync_axi_bus_reg_data2_47_));
DFFPOSX1 DFFPOSX1_287 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__48_), .Q(bus_sync_axi_bus_reg_data2_48_));
DFFPOSX1 DFFPOSX1_288 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__49_), .Q(bus_sync_axi_bus_reg_data2_49_));
DFFPOSX1 DFFPOSX1_289 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__50_), .Q(bus_sync_axi_bus_reg_data2_50_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(SCLK), .D(_0counter_65_0__28_), .Q(counter_28_));
DFFPOSX1 DFFPOSX1_290 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__51_), .Q(bus_sync_axi_bus_reg_data2_51_));
DFFPOSX1 DFFPOSX1_291 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__52_), .Q(bus_sync_axi_bus_reg_data2_52_));
DFFPOSX1 DFFPOSX1_292 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__53_), .Q(bus_sync_axi_bus_reg_data2_53_));
DFFPOSX1 DFFPOSX1_293 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__54_), .Q(bus_sync_axi_bus_reg_data2_54_));
DFFPOSX1 DFFPOSX1_294 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__55_), .Q(bus_sync_axi_bus_reg_data2_55_));
DFFPOSX1 DFFPOSX1_295 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__56_), .Q(bus_sync_axi_bus_reg_data2_56_));
DFFPOSX1 DFFPOSX1_296 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__57_), .Q(bus_sync_axi_bus_reg_data2_57_));
DFFPOSX1 DFFPOSX1_297 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__58_), .Q(bus_sync_axi_bus_reg_data2_58_));
DFFPOSX1 DFFPOSX1_298 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__59_), .Q(bus_sync_axi_bus_reg_data2_59_));
DFFPOSX1 DFFPOSX1_299 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__60_), .Q(bus_sync_axi_bus_reg_data2_60_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(SCLK), .D(_0counter_65_0__2_), .Q(counter_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(SCLK), .D(_0counter_65_0__29_), .Q(counter_29_));
DFFPOSX1 DFFPOSX1_300 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__61_), .Q(bus_sync_axi_bus_reg_data2_61_));
DFFPOSX1 DFFPOSX1_301 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__62_), .Q(bus_sync_axi_bus_reg_data2_62_));
DFFPOSX1 DFFPOSX1_302 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data2_63_0__63_), .Q(bus_sync_axi_bus_reg_data2_63_));
DFFPOSX1 DFFPOSX1_303 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__0_), .Q(\axi_wdata[0] ));
DFFPOSX1 DFFPOSX1_304 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__1_), .Q(\axi_wdata[1] ));
DFFPOSX1 DFFPOSX1_305 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__2_), .Q(\axi_wdata[2] ));
DFFPOSX1 DFFPOSX1_306 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__3_), .Q(\axi_wdata[3] ));
DFFPOSX1 DFFPOSX1_307 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__4_), .Q(\axi_wdata[4] ));
DFFPOSX1 DFFPOSX1_308 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__5_), .Q(\axi_wdata[5] ));
DFFPOSX1 DFFPOSX1_309 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__6_), .Q(\axi_wdata[6] ));
DFFPOSX1 DFFPOSX1_31 ( .CLK(SCLK), .D(_0counter_65_0__30_), .Q(counter_30_));
DFFPOSX1 DFFPOSX1_310 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__7_), .Q(\axi_wdata[7] ));
DFFPOSX1 DFFPOSX1_311 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__8_), .Q(\axi_wdata[8] ));
DFFPOSX1 DFFPOSX1_312 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__9_), .Q(\axi_wdata[9] ));
DFFPOSX1 DFFPOSX1_313 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__10_), .Q(\axi_wdata[10] ));
DFFPOSX1 DFFPOSX1_314 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__11_), .Q(\axi_wdata[11] ));
DFFPOSX1 DFFPOSX1_315 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__12_), .Q(\axi_wdata[12] ));
DFFPOSX1 DFFPOSX1_316 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__13_), .Q(\axi_wdata[13] ));
DFFPOSX1 DFFPOSX1_317 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__14_), .Q(\axi_wdata[14] ));
DFFPOSX1 DFFPOSX1_318 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__15_), .Q(\axi_wdata[15] ));
DFFPOSX1 DFFPOSX1_319 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__16_), .Q(\axi_wdata[16] ));
DFFPOSX1 DFFPOSX1_32 ( .CLK(SCLK), .D(_0counter_65_0__31_), .Q(counter_31_));
DFFPOSX1 DFFPOSX1_320 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__17_), .Q(\axi_wdata[17] ));
DFFPOSX1 DFFPOSX1_321 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__18_), .Q(\axi_wdata[18] ));
DFFPOSX1 DFFPOSX1_322 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__19_), .Q(\axi_wdata[19] ));
DFFPOSX1 DFFPOSX1_323 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__20_), .Q(\axi_wdata[20] ));
DFFPOSX1 DFFPOSX1_324 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__21_), .Q(\axi_wdata[21] ));
DFFPOSX1 DFFPOSX1_325 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__22_), .Q(\axi_wdata[22] ));
DFFPOSX1 DFFPOSX1_326 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__23_), .Q(\axi_wdata[23] ));
DFFPOSX1 DFFPOSX1_327 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__24_), .Q(\axi_wdata[24] ));
DFFPOSX1 DFFPOSX1_328 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__25_), .Q(\axi_wdata[25] ));
DFFPOSX1 DFFPOSX1_329 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__26_), .Q(\axi_wdata[26] ));
DFFPOSX1 DFFPOSX1_33 ( .CLK(SCLK), .D(_0counter_65_0__32_), .Q(counter_32_));
DFFPOSX1 DFFPOSX1_330 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__27_), .Q(\axi_wdata[27] ));
DFFPOSX1 DFFPOSX1_331 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__28_), .Q(\axi_wdata[28] ));
DFFPOSX1 DFFPOSX1_332 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__29_), .Q(\axi_wdata[29] ));
DFFPOSX1 DFFPOSX1_333 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__30_), .Q(\axi_wdata[30] ));
DFFPOSX1 DFFPOSX1_334 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__31_), .Q(\axi_wdata[31] ));
DFFPOSX1 DFFPOSX1_335 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__32_), .Q(\axi_araddr[0] ));
DFFPOSX1 DFFPOSX1_336 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__33_), .Q(\axi_araddr[1] ));
DFFPOSX1 DFFPOSX1_337 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__34_), .Q(\axi_araddr[2] ));
DFFPOSX1 DFFPOSX1_338 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__35_), .Q(\axi_araddr[3] ));
DFFPOSX1 DFFPOSX1_339 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__36_), .Q(\axi_araddr[4] ));
DFFPOSX1 DFFPOSX1_34 ( .CLK(SCLK), .D(_0counter_65_0__33_), .Q(counter_33_));
DFFPOSX1 DFFPOSX1_340 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__37_), .Q(\axi_araddr[5] ));
DFFPOSX1 DFFPOSX1_341 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__38_), .Q(\axi_araddr[6] ));
DFFPOSX1 DFFPOSX1_342 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__39_), .Q(\axi_araddr[7] ));
DFFPOSX1 DFFPOSX1_343 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__40_), .Q(\axi_araddr[8] ));
DFFPOSX1 DFFPOSX1_344 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__41_), .Q(\axi_araddr[9] ));
DFFPOSX1 DFFPOSX1_345 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__42_), .Q(\axi_araddr[10] ));
DFFPOSX1 DFFPOSX1_346 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__43_), .Q(\axi_araddr[11] ));
DFFPOSX1 DFFPOSX1_347 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__44_), .Q(\axi_araddr[12] ));
DFFPOSX1 DFFPOSX1_348 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__45_), .Q(\axi_araddr[13] ));
DFFPOSX1 DFFPOSX1_349 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__46_), .Q(\axi_araddr[14] ));
DFFPOSX1 DFFPOSX1_35 ( .CLK(SCLK), .D(_0counter_65_0__34_), .Q(counter_34_));
DFFPOSX1 DFFPOSX1_350 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__47_), .Q(\axi_araddr[15] ));
DFFPOSX1 DFFPOSX1_351 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__48_), .Q(\axi_araddr[16] ));
DFFPOSX1 DFFPOSX1_352 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__49_), .Q(\axi_araddr[17] ));
DFFPOSX1 DFFPOSX1_353 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__50_), .Q(\axi_araddr[18] ));
DFFPOSX1 DFFPOSX1_354 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__51_), .Q(\axi_araddr[19] ));
DFFPOSX1 DFFPOSX1_355 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__52_), .Q(\axi_araddr[20] ));
DFFPOSX1 DFFPOSX1_356 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__53_), .Q(\axi_araddr[21] ));
DFFPOSX1 DFFPOSX1_357 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__54_), .Q(\axi_araddr[22] ));
DFFPOSX1 DFFPOSX1_358 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__55_), .Q(\axi_araddr[23] ));
DFFPOSX1 DFFPOSX1_359 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__56_), .Q(\axi_araddr[24] ));
DFFPOSX1 DFFPOSX1_36 ( .CLK(SCLK), .D(_0counter_65_0__35_), .Q(counter_35_));
DFFPOSX1 DFFPOSX1_360 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__57_), .Q(\axi_araddr[25] ));
DFFPOSX1 DFFPOSX1_361 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__58_), .Q(\axi_araddr[26] ));
DFFPOSX1 DFFPOSX1_362 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__59_), .Q(\axi_araddr[27] ));
DFFPOSX1 DFFPOSX1_363 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__60_), .Q(\axi_araddr[28] ));
DFFPOSX1 DFFPOSX1_364 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__61_), .Q(\axi_araddr[29] ));
DFFPOSX1 DFFPOSX1_365 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__62_), .Q(\axi_araddr[30] ));
DFFPOSX1 DFFPOSX1_366 ( .CLK(CLK), .D(bus_sync_axi_bus__0reg_data3_63_0__63_), .Q(\axi_araddr[31] ));
DFFPOSX1 DFFPOSX1_367 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__0_), .Q(bus_sync_axi_bus_reg_data1_0_));
DFFPOSX1 DFFPOSX1_368 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__1_), .Q(bus_sync_axi_bus_reg_data1_1_));
DFFPOSX1 DFFPOSX1_369 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__2_), .Q(bus_sync_axi_bus_reg_data1_2_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(SCLK), .D(_0counter_65_0__36_), .Q(counter_36_));
DFFPOSX1 DFFPOSX1_370 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__3_), .Q(bus_sync_axi_bus_reg_data1_3_));
DFFPOSX1 DFFPOSX1_371 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__4_), .Q(bus_sync_axi_bus_reg_data1_4_));
DFFPOSX1 DFFPOSX1_372 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__5_), .Q(bus_sync_axi_bus_reg_data1_5_));
DFFPOSX1 DFFPOSX1_373 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__6_), .Q(bus_sync_axi_bus_reg_data1_6_));
DFFPOSX1 DFFPOSX1_374 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__7_), .Q(bus_sync_axi_bus_reg_data1_7_));
DFFPOSX1 DFFPOSX1_375 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__8_), .Q(bus_sync_axi_bus_reg_data1_8_));
DFFPOSX1 DFFPOSX1_376 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__9_), .Q(bus_sync_axi_bus_reg_data1_9_));
DFFPOSX1 DFFPOSX1_377 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__10_), .Q(bus_sync_axi_bus_reg_data1_10_));
DFFPOSX1 DFFPOSX1_378 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__11_), .Q(bus_sync_axi_bus_reg_data1_11_));
DFFPOSX1 DFFPOSX1_379 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__12_), .Q(bus_sync_axi_bus_reg_data1_12_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(SCLK), .D(_0counter_65_0__37_), .Q(counter_37_));
DFFPOSX1 DFFPOSX1_380 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__13_), .Q(bus_sync_axi_bus_reg_data1_13_));
DFFPOSX1 DFFPOSX1_381 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__14_), .Q(bus_sync_axi_bus_reg_data1_14_));
DFFPOSX1 DFFPOSX1_382 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__15_), .Q(bus_sync_axi_bus_reg_data1_15_));
DFFPOSX1 DFFPOSX1_383 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__16_), .Q(bus_sync_axi_bus_reg_data1_16_));
DFFPOSX1 DFFPOSX1_384 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__17_), .Q(bus_sync_axi_bus_reg_data1_17_));
DFFPOSX1 DFFPOSX1_385 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__18_), .Q(bus_sync_axi_bus_reg_data1_18_));
DFFPOSX1 DFFPOSX1_386 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__19_), .Q(bus_sync_axi_bus_reg_data1_19_));
DFFPOSX1 DFFPOSX1_387 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__20_), .Q(bus_sync_axi_bus_reg_data1_20_));
DFFPOSX1 DFFPOSX1_388 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__21_), .Q(bus_sync_axi_bus_reg_data1_21_));
DFFPOSX1 DFFPOSX1_389 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__22_), .Q(bus_sync_axi_bus_reg_data1_22_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(SCLK), .D(_0counter_65_0__38_), .Q(counter_38_));
DFFPOSX1 DFFPOSX1_390 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__23_), .Q(bus_sync_axi_bus_reg_data1_23_));
DFFPOSX1 DFFPOSX1_391 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__24_), .Q(bus_sync_axi_bus_reg_data1_24_));
DFFPOSX1 DFFPOSX1_392 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__25_), .Q(bus_sync_axi_bus_reg_data1_25_));
DFFPOSX1 DFFPOSX1_393 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__26_), .Q(bus_sync_axi_bus_reg_data1_26_));
DFFPOSX1 DFFPOSX1_394 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__27_), .Q(bus_sync_axi_bus_reg_data1_27_));
DFFPOSX1 DFFPOSX1_395 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__28_), .Q(bus_sync_axi_bus_reg_data1_28_));
DFFPOSX1 DFFPOSX1_396 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__29_), .Q(bus_sync_axi_bus_reg_data1_29_));
DFFPOSX1 DFFPOSX1_397 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__30_), .Q(bus_sync_axi_bus_reg_data1_30_));
DFFPOSX1 DFFPOSX1_398 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__31_), .Q(bus_sync_axi_bus_reg_data1_31_));
DFFPOSX1 DFFPOSX1_399 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__32_), .Q(bus_sync_axi_bus_reg_data1_32_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(SCLK), .D(_0counter_65_0__3_), .Q(counter_3_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(SCLK), .D(_0counter_65_0__39_), .Q(counter_39_));
DFFPOSX1 DFFPOSX1_400 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__33_), .Q(bus_sync_axi_bus_reg_data1_33_));
DFFPOSX1 DFFPOSX1_401 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__34_), .Q(bus_sync_axi_bus_reg_data1_34_));
DFFPOSX1 DFFPOSX1_402 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__35_), .Q(bus_sync_axi_bus_reg_data1_35_));
DFFPOSX1 DFFPOSX1_403 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__36_), .Q(bus_sync_axi_bus_reg_data1_36_));
DFFPOSX1 DFFPOSX1_404 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__37_), .Q(bus_sync_axi_bus_reg_data1_37_));
DFFPOSX1 DFFPOSX1_405 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__38_), .Q(bus_sync_axi_bus_reg_data1_38_));
DFFPOSX1 DFFPOSX1_406 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__39_), .Q(bus_sync_axi_bus_reg_data1_39_));
DFFPOSX1 DFFPOSX1_407 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__40_), .Q(bus_sync_axi_bus_reg_data1_40_));
DFFPOSX1 DFFPOSX1_408 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__41_), .Q(bus_sync_axi_bus_reg_data1_41_));
DFFPOSX1 DFFPOSX1_409 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__42_), .Q(bus_sync_axi_bus_reg_data1_42_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(SCLK), .D(_0counter_65_0__40_), .Q(counter_40_));
DFFPOSX1 DFFPOSX1_410 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__43_), .Q(bus_sync_axi_bus_reg_data1_43_));
DFFPOSX1 DFFPOSX1_411 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__44_), .Q(bus_sync_axi_bus_reg_data1_44_));
DFFPOSX1 DFFPOSX1_412 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__45_), .Q(bus_sync_axi_bus_reg_data1_45_));
DFFPOSX1 DFFPOSX1_413 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__46_), .Q(bus_sync_axi_bus_reg_data1_46_));
DFFPOSX1 DFFPOSX1_414 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__47_), .Q(bus_sync_axi_bus_reg_data1_47_));
DFFPOSX1 DFFPOSX1_415 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__48_), .Q(bus_sync_axi_bus_reg_data1_48_));
DFFPOSX1 DFFPOSX1_416 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__49_), .Q(bus_sync_axi_bus_reg_data1_49_));
DFFPOSX1 DFFPOSX1_417 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__50_), .Q(bus_sync_axi_bus_reg_data1_50_));
DFFPOSX1 DFFPOSX1_418 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__51_), .Q(bus_sync_axi_bus_reg_data1_51_));
DFFPOSX1 DFFPOSX1_419 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__52_), .Q(bus_sync_axi_bus_reg_data1_52_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(SCLK), .D(_0counter_65_0__41_), .Q(counter_41_));
DFFPOSX1 DFFPOSX1_420 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__53_), .Q(bus_sync_axi_bus_reg_data1_53_));
DFFPOSX1 DFFPOSX1_421 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__54_), .Q(bus_sync_axi_bus_reg_data1_54_));
DFFPOSX1 DFFPOSX1_422 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__55_), .Q(bus_sync_axi_bus_reg_data1_55_));
DFFPOSX1 DFFPOSX1_423 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__56_), .Q(bus_sync_axi_bus_reg_data1_56_));
DFFPOSX1 DFFPOSX1_424 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__57_), .Q(bus_sync_axi_bus_reg_data1_57_));
DFFPOSX1 DFFPOSX1_425 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__58_), .Q(bus_sync_axi_bus_reg_data1_58_));
DFFPOSX1 DFFPOSX1_426 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__59_), .Q(bus_sync_axi_bus_reg_data1_59_));
DFFPOSX1 DFFPOSX1_427 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__60_), .Q(bus_sync_axi_bus_reg_data1_60_));
DFFPOSX1 DFFPOSX1_428 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__61_), .Q(bus_sync_axi_bus_reg_data1_61_));
DFFPOSX1 DFFPOSX1_429 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__62_), .Q(bus_sync_axi_bus_reg_data1_62_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(SCLK), .D(_0counter_65_0__42_), .Q(counter_42_));
DFFPOSX1 DFFPOSX1_430 ( .CLK(SCLK), .D(bus_sync_axi_bus__0reg_data1_63_0__63_), .Q(bus_sync_axi_bus_reg_data1_63_));
DFFPOSX1 DFFPOSX1_431 ( .CLK(bus_sync_axi_bus_NCLK2), .D(bus_sync_axi_bus__0ECLK1_0_0_), .Q(bus_sync_axi_bus_ECLK1));
DFFPOSX1 DFFPOSX1_432 ( .CLK(bus_sync_axi_bus_NCLK2), .D(bus_sync_axi_bus__0EECLK1_0_0_), .Q(bus_sync_axi_bus_EECLK1));
DFFPOSX1 DFFPOSX1_433 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__0_), .Q(bus_sync_rdata_data_out_0_));
DFFPOSX1 DFFPOSX1_434 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__1_), .Q(bus_sync_rdata_data_out_1_));
DFFPOSX1 DFFPOSX1_435 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__2_), .Q(bus_sync_rdata_data_out_2_));
DFFPOSX1 DFFPOSX1_436 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__3_), .Q(bus_sync_rdata_data_out_3_));
DFFPOSX1 DFFPOSX1_437 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__4_), .Q(bus_sync_rdata_data_out_4_));
DFFPOSX1 DFFPOSX1_438 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__5_), .Q(bus_sync_rdata_data_out_5_));
DFFPOSX1 DFFPOSX1_439 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__6_), .Q(bus_sync_rdata_data_out_6_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(SCLK), .D(_0counter_65_0__43_), .Q(counter_43_));
DFFPOSX1 DFFPOSX1_440 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__7_), .Q(bus_sync_rdata_data_out_7_));
DFFPOSX1 DFFPOSX1_441 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__8_), .Q(bus_sync_rdata_data_out_8_));
DFFPOSX1 DFFPOSX1_442 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__9_), .Q(bus_sync_rdata_data_out_9_));
DFFPOSX1 DFFPOSX1_443 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__10_), .Q(bus_sync_rdata_data_out_10_));
DFFPOSX1 DFFPOSX1_444 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__11_), .Q(bus_sync_rdata_data_out_11_));
DFFPOSX1 DFFPOSX1_445 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__12_), .Q(bus_sync_rdata_data_out_12_));
DFFPOSX1 DFFPOSX1_446 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__13_), .Q(bus_sync_rdata_data_out_13_));
DFFPOSX1 DFFPOSX1_447 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__14_), .Q(bus_sync_rdata_data_out_14_));
DFFPOSX1 DFFPOSX1_448 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__15_), .Q(bus_sync_rdata_data_out_15_));
DFFPOSX1 DFFPOSX1_449 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__16_), .Q(bus_sync_rdata_data_out_16_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(SCLK), .D(_0counter_65_0__44_), .Q(counter_44_));
DFFPOSX1 DFFPOSX1_450 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__17_), .Q(bus_sync_rdata_data_out_17_));
DFFPOSX1 DFFPOSX1_451 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__18_), .Q(bus_sync_rdata_data_out_18_));
DFFPOSX1 DFFPOSX1_452 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__19_), .Q(bus_sync_rdata_data_out_19_));
DFFPOSX1 DFFPOSX1_453 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__20_), .Q(bus_sync_rdata_data_out_20_));
DFFPOSX1 DFFPOSX1_454 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__21_), .Q(bus_sync_rdata_data_out_21_));
DFFPOSX1 DFFPOSX1_455 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__22_), .Q(bus_sync_rdata_data_out_22_));
DFFPOSX1 DFFPOSX1_456 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__23_), .Q(bus_sync_rdata_data_out_23_));
DFFPOSX1 DFFPOSX1_457 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__24_), .Q(bus_sync_rdata_data_out_24_));
DFFPOSX1 DFFPOSX1_458 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__25_), .Q(bus_sync_rdata_data_out_25_));
DFFPOSX1 DFFPOSX1_459 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__26_), .Q(bus_sync_rdata_data_out_26_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(SCLK), .D(_0counter_65_0__45_), .Q(counter_45_));
DFFPOSX1 DFFPOSX1_460 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__27_), .Q(bus_sync_rdata_data_out_27_));
DFFPOSX1 DFFPOSX1_461 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__28_), .Q(bus_sync_rdata_data_out_28_));
DFFPOSX1 DFFPOSX1_462 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__29_), .Q(bus_sync_rdata_data_out_29_));
DFFPOSX1 DFFPOSX1_463 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__30_), .Q(bus_sync_rdata_data_out_30_));
DFFPOSX1 DFFPOSX1_464 ( .CLK(SCLK), .D(bus_sync_rdata__0reg_data3_31_0__31_), .Q(bus_sync_rdata_data_out_31_));
DFFPOSX1 DFFPOSX1_465 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__0_), .Q(bus_sync_rdata_reg_data1_0_));
DFFPOSX1 DFFPOSX1_466 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__1_), .Q(bus_sync_rdata_reg_data1_1_));
DFFPOSX1 DFFPOSX1_467 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__2_), .Q(bus_sync_rdata_reg_data1_2_));
DFFPOSX1 DFFPOSX1_468 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__3_), .Q(bus_sync_rdata_reg_data1_3_));
DFFPOSX1 DFFPOSX1_469 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__4_), .Q(bus_sync_rdata_reg_data1_4_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(SCLK), .D(_0counter_65_0__46_), .Q(counter_46_));
DFFPOSX1 DFFPOSX1_470 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__5_), .Q(bus_sync_rdata_reg_data1_5_));
DFFPOSX1 DFFPOSX1_471 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__6_), .Q(bus_sync_rdata_reg_data1_6_));
DFFPOSX1 DFFPOSX1_472 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__7_), .Q(bus_sync_rdata_reg_data1_7_));
DFFPOSX1 DFFPOSX1_473 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__8_), .Q(bus_sync_rdata_reg_data1_8_));
DFFPOSX1 DFFPOSX1_474 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__9_), .Q(bus_sync_rdata_reg_data1_9_));
DFFPOSX1 DFFPOSX1_475 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__10_), .Q(bus_sync_rdata_reg_data1_10_));
DFFPOSX1 DFFPOSX1_476 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__11_), .Q(bus_sync_rdata_reg_data1_11_));
DFFPOSX1 DFFPOSX1_477 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__12_), .Q(bus_sync_rdata_reg_data1_12_));
DFFPOSX1 DFFPOSX1_478 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__13_), .Q(bus_sync_rdata_reg_data1_13_));
DFFPOSX1 DFFPOSX1_479 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__14_), .Q(bus_sync_rdata_reg_data1_14_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(SCLK), .D(_0counter_65_0__47_), .Q(counter_47_));
DFFPOSX1 DFFPOSX1_480 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__15_), .Q(bus_sync_rdata_reg_data1_15_));
DFFPOSX1 DFFPOSX1_481 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__16_), .Q(bus_sync_rdata_reg_data1_16_));
DFFPOSX1 DFFPOSX1_482 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__17_), .Q(bus_sync_rdata_reg_data1_17_));
DFFPOSX1 DFFPOSX1_483 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__18_), .Q(bus_sync_rdata_reg_data1_18_));
DFFPOSX1 DFFPOSX1_484 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__19_), .Q(bus_sync_rdata_reg_data1_19_));
DFFPOSX1 DFFPOSX1_485 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__20_), .Q(bus_sync_rdata_reg_data1_20_));
DFFPOSX1 DFFPOSX1_486 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__21_), .Q(bus_sync_rdata_reg_data1_21_));
DFFPOSX1 DFFPOSX1_487 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__22_), .Q(bus_sync_rdata_reg_data1_22_));
DFFPOSX1 DFFPOSX1_488 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__23_), .Q(bus_sync_rdata_reg_data1_23_));
DFFPOSX1 DFFPOSX1_489 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__24_), .Q(bus_sync_rdata_reg_data1_24_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(SCLK), .D(_0counter_65_0__48_), .Q(counter_48_));
DFFPOSX1 DFFPOSX1_490 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__25_), .Q(bus_sync_rdata_reg_data1_25_));
DFFPOSX1 DFFPOSX1_491 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__26_), .Q(bus_sync_rdata_reg_data1_26_));
DFFPOSX1 DFFPOSX1_492 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__27_), .Q(bus_sync_rdata_reg_data1_27_));
DFFPOSX1 DFFPOSX1_493 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__28_), .Q(bus_sync_rdata_reg_data1_28_));
DFFPOSX1 DFFPOSX1_494 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__29_), .Q(bus_sync_rdata_reg_data1_29_));
DFFPOSX1 DFFPOSX1_495 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__30_), .Q(bus_sync_rdata_reg_data1_30_));
DFFPOSX1 DFFPOSX1_496 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data1_31_0__31_), .Q(bus_sync_rdata_reg_data1_31_));
DFFPOSX1 DFFPOSX1_497 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__0_), .Q(bus_sync_rdata_reg_data2_0_));
DFFPOSX1 DFFPOSX1_498 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__1_), .Q(bus_sync_rdata_reg_data2_1_));
DFFPOSX1 DFFPOSX1_499 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__2_), .Q(bus_sync_rdata_reg_data2_2_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(SCLK), .D(_0counter_65_0__4_), .Q(counter_4_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(SCLK), .D(_0counter_65_0__49_), .Q(counter_49_));
DFFPOSX1 DFFPOSX1_500 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__3_), .Q(bus_sync_rdata_reg_data2_3_));
DFFPOSX1 DFFPOSX1_501 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__4_), .Q(bus_sync_rdata_reg_data2_4_));
DFFPOSX1 DFFPOSX1_502 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__5_), .Q(bus_sync_rdata_reg_data2_5_));
DFFPOSX1 DFFPOSX1_503 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__6_), .Q(bus_sync_rdata_reg_data2_6_));
DFFPOSX1 DFFPOSX1_504 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__7_), .Q(bus_sync_rdata_reg_data2_7_));
DFFPOSX1 DFFPOSX1_505 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__8_), .Q(bus_sync_rdata_reg_data2_8_));
DFFPOSX1 DFFPOSX1_506 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__9_), .Q(bus_sync_rdata_reg_data2_9_));
DFFPOSX1 DFFPOSX1_507 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__10_), .Q(bus_sync_rdata_reg_data2_10_));
DFFPOSX1 DFFPOSX1_508 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__11_), .Q(bus_sync_rdata_reg_data2_11_));
DFFPOSX1 DFFPOSX1_509 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__12_), .Q(bus_sync_rdata_reg_data2_12_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(SCLK), .D(_0counter_65_0__50_), .Q(counter_50_));
DFFPOSX1 DFFPOSX1_510 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__13_), .Q(bus_sync_rdata_reg_data2_13_));
DFFPOSX1 DFFPOSX1_511 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__14_), .Q(bus_sync_rdata_reg_data2_14_));
DFFPOSX1 DFFPOSX1_512 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__15_), .Q(bus_sync_rdata_reg_data2_15_));
DFFPOSX1 DFFPOSX1_513 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__16_), .Q(bus_sync_rdata_reg_data2_16_));
DFFPOSX1 DFFPOSX1_514 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__17_), .Q(bus_sync_rdata_reg_data2_17_));
DFFPOSX1 DFFPOSX1_515 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__18_), .Q(bus_sync_rdata_reg_data2_18_));
DFFPOSX1 DFFPOSX1_516 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__19_), .Q(bus_sync_rdata_reg_data2_19_));
DFFPOSX1 DFFPOSX1_517 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__20_), .Q(bus_sync_rdata_reg_data2_20_));
DFFPOSX1 DFFPOSX1_518 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__21_), .Q(bus_sync_rdata_reg_data2_21_));
DFFPOSX1 DFFPOSX1_519 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__22_), .Q(bus_sync_rdata_reg_data2_22_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(SCLK), .D(_0counter_65_0__51_), .Q(counter_51_));
DFFPOSX1 DFFPOSX1_520 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__23_), .Q(bus_sync_rdata_reg_data2_23_));
DFFPOSX1 DFFPOSX1_521 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__24_), .Q(bus_sync_rdata_reg_data2_24_));
DFFPOSX1 DFFPOSX1_522 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__25_), .Q(bus_sync_rdata_reg_data2_25_));
DFFPOSX1 DFFPOSX1_523 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__26_), .Q(bus_sync_rdata_reg_data2_26_));
DFFPOSX1 DFFPOSX1_524 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__27_), .Q(bus_sync_rdata_reg_data2_27_));
DFFPOSX1 DFFPOSX1_525 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__28_), .Q(bus_sync_rdata_reg_data2_28_));
DFFPOSX1 DFFPOSX1_526 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__29_), .Q(bus_sync_rdata_reg_data2_29_));
DFFPOSX1 DFFPOSX1_527 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__30_), .Q(bus_sync_rdata_reg_data2_30_));
DFFPOSX1 DFFPOSX1_528 ( .CLK(CLK), .D(bus_sync_rdata__0reg_data2_31_0__31_), .Q(bus_sync_rdata_reg_data2_31_));
DFFPOSX1 DFFPOSX1_529 ( .CLK(bus_sync_rdata_NCLK1), .D(bus_sync_rdata__0EECLK2_0_0_), .Q(bus_sync_rdata_EECLK2));
DFFPOSX1 DFFPOSX1_53 ( .CLK(SCLK), .D(_0counter_65_0__52_), .Q(counter_52_));
DFFPOSX1 DFFPOSX1_530 ( .CLK(bus_sync_rdata_NCLK1), .D(bus_sync_rdata__0ECLK2_0_0_), .Q(bus_sync_rdata_ECLK2));
DFFPOSX1 DFFPOSX1_531 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data2_3_0__0_), .Q(bus_sync_state_machine_reg_data2_0_));
DFFPOSX1 DFFPOSX1_532 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data2_3_0__1_), .Q(bus_sync_state_machine_reg_data2_1_));
DFFPOSX1 DFFPOSX1_533 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data2_3_0__2_), .Q(bus_sync_state_machine_reg_data2_2_));
DFFPOSX1 DFFPOSX1_534 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data2_3_0__3_), .Q(bus_sync_state_machine_reg_data2_3_));
DFFPOSX1 DFFPOSX1_535 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data3_3_0__0_), .Q(fini_spi_clk));
DFFPOSX1 DFFPOSX1_536 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data3_3_0__1_), .Q(re_clk));
DFFPOSX1 DFFPOSX1_537 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data3_3_0__2_), .Q(we_clk));
DFFPOSX1 DFFPOSX1_538 ( .CLK(CLK), .D(bus_sync_state_machine__0reg_data3_3_0__3_), .Q(PICORV_RST));
DFFPOSX1 DFFPOSX1_539 ( .CLK(SCLK), .D(bus_sync_state_machine__0reg_data1_3_0__0_), .Q(bus_sync_state_machine_reg_data1_0_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(SCLK), .D(_0counter_65_0__53_), .Q(counter_53_));
DFFPOSX1 DFFPOSX1_540 ( .CLK(SCLK), .D(bus_sync_state_machine__0reg_data1_3_0__1_), .Q(bus_sync_state_machine_reg_data1_1_));
DFFPOSX1 DFFPOSX1_541 ( .CLK(SCLK), .D(bus_sync_state_machine__0reg_data1_3_0__2_), .Q(bus_sync_state_machine_reg_data1_2_));
DFFPOSX1 DFFPOSX1_542 ( .CLK(SCLK), .D(bus_sync_state_machine__0reg_data1_3_0__3_), .Q(bus_sync_state_machine_reg_data1_3_));
DFFPOSX1 DFFPOSX1_543 ( .CLK(bus_sync_state_machine_NCLK2), .D(bus_sync_state_machine__0ECLK1_0_0_), .Q(bus_sync_state_machine_ECLK1));
DFFPOSX1 DFFPOSX1_544 ( .CLK(bus_sync_state_machine_NCLK2), .D(bus_sync_state_machine__0EECLK1_0_0_), .Q(bus_sync_state_machine_EECLK1));
DFFPOSX1 DFFPOSX1_545 ( .CLK(SCLK), .D(bus_sync_status__0reg_data3_2_0__0_), .Q(bus_sync_status_data_out_0_));
DFFPOSX1 DFFPOSX1_546 ( .CLK(SCLK), .D(bus_sync_status__0reg_data3_2_0__1_), .Q(bus_sync_status_data_out_1_));
DFFPOSX1 DFFPOSX1_547 ( .CLK(SCLK), .D(bus_sync_status__0reg_data3_2_0__2_), .Q(bus_sync_status_data_out_2_));
DFFPOSX1 DFFPOSX1_548 ( .CLK(CLK), .D(bus_sync_status__0reg_data1_2_0__0_), .Q(bus_sync_status_reg_data1_0_));
DFFPOSX1 DFFPOSX1_549 ( .CLK(CLK), .D(bus_sync_status__0reg_data1_2_0__1_), .Q(bus_sync_status_reg_data1_1_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(SCLK), .D(_0counter_65_0__54_), .Q(counter_54_));
DFFPOSX1 DFFPOSX1_550 ( .CLK(CLK), .D(bus_sync_status__0reg_data1_2_0__2_), .Q(bus_sync_status_reg_data1_2_));
DFFPOSX1 DFFPOSX1_551 ( .CLK(CLK), .D(bus_sync_status__0reg_data2_2_0__0_), .Q(bus_sync_status_reg_data2_0_));
DFFPOSX1 DFFPOSX1_552 ( .CLK(CLK), .D(bus_sync_status__0reg_data2_2_0__1_), .Q(bus_sync_status_reg_data2_1_));
DFFPOSX1 DFFPOSX1_553 ( .CLK(CLK), .D(bus_sync_status__0reg_data2_2_0__2_), .Q(bus_sync_status_reg_data2_2_));
DFFPOSX1 DFFPOSX1_554 ( .CLK(bus_sync_status_NCLK1), .D(bus_sync_status__0EECLK2_0_0_), .Q(bus_sync_status_EECLK2));
DFFPOSX1 DFFPOSX1_555 ( .CLK(bus_sync_status_NCLK1), .D(bus_sync_status__0ECLK2_0_0_), .Q(bus_sync_status_ECLK2));
DFFPOSX1 DFFPOSX1_56 ( .CLK(SCLK), .D(_0counter_65_0__55_), .Q(counter_55_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(SCLK), .D(_0counter_65_0__56_), .Q(counter_56_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(SCLK), .D(_0counter_65_0__57_), .Q(counter_57_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(SCLK), .D(_0counter_65_0__58_), .Q(counter_58_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(SCLK), .D(_0counter_65_0__5_), .Q(counter_5_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(SCLK), .D(_0counter_65_0__59_), .Q(counter_59_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(SCLK), .D(_0counter_65_0__60_), .Q(counter_60_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(SCLK), .D(_0counter_65_0__61_), .Q(counter_61_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(SCLK), .D(_0counter_65_0__62_), .Q(counter_62_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(SCLK), .D(_0counter_65_0__63_), .Q(counter_63_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(SCLK), .D(_0counter_65_0__64_), .Q(counter_64_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(SCLK), .D(_0counter_65_0__65_), .Q(counter_65_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(SCLK), .D(_0fini_spi_0_0_), .Q(fini_spi));
DFFPOSX1 DFFPOSX1_68 ( .CLK(SCLK), .D(_0bus_cap_31_0__0_), .Q(bus_cap_0_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(SCLK), .D(_0bus_cap_31_0__1_), .Q(bus_cap_1_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(SCLK), .D(_0counter_65_0__6_), .Q(counter_6_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(SCLK), .D(_0bus_cap_31_0__2_), .Q(bus_cap_2_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(SCLK), .D(_0bus_cap_31_0__3_), .Q(bus_cap_3_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(SCLK), .D(_0bus_cap_31_0__4_), .Q(bus_cap_4_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(SCLK), .D(_0bus_cap_31_0__5_), .Q(bus_cap_5_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(SCLK), .D(_0bus_cap_31_0__6_), .Q(bus_cap_6_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(SCLK), .D(_0bus_cap_31_0__7_), .Q(bus_cap_7_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(SCLK), .D(_0bus_cap_31_0__8_), .Q(bus_cap_8_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(SCLK), .D(_0bus_cap_31_0__9_), .Q(bus_cap_9_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(SCLK), .D(_0bus_cap_31_0__10_), .Q(bus_cap_10_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(SCLK), .D(_0bus_cap_31_0__11_), .Q(bus_cap_11_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(SCLK), .D(_0counter_65_0__7_), .Q(counter_7_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(SCLK), .D(_0bus_cap_31_0__12_), .Q(bus_cap_12_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(SCLK), .D(_0bus_cap_31_0__13_), .Q(bus_cap_13_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(SCLK), .D(_0bus_cap_31_0__14_), .Q(bus_cap_14_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(SCLK), .D(_0bus_cap_31_0__15_), .Q(bus_cap_15_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(SCLK), .D(_0bus_cap_31_0__16_), .Q(bus_cap_16_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(SCLK), .D(_0bus_cap_31_0__17_), .Q(bus_cap_17_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(SCLK), .D(_0bus_cap_31_0__18_), .Q(bus_cap_18_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(SCLK), .D(_0bus_cap_31_0__19_), .Q(bus_cap_19_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(SCLK), .D(_0bus_cap_31_0__20_), .Q(bus_cap_20_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(SCLK), .D(_0bus_cap_31_0__21_), .Q(bus_cap_21_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(SCLK), .D(_0counter_65_0__8_), .Q(counter_8_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(SCLK), .D(_0bus_cap_31_0__22_), .Q(bus_cap_22_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(SCLK), .D(_0bus_cap_31_0__23_), .Q(bus_cap_23_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(SCLK), .D(_0bus_cap_31_0__24_), .Q(bus_cap_24_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(SCLK), .D(_0bus_cap_31_0__25_), .Q(bus_cap_25_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(SCLK), .D(_0bus_cap_31_0__26_), .Q(bus_cap_26_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(SCLK), .D(_0bus_cap_31_0__27_), .Q(bus_cap_27_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(SCLK), .D(_0bus_cap_31_0__28_), .Q(bus_cap_28_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(SCLK), .D(_0bus_cap_31_0__29_), .Q(bus_cap_29_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(SCLK), .D(_0bus_cap_31_0__30_), .Q(bus_cap_30_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(SCLK), .D(_0bus_cap_31_0__31_), .Q(DOUT));
INVX1 INVX1_1 ( .A(axi_bvalid), .Y(_abc_4268_new_n560_));
INVX1 INVX1_10 ( .A(fini_spi_clk), .Y(_abc_4268_new_n606_));
INVX1 INVX1_11 ( .A(axi_awready), .Y(_abc_4268_new_n610_));
INVX1 INVX1_12 ( .A(_abc_4268_new_n616_), .Y(_abc_4268_new_n617_));
INVX1 INVX1_13 ( .A(counter_1_), .Y(_abc_4268_new_n618_));
INVX1 INVX1_14 ( .A(_abc_4268_new_n621_), .Y(_abc_4268_new_n622_));
INVX1 INVX1_15 ( .A(_abc_4268_new_n624_), .Y(_abc_4268_new_n625_));
INVX1 INVX1_16 ( .A(_abc_4268_new_n626_), .Y(_abc_4268_new_n627_));
INVX1 INVX1_17 ( .A(_abc_4268_new_n628_), .Y(_abc_4268_new_n629_));
INVX1 INVX1_18 ( .A(_abc_4268_new_n630_), .Y(_abc_4268_new_n631_));
INVX1 INVX1_19 ( .A(_abc_4268_new_n633_), .Y(_abc_4268_new_n634_));
INVX1 INVX1_2 ( .A(axi_wready), .Y(_abc_4268_new_n566_));
INVX1 INVX1_20 ( .A(_abc_4268_new_n635_), .Y(_abc_4268_new_n636_));
INVX1 INVX1_21 ( .A(_abc_4268_new_n639_), .Y(_abc_4268_new_n640_));
INVX1 INVX1_22 ( .A(_abc_4268_new_n641_), .Y(_abc_4268_new_n642_));
INVX1 INVX1_23 ( .A(_abc_4268_new_n644_), .Y(_abc_4268_new_n645_));
INVX1 INVX1_24 ( .A(_abc_4268_new_n646_), .Y(_abc_4268_new_n647_));
INVX1 INVX1_25 ( .A(_abc_4268_new_n651_), .Y(_abc_4268_new_n652_));
INVX1 INVX1_26 ( .A(_abc_4268_new_n653_), .Y(_abc_4268_new_n654_));
INVX1 INVX1_27 ( .A(_abc_4268_new_n656_), .Y(_abc_4268_new_n657_));
INVX1 INVX1_28 ( .A(_abc_4268_new_n658_), .Y(_abc_4268_new_n659_));
INVX1 INVX1_29 ( .A(_abc_4268_new_n662_), .Y(_abc_4268_new_n663_));
INVX1 INVX1_3 ( .A(axi_arready), .Y(_abc_4268_new_n575_));
INVX1 INVX1_30 ( .A(_abc_4268_new_n664_), .Y(_abc_4268_new_n665_));
INVX1 INVX1_31 ( .A(_abc_4268_new_n667_), .Y(_abc_4268_new_n668_));
INVX1 INVX1_32 ( .A(counter_18_), .Y(_abc_4268_new_n669_));
INVX1 INVX1_33 ( .A(counter_19_), .Y(_abc_4268_new_n670_));
INVX1 INVX1_34 ( .A(axi_rready), .Y(_abc_4268_new_n955_));
INVX1 INVX1_35 ( .A(CEB), .Y(_abc_4268_new_n1083_));
INVX1 INVX1_36 ( .A(_abc_4268_new_n1085_), .Y(_abc_4268_new_n1087_));
INVX1 INVX1_37 ( .A(_abc_4268_new_n1216_), .Y(_abc_4268_new_n1218_));
INVX1 INVX1_38 ( .A(_abc_4268_new_n1470_), .Y(_0counter_65_0__0_));
INVX1 INVX1_39 ( .A(_abc_4268_new_n1537_), .Y(_abc_4268_new_n1538_));
INVX1 INVX1_4 ( .A(re_clk), .Y(_abc_4268_new_n578_));
INVX1 INVX1_40 ( .A(counter_0_), .Y(_abc_4268_new_n1547_));
INVX1 INVX1_41 ( .A(bus_sync_axi_bus_EECLK1), .Y(bus_sync_axi_bus__abc_3879_new_n393_));
INVX1 INVX1_42 ( .A(CLK), .Y(bus_sync_axi_bus_NCLK2));
INVX1 INVX1_43 ( .A(bus_sync_rdata_EECLK2), .Y(bus_sync_rdata__abc_3653_new_n265_));
INVX1 INVX1_44 ( .A(CLK), .Y(bus_sync_rdata_NCLK1));
INVX1 INVX1_45 ( .A(bus_sync_state_machine_EECLK1), .Y(bus_sync_state_machine__abc_3850_new_n33_));
INVX1 INVX1_46 ( .A(CLK), .Y(bus_sync_state_machine_NCLK2));
INVX1 INVX1_47 ( .A(bus_sync_status_EECLK2), .Y(bus_sync_status__abc_3630_new_n27_));
INVX1 INVX1_48 ( .A(CLK), .Y(bus_sync_status_NCLK1));
INVX1 INVX1_5 ( .A(_abc_4268_new_n580_), .Y(_abc_4268_new_n581_));
INVX1 INVX1_6 ( .A(we_clk), .Y(_abc_4268_new_n583_));
INVX1 INVX1_7 ( .A(axi_rvalid), .Y(_abc_4268_new_n590_));
INVX1 INVX1_8 ( .A(_abc_4268_new_n585_), .Y(_abc_4268_new_n602_));
INVX1 INVX1_9 ( .A(RST), .Y(_abc_4268_new_n605_));
OR2X2 OR2X2_1 ( .A(_abc_4268_new_n559_), .B(_abc_4268_new_n562_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_7_));
OR2X2 OR2X2_10 ( .A(_abc_4268_new_n594_), .B(state_4_), .Y(axi_arvalid));
OR2X2 OR2X2_100 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n782_), .Y(_abc_4268_new_n783_));
OR2X2 OR2X2_101 ( .A(_abc_4268_new_n701_), .B(bus_cap_11_), .Y(_abc_4268_new_n786_));
OR2X2 OR2X2_102 ( .A(_abc_4268_new_n676_), .B(bus_cap_10_), .Y(_abc_4268_new_n787_));
OR2X2 OR2X2_103 ( .A(_abc_4268_new_n788_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n789_));
OR2X2 OR2X2_104 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n790_), .Y(_abc_4268_new_n791_));
OR2X2 OR2X2_105 ( .A(_abc_4268_new_n701_), .B(bus_cap_12_), .Y(_abc_4268_new_n794_));
OR2X2 OR2X2_106 ( .A(_abc_4268_new_n676_), .B(bus_cap_11_), .Y(_abc_4268_new_n795_));
OR2X2 OR2X2_107 ( .A(_abc_4268_new_n796_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n797_));
OR2X2 OR2X2_108 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n798_), .Y(_abc_4268_new_n799_));
OR2X2 OR2X2_109 ( .A(_abc_4268_new_n701_), .B(bus_cap_13_), .Y(_abc_4268_new_n802_));
OR2X2 OR2X2_11 ( .A(state_7_), .B(state_5_), .Y(_abc_4268_new_n596_));
OR2X2 OR2X2_110 ( .A(_abc_4268_new_n676_), .B(bus_cap_12_), .Y(_abc_4268_new_n803_));
OR2X2 OR2X2_111 ( .A(_abc_4268_new_n804_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n805_));
OR2X2 OR2X2_112 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n806_), .Y(_abc_4268_new_n807_));
OR2X2 OR2X2_113 ( .A(_abc_4268_new_n701_), .B(bus_cap_14_), .Y(_abc_4268_new_n810_));
OR2X2 OR2X2_114 ( .A(_abc_4268_new_n676_), .B(bus_cap_13_), .Y(_abc_4268_new_n811_));
OR2X2 OR2X2_115 ( .A(_abc_4268_new_n812_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n813_));
OR2X2 OR2X2_116 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n814_), .Y(_abc_4268_new_n815_));
OR2X2 OR2X2_117 ( .A(_abc_4268_new_n701_), .B(bus_cap_15_), .Y(_abc_4268_new_n818_));
OR2X2 OR2X2_118 ( .A(_abc_4268_new_n676_), .B(bus_cap_14_), .Y(_abc_4268_new_n819_));
OR2X2 OR2X2_119 ( .A(_abc_4268_new_n820_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n821_));
OR2X2 OR2X2_12 ( .A(_abc_4268_new_n564_), .B(_abc_4268_new_n596_), .Y(axi_awvalid));
OR2X2 OR2X2_120 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n822_), .Y(_abc_4268_new_n823_));
OR2X2 OR2X2_121 ( .A(_abc_4268_new_n701_), .B(bus_cap_16_), .Y(_abc_4268_new_n826_));
OR2X2 OR2X2_122 ( .A(_abc_4268_new_n676_), .B(bus_cap_15_), .Y(_abc_4268_new_n827_));
OR2X2 OR2X2_123 ( .A(_abc_4268_new_n828_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n829_));
OR2X2 OR2X2_124 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n830_), .Y(_abc_4268_new_n831_));
OR2X2 OR2X2_125 ( .A(_abc_4268_new_n701_), .B(bus_cap_17_), .Y(_abc_4268_new_n834_));
OR2X2 OR2X2_126 ( .A(_abc_4268_new_n676_), .B(bus_cap_16_), .Y(_abc_4268_new_n835_));
OR2X2 OR2X2_127 ( .A(_abc_4268_new_n836_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n837_));
OR2X2 OR2X2_128 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n838_), .Y(_abc_4268_new_n839_));
OR2X2 OR2X2_129 ( .A(_abc_4268_new_n701_), .B(bus_cap_18_), .Y(_abc_4268_new_n842_));
OR2X2 OR2X2_13 ( .A(state_1_), .B(state_4_), .Y(_abc_4268_new_n598_));
OR2X2 OR2X2_130 ( .A(_abc_4268_new_n676_), .B(bus_cap_17_), .Y(_abc_4268_new_n843_));
OR2X2 OR2X2_131 ( .A(_abc_4268_new_n844_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n845_));
OR2X2 OR2X2_132 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n846_), .Y(_abc_4268_new_n847_));
OR2X2 OR2X2_133 ( .A(_abc_4268_new_n701_), .B(bus_cap_19_), .Y(_abc_4268_new_n850_));
OR2X2 OR2X2_134 ( .A(_abc_4268_new_n676_), .B(bus_cap_18_), .Y(_abc_4268_new_n851_));
OR2X2 OR2X2_135 ( .A(_abc_4268_new_n852_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n853_));
OR2X2 OR2X2_136 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n854_), .Y(_abc_4268_new_n855_));
OR2X2 OR2X2_137 ( .A(_abc_4268_new_n701_), .B(bus_cap_20_), .Y(_abc_4268_new_n858_));
OR2X2 OR2X2_138 ( .A(_abc_4268_new_n676_), .B(bus_cap_19_), .Y(_abc_4268_new_n859_));
OR2X2 OR2X2_139 ( .A(_abc_4268_new_n860_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n861_));
OR2X2 OR2X2_14 ( .A(_abc_4268_new_n596_), .B(_abc_4268_new_n598_), .Y(_abc_4268_new_n599_));
OR2X2 OR2X2_140 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n862_), .Y(_abc_4268_new_n863_));
OR2X2 OR2X2_141 ( .A(_abc_4268_new_n701_), .B(bus_cap_21_), .Y(_abc_4268_new_n866_));
OR2X2 OR2X2_142 ( .A(_abc_4268_new_n676_), .B(bus_cap_20_), .Y(_abc_4268_new_n867_));
OR2X2 OR2X2_143 ( .A(_abc_4268_new_n868_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n869_));
OR2X2 OR2X2_144 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n870_), .Y(_abc_4268_new_n871_));
OR2X2 OR2X2_145 ( .A(_abc_4268_new_n701_), .B(bus_cap_22_), .Y(_abc_4268_new_n874_));
OR2X2 OR2X2_146 ( .A(_abc_4268_new_n676_), .B(bus_cap_21_), .Y(_abc_4268_new_n875_));
OR2X2 OR2X2_147 ( .A(_abc_4268_new_n876_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n877_));
OR2X2 OR2X2_148 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n878_), .Y(_abc_4268_new_n879_));
OR2X2 OR2X2_149 ( .A(_abc_4268_new_n701_), .B(bus_cap_23_), .Y(_abc_4268_new_n882_));
OR2X2 OR2X2_15 ( .A(_abc_4268_new_n564_), .B(_abc_4268_new_n594_), .Y(_abc_4268_new_n600_));
OR2X2 OR2X2_150 ( .A(_abc_4268_new_n676_), .B(bus_cap_22_), .Y(_abc_4268_new_n883_));
OR2X2 OR2X2_151 ( .A(_abc_4268_new_n884_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n885_));
OR2X2 OR2X2_152 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n886_), .Y(_abc_4268_new_n887_));
OR2X2 OR2X2_153 ( .A(_abc_4268_new_n701_), .B(bus_cap_24_), .Y(_abc_4268_new_n890_));
OR2X2 OR2X2_154 ( .A(_abc_4268_new_n676_), .B(bus_cap_23_), .Y(_abc_4268_new_n891_));
OR2X2 OR2X2_155 ( .A(_abc_4268_new_n892_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n893_));
OR2X2 OR2X2_156 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n894_), .Y(_abc_4268_new_n895_));
OR2X2 OR2X2_157 ( .A(_abc_4268_new_n701_), .B(bus_cap_25_), .Y(_abc_4268_new_n898_));
OR2X2 OR2X2_158 ( .A(_abc_4268_new_n676_), .B(bus_cap_24_), .Y(_abc_4268_new_n899_));
OR2X2 OR2X2_159 ( .A(_abc_4268_new_n900_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n901_));
OR2X2 OR2X2_16 ( .A(_abc_4268_new_n599_), .B(_abc_4268_new_n600_), .Y(busy));
OR2X2 OR2X2_160 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n902_), .Y(_abc_4268_new_n903_));
OR2X2 OR2X2_161 ( .A(_abc_4268_new_n701_), .B(bus_cap_26_), .Y(_abc_4268_new_n906_));
OR2X2 OR2X2_162 ( .A(_abc_4268_new_n676_), .B(bus_cap_25_), .Y(_abc_4268_new_n907_));
OR2X2 OR2X2_163 ( .A(_abc_4268_new_n908_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n909_));
OR2X2 OR2X2_164 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n910_), .Y(_abc_4268_new_n911_));
OR2X2 OR2X2_165 ( .A(_abc_4268_new_n701_), .B(bus_cap_27_), .Y(_abc_4268_new_n914_));
OR2X2 OR2X2_166 ( .A(_abc_4268_new_n676_), .B(bus_cap_26_), .Y(_abc_4268_new_n915_));
OR2X2 OR2X2_167 ( .A(_abc_4268_new_n916_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n917_));
OR2X2 OR2X2_168 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n918_), .Y(_abc_4268_new_n919_));
OR2X2 OR2X2_169 ( .A(_abc_4268_new_n701_), .B(bus_cap_28_), .Y(_abc_4268_new_n922_));
OR2X2 OR2X2_17 ( .A(_abc_4268_new_n607_), .B(_abc_4268_new_n605_), .Y(_abc_4268_new_n608_));
OR2X2 OR2X2_170 ( .A(_abc_4268_new_n676_), .B(bus_cap_27_), .Y(_abc_4268_new_n923_));
OR2X2 OR2X2_171 ( .A(_abc_4268_new_n924_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n925_));
OR2X2 OR2X2_172 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n926_), .Y(_abc_4268_new_n927_));
OR2X2 OR2X2_173 ( .A(_abc_4268_new_n701_), .B(bus_cap_29_), .Y(_abc_4268_new_n930_));
OR2X2 OR2X2_174 ( .A(_abc_4268_new_n676_), .B(bus_cap_28_), .Y(_abc_4268_new_n931_));
OR2X2 OR2X2_175 ( .A(_abc_4268_new_n932_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n933_));
OR2X2 OR2X2_176 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n934_), .Y(_abc_4268_new_n935_));
OR2X2 OR2X2_177 ( .A(_abc_4268_new_n701_), .B(bus_cap_30_), .Y(_abc_4268_new_n938_));
OR2X2 OR2X2_178 ( .A(_abc_4268_new_n676_), .B(bus_cap_29_), .Y(_abc_4268_new_n939_));
OR2X2 OR2X2_179 ( .A(_abc_4268_new_n940_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n941_));
OR2X2 OR2X2_18 ( .A(_abc_4268_new_n604_), .B(_abc_4268_new_n608_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_0_));
OR2X2 OR2X2_180 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n942_), .Y(_abc_4268_new_n943_));
OR2X2 OR2X2_181 ( .A(_abc_4268_new_n701_), .B(DOUT), .Y(_abc_4268_new_n946_));
OR2X2 OR2X2_182 ( .A(_abc_4268_new_n676_), .B(bus_cap_30_), .Y(_abc_4268_new_n947_));
OR2X2 OR2X2_183 ( .A(_abc_4268_new_n948_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n949_));
OR2X2 OR2X2_184 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n950_), .Y(_abc_4268_new_n951_));
OR2X2 OR2X2_185 ( .A(_abc_4268_new_n956_), .B(_abc_4268_new_n954_), .Y(_abc_4268_new_n957_));
OR2X2 OR2X2_186 ( .A(_abc_4268_new_n960_), .B(_abc_4268_new_n959_), .Y(_abc_4268_new_n961_));
OR2X2 OR2X2_187 ( .A(_abc_4268_new_n964_), .B(_abc_4268_new_n963_), .Y(_abc_4268_new_n965_));
OR2X2 OR2X2_188 ( .A(_abc_4268_new_n968_), .B(_abc_4268_new_n967_), .Y(_abc_4268_new_n969_));
OR2X2 OR2X2_189 ( .A(_abc_4268_new_n972_), .B(_abc_4268_new_n971_), .Y(_abc_4268_new_n973_));
OR2X2 OR2X2_19 ( .A(_abc_4268_new_n612_), .B(_abc_4268_new_n611_), .Y(_abc_4268_new_n613_));
OR2X2 OR2X2_190 ( .A(_abc_4268_new_n976_), .B(_abc_4268_new_n975_), .Y(_abc_4268_new_n977_));
OR2X2 OR2X2_191 ( .A(_abc_4268_new_n980_), .B(_abc_4268_new_n979_), .Y(_abc_4268_new_n981_));
OR2X2 OR2X2_192 ( .A(_abc_4268_new_n984_), .B(_abc_4268_new_n983_), .Y(_abc_4268_new_n985_));
OR2X2 OR2X2_193 ( .A(_abc_4268_new_n988_), .B(_abc_4268_new_n987_), .Y(_abc_4268_new_n989_));
OR2X2 OR2X2_194 ( .A(_abc_4268_new_n992_), .B(_abc_4268_new_n991_), .Y(_abc_4268_new_n993_));
OR2X2 OR2X2_195 ( .A(_abc_4268_new_n996_), .B(_abc_4268_new_n995_), .Y(_abc_4268_new_n997_));
OR2X2 OR2X2_196 ( .A(_abc_4268_new_n1000_), .B(_abc_4268_new_n999_), .Y(_abc_4268_new_n1001_));
OR2X2 OR2X2_197 ( .A(_abc_4268_new_n1004_), .B(_abc_4268_new_n1003_), .Y(_abc_4268_new_n1005_));
OR2X2 OR2X2_198 ( .A(_abc_4268_new_n1008_), .B(_abc_4268_new_n1007_), .Y(_abc_4268_new_n1009_));
OR2X2 OR2X2_199 ( .A(_abc_4268_new_n1012_), .B(_abc_4268_new_n1011_), .Y(_abc_4268_new_n1013_));
OR2X2 OR2X2_2 ( .A(state_3_), .B(axi_bready), .Y(_abc_4268_new_n564_));
OR2X2 OR2X2_20 ( .A(we), .B(DATA), .Y(_abc_4268_new_n619_));
OR2X2 OR2X2_200 ( .A(_abc_4268_new_n1016_), .B(_abc_4268_new_n1015_), .Y(_abc_4268_new_n1017_));
OR2X2 OR2X2_201 ( .A(_abc_4268_new_n1020_), .B(_abc_4268_new_n1019_), .Y(_abc_4268_new_n1021_));
OR2X2 OR2X2_202 ( .A(_abc_4268_new_n1024_), .B(_abc_4268_new_n1023_), .Y(_abc_4268_new_n1025_));
OR2X2 OR2X2_203 ( .A(_abc_4268_new_n1028_), .B(_abc_4268_new_n1027_), .Y(_abc_4268_new_n1029_));
OR2X2 OR2X2_204 ( .A(_abc_4268_new_n1032_), .B(_abc_4268_new_n1031_), .Y(_abc_4268_new_n1033_));
OR2X2 OR2X2_205 ( .A(_abc_4268_new_n1036_), .B(_abc_4268_new_n1035_), .Y(_abc_4268_new_n1037_));
OR2X2 OR2X2_206 ( .A(_abc_4268_new_n1040_), .B(_abc_4268_new_n1039_), .Y(_abc_4268_new_n1041_));
OR2X2 OR2X2_207 ( .A(_abc_4268_new_n1044_), .B(_abc_4268_new_n1043_), .Y(_abc_4268_new_n1045_));
OR2X2 OR2X2_208 ( .A(_abc_4268_new_n1048_), .B(_abc_4268_new_n1047_), .Y(_abc_4268_new_n1049_));
OR2X2 OR2X2_209 ( .A(_abc_4268_new_n1052_), .B(_abc_4268_new_n1051_), .Y(_abc_4268_new_n1053_));
OR2X2 OR2X2_21 ( .A(_abc_4268_new_n619_), .B(_abc_4268_new_n618_), .Y(_abc_4268_new_n620_));
OR2X2 OR2X2_210 ( .A(_abc_4268_new_n1056_), .B(_abc_4268_new_n1055_), .Y(_abc_4268_new_n1057_));
OR2X2 OR2X2_211 ( .A(_abc_4268_new_n1060_), .B(_abc_4268_new_n1059_), .Y(_abc_4268_new_n1061_));
OR2X2 OR2X2_212 ( .A(_abc_4268_new_n1064_), .B(_abc_4268_new_n1063_), .Y(_abc_4268_new_n1065_));
OR2X2 OR2X2_213 ( .A(_abc_4268_new_n1068_), .B(_abc_4268_new_n1067_), .Y(_abc_4268_new_n1069_));
OR2X2 OR2X2_214 ( .A(_abc_4268_new_n1072_), .B(_abc_4268_new_n1071_), .Y(_abc_4268_new_n1073_));
OR2X2 OR2X2_215 ( .A(_abc_4268_new_n1076_), .B(_abc_4268_new_n1075_), .Y(_abc_4268_new_n1077_));
OR2X2 OR2X2_216 ( .A(_abc_4268_new_n1080_), .B(_abc_4268_new_n1079_), .Y(_abc_4268_new_n1081_));
OR2X2 OR2X2_217 ( .A(_abc_4268_new_n1088_), .B(_abc_4268_new_n1086_), .Y(_abc_4268_new_n1089_));
OR2X2 OR2X2_218 ( .A(_abc_4268_new_n1092_), .B(_abc_4268_new_n1091_), .Y(_abc_4268_new_n1093_));
OR2X2 OR2X2_219 ( .A(_abc_4268_new_n1096_), .B(_abc_4268_new_n1095_), .Y(_abc_4268_new_n1097_));
OR2X2 OR2X2_22 ( .A(re), .B(we), .Y(_abc_4268_new_n624_));
OR2X2 OR2X2_220 ( .A(_abc_4268_new_n1100_), .B(_abc_4268_new_n1099_), .Y(_abc_4268_new_n1101_));
OR2X2 OR2X2_221 ( .A(_abc_4268_new_n1104_), .B(_abc_4268_new_n1103_), .Y(_abc_4268_new_n1105_));
OR2X2 OR2X2_222 ( .A(_abc_4268_new_n1108_), .B(_abc_4268_new_n1107_), .Y(_abc_4268_new_n1109_));
OR2X2 OR2X2_223 ( .A(_abc_4268_new_n1112_), .B(_abc_4268_new_n1111_), .Y(_abc_4268_new_n1113_));
OR2X2 OR2X2_224 ( .A(_abc_4268_new_n1116_), .B(_abc_4268_new_n1115_), .Y(_abc_4268_new_n1117_));
OR2X2 OR2X2_225 ( .A(_abc_4268_new_n1120_), .B(_abc_4268_new_n1119_), .Y(_abc_4268_new_n1121_));
OR2X2 OR2X2_226 ( .A(_abc_4268_new_n1124_), .B(_abc_4268_new_n1123_), .Y(_abc_4268_new_n1125_));
OR2X2 OR2X2_227 ( .A(_abc_4268_new_n1128_), .B(_abc_4268_new_n1127_), .Y(_abc_4268_new_n1129_));
OR2X2 OR2X2_228 ( .A(_abc_4268_new_n1132_), .B(_abc_4268_new_n1131_), .Y(_abc_4268_new_n1133_));
OR2X2 OR2X2_229 ( .A(_abc_4268_new_n1136_), .B(_abc_4268_new_n1135_), .Y(_abc_4268_new_n1137_));
OR2X2 OR2X2_23 ( .A(_abc_4268_new_n625_), .B(_abc_4268_new_n623_), .Y(_abc_4268_new_n626_));
OR2X2 OR2X2_230 ( .A(_abc_4268_new_n1140_), .B(_abc_4268_new_n1139_), .Y(_abc_4268_new_n1141_));
OR2X2 OR2X2_231 ( .A(_abc_4268_new_n1144_), .B(_abc_4268_new_n1143_), .Y(_abc_4268_new_n1145_));
OR2X2 OR2X2_232 ( .A(_abc_4268_new_n1148_), .B(_abc_4268_new_n1147_), .Y(_abc_4268_new_n1149_));
OR2X2 OR2X2_233 ( .A(_abc_4268_new_n1152_), .B(_abc_4268_new_n1151_), .Y(_abc_4268_new_n1153_));
OR2X2 OR2X2_234 ( .A(_abc_4268_new_n1156_), .B(_abc_4268_new_n1155_), .Y(_abc_4268_new_n1157_));
OR2X2 OR2X2_235 ( .A(_abc_4268_new_n1160_), .B(_abc_4268_new_n1159_), .Y(_abc_4268_new_n1161_));
OR2X2 OR2X2_236 ( .A(_abc_4268_new_n1164_), .B(_abc_4268_new_n1163_), .Y(_abc_4268_new_n1165_));
OR2X2 OR2X2_237 ( .A(_abc_4268_new_n1168_), .B(_abc_4268_new_n1167_), .Y(_abc_4268_new_n1169_));
OR2X2 OR2X2_238 ( .A(_abc_4268_new_n1172_), .B(_abc_4268_new_n1171_), .Y(_abc_4268_new_n1173_));
OR2X2 OR2X2_239 ( .A(_abc_4268_new_n1176_), .B(_abc_4268_new_n1175_), .Y(_abc_4268_new_n1177_));
OR2X2 OR2X2_24 ( .A(counter_16_), .B(counter_17_), .Y(_abc_4268_new_n628_));
OR2X2 OR2X2_240 ( .A(_abc_4268_new_n1180_), .B(_abc_4268_new_n1179_), .Y(_abc_4268_new_n1181_));
OR2X2 OR2X2_241 ( .A(_abc_4268_new_n1184_), .B(_abc_4268_new_n1183_), .Y(_abc_4268_new_n1185_));
OR2X2 OR2X2_242 ( .A(_abc_4268_new_n1188_), .B(_abc_4268_new_n1187_), .Y(_abc_4268_new_n1189_));
OR2X2 OR2X2_243 ( .A(_abc_4268_new_n1192_), .B(_abc_4268_new_n1191_), .Y(_abc_4268_new_n1193_));
OR2X2 OR2X2_244 ( .A(_abc_4268_new_n1196_), .B(_abc_4268_new_n1195_), .Y(_abc_4268_new_n1197_));
OR2X2 OR2X2_245 ( .A(_abc_4268_new_n1200_), .B(_abc_4268_new_n1199_), .Y(_abc_4268_new_n1201_));
OR2X2 OR2X2_246 ( .A(_abc_4268_new_n1204_), .B(_abc_4268_new_n1203_), .Y(_abc_4268_new_n1205_));
OR2X2 OR2X2_247 ( .A(_abc_4268_new_n1208_), .B(_abc_4268_new_n1207_), .Y(_abc_4268_new_n1209_));
OR2X2 OR2X2_248 ( .A(_abc_4268_new_n1212_), .B(_abc_4268_new_n1211_), .Y(_abc_4268_new_n1213_));
OR2X2 OR2X2_249 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_0_), .Y(_abc_4268_new_n1217_));
OR2X2 OR2X2_25 ( .A(counter_14_), .B(counter_15_), .Y(_abc_4268_new_n630_));
OR2X2 OR2X2_250 ( .A(_abc_4268_new_n1218_), .B(DATA), .Y(_abc_4268_new_n1219_));
OR2X2 OR2X2_251 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_1_), .Y(_abc_4268_new_n1222_));
OR2X2 OR2X2_252 ( .A(_abc_4268_new_n1218_), .B(sft_reg_0_), .Y(_abc_4268_new_n1223_));
OR2X2 OR2X2_253 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_2_), .Y(_abc_4268_new_n1226_));
OR2X2 OR2X2_254 ( .A(_abc_4268_new_n1218_), .B(sft_reg_1_), .Y(_abc_4268_new_n1227_));
OR2X2 OR2X2_255 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_3_), .Y(_abc_4268_new_n1230_));
OR2X2 OR2X2_256 ( .A(_abc_4268_new_n1218_), .B(sft_reg_2_), .Y(_abc_4268_new_n1231_));
OR2X2 OR2X2_257 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_4_), .Y(_abc_4268_new_n1234_));
OR2X2 OR2X2_258 ( .A(_abc_4268_new_n1218_), .B(sft_reg_3_), .Y(_abc_4268_new_n1235_));
OR2X2 OR2X2_259 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_5_), .Y(_abc_4268_new_n1238_));
OR2X2 OR2X2_26 ( .A(counter_12_), .B(counter_13_), .Y(_abc_4268_new_n633_));
OR2X2 OR2X2_260 ( .A(_abc_4268_new_n1218_), .B(sft_reg_4_), .Y(_abc_4268_new_n1239_));
OR2X2 OR2X2_261 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_6_), .Y(_abc_4268_new_n1242_));
OR2X2 OR2X2_262 ( .A(_abc_4268_new_n1218_), .B(sft_reg_5_), .Y(_abc_4268_new_n1243_));
OR2X2 OR2X2_263 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_7_), .Y(_abc_4268_new_n1246_));
OR2X2 OR2X2_264 ( .A(_abc_4268_new_n1218_), .B(sft_reg_6_), .Y(_abc_4268_new_n1247_));
OR2X2 OR2X2_265 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_8_), .Y(_abc_4268_new_n1250_));
OR2X2 OR2X2_266 ( .A(_abc_4268_new_n1218_), .B(sft_reg_7_), .Y(_abc_4268_new_n1251_));
OR2X2 OR2X2_267 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_9_), .Y(_abc_4268_new_n1254_));
OR2X2 OR2X2_268 ( .A(_abc_4268_new_n1218_), .B(sft_reg_8_), .Y(_abc_4268_new_n1255_));
OR2X2 OR2X2_269 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_10_), .Y(_abc_4268_new_n1258_));
OR2X2 OR2X2_27 ( .A(counter_10_), .B(counter_11_), .Y(_abc_4268_new_n635_));
OR2X2 OR2X2_270 ( .A(_abc_4268_new_n1218_), .B(sft_reg_9_), .Y(_abc_4268_new_n1259_));
OR2X2 OR2X2_271 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_11_), .Y(_abc_4268_new_n1262_));
OR2X2 OR2X2_272 ( .A(_abc_4268_new_n1218_), .B(sft_reg_10_), .Y(_abc_4268_new_n1263_));
OR2X2 OR2X2_273 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_12_), .Y(_abc_4268_new_n1266_));
OR2X2 OR2X2_274 ( .A(_abc_4268_new_n1218_), .B(sft_reg_11_), .Y(_abc_4268_new_n1267_));
OR2X2 OR2X2_275 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_13_), .Y(_abc_4268_new_n1270_));
OR2X2 OR2X2_276 ( .A(_abc_4268_new_n1218_), .B(sft_reg_12_), .Y(_abc_4268_new_n1271_));
OR2X2 OR2X2_277 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_14_), .Y(_abc_4268_new_n1274_));
OR2X2 OR2X2_278 ( .A(_abc_4268_new_n1218_), .B(sft_reg_13_), .Y(_abc_4268_new_n1275_));
OR2X2 OR2X2_279 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_15_), .Y(_abc_4268_new_n1278_));
OR2X2 OR2X2_28 ( .A(counter_4_), .B(counter_5_), .Y(_abc_4268_new_n639_));
OR2X2 OR2X2_280 ( .A(_abc_4268_new_n1218_), .B(sft_reg_14_), .Y(_abc_4268_new_n1279_));
OR2X2 OR2X2_281 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_16_), .Y(_abc_4268_new_n1282_));
OR2X2 OR2X2_282 ( .A(_abc_4268_new_n1218_), .B(sft_reg_15_), .Y(_abc_4268_new_n1283_));
OR2X2 OR2X2_283 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_17_), .Y(_abc_4268_new_n1286_));
OR2X2 OR2X2_284 ( .A(_abc_4268_new_n1218_), .B(sft_reg_16_), .Y(_abc_4268_new_n1287_));
OR2X2 OR2X2_285 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_18_), .Y(_abc_4268_new_n1290_));
OR2X2 OR2X2_286 ( .A(_abc_4268_new_n1218_), .B(sft_reg_17_), .Y(_abc_4268_new_n1291_));
OR2X2 OR2X2_287 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_19_), .Y(_abc_4268_new_n1294_));
OR2X2 OR2X2_288 ( .A(_abc_4268_new_n1218_), .B(sft_reg_18_), .Y(_abc_4268_new_n1295_));
OR2X2 OR2X2_289 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_20_), .Y(_abc_4268_new_n1298_));
OR2X2 OR2X2_29 ( .A(counter_2_), .B(counter_3_), .Y(_abc_4268_new_n641_));
OR2X2 OR2X2_290 ( .A(_abc_4268_new_n1218_), .B(sft_reg_19_), .Y(_abc_4268_new_n1299_));
OR2X2 OR2X2_291 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_21_), .Y(_abc_4268_new_n1302_));
OR2X2 OR2X2_292 ( .A(_abc_4268_new_n1218_), .B(sft_reg_20_), .Y(_abc_4268_new_n1303_));
OR2X2 OR2X2_293 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_22_), .Y(_abc_4268_new_n1306_));
OR2X2 OR2X2_294 ( .A(_abc_4268_new_n1218_), .B(sft_reg_21_), .Y(_abc_4268_new_n1307_));
OR2X2 OR2X2_295 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_23_), .Y(_abc_4268_new_n1310_));
OR2X2 OR2X2_296 ( .A(_abc_4268_new_n1218_), .B(sft_reg_22_), .Y(_abc_4268_new_n1311_));
OR2X2 OR2X2_297 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_24_), .Y(_abc_4268_new_n1314_));
OR2X2 OR2X2_298 ( .A(_abc_4268_new_n1218_), .B(sft_reg_23_), .Y(_abc_4268_new_n1315_));
OR2X2 OR2X2_299 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_25_), .Y(_abc_4268_new_n1318_));
OR2X2 OR2X2_3 ( .A(_abc_4268_new_n564_), .B(state_7_), .Y(axi_wvalid));
OR2X2 OR2X2_30 ( .A(counter_8_), .B(counter_9_), .Y(_abc_4268_new_n644_));
OR2X2 OR2X2_300 ( .A(_abc_4268_new_n1218_), .B(sft_reg_24_), .Y(_abc_4268_new_n1319_));
OR2X2 OR2X2_301 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_26_), .Y(_abc_4268_new_n1322_));
OR2X2 OR2X2_302 ( .A(_abc_4268_new_n1218_), .B(sft_reg_25_), .Y(_abc_4268_new_n1323_));
OR2X2 OR2X2_303 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_27_), .Y(_abc_4268_new_n1326_));
OR2X2 OR2X2_304 ( .A(_abc_4268_new_n1218_), .B(sft_reg_26_), .Y(_abc_4268_new_n1327_));
OR2X2 OR2X2_305 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_28_), .Y(_abc_4268_new_n1330_));
OR2X2 OR2X2_306 ( .A(_abc_4268_new_n1218_), .B(sft_reg_27_), .Y(_abc_4268_new_n1331_));
OR2X2 OR2X2_307 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_29_), .Y(_abc_4268_new_n1334_));
OR2X2 OR2X2_308 ( .A(_abc_4268_new_n1218_), .B(sft_reg_28_), .Y(_abc_4268_new_n1335_));
OR2X2 OR2X2_309 ( .A(_abc_4268_new_n1216_), .B(A_ADDR_30_), .Y(_abc_4268_new_n1338_));
OR2X2 OR2X2_31 ( .A(counter_6_), .B(counter_7_), .Y(_abc_4268_new_n646_));
OR2X2 OR2X2_310 ( .A(_abc_4268_new_n1218_), .B(sft_reg_29_), .Y(_abc_4268_new_n1339_));
OR2X2 OR2X2_311 ( .A(_abc_4268_new_n1343_), .B(_abc_4268_new_n1342_), .Y(_abc_4268_new_n1344_));
OR2X2 OR2X2_312 ( .A(_abc_4268_new_n1083_), .B(sft_reg_0_), .Y(_abc_4268_new_n1346_));
OR2X2 OR2X2_313 ( .A(DATA), .B(CEB), .Y(_abc_4268_new_n1347_));
OR2X2 OR2X2_314 ( .A(_abc_4268_new_n1083_), .B(sft_reg_1_), .Y(_abc_4268_new_n1350_));
OR2X2 OR2X2_315 ( .A(CEB), .B(sft_reg_0_), .Y(_abc_4268_new_n1351_));
OR2X2 OR2X2_316 ( .A(_abc_4268_new_n1083_), .B(sft_reg_2_), .Y(_abc_4268_new_n1354_));
OR2X2 OR2X2_317 ( .A(CEB), .B(sft_reg_1_), .Y(_abc_4268_new_n1355_));
OR2X2 OR2X2_318 ( .A(_abc_4268_new_n1083_), .B(sft_reg_3_), .Y(_abc_4268_new_n1358_));
OR2X2 OR2X2_319 ( .A(CEB), .B(sft_reg_2_), .Y(_abc_4268_new_n1359_));
OR2X2 OR2X2_32 ( .A(counter_28_), .B(counter_29_), .Y(_abc_4268_new_n651_));
OR2X2 OR2X2_320 ( .A(_abc_4268_new_n1083_), .B(sft_reg_4_), .Y(_abc_4268_new_n1362_));
OR2X2 OR2X2_321 ( .A(CEB), .B(sft_reg_3_), .Y(_abc_4268_new_n1363_));
OR2X2 OR2X2_322 ( .A(_abc_4268_new_n1083_), .B(sft_reg_5_), .Y(_abc_4268_new_n1366_));
OR2X2 OR2X2_323 ( .A(CEB), .B(sft_reg_4_), .Y(_abc_4268_new_n1367_));
OR2X2 OR2X2_324 ( .A(_abc_4268_new_n1083_), .B(sft_reg_6_), .Y(_abc_4268_new_n1370_));
OR2X2 OR2X2_325 ( .A(CEB), .B(sft_reg_5_), .Y(_abc_4268_new_n1371_));
OR2X2 OR2X2_326 ( .A(_abc_4268_new_n1083_), .B(sft_reg_7_), .Y(_abc_4268_new_n1374_));
OR2X2 OR2X2_327 ( .A(CEB), .B(sft_reg_6_), .Y(_abc_4268_new_n1375_));
OR2X2 OR2X2_328 ( .A(_abc_4268_new_n1083_), .B(sft_reg_8_), .Y(_abc_4268_new_n1378_));
OR2X2 OR2X2_329 ( .A(CEB), .B(sft_reg_7_), .Y(_abc_4268_new_n1379_));
OR2X2 OR2X2_33 ( .A(counter_26_), .B(counter_27_), .Y(_abc_4268_new_n653_));
OR2X2 OR2X2_330 ( .A(_abc_4268_new_n1083_), .B(sft_reg_9_), .Y(_abc_4268_new_n1382_));
OR2X2 OR2X2_331 ( .A(CEB), .B(sft_reg_8_), .Y(_abc_4268_new_n1383_));
OR2X2 OR2X2_332 ( .A(_abc_4268_new_n1083_), .B(sft_reg_10_), .Y(_abc_4268_new_n1386_));
OR2X2 OR2X2_333 ( .A(CEB), .B(sft_reg_9_), .Y(_abc_4268_new_n1387_));
OR2X2 OR2X2_334 ( .A(_abc_4268_new_n1083_), .B(sft_reg_11_), .Y(_abc_4268_new_n1390_));
OR2X2 OR2X2_335 ( .A(CEB), .B(sft_reg_10_), .Y(_abc_4268_new_n1391_));
OR2X2 OR2X2_336 ( .A(_abc_4268_new_n1083_), .B(sft_reg_12_), .Y(_abc_4268_new_n1394_));
OR2X2 OR2X2_337 ( .A(CEB), .B(sft_reg_11_), .Y(_abc_4268_new_n1395_));
OR2X2 OR2X2_338 ( .A(_abc_4268_new_n1083_), .B(sft_reg_13_), .Y(_abc_4268_new_n1398_));
OR2X2 OR2X2_339 ( .A(CEB), .B(sft_reg_12_), .Y(_abc_4268_new_n1399_));
OR2X2 OR2X2_34 ( .A(counter_32_), .B(counter_33_), .Y(_abc_4268_new_n656_));
OR2X2 OR2X2_340 ( .A(_abc_4268_new_n1083_), .B(sft_reg_14_), .Y(_abc_4268_new_n1402_));
OR2X2 OR2X2_341 ( .A(CEB), .B(sft_reg_13_), .Y(_abc_4268_new_n1403_));
OR2X2 OR2X2_342 ( .A(_abc_4268_new_n1083_), .B(sft_reg_15_), .Y(_abc_4268_new_n1406_));
OR2X2 OR2X2_343 ( .A(CEB), .B(sft_reg_14_), .Y(_abc_4268_new_n1407_));
OR2X2 OR2X2_344 ( .A(_abc_4268_new_n1083_), .B(sft_reg_16_), .Y(_abc_4268_new_n1410_));
OR2X2 OR2X2_345 ( .A(CEB), .B(sft_reg_15_), .Y(_abc_4268_new_n1411_));
OR2X2 OR2X2_346 ( .A(_abc_4268_new_n1083_), .B(sft_reg_17_), .Y(_abc_4268_new_n1414_));
OR2X2 OR2X2_347 ( .A(CEB), .B(sft_reg_16_), .Y(_abc_4268_new_n1415_));
OR2X2 OR2X2_348 ( .A(_abc_4268_new_n1083_), .B(sft_reg_18_), .Y(_abc_4268_new_n1418_));
OR2X2 OR2X2_349 ( .A(CEB), .B(sft_reg_17_), .Y(_abc_4268_new_n1419_));
OR2X2 OR2X2_35 ( .A(counter_30_), .B(counter_31_), .Y(_abc_4268_new_n658_));
OR2X2 OR2X2_350 ( .A(_abc_4268_new_n1083_), .B(sft_reg_19_), .Y(_abc_4268_new_n1422_));
OR2X2 OR2X2_351 ( .A(CEB), .B(sft_reg_18_), .Y(_abc_4268_new_n1423_));
OR2X2 OR2X2_352 ( .A(_abc_4268_new_n1083_), .B(sft_reg_20_), .Y(_abc_4268_new_n1426_));
OR2X2 OR2X2_353 ( .A(CEB), .B(sft_reg_19_), .Y(_abc_4268_new_n1427_));
OR2X2 OR2X2_354 ( .A(_abc_4268_new_n1083_), .B(sft_reg_21_), .Y(_abc_4268_new_n1430_));
OR2X2 OR2X2_355 ( .A(CEB), .B(sft_reg_20_), .Y(_abc_4268_new_n1431_));
OR2X2 OR2X2_356 ( .A(_abc_4268_new_n1083_), .B(sft_reg_22_), .Y(_abc_4268_new_n1434_));
OR2X2 OR2X2_357 ( .A(CEB), .B(sft_reg_21_), .Y(_abc_4268_new_n1435_));
OR2X2 OR2X2_358 ( .A(_abc_4268_new_n1083_), .B(sft_reg_23_), .Y(_abc_4268_new_n1438_));
OR2X2 OR2X2_359 ( .A(CEB), .B(sft_reg_22_), .Y(_abc_4268_new_n1439_));
OR2X2 OR2X2_36 ( .A(counter_24_), .B(counter_25_), .Y(_abc_4268_new_n662_));
OR2X2 OR2X2_360 ( .A(_abc_4268_new_n1083_), .B(sft_reg_24_), .Y(_abc_4268_new_n1442_));
OR2X2 OR2X2_361 ( .A(CEB), .B(sft_reg_23_), .Y(_abc_4268_new_n1443_));
OR2X2 OR2X2_362 ( .A(_abc_4268_new_n1083_), .B(sft_reg_25_), .Y(_abc_4268_new_n1446_));
OR2X2 OR2X2_363 ( .A(CEB), .B(sft_reg_24_), .Y(_abc_4268_new_n1447_));
OR2X2 OR2X2_364 ( .A(_abc_4268_new_n1083_), .B(sft_reg_26_), .Y(_abc_4268_new_n1450_));
OR2X2 OR2X2_365 ( .A(CEB), .B(sft_reg_25_), .Y(_abc_4268_new_n1451_));
OR2X2 OR2X2_366 ( .A(_abc_4268_new_n1083_), .B(sft_reg_27_), .Y(_abc_4268_new_n1454_));
OR2X2 OR2X2_367 ( .A(CEB), .B(sft_reg_26_), .Y(_abc_4268_new_n1455_));
OR2X2 OR2X2_368 ( .A(_abc_4268_new_n1083_), .B(sft_reg_28_), .Y(_abc_4268_new_n1458_));
OR2X2 OR2X2_369 ( .A(CEB), .B(sft_reg_27_), .Y(_abc_4268_new_n1459_));
OR2X2 OR2X2_37 ( .A(counter_22_), .B(counter_23_), .Y(_abc_4268_new_n664_));
OR2X2 OR2X2_370 ( .A(_abc_4268_new_n1083_), .B(sft_reg_29_), .Y(_abc_4268_new_n1462_));
OR2X2 OR2X2_371 ( .A(CEB), .B(sft_reg_28_), .Y(_abc_4268_new_n1463_));
OR2X2 OR2X2_372 ( .A(_abc_4268_new_n1083_), .B(sft_reg_30_), .Y(_abc_4268_new_n1466_));
OR2X2 OR2X2_373 ( .A(CEB), .B(sft_reg_29_), .Y(_abc_4268_new_n1467_));
OR2X2 OR2X2_374 ( .A(_abc_4268_new_n1538_), .B(DATA), .Y(_abc_4268_new_n1539_));
OR2X2 OR2X2_375 ( .A(_abc_4268_new_n1537_), .B(PICORV_RST_SPI), .Y(_abc_4268_new_n1540_));
OR2X2 OR2X2_376 ( .A(_abc_4268_new_n1347_), .B(_abc_4268_new_n618_), .Y(_abc_4268_new_n1543_));
OR2X2 OR2X2_377 ( .A(_0counter_65_0__2_), .B(_abc_4268_new_n1544_), .Y(_abc_4268_new_n1545_));
OR2X2 OR2X2_378 ( .A(_abc_4268_new_n1347_), .B(_abc_4268_new_n1547_), .Y(_abc_4268_new_n1548_));
OR2X2 OR2X2_379 ( .A(_0counter_65_0__1_), .B(_abc_4268_new_n1549_), .Y(_abc_4268_new_n1550_));
OR2X2 OR2X2_38 ( .A(counter_20_), .B(counter_21_), .Y(_abc_4268_new_n667_));
OR2X2 OR2X2_380 ( .A(bus_sync_axi_bus__abc_3879_new_n394_), .B(bus_sync_axi_bus__abc_3879_new_n395_), .Y(bus_sync_axi_bus__abc_3879_new_n396_));
OR2X2 OR2X2_381 ( .A(bus_sync_axi_bus__abc_3879_new_n398_), .B(bus_sync_axi_bus__abc_3879_new_n399_), .Y(bus_sync_axi_bus__abc_3879_new_n400_));
OR2X2 OR2X2_382 ( .A(bus_sync_axi_bus__abc_3879_new_n402_), .B(bus_sync_axi_bus__abc_3879_new_n403_), .Y(bus_sync_axi_bus__abc_3879_new_n404_));
OR2X2 OR2X2_383 ( .A(bus_sync_axi_bus__abc_3879_new_n406_), .B(bus_sync_axi_bus__abc_3879_new_n407_), .Y(bus_sync_axi_bus__abc_3879_new_n408_));
OR2X2 OR2X2_384 ( .A(bus_sync_axi_bus__abc_3879_new_n410_), .B(bus_sync_axi_bus__abc_3879_new_n411_), .Y(bus_sync_axi_bus__abc_3879_new_n412_));
OR2X2 OR2X2_385 ( .A(bus_sync_axi_bus__abc_3879_new_n414_), .B(bus_sync_axi_bus__abc_3879_new_n415_), .Y(bus_sync_axi_bus__abc_3879_new_n416_));
OR2X2 OR2X2_386 ( .A(bus_sync_axi_bus__abc_3879_new_n418_), .B(bus_sync_axi_bus__abc_3879_new_n419_), .Y(bus_sync_axi_bus__abc_3879_new_n420_));
OR2X2 OR2X2_387 ( .A(bus_sync_axi_bus__abc_3879_new_n422_), .B(bus_sync_axi_bus__abc_3879_new_n423_), .Y(bus_sync_axi_bus__abc_3879_new_n424_));
OR2X2 OR2X2_388 ( .A(bus_sync_axi_bus__abc_3879_new_n426_), .B(bus_sync_axi_bus__abc_3879_new_n427_), .Y(bus_sync_axi_bus__abc_3879_new_n428_));
OR2X2 OR2X2_389 ( .A(bus_sync_axi_bus__abc_3879_new_n430_), .B(bus_sync_axi_bus__abc_3879_new_n431_), .Y(bus_sync_axi_bus__abc_3879_new_n432_));
OR2X2 OR2X2_39 ( .A(_abc_4268_new_n675_), .B(_abc_4268_new_n627_), .Y(_abc_4268_new_n676_));
OR2X2 OR2X2_390 ( .A(bus_sync_axi_bus__abc_3879_new_n434_), .B(bus_sync_axi_bus__abc_3879_new_n435_), .Y(bus_sync_axi_bus__abc_3879_new_n436_));
OR2X2 OR2X2_391 ( .A(bus_sync_axi_bus__abc_3879_new_n438_), .B(bus_sync_axi_bus__abc_3879_new_n439_), .Y(bus_sync_axi_bus__abc_3879_new_n440_));
OR2X2 OR2X2_392 ( .A(bus_sync_axi_bus__abc_3879_new_n442_), .B(bus_sync_axi_bus__abc_3879_new_n443_), .Y(bus_sync_axi_bus__abc_3879_new_n444_));
OR2X2 OR2X2_393 ( .A(bus_sync_axi_bus__abc_3879_new_n446_), .B(bus_sync_axi_bus__abc_3879_new_n447_), .Y(bus_sync_axi_bus__abc_3879_new_n448_));
OR2X2 OR2X2_394 ( .A(bus_sync_axi_bus__abc_3879_new_n450_), .B(bus_sync_axi_bus__abc_3879_new_n451_), .Y(bus_sync_axi_bus__abc_3879_new_n452_));
OR2X2 OR2X2_395 ( .A(bus_sync_axi_bus__abc_3879_new_n454_), .B(bus_sync_axi_bus__abc_3879_new_n455_), .Y(bus_sync_axi_bus__abc_3879_new_n456_));
OR2X2 OR2X2_396 ( .A(bus_sync_axi_bus__abc_3879_new_n458_), .B(bus_sync_axi_bus__abc_3879_new_n459_), .Y(bus_sync_axi_bus__abc_3879_new_n460_));
OR2X2 OR2X2_397 ( .A(bus_sync_axi_bus__abc_3879_new_n462_), .B(bus_sync_axi_bus__abc_3879_new_n463_), .Y(bus_sync_axi_bus__abc_3879_new_n464_));
OR2X2 OR2X2_398 ( .A(bus_sync_axi_bus__abc_3879_new_n466_), .B(bus_sync_axi_bus__abc_3879_new_n467_), .Y(bus_sync_axi_bus__abc_3879_new_n468_));
OR2X2 OR2X2_399 ( .A(bus_sync_axi_bus__abc_3879_new_n470_), .B(bus_sync_axi_bus__abc_3879_new_n471_), .Y(bus_sync_axi_bus__abc_3879_new_n472_));
OR2X2 OR2X2_4 ( .A(_abc_4268_new_n567_), .B(_abc_4268_new_n568_), .Y(_abc_4268_new_n569_));
OR2X2 OR2X2_40 ( .A(_abc_4268_new_n677_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n678_));
OR2X2 OR2X2_400 ( .A(bus_sync_axi_bus__abc_3879_new_n474_), .B(bus_sync_axi_bus__abc_3879_new_n475_), .Y(bus_sync_axi_bus__abc_3879_new_n476_));
OR2X2 OR2X2_401 ( .A(bus_sync_axi_bus__abc_3879_new_n478_), .B(bus_sync_axi_bus__abc_3879_new_n479_), .Y(bus_sync_axi_bus__abc_3879_new_n480_));
OR2X2 OR2X2_402 ( .A(bus_sync_axi_bus__abc_3879_new_n482_), .B(bus_sync_axi_bus__abc_3879_new_n483_), .Y(bus_sync_axi_bus__abc_3879_new_n484_));
OR2X2 OR2X2_403 ( .A(bus_sync_axi_bus__abc_3879_new_n486_), .B(bus_sync_axi_bus__abc_3879_new_n487_), .Y(bus_sync_axi_bus__abc_3879_new_n488_));
OR2X2 OR2X2_404 ( .A(bus_sync_axi_bus__abc_3879_new_n490_), .B(bus_sync_axi_bus__abc_3879_new_n491_), .Y(bus_sync_axi_bus__abc_3879_new_n492_));
OR2X2 OR2X2_405 ( .A(bus_sync_axi_bus__abc_3879_new_n494_), .B(bus_sync_axi_bus__abc_3879_new_n495_), .Y(bus_sync_axi_bus__abc_3879_new_n496_));
OR2X2 OR2X2_406 ( .A(bus_sync_axi_bus__abc_3879_new_n498_), .B(bus_sync_axi_bus__abc_3879_new_n499_), .Y(bus_sync_axi_bus__abc_3879_new_n500_));
OR2X2 OR2X2_407 ( .A(bus_sync_axi_bus__abc_3879_new_n502_), .B(bus_sync_axi_bus__abc_3879_new_n503_), .Y(bus_sync_axi_bus__abc_3879_new_n504_));
OR2X2 OR2X2_408 ( .A(bus_sync_axi_bus__abc_3879_new_n506_), .B(bus_sync_axi_bus__abc_3879_new_n507_), .Y(bus_sync_axi_bus__abc_3879_new_n508_));
OR2X2 OR2X2_409 ( .A(bus_sync_axi_bus__abc_3879_new_n510_), .B(bus_sync_axi_bus__abc_3879_new_n511_), .Y(bus_sync_axi_bus__abc_3879_new_n512_));
OR2X2 OR2X2_41 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n680_), .Y(_abc_4268_new_n681_));
OR2X2 OR2X2_410 ( .A(bus_sync_axi_bus__abc_3879_new_n514_), .B(bus_sync_axi_bus__abc_3879_new_n515_), .Y(bus_sync_axi_bus__abc_3879_new_n516_));
OR2X2 OR2X2_411 ( .A(bus_sync_axi_bus__abc_3879_new_n518_), .B(bus_sync_axi_bus__abc_3879_new_n519_), .Y(bus_sync_axi_bus__abc_3879_new_n520_));
OR2X2 OR2X2_412 ( .A(bus_sync_axi_bus__abc_3879_new_n522_), .B(bus_sync_axi_bus__abc_3879_new_n523_), .Y(bus_sync_axi_bus__abc_3879_new_n524_));
OR2X2 OR2X2_413 ( .A(bus_sync_axi_bus__abc_3879_new_n526_), .B(bus_sync_axi_bus__abc_3879_new_n527_), .Y(bus_sync_axi_bus__abc_3879_new_n528_));
OR2X2 OR2X2_414 ( .A(bus_sync_axi_bus__abc_3879_new_n530_), .B(bus_sync_axi_bus__abc_3879_new_n531_), .Y(bus_sync_axi_bus__abc_3879_new_n532_));
OR2X2 OR2X2_415 ( .A(bus_sync_axi_bus__abc_3879_new_n534_), .B(bus_sync_axi_bus__abc_3879_new_n535_), .Y(bus_sync_axi_bus__abc_3879_new_n536_));
OR2X2 OR2X2_416 ( .A(bus_sync_axi_bus__abc_3879_new_n538_), .B(bus_sync_axi_bus__abc_3879_new_n539_), .Y(bus_sync_axi_bus__abc_3879_new_n540_));
OR2X2 OR2X2_417 ( .A(bus_sync_axi_bus__abc_3879_new_n542_), .B(bus_sync_axi_bus__abc_3879_new_n543_), .Y(bus_sync_axi_bus__abc_3879_new_n544_));
OR2X2 OR2X2_418 ( .A(bus_sync_axi_bus__abc_3879_new_n546_), .B(bus_sync_axi_bus__abc_3879_new_n547_), .Y(bus_sync_axi_bus__abc_3879_new_n548_));
OR2X2 OR2X2_419 ( .A(bus_sync_axi_bus__abc_3879_new_n550_), .B(bus_sync_axi_bus__abc_3879_new_n551_), .Y(bus_sync_axi_bus__abc_3879_new_n552_));
OR2X2 OR2X2_42 ( .A(_abc_4268_new_n681_), .B(_abc_4268_new_n679_), .Y(_abc_4268_new_n682_));
OR2X2 OR2X2_420 ( .A(bus_sync_axi_bus__abc_3879_new_n554_), .B(bus_sync_axi_bus__abc_3879_new_n555_), .Y(bus_sync_axi_bus__abc_3879_new_n556_));
OR2X2 OR2X2_421 ( .A(bus_sync_axi_bus__abc_3879_new_n558_), .B(bus_sync_axi_bus__abc_3879_new_n559_), .Y(bus_sync_axi_bus__abc_3879_new_n560_));
OR2X2 OR2X2_422 ( .A(bus_sync_axi_bus__abc_3879_new_n562_), .B(bus_sync_axi_bus__abc_3879_new_n563_), .Y(bus_sync_axi_bus__abc_3879_new_n564_));
OR2X2 OR2X2_423 ( .A(bus_sync_axi_bus__abc_3879_new_n566_), .B(bus_sync_axi_bus__abc_3879_new_n567_), .Y(bus_sync_axi_bus__abc_3879_new_n568_));
OR2X2 OR2X2_424 ( .A(bus_sync_axi_bus__abc_3879_new_n570_), .B(bus_sync_axi_bus__abc_3879_new_n571_), .Y(bus_sync_axi_bus__abc_3879_new_n572_));
OR2X2 OR2X2_425 ( .A(bus_sync_axi_bus__abc_3879_new_n574_), .B(bus_sync_axi_bus__abc_3879_new_n575_), .Y(bus_sync_axi_bus__abc_3879_new_n576_));
OR2X2 OR2X2_426 ( .A(bus_sync_axi_bus__abc_3879_new_n578_), .B(bus_sync_axi_bus__abc_3879_new_n579_), .Y(bus_sync_axi_bus__abc_3879_new_n580_));
OR2X2 OR2X2_427 ( .A(bus_sync_axi_bus__abc_3879_new_n582_), .B(bus_sync_axi_bus__abc_3879_new_n583_), .Y(bus_sync_axi_bus__abc_3879_new_n584_));
OR2X2 OR2X2_428 ( .A(bus_sync_axi_bus__abc_3879_new_n586_), .B(bus_sync_axi_bus__abc_3879_new_n587_), .Y(bus_sync_axi_bus__abc_3879_new_n588_));
OR2X2 OR2X2_429 ( .A(bus_sync_axi_bus__abc_3879_new_n590_), .B(bus_sync_axi_bus__abc_3879_new_n591_), .Y(bus_sync_axi_bus__abc_3879_new_n592_));
OR2X2 OR2X2_43 ( .A(_abc_4268_new_n628_), .B(_abc_4268_new_n630_), .Y(_abc_4268_new_n685_));
OR2X2 OR2X2_430 ( .A(bus_sync_axi_bus__abc_3879_new_n594_), .B(bus_sync_axi_bus__abc_3879_new_n595_), .Y(bus_sync_axi_bus__abc_3879_new_n596_));
OR2X2 OR2X2_431 ( .A(bus_sync_axi_bus__abc_3879_new_n598_), .B(bus_sync_axi_bus__abc_3879_new_n599_), .Y(bus_sync_axi_bus__abc_3879_new_n600_));
OR2X2 OR2X2_432 ( .A(bus_sync_axi_bus__abc_3879_new_n602_), .B(bus_sync_axi_bus__abc_3879_new_n603_), .Y(bus_sync_axi_bus__abc_3879_new_n604_));
OR2X2 OR2X2_433 ( .A(bus_sync_axi_bus__abc_3879_new_n606_), .B(bus_sync_axi_bus__abc_3879_new_n607_), .Y(bus_sync_axi_bus__abc_3879_new_n608_));
OR2X2 OR2X2_434 ( .A(bus_sync_axi_bus__abc_3879_new_n610_), .B(bus_sync_axi_bus__abc_3879_new_n611_), .Y(bus_sync_axi_bus__abc_3879_new_n612_));
OR2X2 OR2X2_435 ( .A(bus_sync_axi_bus__abc_3879_new_n614_), .B(bus_sync_axi_bus__abc_3879_new_n615_), .Y(bus_sync_axi_bus__abc_3879_new_n616_));
OR2X2 OR2X2_436 ( .A(bus_sync_axi_bus__abc_3879_new_n618_), .B(bus_sync_axi_bus__abc_3879_new_n619_), .Y(bus_sync_axi_bus__abc_3879_new_n620_));
OR2X2 OR2X2_437 ( .A(bus_sync_axi_bus__abc_3879_new_n622_), .B(bus_sync_axi_bus__abc_3879_new_n623_), .Y(bus_sync_axi_bus__abc_3879_new_n624_));
OR2X2 OR2X2_438 ( .A(bus_sync_axi_bus__abc_3879_new_n626_), .B(bus_sync_axi_bus__abc_3879_new_n627_), .Y(bus_sync_axi_bus__abc_3879_new_n628_));
OR2X2 OR2X2_439 ( .A(bus_sync_axi_bus__abc_3879_new_n630_), .B(bus_sync_axi_bus__abc_3879_new_n631_), .Y(bus_sync_axi_bus__abc_3879_new_n632_));
OR2X2 OR2X2_44 ( .A(_abc_4268_new_n633_), .B(_abc_4268_new_n635_), .Y(_abc_4268_new_n686_));
OR2X2 OR2X2_440 ( .A(bus_sync_axi_bus__abc_3879_new_n634_), .B(bus_sync_axi_bus__abc_3879_new_n635_), .Y(bus_sync_axi_bus__abc_3879_new_n636_));
OR2X2 OR2X2_441 ( .A(bus_sync_axi_bus__abc_3879_new_n638_), .B(bus_sync_axi_bus__abc_3879_new_n639_), .Y(bus_sync_axi_bus__abc_3879_new_n640_));
OR2X2 OR2X2_442 ( .A(bus_sync_axi_bus__abc_3879_new_n642_), .B(bus_sync_axi_bus__abc_3879_new_n643_), .Y(bus_sync_axi_bus__abc_3879_new_n644_));
OR2X2 OR2X2_443 ( .A(bus_sync_axi_bus__abc_3879_new_n646_), .B(bus_sync_axi_bus__abc_3879_new_n647_), .Y(bus_sync_axi_bus__abc_3879_new_n648_));
OR2X2 OR2X2_444 ( .A(bus_sync_rdata__abc_3653_new_n266_), .B(bus_sync_rdata__abc_3653_new_n267_), .Y(bus_sync_rdata__abc_3653_new_n268_));
OR2X2 OR2X2_445 ( .A(bus_sync_rdata__abc_3653_new_n270_), .B(bus_sync_rdata__abc_3653_new_n271_), .Y(bus_sync_rdata__abc_3653_new_n272_));
OR2X2 OR2X2_446 ( .A(bus_sync_rdata__abc_3653_new_n274_), .B(bus_sync_rdata__abc_3653_new_n275_), .Y(bus_sync_rdata__abc_3653_new_n276_));
OR2X2 OR2X2_447 ( .A(bus_sync_rdata__abc_3653_new_n278_), .B(bus_sync_rdata__abc_3653_new_n279_), .Y(bus_sync_rdata__abc_3653_new_n280_));
OR2X2 OR2X2_448 ( .A(bus_sync_rdata__abc_3653_new_n282_), .B(bus_sync_rdata__abc_3653_new_n283_), .Y(bus_sync_rdata__abc_3653_new_n284_));
OR2X2 OR2X2_449 ( .A(bus_sync_rdata__abc_3653_new_n286_), .B(bus_sync_rdata__abc_3653_new_n287_), .Y(bus_sync_rdata__abc_3653_new_n288_));
OR2X2 OR2X2_45 ( .A(_abc_4268_new_n685_), .B(_abc_4268_new_n686_), .Y(_abc_4268_new_n687_));
OR2X2 OR2X2_450 ( .A(bus_sync_rdata__abc_3653_new_n290_), .B(bus_sync_rdata__abc_3653_new_n291_), .Y(bus_sync_rdata__abc_3653_new_n292_));
OR2X2 OR2X2_451 ( .A(bus_sync_rdata__abc_3653_new_n294_), .B(bus_sync_rdata__abc_3653_new_n295_), .Y(bus_sync_rdata__abc_3653_new_n296_));
OR2X2 OR2X2_452 ( .A(bus_sync_rdata__abc_3653_new_n298_), .B(bus_sync_rdata__abc_3653_new_n299_), .Y(bus_sync_rdata__abc_3653_new_n300_));
OR2X2 OR2X2_453 ( .A(bus_sync_rdata__abc_3653_new_n302_), .B(bus_sync_rdata__abc_3653_new_n303_), .Y(bus_sync_rdata__abc_3653_new_n304_));
OR2X2 OR2X2_454 ( .A(bus_sync_rdata__abc_3653_new_n306_), .B(bus_sync_rdata__abc_3653_new_n307_), .Y(bus_sync_rdata__abc_3653_new_n308_));
OR2X2 OR2X2_455 ( .A(bus_sync_rdata__abc_3653_new_n310_), .B(bus_sync_rdata__abc_3653_new_n311_), .Y(bus_sync_rdata__abc_3653_new_n312_));
OR2X2 OR2X2_456 ( .A(bus_sync_rdata__abc_3653_new_n314_), .B(bus_sync_rdata__abc_3653_new_n315_), .Y(bus_sync_rdata__abc_3653_new_n316_));
OR2X2 OR2X2_457 ( .A(bus_sync_rdata__abc_3653_new_n318_), .B(bus_sync_rdata__abc_3653_new_n319_), .Y(bus_sync_rdata__abc_3653_new_n320_));
OR2X2 OR2X2_458 ( .A(bus_sync_rdata__abc_3653_new_n322_), .B(bus_sync_rdata__abc_3653_new_n323_), .Y(bus_sync_rdata__abc_3653_new_n324_));
OR2X2 OR2X2_459 ( .A(bus_sync_rdata__abc_3653_new_n326_), .B(bus_sync_rdata__abc_3653_new_n327_), .Y(bus_sync_rdata__abc_3653_new_n328_));
OR2X2 OR2X2_46 ( .A(_abc_4268_new_n639_), .B(_abc_4268_new_n641_), .Y(_abc_4268_new_n688_));
OR2X2 OR2X2_460 ( .A(bus_sync_rdata__abc_3653_new_n330_), .B(bus_sync_rdata__abc_3653_new_n331_), .Y(bus_sync_rdata__abc_3653_new_n332_));
OR2X2 OR2X2_461 ( .A(bus_sync_rdata__abc_3653_new_n334_), .B(bus_sync_rdata__abc_3653_new_n335_), .Y(bus_sync_rdata__abc_3653_new_n336_));
OR2X2 OR2X2_462 ( .A(bus_sync_rdata__abc_3653_new_n338_), .B(bus_sync_rdata__abc_3653_new_n339_), .Y(bus_sync_rdata__abc_3653_new_n340_));
OR2X2 OR2X2_463 ( .A(bus_sync_rdata__abc_3653_new_n342_), .B(bus_sync_rdata__abc_3653_new_n343_), .Y(bus_sync_rdata__abc_3653_new_n344_));
OR2X2 OR2X2_464 ( .A(bus_sync_rdata__abc_3653_new_n346_), .B(bus_sync_rdata__abc_3653_new_n347_), .Y(bus_sync_rdata__abc_3653_new_n348_));
OR2X2 OR2X2_465 ( .A(bus_sync_rdata__abc_3653_new_n350_), .B(bus_sync_rdata__abc_3653_new_n351_), .Y(bus_sync_rdata__abc_3653_new_n352_));
OR2X2 OR2X2_466 ( .A(bus_sync_rdata__abc_3653_new_n354_), .B(bus_sync_rdata__abc_3653_new_n355_), .Y(bus_sync_rdata__abc_3653_new_n356_));
OR2X2 OR2X2_467 ( .A(bus_sync_rdata__abc_3653_new_n358_), .B(bus_sync_rdata__abc_3653_new_n359_), .Y(bus_sync_rdata__abc_3653_new_n360_));
OR2X2 OR2X2_468 ( .A(bus_sync_rdata__abc_3653_new_n362_), .B(bus_sync_rdata__abc_3653_new_n363_), .Y(bus_sync_rdata__abc_3653_new_n364_));
OR2X2 OR2X2_469 ( .A(bus_sync_rdata__abc_3653_new_n366_), .B(bus_sync_rdata__abc_3653_new_n367_), .Y(bus_sync_rdata__abc_3653_new_n368_));
OR2X2 OR2X2_47 ( .A(_abc_4268_new_n644_), .B(_abc_4268_new_n646_), .Y(_abc_4268_new_n689_));
OR2X2 OR2X2_470 ( .A(bus_sync_rdata__abc_3653_new_n370_), .B(bus_sync_rdata__abc_3653_new_n371_), .Y(bus_sync_rdata__abc_3653_new_n372_));
OR2X2 OR2X2_471 ( .A(bus_sync_rdata__abc_3653_new_n374_), .B(bus_sync_rdata__abc_3653_new_n375_), .Y(bus_sync_rdata__abc_3653_new_n376_));
OR2X2 OR2X2_472 ( .A(bus_sync_rdata__abc_3653_new_n378_), .B(bus_sync_rdata__abc_3653_new_n379_), .Y(bus_sync_rdata__abc_3653_new_n380_));
OR2X2 OR2X2_473 ( .A(bus_sync_rdata__abc_3653_new_n382_), .B(bus_sync_rdata__abc_3653_new_n383_), .Y(bus_sync_rdata__abc_3653_new_n384_));
OR2X2 OR2X2_474 ( .A(bus_sync_rdata__abc_3653_new_n386_), .B(bus_sync_rdata__abc_3653_new_n387_), .Y(bus_sync_rdata__abc_3653_new_n388_));
OR2X2 OR2X2_475 ( .A(bus_sync_rdata__abc_3653_new_n390_), .B(bus_sync_rdata__abc_3653_new_n391_), .Y(bus_sync_rdata__abc_3653_new_n392_));
OR2X2 OR2X2_476 ( .A(bus_sync_state_machine__abc_3850_new_n34_), .B(bus_sync_state_machine__abc_3850_new_n35_), .Y(bus_sync_state_machine__abc_3850_new_n36_));
OR2X2 OR2X2_477 ( .A(bus_sync_state_machine__abc_3850_new_n38_), .B(bus_sync_state_machine__abc_3850_new_n39_), .Y(bus_sync_state_machine__abc_3850_new_n40_));
OR2X2 OR2X2_478 ( .A(bus_sync_state_machine__abc_3850_new_n42_), .B(bus_sync_state_machine__abc_3850_new_n43_), .Y(bus_sync_state_machine__abc_3850_new_n44_));
OR2X2 OR2X2_479 ( .A(bus_sync_state_machine__abc_3850_new_n46_), .B(bus_sync_state_machine__abc_3850_new_n47_), .Y(bus_sync_state_machine__abc_3850_new_n48_));
OR2X2 OR2X2_48 ( .A(_abc_4268_new_n688_), .B(_abc_4268_new_n689_), .Y(_abc_4268_new_n690_));
OR2X2 OR2X2_480 ( .A(bus_sync_status__abc_3630_new_n28_), .B(bus_sync_status__abc_3630_new_n29_), .Y(bus_sync_status__abc_3630_new_n30_));
OR2X2 OR2X2_481 ( .A(bus_sync_status__abc_3630_new_n32_), .B(bus_sync_status__abc_3630_new_n33_), .Y(bus_sync_status__abc_3630_new_n34_));
OR2X2 OR2X2_482 ( .A(bus_sync_status__abc_3630_new_n36_), .B(bus_sync_status__abc_3630_new_n37_), .Y(bus_sync_status__abc_3630_new_n38_));
OR2X2 OR2X2_49 ( .A(_abc_4268_new_n687_), .B(_abc_4268_new_n690_), .Y(_abc_4268_new_n691_));
OR2X2 OR2X2_5 ( .A(axi_bready), .B(axi_rready), .Y(_abc_4268_new_n571_));
OR2X2 OR2X2_50 ( .A(_abc_4268_new_n651_), .B(_abc_4268_new_n653_), .Y(_abc_4268_new_n692_));
OR2X2 OR2X2_51 ( .A(_abc_4268_new_n656_), .B(_abc_4268_new_n658_), .Y(_abc_4268_new_n693_));
OR2X2 OR2X2_52 ( .A(_abc_4268_new_n692_), .B(_abc_4268_new_n693_), .Y(_abc_4268_new_n694_));
OR2X2 OR2X2_53 ( .A(_abc_4268_new_n662_), .B(_abc_4268_new_n664_), .Y(_abc_4268_new_n695_));
OR2X2 OR2X2_54 ( .A(counter_18_), .B(counter_19_), .Y(_abc_4268_new_n696_));
OR2X2 OR2X2_55 ( .A(_abc_4268_new_n667_), .B(_abc_4268_new_n696_), .Y(_abc_4268_new_n697_));
OR2X2 OR2X2_56 ( .A(_abc_4268_new_n695_), .B(_abc_4268_new_n697_), .Y(_abc_4268_new_n698_));
OR2X2 OR2X2_57 ( .A(_abc_4268_new_n694_), .B(_abc_4268_new_n698_), .Y(_abc_4268_new_n699_));
OR2X2 OR2X2_58 ( .A(_abc_4268_new_n691_), .B(_abc_4268_new_n699_), .Y(_abc_4268_new_n700_));
OR2X2 OR2X2_59 ( .A(_abc_4268_new_n701_), .B(bus_cap_1_), .Y(_abc_4268_new_n702_));
OR2X2 OR2X2_6 ( .A(_abc_4268_new_n571_), .B(_abc_4268_new_n572_), .Y(_abc_4268_new_n573_));
OR2X2 OR2X2_60 ( .A(_abc_4268_new_n676_), .B(bus_cap_0_), .Y(_abc_4268_new_n703_));
OR2X2 OR2X2_61 ( .A(_abc_4268_new_n704_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n705_));
OR2X2 OR2X2_62 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n707_), .Y(_abc_4268_new_n708_));
OR2X2 OR2X2_63 ( .A(_abc_4268_new_n708_), .B(_abc_4268_new_n706_), .Y(_abc_4268_new_n709_));
OR2X2 OR2X2_64 ( .A(_abc_4268_new_n701_), .B(bus_cap_2_), .Y(_abc_4268_new_n712_));
OR2X2 OR2X2_65 ( .A(_abc_4268_new_n676_), .B(bus_cap_1_), .Y(_abc_4268_new_n713_));
OR2X2 OR2X2_66 ( .A(_abc_4268_new_n714_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n715_));
OR2X2 OR2X2_67 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n717_), .Y(_abc_4268_new_n718_));
OR2X2 OR2X2_68 ( .A(_abc_4268_new_n718_), .B(_abc_4268_new_n716_), .Y(_abc_4268_new_n719_));
OR2X2 OR2X2_69 ( .A(_abc_4268_new_n701_), .B(bus_cap_3_), .Y(_abc_4268_new_n722_));
OR2X2 OR2X2_7 ( .A(_abc_4268_new_n587_), .B(_abc_4268_new_n577_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_6_));
OR2X2 OR2X2_70 ( .A(_abc_4268_new_n676_), .B(bus_cap_2_), .Y(_abc_4268_new_n723_));
OR2X2 OR2X2_71 ( .A(_abc_4268_new_n724_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n725_));
OR2X2 OR2X2_72 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n726_), .Y(_abc_4268_new_n727_));
OR2X2 OR2X2_73 ( .A(_abc_4268_new_n701_), .B(bus_cap_4_), .Y(_abc_4268_new_n730_));
OR2X2 OR2X2_74 ( .A(_abc_4268_new_n676_), .B(bus_cap_3_), .Y(_abc_4268_new_n731_));
OR2X2 OR2X2_75 ( .A(_abc_4268_new_n732_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n733_));
OR2X2 OR2X2_76 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n734_), .Y(_abc_4268_new_n735_));
OR2X2 OR2X2_77 ( .A(_abc_4268_new_n701_), .B(bus_cap_5_), .Y(_abc_4268_new_n738_));
OR2X2 OR2X2_78 ( .A(_abc_4268_new_n676_), .B(bus_cap_4_), .Y(_abc_4268_new_n739_));
OR2X2 OR2X2_79 ( .A(_abc_4268_new_n740_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n741_));
OR2X2 OR2X2_8 ( .A(_abc_4268_new_n589_), .B(_abc_4268_new_n592_), .Y(_abc_2903_auto_fsm_map_cc_170_map_fsm_402_4_));
OR2X2 OR2X2_80 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n742_), .Y(_abc_4268_new_n743_));
OR2X2 OR2X2_81 ( .A(_abc_4268_new_n701_), .B(bus_cap_6_), .Y(_abc_4268_new_n746_));
OR2X2 OR2X2_82 ( .A(_abc_4268_new_n676_), .B(bus_cap_5_), .Y(_abc_4268_new_n747_));
OR2X2 OR2X2_83 ( .A(_abc_4268_new_n748_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n749_));
OR2X2 OR2X2_84 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n750_), .Y(_abc_4268_new_n751_));
OR2X2 OR2X2_85 ( .A(_abc_4268_new_n701_), .B(bus_cap_7_), .Y(_abc_4268_new_n754_));
OR2X2 OR2X2_86 ( .A(_abc_4268_new_n676_), .B(bus_cap_6_), .Y(_abc_4268_new_n755_));
OR2X2 OR2X2_87 ( .A(_abc_4268_new_n756_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n757_));
OR2X2 OR2X2_88 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n758_), .Y(_abc_4268_new_n759_));
OR2X2 OR2X2_89 ( .A(_abc_4268_new_n701_), .B(bus_cap_8_), .Y(_abc_4268_new_n762_));
OR2X2 OR2X2_9 ( .A(axi_rready), .B(state_6_), .Y(_abc_4268_new_n594_));
OR2X2 OR2X2_90 ( .A(_abc_4268_new_n676_), .B(bus_cap_7_), .Y(_abc_4268_new_n763_));
OR2X2 OR2X2_91 ( .A(_abc_4268_new_n764_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n765_));
OR2X2 OR2X2_92 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n766_), .Y(_abc_4268_new_n767_));
OR2X2 OR2X2_93 ( .A(_abc_4268_new_n701_), .B(bus_cap_9_), .Y(_abc_4268_new_n770_));
OR2X2 OR2X2_94 ( .A(_abc_4268_new_n676_), .B(bus_cap_8_), .Y(_abc_4268_new_n771_));
OR2X2 OR2X2_95 ( .A(_abc_4268_new_n772_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n773_));
OR2X2 OR2X2_96 ( .A(_abc_4268_new_n621_), .B(_abc_4268_new_n774_), .Y(_abc_4268_new_n775_));
OR2X2 OR2X2_97 ( .A(_abc_4268_new_n701_), .B(bus_cap_10_), .Y(_abc_4268_new_n778_));
OR2X2 OR2X2_98 ( .A(_abc_4268_new_n676_), .B(bus_cap_9_), .Y(_abc_4268_new_n779_));
OR2X2 OR2X2_99 ( .A(_abc_4268_new_n780_), .B(_abc_4268_new_n622_), .Y(_abc_4268_new_n781_));

assign \axi_arprot[0]  = 1'h0;
assign \axi_arprot[1]  = 1'h0;
assign \axi_arprot[2]  = 1'h0;
assign \axi_awprot[0]  = 1'h0;
assign \axi_awprot[1]  = 1'h0;
assign \axi_awprot[2]  = 1'h0;
assign \axi_wstrb[0]  = 1'h1;
assign \axi_wstrb[1]  = 1'h1;
assign \axi_wstrb[2]  = 1'h1;
assign \axi_wstrb[3]  = 1'h1;

endmodule