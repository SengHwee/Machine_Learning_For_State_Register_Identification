
module altor32_lite(clk_i, rst_i, intr_i, nmi_i, enable_i, \mem_dat_i[0] , \mem_dat_i[1] , \mem_dat_i[2] , \mem_dat_i[3] , \mem_dat_i[4] , \mem_dat_i[5] , \mem_dat_i[6] , \mem_dat_i[7] , \mem_dat_i[8] , \mem_dat_i[9] , \mem_dat_i[10] , \mem_dat_i[11] , \mem_dat_i[12] , \mem_dat_i[13] , \mem_dat_i[14] , \mem_dat_i[15] , \mem_dat_i[16] , \mem_dat_i[17] , \mem_dat_i[18] , \mem_dat_i[19] , \mem_dat_i[20] , \mem_dat_i[21] , \mem_dat_i[22] , \mem_dat_i[23] , \mem_dat_i[24] , \mem_dat_i[25] , \mem_dat_i[26] , \mem_dat_i[27] , \mem_dat_i[28] , \mem_dat_i[29] , \mem_dat_i[30] , \mem_dat_i[31] , mem_stall_i, mem_ack_i, fault_o, break_o, \mem_addr_o[0] , \mem_addr_o[1] , \mem_addr_o[2] , \mem_addr_o[3] , \mem_addr_o[4] , \mem_addr_o[5] , \mem_addr_o[6] , \mem_addr_o[7] , \mem_addr_o[8] , \mem_addr_o[9] , \mem_addr_o[10] , \mem_addr_o[11] , \mem_addr_o[12] , \mem_addr_o[13] , \mem_addr_o[14] , \mem_addr_o[15] , \mem_addr_o[16] , \mem_addr_o[17] , \mem_addr_o[18] , \mem_addr_o[19] , \mem_addr_o[20] , \mem_addr_o[21] , \mem_addr_o[22] , \mem_addr_o[23] , \mem_addr_o[24] , \mem_addr_o[25] , \mem_addr_o[26] , \mem_addr_o[27] , \mem_addr_o[28] , \mem_addr_o[29] , \mem_addr_o[30] , \mem_addr_o[31] , \mem_dat_o[0] , \mem_dat_o[1] , \mem_dat_o[2] , \mem_dat_o[3] , \mem_dat_o[4] , \mem_dat_o[5] , \mem_dat_o[6] , \mem_dat_o[7] , \mem_dat_o[8] , \mem_dat_o[9] , \mem_dat_o[10] , \mem_dat_o[11] , \mem_dat_o[12] , \mem_dat_o[13] , \mem_dat_o[14] , \mem_dat_o[15] , \mem_dat_o[16] , \mem_dat_o[17] , \mem_dat_o[18] , \mem_dat_o[19] , \mem_dat_o[20] , \mem_dat_o[21] , \mem_dat_o[22] , \mem_dat_o[23] , \mem_dat_o[24] , \mem_dat_o[25] , \mem_dat_o[26] , \mem_dat_o[27] , \mem_dat_o[28] , \mem_dat_o[29] , \mem_dat_o[30] , \mem_dat_o[31] , \mem_cti_o[0] , \mem_cti_o[1] , \mem_cti_o[2] , mem_cyc_o, mem_stb_o, mem_we_o, \mem_sel_o[0] , \mem_sel_o[1] , \mem_sel_o[2] , \mem_sel_o[3] );
  wire REGFILE_SIM_reg_bank__abc_33898_n2099_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2100;
  wire REGFILE_SIM_reg_bank__abc_33898_n2101_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2102;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n2104;
  wire REGFILE_SIM_reg_bank__abc_33898_n2105_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2106_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2107;
  wire REGFILE_SIM_reg_bank__abc_33898_n2109_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2110;
  wire REGFILE_SIM_reg_bank__abc_33898_n2111_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2112_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2114_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2115_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2116;
  wire REGFILE_SIM_reg_bank__abc_33898_n2117_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2119;
  wire REGFILE_SIM_reg_bank__abc_33898_n2120_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2121_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2122;
  wire REGFILE_SIM_reg_bank__abc_33898_n2124_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2125;
  wire REGFILE_SIM_reg_bank__abc_33898_n2126_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2127_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2129_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2130_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2131;
  wire REGFILE_SIM_reg_bank__abc_33898_n2132_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2134;
  wire REGFILE_SIM_reg_bank__abc_33898_n2135_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2136_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2137;
  wire REGFILE_SIM_reg_bank__abc_33898_n2139_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2140;
  wire REGFILE_SIM_reg_bank__abc_33898_n2141_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2142_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2144_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2145_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2146;
  wire REGFILE_SIM_reg_bank__abc_33898_n2147_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2149;
  wire REGFILE_SIM_reg_bank__abc_33898_n2150_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2151_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2152;
  wire REGFILE_SIM_reg_bank__abc_33898_n2154_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2155;
  wire REGFILE_SIM_reg_bank__abc_33898_n2156_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2157_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2159_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2160_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2161;
  wire REGFILE_SIM_reg_bank__abc_33898_n2162_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2164;
  wire REGFILE_SIM_reg_bank__abc_33898_n2165_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2166_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2167;
  wire REGFILE_SIM_reg_bank__abc_33898_n2169_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2170;
  wire REGFILE_SIM_reg_bank__abc_33898_n2171_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2172_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2174_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2175_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2176;
  wire REGFILE_SIM_reg_bank__abc_33898_n2177_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2179;
  wire REGFILE_SIM_reg_bank__abc_33898_n2180_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2181_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2182;
  wire REGFILE_SIM_reg_bank__abc_33898_n2184_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2185;
  wire REGFILE_SIM_reg_bank__abc_33898_n2186_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2187_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2189_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2190_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2191;
  wire REGFILE_SIM_reg_bank__abc_33898_n2192_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2194;
  wire REGFILE_SIM_reg_bank__abc_33898_n2195_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2196_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2197;
  wire REGFILE_SIM_reg_bank__abc_33898_n2199;
  wire REGFILE_SIM_reg_bank__abc_33898_n2200_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2201;
  wire REGFILE_SIM_reg_bank__abc_33898_n2202_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2204;
  wire REGFILE_SIM_reg_bank__abc_33898_n2205_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2206_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2207;
  wire REGFILE_SIM_reg_bank__abc_33898_n2209_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2210;
  wire REGFILE_SIM_reg_bank__abc_33898_n2211_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2212_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2214_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2215_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2216;
  wire REGFILE_SIM_reg_bank__abc_33898_n2217_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2219;
  wire REGFILE_SIM_reg_bank__abc_33898_n2220_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2221_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2222;
  wire REGFILE_SIM_reg_bank__abc_33898_n2224_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2225;
  wire REGFILE_SIM_reg_bank__abc_33898_n2226_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2227_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2229_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2230_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2231;
  wire REGFILE_SIM_reg_bank__abc_33898_n2232_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2234;
  wire REGFILE_SIM_reg_bank__abc_33898_n2235_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2236_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2237;
  wire REGFILE_SIM_reg_bank__abc_33898_n2239_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2240;
  wire REGFILE_SIM_reg_bank__abc_33898_n2241_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2242_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2244_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2245_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2246;
  wire REGFILE_SIM_reg_bank__abc_33898_n2247_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2249;
  wire REGFILE_SIM_reg_bank__abc_33898_n2250_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2251_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2252;
  wire REGFILE_SIM_reg_bank__abc_33898_n2254_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2255;
  wire REGFILE_SIM_reg_bank__abc_33898_n2256_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2257_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2259_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2260_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2261;
  wire REGFILE_SIM_reg_bank__abc_33898_n2262_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2264;
  wire REGFILE_SIM_reg_bank__abc_33898_n2265_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2266_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2267;
  wire REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2268_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2269_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2270;
  wire REGFILE_SIM_reg_bank__abc_33898_n2272_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2273;
  wire REGFILE_SIM_reg_bank__abc_33898_n2275_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2276;
  wire REGFILE_SIM_reg_bank__abc_33898_n2278_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2279;
  wire REGFILE_SIM_reg_bank__abc_33898_n2281_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2282;
  wire REGFILE_SIM_reg_bank__abc_33898_n2284_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2285;
  wire REGFILE_SIM_reg_bank__abc_33898_n2287_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2288;
  wire REGFILE_SIM_reg_bank__abc_33898_n2290_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2291;
  wire REGFILE_SIM_reg_bank__abc_33898_n2293_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2294;
  wire REGFILE_SIM_reg_bank__abc_33898_n2296;
  wire REGFILE_SIM_reg_bank__abc_33898_n2297_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2299_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2300_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2302_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2303_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2305_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2306_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2308_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2309_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2311_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2312_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2314_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2315_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2317_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2318_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2320_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2321_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2323_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2324_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2326_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2327_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2329_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2330_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2332_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2333_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2335_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2336_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2338_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2339_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2341_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2342_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2344_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2345_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2347_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2348_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2350_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2351_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2353_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2354_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2356_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2357_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2359_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2360_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2362_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2363_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2365_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2366_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2367;
  wire REGFILE_SIM_reg_bank__abc_33898_n2368_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2369_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2370;
  wire REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2371_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2373;
  wire REGFILE_SIM_reg_bank__abc_33898_n2374_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2376;
  wire REGFILE_SIM_reg_bank__abc_33898_n2377_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2379;
  wire REGFILE_SIM_reg_bank__abc_33898_n2380_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2382;
  wire REGFILE_SIM_reg_bank__abc_33898_n2383_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2385;
  wire REGFILE_SIM_reg_bank__abc_33898_n2386_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2388;
  wire REGFILE_SIM_reg_bank__abc_33898_n2389_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2391;
  wire REGFILE_SIM_reg_bank__abc_33898_n2392_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2394_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2395;
  wire REGFILE_SIM_reg_bank__abc_33898_n2397_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2398;
  wire REGFILE_SIM_reg_bank__abc_33898_n2400_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2401;
  wire REGFILE_SIM_reg_bank__abc_33898_n2403_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2404;
  wire REGFILE_SIM_reg_bank__abc_33898_n2406_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2407;
  wire REGFILE_SIM_reg_bank__abc_33898_n2409_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2410;
  wire REGFILE_SIM_reg_bank__abc_33898_n2412_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2413;
  wire REGFILE_SIM_reg_bank__abc_33898_n2415_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2416;
  wire REGFILE_SIM_reg_bank__abc_33898_n2418_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2419;
  wire REGFILE_SIM_reg_bank__abc_33898_n2421_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2422;
  wire REGFILE_SIM_reg_bank__abc_33898_n2424_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2425;
  wire REGFILE_SIM_reg_bank__abc_33898_n2427_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2428;
  wire REGFILE_SIM_reg_bank__abc_33898_n2430_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2431;
  wire REGFILE_SIM_reg_bank__abc_33898_n2433_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2434;
  wire REGFILE_SIM_reg_bank__abc_33898_n2436_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2437;
  wire REGFILE_SIM_reg_bank__abc_33898_n2439_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2440;
  wire REGFILE_SIM_reg_bank__abc_33898_n2442_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2443;
  wire REGFILE_SIM_reg_bank__abc_33898_n2445_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2446;
  wire REGFILE_SIM_reg_bank__abc_33898_n2448_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2449;
  wire REGFILE_SIM_reg_bank__abc_33898_n2451_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2452;
  wire REGFILE_SIM_reg_bank__abc_33898_n2454_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2455;
  wire REGFILE_SIM_reg_bank__abc_33898_n2457_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2458;
  wire REGFILE_SIM_reg_bank__abc_33898_n2460_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2461;
  wire REGFILE_SIM_reg_bank__abc_33898_n2463_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2464;
  wire REGFILE_SIM_reg_bank__abc_33898_n2466_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2467;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n2469_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2470;
  wire REGFILE_SIM_reg_bank__abc_33898_n2471_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2473;
  wire REGFILE_SIM_reg_bank__abc_33898_n2474_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2475_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2477_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2478_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2479;
  wire REGFILE_SIM_reg_bank__abc_33898_n2481_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2482;
  wire REGFILE_SIM_reg_bank__abc_33898_n2483_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2485;
  wire REGFILE_SIM_reg_bank__abc_33898_n2486_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2487_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2489_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2490;
  wire REGFILE_SIM_reg_bank__abc_33898_n2491_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2493_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2494_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2495;
  wire REGFILE_SIM_reg_bank__abc_33898_n2497_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2498;
  wire REGFILE_SIM_reg_bank__abc_33898_n2499_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2501;
  wire REGFILE_SIM_reg_bank__abc_33898_n2502_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2503_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2505_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2506_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2507;
  wire REGFILE_SIM_reg_bank__abc_33898_n2509_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2510;
  wire REGFILE_SIM_reg_bank__abc_33898_n2511_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2513;
  wire REGFILE_SIM_reg_bank__abc_33898_n2514_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2515_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2517_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2518_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2519;
  wire REGFILE_SIM_reg_bank__abc_33898_n2521_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2522;
  wire REGFILE_SIM_reg_bank__abc_33898_n2523_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2525;
  wire REGFILE_SIM_reg_bank__abc_33898_n2526_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2527_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2529_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2530_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2531;
  wire REGFILE_SIM_reg_bank__abc_33898_n2533_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2534;
  wire REGFILE_SIM_reg_bank__abc_33898_n2535_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2537;
  wire REGFILE_SIM_reg_bank__abc_33898_n2538_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2539_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2541_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2542_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2543;
  wire REGFILE_SIM_reg_bank__abc_33898_n2545_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2546;
  wire REGFILE_SIM_reg_bank__abc_33898_n2547_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2549;
  wire REGFILE_SIM_reg_bank__abc_33898_n2550_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2551_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2553_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2554_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2555;
  wire REGFILE_SIM_reg_bank__abc_33898_n2557_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2558;
  wire REGFILE_SIM_reg_bank__abc_33898_n2559_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2561;
  wire REGFILE_SIM_reg_bank__abc_33898_n2562_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2563_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2565_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2566_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2567;
  wire REGFILE_SIM_reg_bank__abc_33898_n2569_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2570;
  wire REGFILE_SIM_reg_bank__abc_33898_n2571_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2573;
  wire REGFILE_SIM_reg_bank__abc_33898_n2574_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2575_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2577_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2578_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2579;
  wire REGFILE_SIM_reg_bank__abc_33898_n2581_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2582;
  wire REGFILE_SIM_reg_bank__abc_33898_n2583_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2585;
  wire REGFILE_SIM_reg_bank__abc_33898_n2586_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2587;
  wire REGFILE_SIM_reg_bank__abc_33898_n2589;
  wire REGFILE_SIM_reg_bank__abc_33898_n2590_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2591_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2593_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2594_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2595;
  wire REGFILE_SIM_reg_bank__abc_33898_n2597_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2598;
  wire REGFILE_SIM_reg_bank__abc_33898_n2599_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2600_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2601;
  wire REGFILE_SIM_reg_bank__abc_33898_n2602_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2603_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2605_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2606_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2608_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2609_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2611_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2612_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2614_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2615_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2617_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2618_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2620_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2621_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2623_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2624_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2626_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2627_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2629_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2630_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2632_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2633_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2635_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2636_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2638_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2639_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2641_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2642_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2644_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2645_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2647_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2648_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2650_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2651_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2653_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2654_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2656_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2657_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2659_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2660_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2662_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2663_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2665_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2666_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2668_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2669_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2671_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2672_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2674_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2675_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2677_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2678_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2680_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2681_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2683_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2684;
  wire REGFILE_SIM_reg_bank__abc_33898_n2686;
  wire REGFILE_SIM_reg_bank__abc_33898_n2687_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2689;
  wire REGFILE_SIM_reg_bank__abc_33898_n2690_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2692;
  wire REGFILE_SIM_reg_bank__abc_33898_n2693_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2695;
  wire REGFILE_SIM_reg_bank__abc_33898_n2696_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2698;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n2700_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2701;
  wire REGFILE_SIM_reg_bank__abc_33898_n2702_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2704;
  wire REGFILE_SIM_reg_bank__abc_33898_n2705_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2706_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2708_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2709_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2710;
  wire REGFILE_SIM_reg_bank__abc_33898_n2712_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2713;
  wire REGFILE_SIM_reg_bank__abc_33898_n2714_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2716;
  wire REGFILE_SIM_reg_bank__abc_33898_n2717_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2718_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2720_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2721_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2722;
  wire REGFILE_SIM_reg_bank__abc_33898_n2724_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2725;
  wire REGFILE_SIM_reg_bank__abc_33898_n2726_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2728;
  wire REGFILE_SIM_reg_bank__abc_33898_n2729_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2730_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2732_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2733_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2734;
  wire REGFILE_SIM_reg_bank__abc_33898_n2736_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2737;
  wire REGFILE_SIM_reg_bank__abc_33898_n2738_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2740;
  wire REGFILE_SIM_reg_bank__abc_33898_n2741_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2742_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2744_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2745_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2746;
  wire REGFILE_SIM_reg_bank__abc_33898_n2748_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2749;
  wire REGFILE_SIM_reg_bank__abc_33898_n2750_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2752;
  wire REGFILE_SIM_reg_bank__abc_33898_n2753_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2754_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2756_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2757_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2758;
  wire REGFILE_SIM_reg_bank__abc_33898_n2760_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2761;
  wire REGFILE_SIM_reg_bank__abc_33898_n2762_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2764;
  wire REGFILE_SIM_reg_bank__abc_33898_n2765_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2766_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2768_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2769_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2770;
  wire REGFILE_SIM_reg_bank__abc_33898_n2772_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2773;
  wire REGFILE_SIM_reg_bank__abc_33898_n2774_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2776;
  wire REGFILE_SIM_reg_bank__abc_33898_n2777_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2778_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2780_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2781;
  wire REGFILE_SIM_reg_bank__abc_33898_n2782_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2784_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2785_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2786;
  wire REGFILE_SIM_reg_bank__abc_33898_n2788_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2789;
  wire REGFILE_SIM_reg_bank__abc_33898_n2790_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2792;
  wire REGFILE_SIM_reg_bank__abc_33898_n2793_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2794_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2796_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2797_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2798;
  wire REGFILE_SIM_reg_bank__abc_33898_n2800_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2801;
  wire REGFILE_SIM_reg_bank__abc_33898_n2802_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2804;
  wire REGFILE_SIM_reg_bank__abc_33898_n2805_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2806_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2808_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2809_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2810;
  wire REGFILE_SIM_reg_bank__abc_33898_n2812_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2813;
  wire REGFILE_SIM_reg_bank__abc_33898_n2814_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2816;
  wire REGFILE_SIM_reg_bank__abc_33898_n2817_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2818_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2820_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2821_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2822;
  wire REGFILE_SIM_reg_bank__abc_33898_n2824_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2825;
  wire REGFILE_SIM_reg_bank__abc_33898_n2826_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2828;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n2830_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2831;
  wire REGFILE_SIM_reg_bank__abc_33898_n2832_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2834;
  wire REGFILE_SIM_reg_bank__abc_33898_n2835_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2836_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2838_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2839_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2840;
  wire REGFILE_SIM_reg_bank__abc_33898_n2842_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2843;
  wire REGFILE_SIM_reg_bank__abc_33898_n2844_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2846;
  wire REGFILE_SIM_reg_bank__abc_33898_n2847_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2848_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2850_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2851_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2852;
  wire REGFILE_SIM_reg_bank__abc_33898_n2854_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2855;
  wire REGFILE_SIM_reg_bank__abc_33898_n2856_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2858;
  wire REGFILE_SIM_reg_bank__abc_33898_n2859_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2860_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2862_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2863_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2864;
  wire REGFILE_SIM_reg_bank__abc_33898_n2866_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2867;
  wire REGFILE_SIM_reg_bank__abc_33898_n2868_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2870;
  wire REGFILE_SIM_reg_bank__abc_33898_n2871_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2872_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2874_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2875_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2876;
  wire REGFILE_SIM_reg_bank__abc_33898_n2878;
  wire REGFILE_SIM_reg_bank__abc_33898_n2879_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2880;
  wire REGFILE_SIM_reg_bank__abc_33898_n2882_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2883;
  wire REGFILE_SIM_reg_bank__abc_33898_n2884_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2886;
  wire REGFILE_SIM_reg_bank__abc_33898_n2887_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2888_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2890_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2891_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2892;
  wire REGFILE_SIM_reg_bank__abc_33898_n2894_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2895;
  wire REGFILE_SIM_reg_bank__abc_33898_n2896_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2898;
  wire REGFILE_SIM_reg_bank__abc_33898_n2899_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2900_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2902_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2903_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2904;
  wire REGFILE_SIM_reg_bank__abc_33898_n2906_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2907;
  wire REGFILE_SIM_reg_bank__abc_33898_n2908_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2910;
  wire REGFILE_SIM_reg_bank__abc_33898_n2911_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2912_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2914_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2915_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2916;
  wire REGFILE_SIM_reg_bank__abc_33898_n2918_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2919;
  wire REGFILE_SIM_reg_bank__abc_33898_n2920_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2922;
  wire REGFILE_SIM_reg_bank__abc_33898_n2923_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2924_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2926_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2927_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2928;
  wire REGFILE_SIM_reg_bank__abc_33898_n2930_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2931;
  wire REGFILE_SIM_reg_bank__abc_33898_n2932_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2934;
  wire REGFILE_SIM_reg_bank__abc_33898_n2935_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2936_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2938_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2939_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2940;
  wire REGFILE_SIM_reg_bank__abc_33898_n2942_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2943;
  wire REGFILE_SIM_reg_bank__abc_33898_n2944_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2946;
  wire REGFILE_SIM_reg_bank__abc_33898_n2947_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2948_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2950_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2951_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2952;
  wire REGFILE_SIM_reg_bank__abc_33898_n2954_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2955;
  wire REGFILE_SIM_reg_bank__abc_33898_n2956_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2958;
  wire REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2959_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2960_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n2961;
  wire REGFILE_SIM_reg_bank__abc_33898_n2963_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2964;
  wire REGFILE_SIM_reg_bank__abc_33898_n2966_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2967;
  wire REGFILE_SIM_reg_bank__abc_33898_n2969_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2970;
  wire REGFILE_SIM_reg_bank__abc_33898_n2972_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2973;
  wire REGFILE_SIM_reg_bank__abc_33898_n2975;
  wire REGFILE_SIM_reg_bank__abc_33898_n2976_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2978_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2979_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2981_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2982_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2984_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2985_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2987_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2988_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2990_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2991_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2993_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2994_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2996_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2997_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n2999_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3000_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3002_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3003_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3005_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3006_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3008_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3009_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3011_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3012_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3014_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3015_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3017_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3018_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3020_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3021_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3023_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3024_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3026_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3027_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3029_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3030_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3032_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3033_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3035_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3036_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3038_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3039_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3041_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3042_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3044_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3045_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3047_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3048_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3050_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3051_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3053_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3054_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3056_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3057_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3058;
  wire REGFILE_SIM_reg_bank__abc_33898_n3059_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3060_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3061;
  wire REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3062_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3064;
  wire REGFILE_SIM_reg_bank__abc_33898_n3065_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3067;
  wire REGFILE_SIM_reg_bank__abc_33898_n3068_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3070;
  wire REGFILE_SIM_reg_bank__abc_33898_n3071_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3073;
  wire REGFILE_SIM_reg_bank__abc_33898_n3074_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3076;
  wire REGFILE_SIM_reg_bank__abc_33898_n3077_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3079_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3080;
  wire REGFILE_SIM_reg_bank__abc_33898_n3082;
  wire REGFILE_SIM_reg_bank__abc_33898_n3083;
  wire REGFILE_SIM_reg_bank__abc_33898_n3085;
  wire REGFILE_SIM_reg_bank__abc_33898_n3086;
  wire REGFILE_SIM_reg_bank__abc_33898_n3088;
  wire REGFILE_SIM_reg_bank__abc_33898_n3089;
  wire REGFILE_SIM_reg_bank__abc_33898_n3091;
  wire REGFILE_SIM_reg_bank__abc_33898_n3092;
  wire REGFILE_SIM_reg_bank__abc_33898_n3094;
  wire REGFILE_SIM_reg_bank__abc_33898_n3095;
  wire REGFILE_SIM_reg_bank__abc_33898_n3097;
  wire REGFILE_SIM_reg_bank__abc_33898_n3098;
  wire REGFILE_SIM_reg_bank__abc_33898_n3100;
  wire REGFILE_SIM_reg_bank__abc_33898_n3101;
  wire REGFILE_SIM_reg_bank__abc_33898_n3103;
  wire REGFILE_SIM_reg_bank__abc_33898_n3104;
  wire REGFILE_SIM_reg_bank__abc_33898_n3106;
  wire REGFILE_SIM_reg_bank__abc_33898_n3107;
  wire REGFILE_SIM_reg_bank__abc_33898_n3109;
  wire REGFILE_SIM_reg_bank__abc_33898_n3110;
  wire REGFILE_SIM_reg_bank__abc_33898_n3112;
  wire REGFILE_SIM_reg_bank__abc_33898_n3113;
  wire REGFILE_SIM_reg_bank__abc_33898_n3115;
  wire REGFILE_SIM_reg_bank__abc_33898_n3116;
  wire REGFILE_SIM_reg_bank__abc_33898_n3118;
  wire REGFILE_SIM_reg_bank__abc_33898_n3119;
  wire REGFILE_SIM_reg_bank__abc_33898_n3121;
  wire REGFILE_SIM_reg_bank__abc_33898_n3122;
  wire REGFILE_SIM_reg_bank__abc_33898_n3124;
  wire REGFILE_SIM_reg_bank__abc_33898_n3125;
  wire REGFILE_SIM_reg_bank__abc_33898_n3127;
  wire REGFILE_SIM_reg_bank__abc_33898_n3128;
  wire REGFILE_SIM_reg_bank__abc_33898_n3130;
  wire REGFILE_SIM_reg_bank__abc_33898_n3131;
  wire REGFILE_SIM_reg_bank__abc_33898_n3133;
  wire REGFILE_SIM_reg_bank__abc_33898_n3134;
  wire REGFILE_SIM_reg_bank__abc_33898_n3136;
  wire REGFILE_SIM_reg_bank__abc_33898_n3137;
  wire REGFILE_SIM_reg_bank__abc_33898_n3139;
  wire REGFILE_SIM_reg_bank__abc_33898_n3140;
  wire REGFILE_SIM_reg_bank__abc_33898_n3142;
  wire REGFILE_SIM_reg_bank__abc_33898_n3143;
  wire REGFILE_SIM_reg_bank__abc_33898_n3145;
  wire REGFILE_SIM_reg_bank__abc_33898_n3146;
  wire REGFILE_SIM_reg_bank__abc_33898_n3148;
  wire REGFILE_SIM_reg_bank__abc_33898_n3149;
  wire REGFILE_SIM_reg_bank__abc_33898_n3151;
  wire REGFILE_SIM_reg_bank__abc_33898_n3152;
  wire REGFILE_SIM_reg_bank__abc_33898_n3154;
  wire REGFILE_SIM_reg_bank__abc_33898_n3155;
  wire REGFILE_SIM_reg_bank__abc_33898_n3157;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n3159;
  wire REGFILE_SIM_reg_bank__abc_33898_n3160;
  wire REGFILE_SIM_reg_bank__abc_33898_n3161;
  wire REGFILE_SIM_reg_bank__abc_33898_n3163;
  wire REGFILE_SIM_reg_bank__abc_33898_n3164;
  wire REGFILE_SIM_reg_bank__abc_33898_n3165;
  wire REGFILE_SIM_reg_bank__abc_33898_n3167;
  wire REGFILE_SIM_reg_bank__abc_33898_n3168;
  wire REGFILE_SIM_reg_bank__abc_33898_n3169;
  wire REGFILE_SIM_reg_bank__abc_33898_n3171;
  wire REGFILE_SIM_reg_bank__abc_33898_n3172;
  wire REGFILE_SIM_reg_bank__abc_33898_n3173;
  wire REGFILE_SIM_reg_bank__abc_33898_n3175;
  wire REGFILE_SIM_reg_bank__abc_33898_n3176;
  wire REGFILE_SIM_reg_bank__abc_33898_n3177;
  wire REGFILE_SIM_reg_bank__abc_33898_n3179;
  wire REGFILE_SIM_reg_bank__abc_33898_n3180;
  wire REGFILE_SIM_reg_bank__abc_33898_n3181;
  wire REGFILE_SIM_reg_bank__abc_33898_n3183;
  wire REGFILE_SIM_reg_bank__abc_33898_n3184;
  wire REGFILE_SIM_reg_bank__abc_33898_n3185;
  wire REGFILE_SIM_reg_bank__abc_33898_n3187;
  wire REGFILE_SIM_reg_bank__abc_33898_n3188;
  wire REGFILE_SIM_reg_bank__abc_33898_n3189;
  wire REGFILE_SIM_reg_bank__abc_33898_n3191;
  wire REGFILE_SIM_reg_bank__abc_33898_n3192;
  wire REGFILE_SIM_reg_bank__abc_33898_n3193;
  wire REGFILE_SIM_reg_bank__abc_33898_n3195;
  wire REGFILE_SIM_reg_bank__abc_33898_n3196;
  wire REGFILE_SIM_reg_bank__abc_33898_n3197_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3199;
  wire REGFILE_SIM_reg_bank__abc_33898_n3200;
  wire REGFILE_SIM_reg_bank__abc_33898_n3201;
  wire REGFILE_SIM_reg_bank__abc_33898_n3203;
  wire REGFILE_SIM_reg_bank__abc_33898_n3204;
  wire REGFILE_SIM_reg_bank__abc_33898_n3205;
  wire REGFILE_SIM_reg_bank__abc_33898_n3207;
  wire REGFILE_SIM_reg_bank__abc_33898_n3208;
  wire REGFILE_SIM_reg_bank__abc_33898_n3209;
  wire REGFILE_SIM_reg_bank__abc_33898_n3211;
  wire REGFILE_SIM_reg_bank__abc_33898_n3212;
  wire REGFILE_SIM_reg_bank__abc_33898_n3213;
  wire REGFILE_SIM_reg_bank__abc_33898_n3215;
  wire REGFILE_SIM_reg_bank__abc_33898_n3216;
  wire REGFILE_SIM_reg_bank__abc_33898_n3217;
  wire REGFILE_SIM_reg_bank__abc_33898_n3219;
  wire REGFILE_SIM_reg_bank__abc_33898_n3220;
  wire REGFILE_SIM_reg_bank__abc_33898_n3221;
  wire REGFILE_SIM_reg_bank__abc_33898_n3223;
  wire REGFILE_SIM_reg_bank__abc_33898_n3224;
  wire REGFILE_SIM_reg_bank__abc_33898_n3225;
  wire REGFILE_SIM_reg_bank__abc_33898_n3227;
  wire REGFILE_SIM_reg_bank__abc_33898_n3228;
  wire REGFILE_SIM_reg_bank__abc_33898_n3229_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3231;
  wire REGFILE_SIM_reg_bank__abc_33898_n3232;
  wire REGFILE_SIM_reg_bank__abc_33898_n3233;
  wire REGFILE_SIM_reg_bank__abc_33898_n3235;
  wire REGFILE_SIM_reg_bank__abc_33898_n3236;
  wire REGFILE_SIM_reg_bank__abc_33898_n3237;
  wire REGFILE_SIM_reg_bank__abc_33898_n3239;
  wire REGFILE_SIM_reg_bank__abc_33898_n3240;
  wire REGFILE_SIM_reg_bank__abc_33898_n3241;
  wire REGFILE_SIM_reg_bank__abc_33898_n3243;
  wire REGFILE_SIM_reg_bank__abc_33898_n3244;
  wire REGFILE_SIM_reg_bank__abc_33898_n3245;
  wire REGFILE_SIM_reg_bank__abc_33898_n3247;
  wire REGFILE_SIM_reg_bank__abc_33898_n3248;
  wire REGFILE_SIM_reg_bank__abc_33898_n3249;
  wire REGFILE_SIM_reg_bank__abc_33898_n3251;
  wire REGFILE_SIM_reg_bank__abc_33898_n3252;
  wire REGFILE_SIM_reg_bank__abc_33898_n3253;
  wire REGFILE_SIM_reg_bank__abc_33898_n3255;
  wire REGFILE_SIM_reg_bank__abc_33898_n3256;
  wire REGFILE_SIM_reg_bank__abc_33898_n3257;
  wire REGFILE_SIM_reg_bank__abc_33898_n3259;
  wire REGFILE_SIM_reg_bank__abc_33898_n3260;
  wire REGFILE_SIM_reg_bank__abc_33898_n3261_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3263;
  wire REGFILE_SIM_reg_bank__abc_33898_n3264;
  wire REGFILE_SIM_reg_bank__abc_33898_n3265;
  wire REGFILE_SIM_reg_bank__abc_33898_n3267;
  wire REGFILE_SIM_reg_bank__abc_33898_n3268;
  wire REGFILE_SIM_reg_bank__abc_33898_n3269;
  wire REGFILE_SIM_reg_bank__abc_33898_n3271;
  wire REGFILE_SIM_reg_bank__abc_33898_n3272;
  wire REGFILE_SIM_reg_bank__abc_33898_n3273;
  wire REGFILE_SIM_reg_bank__abc_33898_n3275;
  wire REGFILE_SIM_reg_bank__abc_33898_n3276;
  wire REGFILE_SIM_reg_bank__abc_33898_n3277;
  wire REGFILE_SIM_reg_bank__abc_33898_n3279;
  wire REGFILE_SIM_reg_bank__abc_33898_n3280;
  wire REGFILE_SIM_reg_bank__abc_33898_n3281;
  wire REGFILE_SIM_reg_bank__abc_33898_n3283;
  wire REGFILE_SIM_reg_bank__abc_33898_n3284;
  wire REGFILE_SIM_reg_bank__abc_33898_n3285;
  wire REGFILE_SIM_reg_bank__abc_33898_n3287;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n3289;
  wire REGFILE_SIM_reg_bank__abc_33898_n3290;
  wire REGFILE_SIM_reg_bank__abc_33898_n3291;
  wire REGFILE_SIM_reg_bank__abc_33898_n3293_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3294;
  wire REGFILE_SIM_reg_bank__abc_33898_n3295;
  wire REGFILE_SIM_reg_bank__abc_33898_n3297;
  wire REGFILE_SIM_reg_bank__abc_33898_n3298;
  wire REGFILE_SIM_reg_bank__abc_33898_n3299;
  wire REGFILE_SIM_reg_bank__abc_33898_n3301;
  wire REGFILE_SIM_reg_bank__abc_33898_n3302;
  wire REGFILE_SIM_reg_bank__abc_33898_n3303;
  wire REGFILE_SIM_reg_bank__abc_33898_n3305;
  wire REGFILE_SIM_reg_bank__abc_33898_n3306;
  wire REGFILE_SIM_reg_bank__abc_33898_n3307;
  wire REGFILE_SIM_reg_bank__abc_33898_n3309;
  wire REGFILE_SIM_reg_bank__abc_33898_n3310;
  wire REGFILE_SIM_reg_bank__abc_33898_n3311;
  wire REGFILE_SIM_reg_bank__abc_33898_n3313;
  wire REGFILE_SIM_reg_bank__abc_33898_n3314;
  wire REGFILE_SIM_reg_bank__abc_33898_n3315;
  wire REGFILE_SIM_reg_bank__abc_33898_n3317;
  wire REGFILE_SIM_reg_bank__abc_33898_n3318;
  wire REGFILE_SIM_reg_bank__abc_33898_n3319;
  wire REGFILE_SIM_reg_bank__abc_33898_n3321;
  wire REGFILE_SIM_reg_bank__abc_33898_n3322;
  wire REGFILE_SIM_reg_bank__abc_33898_n3323;
  wire REGFILE_SIM_reg_bank__abc_33898_n3325_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3326;
  wire REGFILE_SIM_reg_bank__abc_33898_n3327;
  wire REGFILE_SIM_reg_bank__abc_33898_n3329;
  wire REGFILE_SIM_reg_bank__abc_33898_n3330;
  wire REGFILE_SIM_reg_bank__abc_33898_n3331;
  wire REGFILE_SIM_reg_bank__abc_33898_n3333;
  wire REGFILE_SIM_reg_bank__abc_33898_n3334;
  wire REGFILE_SIM_reg_bank__abc_33898_n3335;
  wire REGFILE_SIM_reg_bank__abc_33898_n3337;
  wire REGFILE_SIM_reg_bank__abc_33898_n3338;
  wire REGFILE_SIM_reg_bank__abc_33898_n3339;
  wire REGFILE_SIM_reg_bank__abc_33898_n3341;
  wire REGFILE_SIM_reg_bank__abc_33898_n3342;
  wire REGFILE_SIM_reg_bank__abc_33898_n3343;
  wire REGFILE_SIM_reg_bank__abc_33898_n3345;
  wire REGFILE_SIM_reg_bank__abc_33898_n3346;
  wire REGFILE_SIM_reg_bank__abc_33898_n3347;
  wire REGFILE_SIM_reg_bank__abc_33898_n3349;
  wire REGFILE_SIM_reg_bank__abc_33898_n3350;
  wire REGFILE_SIM_reg_bank__abc_33898_n3351;
  wire REGFILE_SIM_reg_bank__abc_33898_n3353;
  wire REGFILE_SIM_reg_bank__abc_33898_n3354;
  wire REGFILE_SIM_reg_bank__abc_33898_n3355;
  wire REGFILE_SIM_reg_bank__abc_33898_n3357_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3358;
  wire REGFILE_SIM_reg_bank__abc_33898_n3359;
  wire REGFILE_SIM_reg_bank__abc_33898_n3361;
  wire REGFILE_SIM_reg_bank__abc_33898_n3362;
  wire REGFILE_SIM_reg_bank__abc_33898_n3363;
  wire REGFILE_SIM_reg_bank__abc_33898_n3365;
  wire REGFILE_SIM_reg_bank__abc_33898_n3366;
  wire REGFILE_SIM_reg_bank__abc_33898_n3367;
  wire REGFILE_SIM_reg_bank__abc_33898_n3369;
  wire REGFILE_SIM_reg_bank__abc_33898_n3370;
  wire REGFILE_SIM_reg_bank__abc_33898_n3371;
  wire REGFILE_SIM_reg_bank__abc_33898_n3373;
  wire REGFILE_SIM_reg_bank__abc_33898_n3374;
  wire REGFILE_SIM_reg_bank__abc_33898_n3375;
  wire REGFILE_SIM_reg_bank__abc_33898_n3377;
  wire REGFILE_SIM_reg_bank__abc_33898_n3378;
  wire REGFILE_SIM_reg_bank__abc_33898_n3379;
  wire REGFILE_SIM_reg_bank__abc_33898_n3381;
  wire REGFILE_SIM_reg_bank__abc_33898_n3382;
  wire REGFILE_SIM_reg_bank__abc_33898_n3383;
  wire REGFILE_SIM_reg_bank__abc_33898_n3385;
  wire REGFILE_SIM_reg_bank__abc_33898_n3386;
  wire REGFILE_SIM_reg_bank__abc_33898_n3387;
  wire REGFILE_SIM_reg_bank__abc_33898_n3389_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3390;
  wire REGFILE_SIM_reg_bank__abc_33898_n3391;
  wire REGFILE_SIM_reg_bank__abc_33898_n3393;
  wire REGFILE_SIM_reg_bank__abc_33898_n3394;
  wire REGFILE_SIM_reg_bank__abc_33898_n3395;
  wire REGFILE_SIM_reg_bank__abc_33898_n3397;
  wire REGFILE_SIM_reg_bank__abc_33898_n3398;
  wire REGFILE_SIM_reg_bank__abc_33898_n3399;
  wire REGFILE_SIM_reg_bank__abc_33898_n3401;
  wire REGFILE_SIM_reg_bank__abc_33898_n3402;
  wire REGFILE_SIM_reg_bank__abc_33898_n3403;
  wire REGFILE_SIM_reg_bank__abc_33898_n3405;
  wire REGFILE_SIM_reg_bank__abc_33898_n3406;
  wire REGFILE_SIM_reg_bank__abc_33898_n3407;
  wire REGFILE_SIM_reg_bank__abc_33898_n3409;
  wire REGFILE_SIM_reg_bank__abc_33898_n3410;
  wire REGFILE_SIM_reg_bank__abc_33898_n3411;
  wire REGFILE_SIM_reg_bank__abc_33898_n3413;
  wire REGFILE_SIM_reg_bank__abc_33898_n3414;
  wire REGFILE_SIM_reg_bank__abc_33898_n3415;
  wire REGFILE_SIM_reg_bank__abc_33898_n3417;
  wire REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3418;
  wire REGFILE_SIM_reg_bank__abc_33898_n3419;
  wire REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3420;
  wire REGFILE_SIM_reg_bank__abc_33898_n3422;
  wire REGFILE_SIM_reg_bank__abc_33898_n3423;
  wire REGFILE_SIM_reg_bank__abc_33898_n3425;
  wire REGFILE_SIM_reg_bank__abc_33898_n3426;
  wire REGFILE_SIM_reg_bank__abc_33898_n3428;
  wire REGFILE_SIM_reg_bank__abc_33898_n3429;
  wire REGFILE_SIM_reg_bank__abc_33898_n3431;
  wire REGFILE_SIM_reg_bank__abc_33898_n3432;
  wire REGFILE_SIM_reg_bank__abc_33898_n3434;
  wire REGFILE_SIM_reg_bank__abc_33898_n3435;
  wire REGFILE_SIM_reg_bank__abc_33898_n3437;
  wire REGFILE_SIM_reg_bank__abc_33898_n3438;
  wire REGFILE_SIM_reg_bank__abc_33898_n3440;
  wire REGFILE_SIM_reg_bank__abc_33898_n3441;
  wire REGFILE_SIM_reg_bank__abc_33898_n3443;
  wire REGFILE_SIM_reg_bank__abc_33898_n3444;
  wire REGFILE_SIM_reg_bank__abc_33898_n3446;
  wire REGFILE_SIM_reg_bank__abc_33898_n3447;
  wire REGFILE_SIM_reg_bank__abc_33898_n3449;
  wire REGFILE_SIM_reg_bank__abc_33898_n3450;
  wire REGFILE_SIM_reg_bank__abc_33898_n3452;
  wire REGFILE_SIM_reg_bank__abc_33898_n3453_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3455;
  wire REGFILE_SIM_reg_bank__abc_33898_n3456;
  wire REGFILE_SIM_reg_bank__abc_33898_n3458;
  wire REGFILE_SIM_reg_bank__abc_33898_n3459;
  wire REGFILE_SIM_reg_bank__abc_33898_n3461;
  wire REGFILE_SIM_reg_bank__abc_33898_n3462;
  wire REGFILE_SIM_reg_bank__abc_33898_n3464;
  wire REGFILE_SIM_reg_bank__abc_33898_n3465;
  wire REGFILE_SIM_reg_bank__abc_33898_n3467;
  wire REGFILE_SIM_reg_bank__abc_33898_n3468;
  wire REGFILE_SIM_reg_bank__abc_33898_n3470;
  wire REGFILE_SIM_reg_bank__abc_33898_n3471;
  wire REGFILE_SIM_reg_bank__abc_33898_n3473;
  wire REGFILE_SIM_reg_bank__abc_33898_n3474;
  wire REGFILE_SIM_reg_bank__abc_33898_n3476;
  wire REGFILE_SIM_reg_bank__abc_33898_n3477;
  wire REGFILE_SIM_reg_bank__abc_33898_n3479;
  wire REGFILE_SIM_reg_bank__abc_33898_n3480;
  wire REGFILE_SIM_reg_bank__abc_33898_n3482;
  wire REGFILE_SIM_reg_bank__abc_33898_n3483;
  wire REGFILE_SIM_reg_bank__abc_33898_n3485_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3486;
  wire REGFILE_SIM_reg_bank__abc_33898_n3488;
  wire REGFILE_SIM_reg_bank__abc_33898_n3489;
  wire REGFILE_SIM_reg_bank__abc_33898_n3491;
  wire REGFILE_SIM_reg_bank__abc_33898_n3492;
  wire REGFILE_SIM_reg_bank__abc_33898_n3494;
  wire REGFILE_SIM_reg_bank__abc_33898_n3495;
  wire REGFILE_SIM_reg_bank__abc_33898_n3497;
  wire REGFILE_SIM_reg_bank__abc_33898_n3498;
  wire REGFILE_SIM_reg_bank__abc_33898_n3500;
  wire REGFILE_SIM_reg_bank__abc_33898_n3501;
  wire REGFILE_SIM_reg_bank__abc_33898_n3503;
  wire REGFILE_SIM_reg_bank__abc_33898_n3504;
  wire REGFILE_SIM_reg_bank__abc_33898_n3506;
  wire REGFILE_SIM_reg_bank__abc_33898_n3507;
  wire REGFILE_SIM_reg_bank__abc_33898_n3509;
  wire REGFILE_SIM_reg_bank__abc_33898_n3510;
  wire REGFILE_SIM_reg_bank__abc_33898_n3512;
  wire REGFILE_SIM_reg_bank__abc_33898_n3513;
  wire REGFILE_SIM_reg_bank__abc_33898_n3515;
  wire REGFILE_SIM_reg_bank__abc_33898_n3516;
  wire REGFILE_SIM_reg_bank__abc_33898_n3517_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3518;
  wire REGFILE_SIM_reg_bank__abc_33898_n3519;
  wire REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3520;
  wire REGFILE_SIM_reg_bank__abc_33898_n3522;
  wire REGFILE_SIM_reg_bank__abc_33898_n3523;
  wire REGFILE_SIM_reg_bank__abc_33898_n3525;
  wire REGFILE_SIM_reg_bank__abc_33898_n3526;
  wire REGFILE_SIM_reg_bank__abc_33898_n3528;
  wire REGFILE_SIM_reg_bank__abc_33898_n3529;
  wire REGFILE_SIM_reg_bank__abc_33898_n3531;
  wire REGFILE_SIM_reg_bank__abc_33898_n3532;
  wire REGFILE_SIM_reg_bank__abc_33898_n3534;
  wire REGFILE_SIM_reg_bank__abc_33898_n3535;
  wire REGFILE_SIM_reg_bank__abc_33898_n3537;
  wire REGFILE_SIM_reg_bank__abc_33898_n3538;
  wire REGFILE_SIM_reg_bank__abc_33898_n3540;
  wire REGFILE_SIM_reg_bank__abc_33898_n3541;
  wire REGFILE_SIM_reg_bank__abc_33898_n3543;
  wire REGFILE_SIM_reg_bank__abc_33898_n3544;
  wire REGFILE_SIM_reg_bank__abc_33898_n3546;
  wire REGFILE_SIM_reg_bank__abc_33898_n3547;
  wire REGFILE_SIM_reg_bank__abc_33898_n3549_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3550;
  wire REGFILE_SIM_reg_bank__abc_33898_n3552;
  wire REGFILE_SIM_reg_bank__abc_33898_n3553;
  wire REGFILE_SIM_reg_bank__abc_33898_n3555;
  wire REGFILE_SIM_reg_bank__abc_33898_n3556;
  wire REGFILE_SIM_reg_bank__abc_33898_n3558;
  wire REGFILE_SIM_reg_bank__abc_33898_n3559;
  wire REGFILE_SIM_reg_bank__abc_33898_n3561;
  wire REGFILE_SIM_reg_bank__abc_33898_n3562;
  wire REGFILE_SIM_reg_bank__abc_33898_n3564;
  wire REGFILE_SIM_reg_bank__abc_33898_n3565;
  wire REGFILE_SIM_reg_bank__abc_33898_n3567;
  wire REGFILE_SIM_reg_bank__abc_33898_n3568;
  wire REGFILE_SIM_reg_bank__abc_33898_n3570;
  wire REGFILE_SIM_reg_bank__abc_33898_n3571;
  wire REGFILE_SIM_reg_bank__abc_33898_n3573;
  wire REGFILE_SIM_reg_bank__abc_33898_n3574;
  wire REGFILE_SIM_reg_bank__abc_33898_n3576;
  wire REGFILE_SIM_reg_bank__abc_33898_n3577;
  wire REGFILE_SIM_reg_bank__abc_33898_n3579;
  wire REGFILE_SIM_reg_bank__abc_33898_n3580;
  wire REGFILE_SIM_reg_bank__abc_33898_n3582;
  wire REGFILE_SIM_reg_bank__abc_33898_n3583;
  wire REGFILE_SIM_reg_bank__abc_33898_n3585;
  wire REGFILE_SIM_reg_bank__abc_33898_n3586;
  wire REGFILE_SIM_reg_bank__abc_33898_n3588;
  wire REGFILE_SIM_reg_bank__abc_33898_n3589;
  wire REGFILE_SIM_reg_bank__abc_33898_n3591;
  wire REGFILE_SIM_reg_bank__abc_33898_n3592;
  wire REGFILE_SIM_reg_bank__abc_33898_n3594;
  wire REGFILE_SIM_reg_bank__abc_33898_n3595;
  wire REGFILE_SIM_reg_bank__abc_33898_n3597;
  wire REGFILE_SIM_reg_bank__abc_33898_n3598;
  wire REGFILE_SIM_reg_bank__abc_33898_n3600;
  wire REGFILE_SIM_reg_bank__abc_33898_n3601;
  wire REGFILE_SIM_reg_bank__abc_33898_n3603;
  wire REGFILE_SIM_reg_bank__abc_33898_n3604;
  wire REGFILE_SIM_reg_bank__abc_33898_n3606;
  wire REGFILE_SIM_reg_bank__abc_33898_n3607;
  wire REGFILE_SIM_reg_bank__abc_33898_n3609;
  wire REGFILE_SIM_reg_bank__abc_33898_n3610;
  wire REGFILE_SIM_reg_bank__abc_33898_n3612;
  wire REGFILE_SIM_reg_bank__abc_33898_n3613_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3615;
  wire REGFILE_SIM_reg_bank__abc_33898_n3616;
  wire REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3617;
  wire REGFILE_SIM_reg_bank__abc_33898_n3618;
  wire REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3619;
  wire REGFILE_SIM_reg_bank__abc_33898_n3621;
  wire REGFILE_SIM_reg_bank__abc_33898_n3622;
  wire REGFILE_SIM_reg_bank__abc_33898_n3624;
  wire REGFILE_SIM_reg_bank__abc_33898_n3625;
  wire REGFILE_SIM_reg_bank__abc_33898_n3627;
  wire REGFILE_SIM_reg_bank__abc_33898_n3628;
  wire REGFILE_SIM_reg_bank__abc_33898_n3630;
  wire REGFILE_SIM_reg_bank__abc_33898_n3631;
  wire REGFILE_SIM_reg_bank__abc_33898_n3633;
  wire REGFILE_SIM_reg_bank__abc_33898_n3634;
  wire REGFILE_SIM_reg_bank__abc_33898_n3636;
  wire REGFILE_SIM_reg_bank__abc_33898_n3637;
  wire REGFILE_SIM_reg_bank__abc_33898_n3639;
  wire REGFILE_SIM_reg_bank__abc_33898_n3640;
  wire REGFILE_SIM_reg_bank__abc_33898_n3642;
  wire REGFILE_SIM_reg_bank__abc_33898_n3643;
  wire REGFILE_SIM_reg_bank__abc_33898_n3645_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3646;
  wire REGFILE_SIM_reg_bank__abc_33898_n3648;
  wire REGFILE_SIM_reg_bank__abc_33898_n3649;
  wire REGFILE_SIM_reg_bank__abc_33898_n3651;
  wire REGFILE_SIM_reg_bank__abc_33898_n3652;
  wire REGFILE_SIM_reg_bank__abc_33898_n3654;
  wire REGFILE_SIM_reg_bank__abc_33898_n3655;
  wire REGFILE_SIM_reg_bank__abc_33898_n3657;
  wire REGFILE_SIM_reg_bank__abc_33898_n3658;
  wire REGFILE_SIM_reg_bank__abc_33898_n3660;
  wire REGFILE_SIM_reg_bank__abc_33898_n3661;
  wire REGFILE_SIM_reg_bank__abc_33898_n3663;
  wire REGFILE_SIM_reg_bank__abc_33898_n3664;
  wire REGFILE_SIM_reg_bank__abc_33898_n3666;
  wire REGFILE_SIM_reg_bank__abc_33898_n3667;
  wire REGFILE_SIM_reg_bank__abc_33898_n3669;
  wire REGFILE_SIM_reg_bank__abc_33898_n3670;
  wire REGFILE_SIM_reg_bank__abc_33898_n3672;
  wire REGFILE_SIM_reg_bank__abc_33898_n3673;
  wire REGFILE_SIM_reg_bank__abc_33898_n3675;
  wire REGFILE_SIM_reg_bank__abc_33898_n3676;
  wire REGFILE_SIM_reg_bank__abc_33898_n3678;
  wire REGFILE_SIM_reg_bank__abc_33898_n3679;
  wire REGFILE_SIM_reg_bank__abc_33898_n3681;
  wire REGFILE_SIM_reg_bank__abc_33898_n3682;
  wire REGFILE_SIM_reg_bank__abc_33898_n3684;
  wire REGFILE_SIM_reg_bank__abc_33898_n3685;
  wire REGFILE_SIM_reg_bank__abc_33898_n3687;
  wire REGFILE_SIM_reg_bank__abc_33898_n3688;
  wire REGFILE_SIM_reg_bank__abc_33898_n3690;
  wire REGFILE_SIM_reg_bank__abc_33898_n3691;
  wire REGFILE_SIM_reg_bank__abc_33898_n3693;
  wire REGFILE_SIM_reg_bank__abc_33898_n3694;
  wire REGFILE_SIM_reg_bank__abc_33898_n3696;
  wire REGFILE_SIM_reg_bank__abc_33898_n3697;
  wire REGFILE_SIM_reg_bank__abc_33898_n3699;
  wire REGFILE_SIM_reg_bank__abc_33898_n3700;
  wire REGFILE_SIM_reg_bank__abc_33898_n3702;
  wire REGFILE_SIM_reg_bank__abc_33898_n3703;
  wire REGFILE_SIM_reg_bank__abc_33898_n3705;
  wire REGFILE_SIM_reg_bank__abc_33898_n3706;
  wire REGFILE_SIM_reg_bank__abc_33898_n3708;
  wire REGFILE_SIM_reg_bank__abc_33898_n3709_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3711;
  wire REGFILE_SIM_reg_bank__abc_33898_n3712;
  wire REGFILE_SIM_reg_bank__abc_33898_n3714;
  wire REGFILE_SIM_reg_bank__abc_33898_n3715;
  wire REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3716;
  wire REGFILE_SIM_reg_bank__abc_33898_n3717;
  wire REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3718;
  wire REGFILE_SIM_reg_bank__abc_33898_n3720;
  wire REGFILE_SIM_reg_bank__abc_33898_n3721;
  wire REGFILE_SIM_reg_bank__abc_33898_n3723;
  wire REGFILE_SIM_reg_bank__abc_33898_n3724;
  wire REGFILE_SIM_reg_bank__abc_33898_n3726;
  wire REGFILE_SIM_reg_bank__abc_33898_n3727;
  wire REGFILE_SIM_reg_bank__abc_33898_n3729;
  wire REGFILE_SIM_reg_bank__abc_33898_n3730;
  wire REGFILE_SIM_reg_bank__abc_33898_n3732;
  wire REGFILE_SIM_reg_bank__abc_33898_n3733;
  wire REGFILE_SIM_reg_bank__abc_33898_n3735;
  wire REGFILE_SIM_reg_bank__abc_33898_n3736;
  wire REGFILE_SIM_reg_bank__abc_33898_n3738;
  wire REGFILE_SIM_reg_bank__abc_33898_n3739;
  wire REGFILE_SIM_reg_bank__abc_33898_n3741_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3742;
  wire REGFILE_SIM_reg_bank__abc_33898_n3744;
  wire REGFILE_SIM_reg_bank__abc_33898_n3745;
  wire REGFILE_SIM_reg_bank__abc_33898_n3747;
  wire REGFILE_SIM_reg_bank__abc_33898_n3748;
  wire REGFILE_SIM_reg_bank__abc_33898_n3750;
  wire REGFILE_SIM_reg_bank__abc_33898_n3751;
  wire REGFILE_SIM_reg_bank__abc_33898_n3753;
  wire REGFILE_SIM_reg_bank__abc_33898_n3754;
  wire REGFILE_SIM_reg_bank__abc_33898_n3756;
  wire REGFILE_SIM_reg_bank__abc_33898_n3757;
  wire REGFILE_SIM_reg_bank__abc_33898_n3759;
  wire REGFILE_SIM_reg_bank__abc_33898_n3760;
  wire REGFILE_SIM_reg_bank__abc_33898_n3762;
  wire REGFILE_SIM_reg_bank__abc_33898_n3763;
  wire REGFILE_SIM_reg_bank__abc_33898_n3765;
  wire REGFILE_SIM_reg_bank__abc_33898_n3766;
  wire REGFILE_SIM_reg_bank__abc_33898_n3768;
  wire REGFILE_SIM_reg_bank__abc_33898_n3769;
  wire REGFILE_SIM_reg_bank__abc_33898_n3771;
  wire REGFILE_SIM_reg_bank__abc_33898_n3772;
  wire REGFILE_SIM_reg_bank__abc_33898_n3774;
  wire REGFILE_SIM_reg_bank__abc_33898_n3775;
  wire REGFILE_SIM_reg_bank__abc_33898_n3777;
  wire REGFILE_SIM_reg_bank__abc_33898_n3778;
  wire REGFILE_SIM_reg_bank__abc_33898_n3780;
  wire REGFILE_SIM_reg_bank__abc_33898_n3781;
  wire REGFILE_SIM_reg_bank__abc_33898_n3783;
  wire REGFILE_SIM_reg_bank__abc_33898_n3784;
  wire REGFILE_SIM_reg_bank__abc_33898_n3786;
  wire REGFILE_SIM_reg_bank__abc_33898_n3787;
  wire REGFILE_SIM_reg_bank__abc_33898_n3789;
  wire REGFILE_SIM_reg_bank__abc_33898_n3790;
  wire REGFILE_SIM_reg_bank__abc_33898_n3792;
  wire REGFILE_SIM_reg_bank__abc_33898_n3793;
  wire REGFILE_SIM_reg_bank__abc_33898_n3795;
  wire REGFILE_SIM_reg_bank__abc_33898_n3796;
  wire REGFILE_SIM_reg_bank__abc_33898_n3798;
  wire REGFILE_SIM_reg_bank__abc_33898_n3799;
  wire REGFILE_SIM_reg_bank__abc_33898_n3801;
  wire REGFILE_SIM_reg_bank__abc_33898_n3802;
  wire REGFILE_SIM_reg_bank__abc_33898_n3804;
  wire REGFILE_SIM_reg_bank__abc_33898_n3805_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3807;
  wire REGFILE_SIM_reg_bank__abc_33898_n3808;
  wire REGFILE_SIM_reg_bank__abc_33898_n3810;
  wire REGFILE_SIM_reg_bank__abc_33898_n3811;
  wire REGFILE_SIM_reg_bank__abc_33898_n3813;
  wire REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3814;
  wire REGFILE_SIM_reg_bank__abc_33898_n3815;
  wire REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3816;
  wire REGFILE_SIM_reg_bank__abc_33898_n3818;
  wire REGFILE_SIM_reg_bank__abc_33898_n3819;
  wire REGFILE_SIM_reg_bank__abc_33898_n3821;
  wire REGFILE_SIM_reg_bank__abc_33898_n3822;
  wire REGFILE_SIM_reg_bank__abc_33898_n3824;
  wire REGFILE_SIM_reg_bank__abc_33898_n3825;
  wire REGFILE_SIM_reg_bank__abc_33898_n3827;
  wire REGFILE_SIM_reg_bank__abc_33898_n3828;
  wire REGFILE_SIM_reg_bank__abc_33898_n3830;
  wire REGFILE_SIM_reg_bank__abc_33898_n3831;
  wire REGFILE_SIM_reg_bank__abc_33898_n3833;
  wire REGFILE_SIM_reg_bank__abc_33898_n3834;
  wire REGFILE_SIM_reg_bank__abc_33898_n3836;
  wire REGFILE_SIM_reg_bank__abc_33898_n3837_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3839;
  wire REGFILE_SIM_reg_bank__abc_33898_n3840;
  wire REGFILE_SIM_reg_bank__abc_33898_n3842;
  wire REGFILE_SIM_reg_bank__abc_33898_n3843;
  wire REGFILE_SIM_reg_bank__abc_33898_n3845;
  wire REGFILE_SIM_reg_bank__abc_33898_n3846;
  wire REGFILE_SIM_reg_bank__abc_33898_n3848;
  wire REGFILE_SIM_reg_bank__abc_33898_n3849;
  wire REGFILE_SIM_reg_bank__abc_33898_n3851;
  wire REGFILE_SIM_reg_bank__abc_33898_n3852;
  wire REGFILE_SIM_reg_bank__abc_33898_n3854;
  wire REGFILE_SIM_reg_bank__abc_33898_n3855;
  wire REGFILE_SIM_reg_bank__abc_33898_n3857;
  wire REGFILE_SIM_reg_bank__abc_33898_n3858;
  wire REGFILE_SIM_reg_bank__abc_33898_n3860;
  wire REGFILE_SIM_reg_bank__abc_33898_n3861;
  wire REGFILE_SIM_reg_bank__abc_33898_n3863;
  wire REGFILE_SIM_reg_bank__abc_33898_n3864;
  wire REGFILE_SIM_reg_bank__abc_33898_n3866;
  wire REGFILE_SIM_reg_bank__abc_33898_n3867;
  wire REGFILE_SIM_reg_bank__abc_33898_n3869_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3870;
  wire REGFILE_SIM_reg_bank__abc_33898_n3872;
  wire REGFILE_SIM_reg_bank__abc_33898_n3873;
  wire REGFILE_SIM_reg_bank__abc_33898_n3875;
  wire REGFILE_SIM_reg_bank__abc_33898_n3876;
  wire REGFILE_SIM_reg_bank__abc_33898_n3878;
  wire REGFILE_SIM_reg_bank__abc_33898_n3879;
  wire REGFILE_SIM_reg_bank__abc_33898_n3881;
  wire REGFILE_SIM_reg_bank__abc_33898_n3882;
  wire REGFILE_SIM_reg_bank__abc_33898_n3884;
  wire REGFILE_SIM_reg_bank__abc_33898_n3885;
  wire REGFILE_SIM_reg_bank__abc_33898_n3887;
  wire REGFILE_SIM_reg_bank__abc_33898_n3888;
  wire REGFILE_SIM_reg_bank__abc_33898_n3890;
  wire REGFILE_SIM_reg_bank__abc_33898_n3891;
  wire REGFILE_SIM_reg_bank__abc_33898_n3893;
  wire REGFILE_SIM_reg_bank__abc_33898_n3894;
  wire REGFILE_SIM_reg_bank__abc_33898_n3896;
  wire REGFILE_SIM_reg_bank__abc_33898_n3897;
  wire REGFILE_SIM_reg_bank__abc_33898_n3899;
  wire REGFILE_SIM_reg_bank__abc_33898_n3900;
  wire REGFILE_SIM_reg_bank__abc_33898_n3902;
  wire REGFILE_SIM_reg_bank__abc_33898_n3903;
  wire REGFILE_SIM_reg_bank__abc_33898_n3905;
  wire REGFILE_SIM_reg_bank__abc_33898_n3906;
  wire REGFILE_SIM_reg_bank__abc_33898_n3908;
  wire REGFILE_SIM_reg_bank__abc_33898_n3909;
  wire REGFILE_SIM_reg_bank__abc_33898_n3911;
  wire REGFILE_SIM_reg_bank__abc_33898_n3912;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n3914;
  wire REGFILE_SIM_reg_bank__abc_33898_n3915;
  wire REGFILE_SIM_reg_bank__abc_33898_n3916;
  wire REGFILE_SIM_reg_bank__abc_33898_n3918;
  wire REGFILE_SIM_reg_bank__abc_33898_n3919;
  wire REGFILE_SIM_reg_bank__abc_33898_n3920;
  wire REGFILE_SIM_reg_bank__abc_33898_n3922;
  wire REGFILE_SIM_reg_bank__abc_33898_n3923;
  wire REGFILE_SIM_reg_bank__abc_33898_n3924;
  wire REGFILE_SIM_reg_bank__abc_33898_n3926;
  wire REGFILE_SIM_reg_bank__abc_33898_n3927;
  wire REGFILE_SIM_reg_bank__abc_33898_n3928;
  wire REGFILE_SIM_reg_bank__abc_33898_n3930;
  wire REGFILE_SIM_reg_bank__abc_33898_n3931;
  wire REGFILE_SIM_reg_bank__abc_33898_n3932;
  wire REGFILE_SIM_reg_bank__abc_33898_n3934;
  wire REGFILE_SIM_reg_bank__abc_33898_n3935;
  wire REGFILE_SIM_reg_bank__abc_33898_n3936;
  wire REGFILE_SIM_reg_bank__abc_33898_n3938;
  wire REGFILE_SIM_reg_bank__abc_33898_n3939;
  wire REGFILE_SIM_reg_bank__abc_33898_n3940;
  wire REGFILE_SIM_reg_bank__abc_33898_n3942;
  wire REGFILE_SIM_reg_bank__abc_33898_n3943;
  wire REGFILE_SIM_reg_bank__abc_33898_n3944;
  wire REGFILE_SIM_reg_bank__abc_33898_n3946;
  wire REGFILE_SIM_reg_bank__abc_33898_n3947;
  wire REGFILE_SIM_reg_bank__abc_33898_n3948;
  wire REGFILE_SIM_reg_bank__abc_33898_n3950;
  wire REGFILE_SIM_reg_bank__abc_33898_n3951;
  wire REGFILE_SIM_reg_bank__abc_33898_n3952;
  wire REGFILE_SIM_reg_bank__abc_33898_n3954;
  wire REGFILE_SIM_reg_bank__abc_33898_n3955;
  wire REGFILE_SIM_reg_bank__abc_33898_n3956;
  wire REGFILE_SIM_reg_bank__abc_33898_n3958;
  wire REGFILE_SIM_reg_bank__abc_33898_n3959;
  wire REGFILE_SIM_reg_bank__abc_33898_n3960;
  wire REGFILE_SIM_reg_bank__abc_33898_n3962;
  wire REGFILE_SIM_reg_bank__abc_33898_n3963;
  wire REGFILE_SIM_reg_bank__abc_33898_n3964;
  wire REGFILE_SIM_reg_bank__abc_33898_n3966;
  wire REGFILE_SIM_reg_bank__abc_33898_n3967;
  wire REGFILE_SIM_reg_bank__abc_33898_n3968;
  wire REGFILE_SIM_reg_bank__abc_33898_n3970;
  wire REGFILE_SIM_reg_bank__abc_33898_n3971;
  wire REGFILE_SIM_reg_bank__abc_33898_n3972;
  wire REGFILE_SIM_reg_bank__abc_33898_n3974;
  wire REGFILE_SIM_reg_bank__abc_33898_n3975;
  wire REGFILE_SIM_reg_bank__abc_33898_n3976;
  wire REGFILE_SIM_reg_bank__abc_33898_n3978;
  wire REGFILE_SIM_reg_bank__abc_33898_n3979;
  wire REGFILE_SIM_reg_bank__abc_33898_n3980;
  wire REGFILE_SIM_reg_bank__abc_33898_n3982;
  wire REGFILE_SIM_reg_bank__abc_33898_n3983;
  wire REGFILE_SIM_reg_bank__abc_33898_n3984;
  wire REGFILE_SIM_reg_bank__abc_33898_n3986;
  wire REGFILE_SIM_reg_bank__abc_33898_n3987;
  wire REGFILE_SIM_reg_bank__abc_33898_n3988;
  wire REGFILE_SIM_reg_bank__abc_33898_n3990;
  wire REGFILE_SIM_reg_bank__abc_33898_n3991;
  wire REGFILE_SIM_reg_bank__abc_33898_n3992;
  wire REGFILE_SIM_reg_bank__abc_33898_n3994;
  wire REGFILE_SIM_reg_bank__abc_33898_n3995;
  wire REGFILE_SIM_reg_bank__abc_33898_n3996;
  wire REGFILE_SIM_reg_bank__abc_33898_n3998;
  wire REGFILE_SIM_reg_bank__abc_33898_n3999;
  wire REGFILE_SIM_reg_bank__abc_33898_n4000;
  wire REGFILE_SIM_reg_bank__abc_33898_n4002;
  wire REGFILE_SIM_reg_bank__abc_33898_n4003;
  wire REGFILE_SIM_reg_bank__abc_33898_n4004;
  wire REGFILE_SIM_reg_bank__abc_33898_n4006;
  wire REGFILE_SIM_reg_bank__abc_33898_n4007;
  wire REGFILE_SIM_reg_bank__abc_33898_n4008;
  wire REGFILE_SIM_reg_bank__abc_33898_n4010;
  wire REGFILE_SIM_reg_bank__abc_33898_n4011;
  wire REGFILE_SIM_reg_bank__abc_33898_n4012;
  wire REGFILE_SIM_reg_bank__abc_33898_n4014;
  wire REGFILE_SIM_reg_bank__abc_33898_n4015;
  wire REGFILE_SIM_reg_bank__abc_33898_n4016;
  wire REGFILE_SIM_reg_bank__abc_33898_n4018;
  wire REGFILE_SIM_reg_bank__abc_33898_n4019;
  wire REGFILE_SIM_reg_bank__abc_33898_n4020;
  wire REGFILE_SIM_reg_bank__abc_33898_n4022;
  wire REGFILE_SIM_reg_bank__abc_33898_n4023;
  wire REGFILE_SIM_reg_bank__abc_33898_n4024;
  wire REGFILE_SIM_reg_bank__abc_33898_n4026;
  wire REGFILE_SIM_reg_bank__abc_33898_n4027;
  wire REGFILE_SIM_reg_bank__abc_33898_n4028;
  wire REGFILE_SIM_reg_bank__abc_33898_n4030;
  wire REGFILE_SIM_reg_bank__abc_33898_n4031;
  wire REGFILE_SIM_reg_bank__abc_33898_n4032;
  wire REGFILE_SIM_reg_bank__abc_33898_n4034;
  wire REGFILE_SIM_reg_bank__abc_33898_n4035;
  wire REGFILE_SIM_reg_bank__abc_33898_n4036;
  wire REGFILE_SIM_reg_bank__abc_33898_n4038;
  wire REGFILE_SIM_reg_bank__abc_33898_n4039;
  wire REGFILE_SIM_reg_bank__abc_33898_n4040;
  wire REGFILE_SIM_reg_bank__abc_33898_n4042;
  wire REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4043;
  wire REGFILE_SIM_reg_bank__abc_33898_n4044;
  wire REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4045;
  wire REGFILE_SIM_reg_bank__abc_33898_n4047;
  wire REGFILE_SIM_reg_bank__abc_33898_n4048;
  wire REGFILE_SIM_reg_bank__abc_33898_n4050;
  wire REGFILE_SIM_reg_bank__abc_33898_n4051;
  wire REGFILE_SIM_reg_bank__abc_33898_n4053;
  wire REGFILE_SIM_reg_bank__abc_33898_n4054;
  wire REGFILE_SIM_reg_bank__abc_33898_n4056;
  wire REGFILE_SIM_reg_bank__abc_33898_n4057;
  wire REGFILE_SIM_reg_bank__abc_33898_n4059;
  wire REGFILE_SIM_reg_bank__abc_33898_n4060;
  wire REGFILE_SIM_reg_bank__abc_33898_n4062;
  wire REGFILE_SIM_reg_bank__abc_33898_n4063;
  wire REGFILE_SIM_reg_bank__abc_33898_n4065;
  wire REGFILE_SIM_reg_bank__abc_33898_n4066;
  wire REGFILE_SIM_reg_bank__abc_33898_n4068;
  wire REGFILE_SIM_reg_bank__abc_33898_n4069;
  wire REGFILE_SIM_reg_bank__abc_33898_n4071;
  wire REGFILE_SIM_reg_bank__abc_33898_n4072;
  wire REGFILE_SIM_reg_bank__abc_33898_n4074;
  wire REGFILE_SIM_reg_bank__abc_33898_n4075;
  wire REGFILE_SIM_reg_bank__abc_33898_n4077;
  wire REGFILE_SIM_reg_bank__abc_33898_n4078;
  wire REGFILE_SIM_reg_bank__abc_33898_n4080;
  wire REGFILE_SIM_reg_bank__abc_33898_n4081;
  wire REGFILE_SIM_reg_bank__abc_33898_n4083;
  wire REGFILE_SIM_reg_bank__abc_33898_n4084;
  wire REGFILE_SIM_reg_bank__abc_33898_n4086;
  wire REGFILE_SIM_reg_bank__abc_33898_n4087;
  wire REGFILE_SIM_reg_bank__abc_33898_n4089;
  wire REGFILE_SIM_reg_bank__abc_33898_n4090;
  wire REGFILE_SIM_reg_bank__abc_33898_n4092;
  wire REGFILE_SIM_reg_bank__abc_33898_n4093_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4095;
  wire REGFILE_SIM_reg_bank__abc_33898_n4096;
  wire REGFILE_SIM_reg_bank__abc_33898_n4098;
  wire REGFILE_SIM_reg_bank__abc_33898_n4099;
  wire REGFILE_SIM_reg_bank__abc_33898_n4101;
  wire REGFILE_SIM_reg_bank__abc_33898_n4102;
  wire REGFILE_SIM_reg_bank__abc_33898_n4104;
  wire REGFILE_SIM_reg_bank__abc_33898_n4105;
  wire REGFILE_SIM_reg_bank__abc_33898_n4107;
  wire REGFILE_SIM_reg_bank__abc_33898_n4108;
  wire REGFILE_SIM_reg_bank__abc_33898_n4110;
  wire REGFILE_SIM_reg_bank__abc_33898_n4111;
  wire REGFILE_SIM_reg_bank__abc_33898_n4113;
  wire REGFILE_SIM_reg_bank__abc_33898_n4114;
  wire REGFILE_SIM_reg_bank__abc_33898_n4116;
  wire REGFILE_SIM_reg_bank__abc_33898_n4117;
  wire REGFILE_SIM_reg_bank__abc_33898_n4119;
  wire REGFILE_SIM_reg_bank__abc_33898_n4120;
  wire REGFILE_SIM_reg_bank__abc_33898_n4122;
  wire REGFILE_SIM_reg_bank__abc_33898_n4123;
  wire REGFILE_SIM_reg_bank__abc_33898_n4125_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4126;
  wire REGFILE_SIM_reg_bank__abc_33898_n4128;
  wire REGFILE_SIM_reg_bank__abc_33898_n4129;
  wire REGFILE_SIM_reg_bank__abc_33898_n4131;
  wire REGFILE_SIM_reg_bank__abc_33898_n4132;
  wire REGFILE_SIM_reg_bank__abc_33898_n4134;
  wire REGFILE_SIM_reg_bank__abc_33898_n4135;
  wire REGFILE_SIM_reg_bank__abc_33898_n4137;
  wire REGFILE_SIM_reg_bank__abc_33898_n4138;
  wire REGFILE_SIM_reg_bank__abc_33898_n4140;
  wire REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4141;
  wire REGFILE_SIM_reg_bank__abc_33898_n4142;
  wire REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4143;
  wire REGFILE_SIM_reg_bank__abc_33898_n4145;
  wire REGFILE_SIM_reg_bank__abc_33898_n4146;
  wire REGFILE_SIM_reg_bank__abc_33898_n4148;
  wire REGFILE_SIM_reg_bank__abc_33898_n4149;
  wire REGFILE_SIM_reg_bank__abc_33898_n4151;
  wire REGFILE_SIM_reg_bank__abc_33898_n4152;
  wire REGFILE_SIM_reg_bank__abc_33898_n4154;
  wire REGFILE_SIM_reg_bank__abc_33898_n4155;
  wire REGFILE_SIM_reg_bank__abc_33898_n4157_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4158;
  wire REGFILE_SIM_reg_bank__abc_33898_n4160;
  wire REGFILE_SIM_reg_bank__abc_33898_n4161;
  wire REGFILE_SIM_reg_bank__abc_33898_n4163;
  wire REGFILE_SIM_reg_bank__abc_33898_n4164;
  wire REGFILE_SIM_reg_bank__abc_33898_n4166;
  wire REGFILE_SIM_reg_bank__abc_33898_n4167;
  wire REGFILE_SIM_reg_bank__abc_33898_n4169;
  wire REGFILE_SIM_reg_bank__abc_33898_n4170;
  wire REGFILE_SIM_reg_bank__abc_33898_n4172;
  wire REGFILE_SIM_reg_bank__abc_33898_n4173;
  wire REGFILE_SIM_reg_bank__abc_33898_n4175;
  wire REGFILE_SIM_reg_bank__abc_33898_n4176;
  wire REGFILE_SIM_reg_bank__abc_33898_n4178;
  wire REGFILE_SIM_reg_bank__abc_33898_n4179;
  wire REGFILE_SIM_reg_bank__abc_33898_n4181;
  wire REGFILE_SIM_reg_bank__abc_33898_n4182;
  wire REGFILE_SIM_reg_bank__abc_33898_n4184;
  wire REGFILE_SIM_reg_bank__abc_33898_n4185;
  wire REGFILE_SIM_reg_bank__abc_33898_n4187;
  wire REGFILE_SIM_reg_bank__abc_33898_n4188;
  wire REGFILE_SIM_reg_bank__abc_33898_n4190_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4191;
  wire REGFILE_SIM_reg_bank__abc_33898_n4193_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4194;
  wire REGFILE_SIM_reg_bank__abc_33898_n4196;
  wire REGFILE_SIM_reg_bank__abc_33898_n4197_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4199;
  wire REGFILE_SIM_reg_bank__abc_33898_n4200;
  wire REGFILE_SIM_reg_bank__abc_33898_n4202;
  wire REGFILE_SIM_reg_bank__abc_33898_n4203;
  wire REGFILE_SIM_reg_bank__abc_33898_n4205;
  wire REGFILE_SIM_reg_bank__abc_33898_n4206;
  wire REGFILE_SIM_reg_bank__abc_33898_n4208;
  wire REGFILE_SIM_reg_bank__abc_33898_n4209;
  wire REGFILE_SIM_reg_bank__abc_33898_n4211;
  wire REGFILE_SIM_reg_bank__abc_33898_n4212;
  wire REGFILE_SIM_reg_bank__abc_33898_n4214;
  wire REGFILE_SIM_reg_bank__abc_33898_n4215;
  wire REGFILE_SIM_reg_bank__abc_33898_n4217;
  wire REGFILE_SIM_reg_bank__abc_33898_n4218;
  wire REGFILE_SIM_reg_bank__abc_33898_n4220;
  wire REGFILE_SIM_reg_bank__abc_33898_n4221;
  wire REGFILE_SIM_reg_bank__abc_33898_n4223;
  wire REGFILE_SIM_reg_bank__abc_33898_n4224;
  wire REGFILE_SIM_reg_bank__abc_33898_n4226;
  wire REGFILE_SIM_reg_bank__abc_33898_n4227;
  wire REGFILE_SIM_reg_bank__abc_33898_n4229;
  wire REGFILE_SIM_reg_bank__abc_33898_n4230;
  wire REGFILE_SIM_reg_bank__abc_33898_n4232;
  wire REGFILE_SIM_reg_bank__abc_33898_n4233;
  wire REGFILE_SIM_reg_bank__abc_33898_n4235;
  wire REGFILE_SIM_reg_bank__abc_33898_n4236;
  wire REGFILE_SIM_reg_bank__abc_33898_n4238;
  wire REGFILE_SIM_reg_bank__abc_33898_n4239;
  wire REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4240;
  wire REGFILE_SIM_reg_bank__abc_33898_n4241;
  wire REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4242;
  wire REGFILE_SIM_reg_bank__abc_33898_n4244;
  wire REGFILE_SIM_reg_bank__abc_33898_n4245;
  wire REGFILE_SIM_reg_bank__abc_33898_n4247;
  wire REGFILE_SIM_reg_bank__abc_33898_n4248;
  wire REGFILE_SIM_reg_bank__abc_33898_n4250;
  wire REGFILE_SIM_reg_bank__abc_33898_n4251;
  wire REGFILE_SIM_reg_bank__abc_33898_n4253;
  wire REGFILE_SIM_reg_bank__abc_33898_n4254;
  wire REGFILE_SIM_reg_bank__abc_33898_n4256;
  wire REGFILE_SIM_reg_bank__abc_33898_n4257;
  wire REGFILE_SIM_reg_bank__abc_33898_n4259;
  wire REGFILE_SIM_reg_bank__abc_33898_n4260;
  wire REGFILE_SIM_reg_bank__abc_33898_n4262;
  wire REGFILE_SIM_reg_bank__abc_33898_n4263;
  wire REGFILE_SIM_reg_bank__abc_33898_n4265;
  wire REGFILE_SIM_reg_bank__abc_33898_n4266;
  wire REGFILE_SIM_reg_bank__abc_33898_n4268;
  wire REGFILE_SIM_reg_bank__abc_33898_n4269;
  wire REGFILE_SIM_reg_bank__abc_33898_n4271;
  wire REGFILE_SIM_reg_bank__abc_33898_n4272;
  wire REGFILE_SIM_reg_bank__abc_33898_n4274;
  wire REGFILE_SIM_reg_bank__abc_33898_n4275;
  wire REGFILE_SIM_reg_bank__abc_33898_n4277;
  wire REGFILE_SIM_reg_bank__abc_33898_n4278;
  wire REGFILE_SIM_reg_bank__abc_33898_n4280;
  wire REGFILE_SIM_reg_bank__abc_33898_n4281;
  wire REGFILE_SIM_reg_bank__abc_33898_n4283;
  wire REGFILE_SIM_reg_bank__abc_33898_n4284;
  wire REGFILE_SIM_reg_bank__abc_33898_n4286;
  wire REGFILE_SIM_reg_bank__abc_33898_n4287;
  wire REGFILE_SIM_reg_bank__abc_33898_n4289;
  wire REGFILE_SIM_reg_bank__abc_33898_n4290;
  wire REGFILE_SIM_reg_bank__abc_33898_n4292;
  wire REGFILE_SIM_reg_bank__abc_33898_n4293;
  wire REGFILE_SIM_reg_bank__abc_33898_n4295;
  wire REGFILE_SIM_reg_bank__abc_33898_n4296;
  wire REGFILE_SIM_reg_bank__abc_33898_n4298;
  wire REGFILE_SIM_reg_bank__abc_33898_n4299;
  wire REGFILE_SIM_reg_bank__abc_33898_n4301;
  wire REGFILE_SIM_reg_bank__abc_33898_n4302;
  wire REGFILE_SIM_reg_bank__abc_33898_n4304;
  wire REGFILE_SIM_reg_bank__abc_33898_n4305;
  wire REGFILE_SIM_reg_bank__abc_33898_n4307;
  wire REGFILE_SIM_reg_bank__abc_33898_n4308;
  wire REGFILE_SIM_reg_bank__abc_33898_n4310;
  wire REGFILE_SIM_reg_bank__abc_33898_n4311;
  wire REGFILE_SIM_reg_bank__abc_33898_n4313_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4314;
  wire REGFILE_SIM_reg_bank__abc_33898_n4316;
  wire REGFILE_SIM_reg_bank__abc_33898_n4317;
  wire REGFILE_SIM_reg_bank__abc_33898_n4319;
  wire REGFILE_SIM_reg_bank__abc_33898_n4320;
  wire REGFILE_SIM_reg_bank__abc_33898_n4322;
  wire REGFILE_SIM_reg_bank__abc_33898_n4323;
  wire REGFILE_SIM_reg_bank__abc_33898_n4325;
  wire REGFILE_SIM_reg_bank__abc_33898_n4326;
  wire REGFILE_SIM_reg_bank__abc_33898_n4328;
  wire REGFILE_SIM_reg_bank__abc_33898_n4329;
  wire REGFILE_SIM_reg_bank__abc_33898_n4331;
  wire REGFILE_SIM_reg_bank__abc_33898_n4332;
  wire REGFILE_SIM_reg_bank__abc_33898_n4334;
  wire REGFILE_SIM_reg_bank__abc_33898_n4335;
  wire REGFILE_SIM_reg_bank__abc_33898_n4337;
  wire REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4338;
  wire REGFILE_SIM_reg_bank__abc_33898_n4339;
  wire REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4340;
  wire REGFILE_SIM_reg_bank__abc_33898_n4342;
  wire REGFILE_SIM_reg_bank__abc_33898_n4343_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4345;
  wire REGFILE_SIM_reg_bank__abc_33898_n4346;
  wire REGFILE_SIM_reg_bank__abc_33898_n4348;
  wire REGFILE_SIM_reg_bank__abc_33898_n4349;
  wire REGFILE_SIM_reg_bank__abc_33898_n4351;
  wire REGFILE_SIM_reg_bank__abc_33898_n4352;
  wire REGFILE_SIM_reg_bank__abc_33898_n4354;
  wire REGFILE_SIM_reg_bank__abc_33898_n4355;
  wire REGFILE_SIM_reg_bank__abc_33898_n4357;
  wire REGFILE_SIM_reg_bank__abc_33898_n4358;
  wire REGFILE_SIM_reg_bank__abc_33898_n4360;
  wire REGFILE_SIM_reg_bank__abc_33898_n4361;
  wire REGFILE_SIM_reg_bank__abc_33898_n4363;
  wire REGFILE_SIM_reg_bank__abc_33898_n4364;
  wire REGFILE_SIM_reg_bank__abc_33898_n4366;
  wire REGFILE_SIM_reg_bank__abc_33898_n4367;
  wire REGFILE_SIM_reg_bank__abc_33898_n4369;
  wire REGFILE_SIM_reg_bank__abc_33898_n4370;
  wire REGFILE_SIM_reg_bank__abc_33898_n4372;
  wire REGFILE_SIM_reg_bank__abc_33898_n4373_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4375;
  wire REGFILE_SIM_reg_bank__abc_33898_n4376;
  wire REGFILE_SIM_reg_bank__abc_33898_n4378;
  wire REGFILE_SIM_reg_bank__abc_33898_n4379;
  wire REGFILE_SIM_reg_bank__abc_33898_n4381;
  wire REGFILE_SIM_reg_bank__abc_33898_n4382;
  wire REGFILE_SIM_reg_bank__abc_33898_n4384;
  wire REGFILE_SIM_reg_bank__abc_33898_n4385;
  wire REGFILE_SIM_reg_bank__abc_33898_n4387;
  wire REGFILE_SIM_reg_bank__abc_33898_n4388;
  wire REGFILE_SIM_reg_bank__abc_33898_n4390;
  wire REGFILE_SIM_reg_bank__abc_33898_n4391;
  wire REGFILE_SIM_reg_bank__abc_33898_n4393;
  wire REGFILE_SIM_reg_bank__abc_33898_n4394;
  wire REGFILE_SIM_reg_bank__abc_33898_n4396;
  wire REGFILE_SIM_reg_bank__abc_33898_n4397;
  wire REGFILE_SIM_reg_bank__abc_33898_n4399;
  wire REGFILE_SIM_reg_bank__abc_33898_n4400;
  wire REGFILE_SIM_reg_bank__abc_33898_n4402;
  wire REGFILE_SIM_reg_bank__abc_33898_n4403_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4405;
  wire REGFILE_SIM_reg_bank__abc_33898_n4406;
  wire REGFILE_SIM_reg_bank__abc_33898_n4408;
  wire REGFILE_SIM_reg_bank__abc_33898_n4409;
  wire REGFILE_SIM_reg_bank__abc_33898_n4411;
  wire REGFILE_SIM_reg_bank__abc_33898_n4412;
  wire REGFILE_SIM_reg_bank__abc_33898_n4414;
  wire REGFILE_SIM_reg_bank__abc_33898_n4415;
  wire REGFILE_SIM_reg_bank__abc_33898_n4417;
  wire REGFILE_SIM_reg_bank__abc_33898_n4418;
  wire REGFILE_SIM_reg_bank__abc_33898_n4420;
  wire REGFILE_SIM_reg_bank__abc_33898_n4421;
  wire REGFILE_SIM_reg_bank__abc_33898_n4423;
  wire REGFILE_SIM_reg_bank__abc_33898_n4424;
  wire REGFILE_SIM_reg_bank__abc_33898_n4426;
  wire REGFILE_SIM_reg_bank__abc_33898_n4427;
  wire REGFILE_SIM_reg_bank__abc_33898_n4429;
  wire REGFILE_SIM_reg_bank__abc_33898_n4430;
  wire REGFILE_SIM_reg_bank__abc_33898_n4432;
  wire REGFILE_SIM_reg_bank__abc_33898_n4433_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n4436;
  wire REGFILE_SIM_reg_bank__abc_33898_n4437;
  wire REGFILE_SIM_reg_bank__abc_33898_n4438;
  wire REGFILE_SIM_reg_bank__abc_33898_n4440;
  wire REGFILE_SIM_reg_bank__abc_33898_n4441;
  wire REGFILE_SIM_reg_bank__abc_33898_n4442;
  wire REGFILE_SIM_reg_bank__abc_33898_n4444;
  wire REGFILE_SIM_reg_bank__abc_33898_n4445;
  wire REGFILE_SIM_reg_bank__abc_33898_n4446;
  wire REGFILE_SIM_reg_bank__abc_33898_n4448;
  wire REGFILE_SIM_reg_bank__abc_33898_n4449;
  wire REGFILE_SIM_reg_bank__abc_33898_n4450;
  wire REGFILE_SIM_reg_bank__abc_33898_n4452;
  wire REGFILE_SIM_reg_bank__abc_33898_n4453;
  wire REGFILE_SIM_reg_bank__abc_33898_n4454;
  wire REGFILE_SIM_reg_bank__abc_33898_n4456;
  wire REGFILE_SIM_reg_bank__abc_33898_n4457;
  wire REGFILE_SIM_reg_bank__abc_33898_n4458;
  wire REGFILE_SIM_reg_bank__abc_33898_n4460;
  wire REGFILE_SIM_reg_bank__abc_33898_n4461;
  wire REGFILE_SIM_reg_bank__abc_33898_n4462;
  wire REGFILE_SIM_reg_bank__abc_33898_n4464;
  wire REGFILE_SIM_reg_bank__abc_33898_n4465;
  wire REGFILE_SIM_reg_bank__abc_33898_n4466;
  wire REGFILE_SIM_reg_bank__abc_33898_n4468;
  wire REGFILE_SIM_reg_bank__abc_33898_n4469;
  wire REGFILE_SIM_reg_bank__abc_33898_n4470;
  wire REGFILE_SIM_reg_bank__abc_33898_n4472;
  wire REGFILE_SIM_reg_bank__abc_33898_n4473;
  wire REGFILE_SIM_reg_bank__abc_33898_n4474;
  wire REGFILE_SIM_reg_bank__abc_33898_n4476;
  wire REGFILE_SIM_reg_bank__abc_33898_n4477;
  wire REGFILE_SIM_reg_bank__abc_33898_n4478;
  wire REGFILE_SIM_reg_bank__abc_33898_n4480;
  wire REGFILE_SIM_reg_bank__abc_33898_n4481;
  wire REGFILE_SIM_reg_bank__abc_33898_n4482;
  wire REGFILE_SIM_reg_bank__abc_33898_n4484;
  wire REGFILE_SIM_reg_bank__abc_33898_n4485;
  wire REGFILE_SIM_reg_bank__abc_33898_n4486;
  wire REGFILE_SIM_reg_bank__abc_33898_n4488;
  wire REGFILE_SIM_reg_bank__abc_33898_n4489;
  wire REGFILE_SIM_reg_bank__abc_33898_n4490;
  wire REGFILE_SIM_reg_bank__abc_33898_n4492;
  wire REGFILE_SIM_reg_bank__abc_33898_n4493_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4494;
  wire REGFILE_SIM_reg_bank__abc_33898_n4496;
  wire REGFILE_SIM_reg_bank__abc_33898_n4497;
  wire REGFILE_SIM_reg_bank__abc_33898_n4498;
  wire REGFILE_SIM_reg_bank__abc_33898_n4500;
  wire REGFILE_SIM_reg_bank__abc_33898_n4501;
  wire REGFILE_SIM_reg_bank__abc_33898_n4502;
  wire REGFILE_SIM_reg_bank__abc_33898_n4504;
  wire REGFILE_SIM_reg_bank__abc_33898_n4505;
  wire REGFILE_SIM_reg_bank__abc_33898_n4506;
  wire REGFILE_SIM_reg_bank__abc_33898_n4508;
  wire REGFILE_SIM_reg_bank__abc_33898_n4509;
  wire REGFILE_SIM_reg_bank__abc_33898_n4510;
  wire REGFILE_SIM_reg_bank__abc_33898_n4512;
  wire REGFILE_SIM_reg_bank__abc_33898_n4513;
  wire REGFILE_SIM_reg_bank__abc_33898_n4514;
  wire REGFILE_SIM_reg_bank__abc_33898_n4516;
  wire REGFILE_SIM_reg_bank__abc_33898_n4517;
  wire REGFILE_SIM_reg_bank__abc_33898_n4518;
  wire REGFILE_SIM_reg_bank__abc_33898_n4520;
  wire REGFILE_SIM_reg_bank__abc_33898_n4521;
  wire REGFILE_SIM_reg_bank__abc_33898_n4522;
  wire REGFILE_SIM_reg_bank__abc_33898_n4524;
  wire REGFILE_SIM_reg_bank__abc_33898_n4525;
  wire REGFILE_SIM_reg_bank__abc_33898_n4526;
  wire REGFILE_SIM_reg_bank__abc_33898_n4528;
  wire REGFILE_SIM_reg_bank__abc_33898_n4529;
  wire REGFILE_SIM_reg_bank__abc_33898_n4530;
  wire REGFILE_SIM_reg_bank__abc_33898_n4532;
  wire REGFILE_SIM_reg_bank__abc_33898_n4533;
  wire REGFILE_SIM_reg_bank__abc_33898_n4534;
  wire REGFILE_SIM_reg_bank__abc_33898_n4536;
  wire REGFILE_SIM_reg_bank__abc_33898_n4537;
  wire REGFILE_SIM_reg_bank__abc_33898_n4538;
  wire REGFILE_SIM_reg_bank__abc_33898_n4540;
  wire REGFILE_SIM_reg_bank__abc_33898_n4541;
  wire REGFILE_SIM_reg_bank__abc_33898_n4542;
  wire REGFILE_SIM_reg_bank__abc_33898_n4544;
  wire REGFILE_SIM_reg_bank__abc_33898_n4545;
  wire REGFILE_SIM_reg_bank__abc_33898_n4546;
  wire REGFILE_SIM_reg_bank__abc_33898_n4548;
  wire REGFILE_SIM_reg_bank__abc_33898_n4549;
  wire REGFILE_SIM_reg_bank__abc_33898_n4550;
  wire REGFILE_SIM_reg_bank__abc_33898_n4552;
  wire REGFILE_SIM_reg_bank__abc_33898_n4553_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4554;
  wire REGFILE_SIM_reg_bank__abc_33898_n4556;
  wire REGFILE_SIM_reg_bank__abc_33898_n4557;
  wire REGFILE_SIM_reg_bank__abc_33898_n4558;
  wire REGFILE_SIM_reg_bank__abc_33898_n4560;
  wire REGFILE_SIM_reg_bank__abc_33898_n4561;
  wire REGFILE_SIM_reg_bank__abc_33898_n4562;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n4565;
  wire REGFILE_SIM_reg_bank__abc_33898_n4566;
  wire REGFILE_SIM_reg_bank__abc_33898_n4567;
  wire REGFILE_SIM_reg_bank__abc_33898_n4569;
  wire REGFILE_SIM_reg_bank__abc_33898_n4570;
  wire REGFILE_SIM_reg_bank__abc_33898_n4571;
  wire REGFILE_SIM_reg_bank__abc_33898_n4573;
  wire REGFILE_SIM_reg_bank__abc_33898_n4574;
  wire REGFILE_SIM_reg_bank__abc_33898_n4575;
  wire REGFILE_SIM_reg_bank__abc_33898_n4577;
  wire REGFILE_SIM_reg_bank__abc_33898_n4578;
  wire REGFILE_SIM_reg_bank__abc_33898_n4579;
  wire REGFILE_SIM_reg_bank__abc_33898_n4581;
  wire REGFILE_SIM_reg_bank__abc_33898_n4582;
  wire REGFILE_SIM_reg_bank__abc_33898_n4583_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4585;
  wire REGFILE_SIM_reg_bank__abc_33898_n4586;
  wire REGFILE_SIM_reg_bank__abc_33898_n4587;
  wire REGFILE_SIM_reg_bank__abc_33898_n4589;
  wire REGFILE_SIM_reg_bank__abc_33898_n4590;
  wire REGFILE_SIM_reg_bank__abc_33898_n4591;
  wire REGFILE_SIM_reg_bank__abc_33898_n4593;
  wire REGFILE_SIM_reg_bank__abc_33898_n4594;
  wire REGFILE_SIM_reg_bank__abc_33898_n4595;
  wire REGFILE_SIM_reg_bank__abc_33898_n4597;
  wire REGFILE_SIM_reg_bank__abc_33898_n4598;
  wire REGFILE_SIM_reg_bank__abc_33898_n4599;
  wire REGFILE_SIM_reg_bank__abc_33898_n4601;
  wire REGFILE_SIM_reg_bank__abc_33898_n4602;
  wire REGFILE_SIM_reg_bank__abc_33898_n4603;
  wire REGFILE_SIM_reg_bank__abc_33898_n4605;
  wire REGFILE_SIM_reg_bank__abc_33898_n4606;
  wire REGFILE_SIM_reg_bank__abc_33898_n4607;
  wire REGFILE_SIM_reg_bank__abc_33898_n4609;
  wire REGFILE_SIM_reg_bank__abc_33898_n4610;
  wire REGFILE_SIM_reg_bank__abc_33898_n4611;
  wire REGFILE_SIM_reg_bank__abc_33898_n4613_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4614;
  wire REGFILE_SIM_reg_bank__abc_33898_n4615;
  wire REGFILE_SIM_reg_bank__abc_33898_n4617;
  wire REGFILE_SIM_reg_bank__abc_33898_n4618;
  wire REGFILE_SIM_reg_bank__abc_33898_n4619;
  wire REGFILE_SIM_reg_bank__abc_33898_n4621;
  wire REGFILE_SIM_reg_bank__abc_33898_n4622;
  wire REGFILE_SIM_reg_bank__abc_33898_n4623;
  wire REGFILE_SIM_reg_bank__abc_33898_n4625;
  wire REGFILE_SIM_reg_bank__abc_33898_n4626;
  wire REGFILE_SIM_reg_bank__abc_33898_n4627;
  wire REGFILE_SIM_reg_bank__abc_33898_n4629;
  wire REGFILE_SIM_reg_bank__abc_33898_n4630;
  wire REGFILE_SIM_reg_bank__abc_33898_n4631;
  wire REGFILE_SIM_reg_bank__abc_33898_n4633;
  wire REGFILE_SIM_reg_bank__abc_33898_n4634;
  wire REGFILE_SIM_reg_bank__abc_33898_n4635;
  wire REGFILE_SIM_reg_bank__abc_33898_n4637;
  wire REGFILE_SIM_reg_bank__abc_33898_n4638;
  wire REGFILE_SIM_reg_bank__abc_33898_n4639;
  wire REGFILE_SIM_reg_bank__abc_33898_n4641;
  wire REGFILE_SIM_reg_bank__abc_33898_n4642;
  wire REGFILE_SIM_reg_bank__abc_33898_n4643_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4645;
  wire REGFILE_SIM_reg_bank__abc_33898_n4646;
  wire REGFILE_SIM_reg_bank__abc_33898_n4647;
  wire REGFILE_SIM_reg_bank__abc_33898_n4649;
  wire REGFILE_SIM_reg_bank__abc_33898_n4650;
  wire REGFILE_SIM_reg_bank__abc_33898_n4651;
  wire REGFILE_SIM_reg_bank__abc_33898_n4653;
  wire REGFILE_SIM_reg_bank__abc_33898_n4654;
  wire REGFILE_SIM_reg_bank__abc_33898_n4655;
  wire REGFILE_SIM_reg_bank__abc_33898_n4657;
  wire REGFILE_SIM_reg_bank__abc_33898_n4658;
  wire REGFILE_SIM_reg_bank__abc_33898_n4659;
  wire REGFILE_SIM_reg_bank__abc_33898_n4661;
  wire REGFILE_SIM_reg_bank__abc_33898_n4662;
  wire REGFILE_SIM_reg_bank__abc_33898_n4663;
  wire REGFILE_SIM_reg_bank__abc_33898_n4665;
  wire REGFILE_SIM_reg_bank__abc_33898_n4666;
  wire REGFILE_SIM_reg_bank__abc_33898_n4667;
  wire REGFILE_SIM_reg_bank__abc_33898_n4669;
  wire REGFILE_SIM_reg_bank__abc_33898_n4670;
  wire REGFILE_SIM_reg_bank__abc_33898_n4671;
  wire REGFILE_SIM_reg_bank__abc_33898_n4673_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4674;
  wire REGFILE_SIM_reg_bank__abc_33898_n4675;
  wire REGFILE_SIM_reg_bank__abc_33898_n4677;
  wire REGFILE_SIM_reg_bank__abc_33898_n4678;
  wire REGFILE_SIM_reg_bank__abc_33898_n4679;
  wire REGFILE_SIM_reg_bank__abc_33898_n4681;
  wire REGFILE_SIM_reg_bank__abc_33898_n4682;
  wire REGFILE_SIM_reg_bank__abc_33898_n4683;
  wire REGFILE_SIM_reg_bank__abc_33898_n4685;
  wire REGFILE_SIM_reg_bank__abc_33898_n4686;
  wire REGFILE_SIM_reg_bank__abc_33898_n4687;
  wire REGFILE_SIM_reg_bank__abc_33898_n4689;
  wire REGFILE_SIM_reg_bank__abc_33898_n4690;
  wire REGFILE_SIM_reg_bank__abc_33898_n4691;
  wire REGFILE_SIM_reg_bank__abc_33898_n4693;
  wire REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4694;
  wire REGFILE_SIM_reg_bank__abc_33898_n4695;
  wire REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4696;
  wire REGFILE_SIM_reg_bank__abc_33898_n4698;
  wire REGFILE_SIM_reg_bank__abc_33898_n4699;
  wire REGFILE_SIM_reg_bank__abc_33898_n4701;
  wire REGFILE_SIM_reg_bank__abc_33898_n4702;
  wire REGFILE_SIM_reg_bank__abc_33898_n4704;
  wire REGFILE_SIM_reg_bank__abc_33898_n4705;
  wire REGFILE_SIM_reg_bank__abc_33898_n4707;
  wire REGFILE_SIM_reg_bank__abc_33898_n4708;
  wire REGFILE_SIM_reg_bank__abc_33898_n4710;
  wire REGFILE_SIM_reg_bank__abc_33898_n4711;
  wire REGFILE_SIM_reg_bank__abc_33898_n4713;
  wire REGFILE_SIM_reg_bank__abc_33898_n4714;
  wire REGFILE_SIM_reg_bank__abc_33898_n4716;
  wire REGFILE_SIM_reg_bank__abc_33898_n4717;
  wire REGFILE_SIM_reg_bank__abc_33898_n4719;
  wire REGFILE_SIM_reg_bank__abc_33898_n4720;
  wire REGFILE_SIM_reg_bank__abc_33898_n4722;
  wire REGFILE_SIM_reg_bank__abc_33898_n4723;
  wire REGFILE_SIM_reg_bank__abc_33898_n4725;
  wire REGFILE_SIM_reg_bank__abc_33898_n4726;
  wire REGFILE_SIM_reg_bank__abc_33898_n4728;
  wire REGFILE_SIM_reg_bank__abc_33898_n4729;
  wire REGFILE_SIM_reg_bank__abc_33898_n4731;
  wire REGFILE_SIM_reg_bank__abc_33898_n4732;
  wire REGFILE_SIM_reg_bank__abc_33898_n4734;
  wire REGFILE_SIM_reg_bank__abc_33898_n4735;
  wire REGFILE_SIM_reg_bank__abc_33898_n4737;
  wire REGFILE_SIM_reg_bank__abc_33898_n4738;
  wire REGFILE_SIM_reg_bank__abc_33898_n4740;
  wire REGFILE_SIM_reg_bank__abc_33898_n4741;
  wire REGFILE_SIM_reg_bank__abc_33898_n4743;
  wire REGFILE_SIM_reg_bank__abc_33898_n4744;
  wire REGFILE_SIM_reg_bank__abc_33898_n4746;
  wire REGFILE_SIM_reg_bank__abc_33898_n4747;
  wire REGFILE_SIM_reg_bank__abc_33898_n4749;
  wire REGFILE_SIM_reg_bank__abc_33898_n4750;
  wire REGFILE_SIM_reg_bank__abc_33898_n4752;
  wire REGFILE_SIM_reg_bank__abc_33898_n4753;
  wire REGFILE_SIM_reg_bank__abc_33898_n4755;
  wire REGFILE_SIM_reg_bank__abc_33898_n4756;
  wire REGFILE_SIM_reg_bank__abc_33898_n4758;
  wire REGFILE_SIM_reg_bank__abc_33898_n4759;
  wire REGFILE_SIM_reg_bank__abc_33898_n4761;
  wire REGFILE_SIM_reg_bank__abc_33898_n4762;
  wire REGFILE_SIM_reg_bank__abc_33898_n4764;
  wire REGFILE_SIM_reg_bank__abc_33898_n4765;
  wire REGFILE_SIM_reg_bank__abc_33898_n4767;
  wire REGFILE_SIM_reg_bank__abc_33898_n4768;
  wire REGFILE_SIM_reg_bank__abc_33898_n4770;
  wire REGFILE_SIM_reg_bank__abc_33898_n4771;
  wire REGFILE_SIM_reg_bank__abc_33898_n4773;
  wire REGFILE_SIM_reg_bank__abc_33898_n4774;
  wire REGFILE_SIM_reg_bank__abc_33898_n4776;
  wire REGFILE_SIM_reg_bank__abc_33898_n4777;
  wire REGFILE_SIM_reg_bank__abc_33898_n4779;
  wire REGFILE_SIM_reg_bank__abc_33898_n4780;
  wire REGFILE_SIM_reg_bank__abc_33898_n4782;
  wire REGFILE_SIM_reg_bank__abc_33898_n4783;
  wire REGFILE_SIM_reg_bank__abc_33898_n4785;
  wire REGFILE_SIM_reg_bank__abc_33898_n4786;
  wire REGFILE_SIM_reg_bank__abc_33898_n4788;
  wire REGFILE_SIM_reg_bank__abc_33898_n4789;
  wire REGFILE_SIM_reg_bank__abc_33898_n4791;
  wire REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4792;
  wire REGFILE_SIM_reg_bank__abc_33898_n4793_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4794;
  wire REGFILE_SIM_reg_bank__abc_33898_n4796;
  wire REGFILE_SIM_reg_bank__abc_33898_n4797;
  wire REGFILE_SIM_reg_bank__abc_33898_n4799;
  wire REGFILE_SIM_reg_bank__abc_33898_n4800;
  wire REGFILE_SIM_reg_bank__abc_33898_n4802;
  wire REGFILE_SIM_reg_bank__abc_33898_n4803;
  wire REGFILE_SIM_reg_bank__abc_33898_n4805;
  wire REGFILE_SIM_reg_bank__abc_33898_n4806;
  wire REGFILE_SIM_reg_bank__abc_33898_n4808;
  wire REGFILE_SIM_reg_bank__abc_33898_n4809;
  wire REGFILE_SIM_reg_bank__abc_33898_n4811;
  wire REGFILE_SIM_reg_bank__abc_33898_n4812;
  wire REGFILE_SIM_reg_bank__abc_33898_n4814;
  wire REGFILE_SIM_reg_bank__abc_33898_n4815;
  wire REGFILE_SIM_reg_bank__abc_33898_n4817;
  wire REGFILE_SIM_reg_bank__abc_33898_n4818;
  wire REGFILE_SIM_reg_bank__abc_33898_n4820;
  wire REGFILE_SIM_reg_bank__abc_33898_n4821;
  wire REGFILE_SIM_reg_bank__abc_33898_n4823_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4824;
  wire REGFILE_SIM_reg_bank__abc_33898_n4826;
  wire REGFILE_SIM_reg_bank__abc_33898_n4827;
  wire REGFILE_SIM_reg_bank__abc_33898_n4829;
  wire REGFILE_SIM_reg_bank__abc_33898_n4830;
  wire REGFILE_SIM_reg_bank__abc_33898_n4832;
  wire REGFILE_SIM_reg_bank__abc_33898_n4833;
  wire REGFILE_SIM_reg_bank__abc_33898_n4835;
  wire REGFILE_SIM_reg_bank__abc_33898_n4836;
  wire REGFILE_SIM_reg_bank__abc_33898_n4838;
  wire REGFILE_SIM_reg_bank__abc_33898_n4839;
  wire REGFILE_SIM_reg_bank__abc_33898_n4841;
  wire REGFILE_SIM_reg_bank__abc_33898_n4842;
  wire REGFILE_SIM_reg_bank__abc_33898_n4844;
  wire REGFILE_SIM_reg_bank__abc_33898_n4845;
  wire REGFILE_SIM_reg_bank__abc_33898_n4847;
  wire REGFILE_SIM_reg_bank__abc_33898_n4848;
  wire REGFILE_SIM_reg_bank__abc_33898_n4850;
  wire REGFILE_SIM_reg_bank__abc_33898_n4851;
  wire REGFILE_SIM_reg_bank__abc_33898_n4853_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4854;
  wire REGFILE_SIM_reg_bank__abc_33898_n4856;
  wire REGFILE_SIM_reg_bank__abc_33898_n4857;
  wire REGFILE_SIM_reg_bank__abc_33898_n4859;
  wire REGFILE_SIM_reg_bank__abc_33898_n4860;
  wire REGFILE_SIM_reg_bank__abc_33898_n4862;
  wire REGFILE_SIM_reg_bank__abc_33898_n4863;
  wire REGFILE_SIM_reg_bank__abc_33898_n4865;
  wire REGFILE_SIM_reg_bank__abc_33898_n4866;
  wire REGFILE_SIM_reg_bank__abc_33898_n4868;
  wire REGFILE_SIM_reg_bank__abc_33898_n4869;
  wire REGFILE_SIM_reg_bank__abc_33898_n4871;
  wire REGFILE_SIM_reg_bank__abc_33898_n4872;
  wire REGFILE_SIM_reg_bank__abc_33898_n4874;
  wire REGFILE_SIM_reg_bank__abc_33898_n4875;
  wire REGFILE_SIM_reg_bank__abc_33898_n4877;
  wire REGFILE_SIM_reg_bank__abc_33898_n4878;
  wire REGFILE_SIM_reg_bank__abc_33898_n4880;
  wire REGFILE_SIM_reg_bank__abc_33898_n4881;
  wire REGFILE_SIM_reg_bank__abc_33898_n4883_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4884;
  wire REGFILE_SIM_reg_bank__abc_33898_n4886;
  wire REGFILE_SIM_reg_bank__abc_33898_n4887;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n4890;
  wire REGFILE_SIM_reg_bank__abc_33898_n4891;
  wire REGFILE_SIM_reg_bank__abc_33898_n4892;
  wire REGFILE_SIM_reg_bank__abc_33898_n4894;
  wire REGFILE_SIM_reg_bank__abc_33898_n4895;
  wire REGFILE_SIM_reg_bank__abc_33898_n4896;
  wire REGFILE_SIM_reg_bank__abc_33898_n4898;
  wire REGFILE_SIM_reg_bank__abc_33898_n4899;
  wire REGFILE_SIM_reg_bank__abc_33898_n4900;
  wire REGFILE_SIM_reg_bank__abc_33898_n4902;
  wire REGFILE_SIM_reg_bank__abc_33898_n4903;
  wire REGFILE_SIM_reg_bank__abc_33898_n4904;
  wire REGFILE_SIM_reg_bank__abc_33898_n4906;
  wire REGFILE_SIM_reg_bank__abc_33898_n4907;
  wire REGFILE_SIM_reg_bank__abc_33898_n4908;
  wire REGFILE_SIM_reg_bank__abc_33898_n4910;
  wire REGFILE_SIM_reg_bank__abc_33898_n4911;
  wire REGFILE_SIM_reg_bank__abc_33898_n4912;
  wire REGFILE_SIM_reg_bank__abc_33898_n4914;
  wire REGFILE_SIM_reg_bank__abc_33898_n4915;
  wire REGFILE_SIM_reg_bank__abc_33898_n4916;
  wire REGFILE_SIM_reg_bank__abc_33898_n4918;
  wire REGFILE_SIM_reg_bank__abc_33898_n4919;
  wire REGFILE_SIM_reg_bank__abc_33898_n4920;
  wire REGFILE_SIM_reg_bank__abc_33898_n4922;
  wire REGFILE_SIM_reg_bank__abc_33898_n4923;
  wire REGFILE_SIM_reg_bank__abc_33898_n4924;
  wire REGFILE_SIM_reg_bank__abc_33898_n4926;
  wire REGFILE_SIM_reg_bank__abc_33898_n4927;
  wire REGFILE_SIM_reg_bank__abc_33898_n4928;
  wire REGFILE_SIM_reg_bank__abc_33898_n4930;
  wire REGFILE_SIM_reg_bank__abc_33898_n4931;
  wire REGFILE_SIM_reg_bank__abc_33898_n4932;
  wire REGFILE_SIM_reg_bank__abc_33898_n4934;
  wire REGFILE_SIM_reg_bank__abc_33898_n4935;
  wire REGFILE_SIM_reg_bank__abc_33898_n4936;
  wire REGFILE_SIM_reg_bank__abc_33898_n4938;
  wire REGFILE_SIM_reg_bank__abc_33898_n4939;
  wire REGFILE_SIM_reg_bank__abc_33898_n4940;
  wire REGFILE_SIM_reg_bank__abc_33898_n4942;
  wire REGFILE_SIM_reg_bank__abc_33898_n4943_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n4944;
  wire REGFILE_SIM_reg_bank__abc_33898_n4946;
  wire REGFILE_SIM_reg_bank__abc_33898_n4947;
  wire REGFILE_SIM_reg_bank__abc_33898_n4948;
  wire REGFILE_SIM_reg_bank__abc_33898_n4950;
  wire REGFILE_SIM_reg_bank__abc_33898_n4951;
  wire REGFILE_SIM_reg_bank__abc_33898_n4952;
  wire REGFILE_SIM_reg_bank__abc_33898_n4954;
  wire REGFILE_SIM_reg_bank__abc_33898_n4955;
  wire REGFILE_SIM_reg_bank__abc_33898_n4956;
  wire REGFILE_SIM_reg_bank__abc_33898_n4958;
  wire REGFILE_SIM_reg_bank__abc_33898_n4959;
  wire REGFILE_SIM_reg_bank__abc_33898_n4960;
  wire REGFILE_SIM_reg_bank__abc_33898_n4962;
  wire REGFILE_SIM_reg_bank__abc_33898_n4963;
  wire REGFILE_SIM_reg_bank__abc_33898_n4964;
  wire REGFILE_SIM_reg_bank__abc_33898_n4966;
  wire REGFILE_SIM_reg_bank__abc_33898_n4967;
  wire REGFILE_SIM_reg_bank__abc_33898_n4968;
  wire REGFILE_SIM_reg_bank__abc_33898_n4970;
  wire REGFILE_SIM_reg_bank__abc_33898_n4971;
  wire REGFILE_SIM_reg_bank__abc_33898_n4972;
  wire REGFILE_SIM_reg_bank__abc_33898_n4974;
  wire REGFILE_SIM_reg_bank__abc_33898_n4975;
  wire REGFILE_SIM_reg_bank__abc_33898_n4976;
  wire REGFILE_SIM_reg_bank__abc_33898_n4978;
  wire REGFILE_SIM_reg_bank__abc_33898_n4979;
  wire REGFILE_SIM_reg_bank__abc_33898_n4980;
  wire REGFILE_SIM_reg_bank__abc_33898_n4982;
  wire REGFILE_SIM_reg_bank__abc_33898_n4983;
  wire REGFILE_SIM_reg_bank__abc_33898_n4984;
  wire REGFILE_SIM_reg_bank__abc_33898_n4986;
  wire REGFILE_SIM_reg_bank__abc_33898_n4987;
  wire REGFILE_SIM_reg_bank__abc_33898_n4988;
  wire REGFILE_SIM_reg_bank__abc_33898_n4990;
  wire REGFILE_SIM_reg_bank__abc_33898_n4991;
  wire REGFILE_SIM_reg_bank__abc_33898_n4992;
  wire REGFILE_SIM_reg_bank__abc_33898_n4994;
  wire REGFILE_SIM_reg_bank__abc_33898_n4995;
  wire REGFILE_SIM_reg_bank__abc_33898_n4996;
  wire REGFILE_SIM_reg_bank__abc_33898_n4998;
  wire REGFILE_SIM_reg_bank__abc_33898_n4999;
  wire REGFILE_SIM_reg_bank__abc_33898_n5000;
  wire REGFILE_SIM_reg_bank__abc_33898_n5002;
  wire REGFILE_SIM_reg_bank__abc_33898_n5003_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5004;
  wire REGFILE_SIM_reg_bank__abc_33898_n5006;
  wire REGFILE_SIM_reg_bank__abc_33898_n5007;
  wire REGFILE_SIM_reg_bank__abc_33898_n5008;
  wire REGFILE_SIM_reg_bank__abc_33898_n5010;
  wire REGFILE_SIM_reg_bank__abc_33898_n5011;
  wire REGFILE_SIM_reg_bank__abc_33898_n5012;
  wire REGFILE_SIM_reg_bank__abc_33898_n5014;
  wire REGFILE_SIM_reg_bank__abc_33898_n5015;
  wire REGFILE_SIM_reg_bank__abc_33898_n5016;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n5019;
  wire REGFILE_SIM_reg_bank__abc_33898_n5020;
  wire REGFILE_SIM_reg_bank__abc_33898_n5021;
  wire REGFILE_SIM_reg_bank__abc_33898_n5023;
  wire REGFILE_SIM_reg_bank__abc_33898_n5024;
  wire REGFILE_SIM_reg_bank__abc_33898_n5025;
  wire REGFILE_SIM_reg_bank__abc_33898_n5027;
  wire REGFILE_SIM_reg_bank__abc_33898_n5028;
  wire REGFILE_SIM_reg_bank__abc_33898_n5029;
  wire REGFILE_SIM_reg_bank__abc_33898_n5031;
  wire REGFILE_SIM_reg_bank__abc_33898_n5032;
  wire REGFILE_SIM_reg_bank__abc_33898_n5033_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5035;
  wire REGFILE_SIM_reg_bank__abc_33898_n5036;
  wire REGFILE_SIM_reg_bank__abc_33898_n5037;
  wire REGFILE_SIM_reg_bank__abc_33898_n5039;
  wire REGFILE_SIM_reg_bank__abc_33898_n5040;
  wire REGFILE_SIM_reg_bank__abc_33898_n5041;
  wire REGFILE_SIM_reg_bank__abc_33898_n5043;
  wire REGFILE_SIM_reg_bank__abc_33898_n5044;
  wire REGFILE_SIM_reg_bank__abc_33898_n5045;
  wire REGFILE_SIM_reg_bank__abc_33898_n5047;
  wire REGFILE_SIM_reg_bank__abc_33898_n5048;
  wire REGFILE_SIM_reg_bank__abc_33898_n5049;
  wire REGFILE_SIM_reg_bank__abc_33898_n5051;
  wire REGFILE_SIM_reg_bank__abc_33898_n5052;
  wire REGFILE_SIM_reg_bank__abc_33898_n5053;
  wire REGFILE_SIM_reg_bank__abc_33898_n5055;
  wire REGFILE_SIM_reg_bank__abc_33898_n5056;
  wire REGFILE_SIM_reg_bank__abc_33898_n5057;
  wire REGFILE_SIM_reg_bank__abc_33898_n5059;
  wire REGFILE_SIM_reg_bank__abc_33898_n5060;
  wire REGFILE_SIM_reg_bank__abc_33898_n5061;
  wire REGFILE_SIM_reg_bank__abc_33898_n5063_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5064;
  wire REGFILE_SIM_reg_bank__abc_33898_n5065;
  wire REGFILE_SIM_reg_bank__abc_33898_n5067;
  wire REGFILE_SIM_reg_bank__abc_33898_n5068;
  wire REGFILE_SIM_reg_bank__abc_33898_n5069;
  wire REGFILE_SIM_reg_bank__abc_33898_n5071;
  wire REGFILE_SIM_reg_bank__abc_33898_n5072;
  wire REGFILE_SIM_reg_bank__abc_33898_n5073;
  wire REGFILE_SIM_reg_bank__abc_33898_n5075;
  wire REGFILE_SIM_reg_bank__abc_33898_n5076;
  wire REGFILE_SIM_reg_bank__abc_33898_n5077;
  wire REGFILE_SIM_reg_bank__abc_33898_n5079;
  wire REGFILE_SIM_reg_bank__abc_33898_n5080;
  wire REGFILE_SIM_reg_bank__abc_33898_n5081;
  wire REGFILE_SIM_reg_bank__abc_33898_n5083;
  wire REGFILE_SIM_reg_bank__abc_33898_n5084;
  wire REGFILE_SIM_reg_bank__abc_33898_n5085;
  wire REGFILE_SIM_reg_bank__abc_33898_n5087;
  wire REGFILE_SIM_reg_bank__abc_33898_n5088;
  wire REGFILE_SIM_reg_bank__abc_33898_n5089;
  wire REGFILE_SIM_reg_bank__abc_33898_n5091;
  wire REGFILE_SIM_reg_bank__abc_33898_n5092;
  wire REGFILE_SIM_reg_bank__abc_33898_n5093_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5095;
  wire REGFILE_SIM_reg_bank__abc_33898_n5096;
  wire REGFILE_SIM_reg_bank__abc_33898_n5097;
  wire REGFILE_SIM_reg_bank__abc_33898_n5099;
  wire REGFILE_SIM_reg_bank__abc_33898_n5100;
  wire REGFILE_SIM_reg_bank__abc_33898_n5101;
  wire REGFILE_SIM_reg_bank__abc_33898_n5103;
  wire REGFILE_SIM_reg_bank__abc_33898_n5104;
  wire REGFILE_SIM_reg_bank__abc_33898_n5105;
  wire REGFILE_SIM_reg_bank__abc_33898_n5107;
  wire REGFILE_SIM_reg_bank__abc_33898_n5108;
  wire REGFILE_SIM_reg_bank__abc_33898_n5109;
  wire REGFILE_SIM_reg_bank__abc_33898_n5111;
  wire REGFILE_SIM_reg_bank__abc_33898_n5112;
  wire REGFILE_SIM_reg_bank__abc_33898_n5113;
  wire REGFILE_SIM_reg_bank__abc_33898_n5115;
  wire REGFILE_SIM_reg_bank__abc_33898_n5116;
  wire REGFILE_SIM_reg_bank__abc_33898_n5117;
  wire REGFILE_SIM_reg_bank__abc_33898_n5119;
  wire REGFILE_SIM_reg_bank__abc_33898_n5120;
  wire REGFILE_SIM_reg_bank__abc_33898_n5121;
  wire REGFILE_SIM_reg_bank__abc_33898_n5123_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5124;
  wire REGFILE_SIM_reg_bank__abc_33898_n5125;
  wire REGFILE_SIM_reg_bank__abc_33898_n5127;
  wire REGFILE_SIM_reg_bank__abc_33898_n5128;
  wire REGFILE_SIM_reg_bank__abc_33898_n5129;
  wire REGFILE_SIM_reg_bank__abc_33898_n5131;
  wire REGFILE_SIM_reg_bank__abc_33898_n5132;
  wire REGFILE_SIM_reg_bank__abc_33898_n5133;
  wire REGFILE_SIM_reg_bank__abc_33898_n5135;
  wire REGFILE_SIM_reg_bank__abc_33898_n5136;
  wire REGFILE_SIM_reg_bank__abc_33898_n5137;
  wire REGFILE_SIM_reg_bank__abc_33898_n5139;
  wire REGFILE_SIM_reg_bank__abc_33898_n5140;
  wire REGFILE_SIM_reg_bank__abc_33898_n5141;
  wire REGFILE_SIM_reg_bank__abc_33898_n5143;
  wire REGFILE_SIM_reg_bank__abc_33898_n5144;
  wire REGFILE_SIM_reg_bank__abc_33898_n5145;
  wire REGFILE_SIM_reg_bank__abc_33898_n5147;
  wire REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5148;
  wire REGFILE_SIM_reg_bank__abc_33898_n5149;
  wire REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5150;
  wire REGFILE_SIM_reg_bank__abc_33898_n5152;
  wire REGFILE_SIM_reg_bank__abc_33898_n5153_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5155;
  wire REGFILE_SIM_reg_bank__abc_33898_n5156;
  wire REGFILE_SIM_reg_bank__abc_33898_n5158;
  wire REGFILE_SIM_reg_bank__abc_33898_n5159;
  wire REGFILE_SIM_reg_bank__abc_33898_n5161;
  wire REGFILE_SIM_reg_bank__abc_33898_n5162;
  wire REGFILE_SIM_reg_bank__abc_33898_n5164;
  wire REGFILE_SIM_reg_bank__abc_33898_n5165;
  wire REGFILE_SIM_reg_bank__abc_33898_n5167;
  wire REGFILE_SIM_reg_bank__abc_33898_n5168;
  wire REGFILE_SIM_reg_bank__abc_33898_n5170;
  wire REGFILE_SIM_reg_bank__abc_33898_n5171;
  wire REGFILE_SIM_reg_bank__abc_33898_n5173;
  wire REGFILE_SIM_reg_bank__abc_33898_n5174;
  wire REGFILE_SIM_reg_bank__abc_33898_n5176;
  wire REGFILE_SIM_reg_bank__abc_33898_n5177;
  wire REGFILE_SIM_reg_bank__abc_33898_n5179;
  wire REGFILE_SIM_reg_bank__abc_33898_n5180;
  wire REGFILE_SIM_reg_bank__abc_33898_n5182;
  wire REGFILE_SIM_reg_bank__abc_33898_n5183_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5185;
  wire REGFILE_SIM_reg_bank__abc_33898_n5186;
  wire REGFILE_SIM_reg_bank__abc_33898_n5188;
  wire REGFILE_SIM_reg_bank__abc_33898_n5189;
  wire REGFILE_SIM_reg_bank__abc_33898_n5191;
  wire REGFILE_SIM_reg_bank__abc_33898_n5192;
  wire REGFILE_SIM_reg_bank__abc_33898_n5194;
  wire REGFILE_SIM_reg_bank__abc_33898_n5195;
  wire REGFILE_SIM_reg_bank__abc_33898_n5197;
  wire REGFILE_SIM_reg_bank__abc_33898_n5198;
  wire REGFILE_SIM_reg_bank__abc_33898_n5200;
  wire REGFILE_SIM_reg_bank__abc_33898_n5201;
  wire REGFILE_SIM_reg_bank__abc_33898_n5203;
  wire REGFILE_SIM_reg_bank__abc_33898_n5204;
  wire REGFILE_SIM_reg_bank__abc_33898_n5206;
  wire REGFILE_SIM_reg_bank__abc_33898_n5207;
  wire REGFILE_SIM_reg_bank__abc_33898_n5209;
  wire REGFILE_SIM_reg_bank__abc_33898_n5210;
  wire REGFILE_SIM_reg_bank__abc_33898_n5212;
  wire REGFILE_SIM_reg_bank__abc_33898_n5213_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5215;
  wire REGFILE_SIM_reg_bank__abc_33898_n5216;
  wire REGFILE_SIM_reg_bank__abc_33898_n5218;
  wire REGFILE_SIM_reg_bank__abc_33898_n5219;
  wire REGFILE_SIM_reg_bank__abc_33898_n5221;
  wire REGFILE_SIM_reg_bank__abc_33898_n5222;
  wire REGFILE_SIM_reg_bank__abc_33898_n5224;
  wire REGFILE_SIM_reg_bank__abc_33898_n5225;
  wire REGFILE_SIM_reg_bank__abc_33898_n5227;
  wire REGFILE_SIM_reg_bank__abc_33898_n5228;
  wire REGFILE_SIM_reg_bank__abc_33898_n5230;
  wire REGFILE_SIM_reg_bank__abc_33898_n5231;
  wire REGFILE_SIM_reg_bank__abc_33898_n5233;
  wire REGFILE_SIM_reg_bank__abc_33898_n5234;
  wire REGFILE_SIM_reg_bank__abc_33898_n5236;
  wire REGFILE_SIM_reg_bank__abc_33898_n5237;
  wire REGFILE_SIM_reg_bank__abc_33898_n5239;
  wire REGFILE_SIM_reg_bank__abc_33898_n5240;
  wire REGFILE_SIM_reg_bank__abc_33898_n5242;
  wire REGFILE_SIM_reg_bank__abc_33898_n5243_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7;
  wire REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8;
  wire REGFILE_SIM_reg_bank__abc_33898_n5246;
  wire REGFILE_SIM_reg_bank__abc_33898_n5247;
  wire REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5248;
  wire REGFILE_SIM_reg_bank__abc_33898_n5250;
  wire REGFILE_SIM_reg_bank__abc_33898_n5251;
  wire REGFILE_SIM_reg_bank__abc_33898_n5253;
  wire REGFILE_SIM_reg_bank__abc_33898_n5254;
  wire REGFILE_SIM_reg_bank__abc_33898_n5256;
  wire REGFILE_SIM_reg_bank__abc_33898_n5257;
  wire REGFILE_SIM_reg_bank__abc_33898_n5259;
  wire REGFILE_SIM_reg_bank__abc_33898_n5260;
  wire REGFILE_SIM_reg_bank__abc_33898_n5262;
  wire REGFILE_SIM_reg_bank__abc_33898_n5263;
  wire REGFILE_SIM_reg_bank__abc_33898_n5265;
  wire REGFILE_SIM_reg_bank__abc_33898_n5266;
  wire REGFILE_SIM_reg_bank__abc_33898_n5268;
  wire REGFILE_SIM_reg_bank__abc_33898_n5269;
  wire REGFILE_SIM_reg_bank__abc_33898_n5271;
  wire REGFILE_SIM_reg_bank__abc_33898_n5272;
  wire REGFILE_SIM_reg_bank__abc_33898_n5274;
  wire REGFILE_SIM_reg_bank__abc_33898_n5275;
  wire REGFILE_SIM_reg_bank__abc_33898_n5277;
  wire REGFILE_SIM_reg_bank__abc_33898_n5278;
  wire REGFILE_SIM_reg_bank__abc_33898_n5280;
  wire REGFILE_SIM_reg_bank__abc_33898_n5281;
  wire REGFILE_SIM_reg_bank__abc_33898_n5283;
  wire REGFILE_SIM_reg_bank__abc_33898_n5284;
  wire REGFILE_SIM_reg_bank__abc_33898_n5286;
  wire REGFILE_SIM_reg_bank__abc_33898_n5287;
  wire REGFILE_SIM_reg_bank__abc_33898_n5289;
  wire REGFILE_SIM_reg_bank__abc_33898_n5290;
  wire REGFILE_SIM_reg_bank__abc_33898_n5292;
  wire REGFILE_SIM_reg_bank__abc_33898_n5293;
  wire REGFILE_SIM_reg_bank__abc_33898_n5295;
  wire REGFILE_SIM_reg_bank__abc_33898_n5296;
  wire REGFILE_SIM_reg_bank__abc_33898_n5298;
  wire REGFILE_SIM_reg_bank__abc_33898_n5299;
  wire REGFILE_SIM_reg_bank__abc_33898_n5301;
  wire REGFILE_SIM_reg_bank__abc_33898_n5302;
  wire REGFILE_SIM_reg_bank__abc_33898_n5304;
  wire REGFILE_SIM_reg_bank__abc_33898_n5305;
  wire REGFILE_SIM_reg_bank__abc_33898_n5307;
  wire REGFILE_SIM_reg_bank__abc_33898_n5308;
  wire REGFILE_SIM_reg_bank__abc_33898_n5310;
  wire REGFILE_SIM_reg_bank__abc_33898_n5311;
  wire REGFILE_SIM_reg_bank__abc_33898_n5313;
  wire REGFILE_SIM_reg_bank__abc_33898_n5314;
  wire REGFILE_SIM_reg_bank__abc_33898_n5316;
  wire REGFILE_SIM_reg_bank__abc_33898_n5317;
  wire REGFILE_SIM_reg_bank__abc_33898_n5319;
  wire REGFILE_SIM_reg_bank__abc_33898_n5320;
  wire REGFILE_SIM_reg_bank__abc_33898_n5322;
  wire REGFILE_SIM_reg_bank__abc_33898_n5323;
  wire REGFILE_SIM_reg_bank__abc_33898_n5325;
  wire REGFILE_SIM_reg_bank__abc_33898_n5326;
  wire REGFILE_SIM_reg_bank__abc_33898_n5328;
  wire REGFILE_SIM_reg_bank__abc_33898_n5329;
  wire REGFILE_SIM_reg_bank__abc_33898_n5331;
  wire REGFILE_SIM_reg_bank__abc_33898_n5332;
  wire REGFILE_SIM_reg_bank__abc_33898_n5334;
  wire REGFILE_SIM_reg_bank__abc_33898_n5335;
  wire REGFILE_SIM_reg_bank__abc_33898_n5337;
  wire REGFILE_SIM_reg_bank__abc_33898_n5338;
  wire REGFILE_SIM_reg_bank__abc_33898_n5340;
  wire REGFILE_SIM_reg_bank__abc_33898_n5341;
  wire REGFILE_SIM_reg_bank__abc_33898_n5343;
  wire REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5344;
  wire REGFILE_SIM_reg_bank__abc_33898_n5345;
  wire REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5346;
  wire REGFILE_SIM_reg_bank__abc_33898_n5348;
  wire REGFILE_SIM_reg_bank__abc_33898_n5349;
  wire REGFILE_SIM_reg_bank__abc_33898_n5351;
  wire REGFILE_SIM_reg_bank__abc_33898_n5352;
  wire REGFILE_SIM_reg_bank__abc_33898_n5354;
  wire REGFILE_SIM_reg_bank__abc_33898_n5355;
  wire REGFILE_SIM_reg_bank__abc_33898_n5357;
  wire REGFILE_SIM_reg_bank__abc_33898_n5358;
  wire REGFILE_SIM_reg_bank__abc_33898_n5360;
  wire REGFILE_SIM_reg_bank__abc_33898_n5361;
  wire REGFILE_SIM_reg_bank__abc_33898_n5363;
  wire REGFILE_SIM_reg_bank__abc_33898_n5364;
  wire REGFILE_SIM_reg_bank__abc_33898_n5366;
  wire REGFILE_SIM_reg_bank__abc_33898_n5367;
  wire REGFILE_SIM_reg_bank__abc_33898_n5369;
  wire REGFILE_SIM_reg_bank__abc_33898_n5370;
  wire REGFILE_SIM_reg_bank__abc_33898_n5372;
  wire REGFILE_SIM_reg_bank__abc_33898_n5373;
  wire REGFILE_SIM_reg_bank__abc_33898_n5375;
  wire REGFILE_SIM_reg_bank__abc_33898_n5376;
  wire REGFILE_SIM_reg_bank__abc_33898_n5378;
  wire REGFILE_SIM_reg_bank__abc_33898_n5379;
  wire REGFILE_SIM_reg_bank__abc_33898_n5381;
  wire REGFILE_SIM_reg_bank__abc_33898_n5382;
  wire REGFILE_SIM_reg_bank__abc_33898_n5384;
  wire REGFILE_SIM_reg_bank__abc_33898_n5385;
  wire REGFILE_SIM_reg_bank__abc_33898_n5387;
  wire REGFILE_SIM_reg_bank__abc_33898_n5388;
  wire REGFILE_SIM_reg_bank__abc_33898_n5390;
  wire REGFILE_SIM_reg_bank__abc_33898_n5391;
  wire REGFILE_SIM_reg_bank__abc_33898_n5393;
  wire REGFILE_SIM_reg_bank__abc_33898_n5394;
  wire REGFILE_SIM_reg_bank__abc_33898_n5396;
  wire REGFILE_SIM_reg_bank__abc_33898_n5397;
  wire REGFILE_SIM_reg_bank__abc_33898_n5399;
  wire REGFILE_SIM_reg_bank__abc_33898_n5400;
  wire REGFILE_SIM_reg_bank__abc_33898_n5402;
  wire REGFILE_SIM_reg_bank__abc_33898_n5403;
  wire REGFILE_SIM_reg_bank__abc_33898_n5405;
  wire REGFILE_SIM_reg_bank__abc_33898_n5406;
  wire REGFILE_SIM_reg_bank__abc_33898_n5408;
  wire REGFILE_SIM_reg_bank__abc_33898_n5409;
  wire REGFILE_SIM_reg_bank__abc_33898_n5411;
  wire REGFILE_SIM_reg_bank__abc_33898_n5412;
  wire REGFILE_SIM_reg_bank__abc_33898_n5414;
  wire REGFILE_SIM_reg_bank__abc_33898_n5415;
  wire REGFILE_SIM_reg_bank__abc_33898_n5417;
  wire REGFILE_SIM_reg_bank__abc_33898_n5418;
  wire REGFILE_SIM_reg_bank__abc_33898_n5420;
  wire REGFILE_SIM_reg_bank__abc_33898_n5421;
  wire REGFILE_SIM_reg_bank__abc_33898_n5423;
  wire REGFILE_SIM_reg_bank__abc_33898_n5424;
  wire REGFILE_SIM_reg_bank__abc_33898_n5426;
  wire REGFILE_SIM_reg_bank__abc_33898_n5427;
  wire REGFILE_SIM_reg_bank__abc_33898_n5429;
  wire REGFILE_SIM_reg_bank__abc_33898_n5430;
  wire REGFILE_SIM_reg_bank__abc_33898_n5432;
  wire REGFILE_SIM_reg_bank__abc_33898_n5433;
  wire REGFILE_SIM_reg_bank__abc_33898_n5435;
  wire REGFILE_SIM_reg_bank__abc_33898_n5436;
  wire REGFILE_SIM_reg_bank__abc_33898_n5438;
  wire REGFILE_SIM_reg_bank__abc_33898_n5439;
  wire REGFILE_SIM_reg_bank__abc_33898_n5441;
  wire REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5442;
  wire REGFILE_SIM_reg_bank__abc_33898_n5443;
  wire REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5444;
  wire REGFILE_SIM_reg_bank__abc_33898_n5446;
  wire REGFILE_SIM_reg_bank__abc_33898_n5447;
  wire REGFILE_SIM_reg_bank__abc_33898_n5449;
  wire REGFILE_SIM_reg_bank__abc_33898_n5450;
  wire REGFILE_SIM_reg_bank__abc_33898_n5452;
  wire REGFILE_SIM_reg_bank__abc_33898_n5453;
  wire REGFILE_SIM_reg_bank__abc_33898_n5455;
  wire REGFILE_SIM_reg_bank__abc_33898_n5456;
  wire REGFILE_SIM_reg_bank__abc_33898_n5458;
  wire REGFILE_SIM_reg_bank__abc_33898_n5459;
  wire REGFILE_SIM_reg_bank__abc_33898_n5461;
  wire REGFILE_SIM_reg_bank__abc_33898_n5462;
  wire REGFILE_SIM_reg_bank__abc_33898_n5464;
  wire REGFILE_SIM_reg_bank__abc_33898_n5465;
  wire REGFILE_SIM_reg_bank__abc_33898_n5467;
  wire REGFILE_SIM_reg_bank__abc_33898_n5468;
  wire REGFILE_SIM_reg_bank__abc_33898_n5470;
  wire REGFILE_SIM_reg_bank__abc_33898_n5471;
  wire REGFILE_SIM_reg_bank__abc_33898_n5473;
  wire REGFILE_SIM_reg_bank__abc_33898_n5474;
  wire REGFILE_SIM_reg_bank__abc_33898_n5476;
  wire REGFILE_SIM_reg_bank__abc_33898_n5477;
  wire REGFILE_SIM_reg_bank__abc_33898_n5479;
  wire REGFILE_SIM_reg_bank__abc_33898_n5480;
  wire REGFILE_SIM_reg_bank__abc_33898_n5482;
  wire REGFILE_SIM_reg_bank__abc_33898_n5483;
  wire REGFILE_SIM_reg_bank__abc_33898_n5485;
  wire REGFILE_SIM_reg_bank__abc_33898_n5486;
  wire REGFILE_SIM_reg_bank__abc_33898_n5488;
  wire REGFILE_SIM_reg_bank__abc_33898_n5489;
  wire REGFILE_SIM_reg_bank__abc_33898_n5491;
  wire REGFILE_SIM_reg_bank__abc_33898_n5492;
  wire REGFILE_SIM_reg_bank__abc_33898_n5494;
  wire REGFILE_SIM_reg_bank__abc_33898_n5495;
  wire REGFILE_SIM_reg_bank__abc_33898_n5497;
  wire REGFILE_SIM_reg_bank__abc_33898_n5498;
  wire REGFILE_SIM_reg_bank__abc_33898_n5500;
  wire REGFILE_SIM_reg_bank__abc_33898_n5501;
  wire REGFILE_SIM_reg_bank__abc_33898_n5503;
  wire REGFILE_SIM_reg_bank__abc_33898_n5504;
  wire REGFILE_SIM_reg_bank__abc_33898_n5506;
  wire REGFILE_SIM_reg_bank__abc_33898_n5507;
  wire REGFILE_SIM_reg_bank__abc_33898_n5509;
  wire REGFILE_SIM_reg_bank__abc_33898_n5510;
  wire REGFILE_SIM_reg_bank__abc_33898_n5512;
  wire REGFILE_SIM_reg_bank__abc_33898_n5513;
  wire REGFILE_SIM_reg_bank__abc_33898_n5515;
  wire REGFILE_SIM_reg_bank__abc_33898_n5516;
  wire REGFILE_SIM_reg_bank__abc_33898_n5518;
  wire REGFILE_SIM_reg_bank__abc_33898_n5519;
  wire REGFILE_SIM_reg_bank__abc_33898_n5521;
  wire REGFILE_SIM_reg_bank__abc_33898_n5522;
  wire REGFILE_SIM_reg_bank__abc_33898_n5524;
  wire REGFILE_SIM_reg_bank__abc_33898_n5525;
  wire REGFILE_SIM_reg_bank__abc_33898_n5527;
  wire REGFILE_SIM_reg_bank__abc_33898_n5528;
  wire REGFILE_SIM_reg_bank__abc_33898_n5530;
  wire REGFILE_SIM_reg_bank__abc_33898_n5531;
  wire REGFILE_SIM_reg_bank__abc_33898_n5533;
  wire REGFILE_SIM_reg_bank__abc_33898_n5534;
  wire REGFILE_SIM_reg_bank__abc_33898_n5536;
  wire REGFILE_SIM_reg_bank__abc_33898_n5537;
  wire REGFILE_SIM_reg_bank__abc_33898_n5539;
  wire REGFILE_SIM_reg_bank__abc_33898_n5540;
  wire REGFILE_SIM_reg_bank__abc_33898_n5541;
  wire REGFILE_SIM_reg_bank__abc_33898_n5542;
  wire REGFILE_SIM_reg_bank__abc_33898_n5543;
  wire REGFILE_SIM_reg_bank__abc_33898_n5544;
  wire REGFILE_SIM_reg_bank__abc_33898_n5545;
  wire REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5546;
  wire REGFILE_SIM_reg_bank__abc_33898_n5547;
  wire REGFILE_SIM_reg_bank__abc_33898_n5548;
  wire REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5549;
  wire REGFILE_SIM_reg_bank__abc_33898_n5550;
  wire REGFILE_SIM_reg_bank__abc_33898_n5551;
  wire REGFILE_SIM_reg_bank__abc_33898_n5552;
  wire REGFILE_SIM_reg_bank__abc_33898_n5553;
  wire REGFILE_SIM_reg_bank__abc_33898_n5554;
  wire REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5555;
  wire REGFILE_SIM_reg_bank__abc_33898_n5556;
  wire REGFILE_SIM_reg_bank__abc_33898_n5557;
  wire REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5558;
  wire REGFILE_SIM_reg_bank__abc_33898_n5559;
  wire REGFILE_SIM_reg_bank__abc_33898_n5560;
  wire REGFILE_SIM_reg_bank__abc_33898_n5561;
  wire REGFILE_SIM_reg_bank__abc_33898_n5562;
  wire REGFILE_SIM_reg_bank__abc_33898_n5563;
  wire REGFILE_SIM_reg_bank__abc_33898_n5564;
  wire REGFILE_SIM_reg_bank__abc_33898_n5565;
  wire REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5566;
  wire REGFILE_SIM_reg_bank__abc_33898_n5567;
  wire REGFILE_SIM_reg_bank__abc_33898_n5568;
  wire REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5569;
  wire REGFILE_SIM_reg_bank__abc_33898_n5570;
  wire REGFILE_SIM_reg_bank__abc_33898_n5571;
  wire REGFILE_SIM_reg_bank__abc_33898_n5572;
  wire REGFILE_SIM_reg_bank__abc_33898_n5573;
  wire REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5574;
  wire REGFILE_SIM_reg_bank__abc_33898_n5575;
  wire REGFILE_SIM_reg_bank__abc_33898_n5576;
  wire REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5577;
  wire REGFILE_SIM_reg_bank__abc_33898_n5578;
  wire REGFILE_SIM_reg_bank__abc_33898_n5579;
  wire REGFILE_SIM_reg_bank__abc_33898_n5580;
  wire REGFILE_SIM_reg_bank__abc_33898_n5581;
  wire REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5582;
  wire REGFILE_SIM_reg_bank__abc_33898_n5583;
  wire REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5584;
  wire REGFILE_SIM_reg_bank__abc_33898_n5585;
  wire REGFILE_SIM_reg_bank__abc_33898_n5586;
  wire REGFILE_SIM_reg_bank__abc_33898_n5587;
  wire REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5588;
  wire REGFILE_SIM_reg_bank__abc_33898_n5589;
  wire REGFILE_SIM_reg_bank__abc_33898_n5590;
  wire REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5591;
  wire REGFILE_SIM_reg_bank__abc_33898_n5592;
  wire REGFILE_SIM_reg_bank__abc_33898_n5593;
  wire REGFILE_SIM_reg_bank__abc_33898_n5594;
  wire REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5595;
  wire REGFILE_SIM_reg_bank__abc_33898_n5596;
  wire REGFILE_SIM_reg_bank__abc_33898_n5597;
  wire REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5598;
  wire REGFILE_SIM_reg_bank__abc_33898_n5599;
  wire REGFILE_SIM_reg_bank__abc_33898_n5600;
  wire REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5601;
  wire REGFILE_SIM_reg_bank__abc_33898_n5602;
  wire REGFILE_SIM_reg_bank__abc_33898_n5603;
  wire REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5604;
  wire REGFILE_SIM_reg_bank__abc_33898_n5605;
  wire REGFILE_SIM_reg_bank__abc_33898_n5606;
  wire REGFILE_SIM_reg_bank__abc_33898_n5607;
  wire REGFILE_SIM_reg_bank__abc_33898_n5608;
  wire REGFILE_SIM_reg_bank__abc_33898_n5609;
  wire REGFILE_SIM_reg_bank__abc_33898_n5610;
  wire REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5611;
  wire REGFILE_SIM_reg_bank__abc_33898_n5612;
  wire REGFILE_SIM_reg_bank__abc_33898_n5613;
  wire REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5614;
  wire REGFILE_SIM_reg_bank__abc_33898_n5615;
  wire REGFILE_SIM_reg_bank__abc_33898_n5616;
  wire REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5617;
  wire REGFILE_SIM_reg_bank__abc_33898_n5618;
  wire REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5619;
  wire REGFILE_SIM_reg_bank__abc_33898_n5620;
  wire REGFILE_SIM_reg_bank__abc_33898_n5621;
  wire REGFILE_SIM_reg_bank__abc_33898_n5622;
  wire REGFILE_SIM_reg_bank__abc_33898_n5623;
  wire REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5624;
  wire REGFILE_SIM_reg_bank__abc_33898_n5625;
  wire REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5626;
  wire REGFILE_SIM_reg_bank__abc_33898_n5627;
  wire REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5628;
  wire REGFILE_SIM_reg_bank__abc_33898_n5629;
  wire REGFILE_SIM_reg_bank__abc_33898_n5630;
  wire REGFILE_SIM_reg_bank__abc_33898_n5631;
  wire REGFILE_SIM_reg_bank__abc_33898_n5632;
  wire REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5633;
  wire REGFILE_SIM_reg_bank__abc_33898_n5634;
  wire REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5635;
  wire REGFILE_SIM_reg_bank__abc_33898_n5636;
  wire REGFILE_SIM_reg_bank__abc_33898_n5637;
  wire REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5638;
  wire REGFILE_SIM_reg_bank__abc_33898_n5639;
  wire REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5640;
  wire REGFILE_SIM_reg_bank__abc_33898_n5641;
  wire REGFILE_SIM_reg_bank__abc_33898_n5642;
  wire REGFILE_SIM_reg_bank__abc_33898_n5643;
  wire REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5644;
  wire REGFILE_SIM_reg_bank__abc_33898_n5645;
  wire REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5646;
  wire REGFILE_SIM_reg_bank__abc_33898_n5647;
  wire REGFILE_SIM_reg_bank__abc_33898_n5648;
  wire REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5649;
  wire REGFILE_SIM_reg_bank__abc_33898_n5650;
  wire REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n5651;
  wire REGFILE_SIM_reg_bank__abc_33898_n5652;
  wire REGFILE_SIM_reg_bank__abc_33898_n5653;
  wire REGFILE_SIM_reg_bank__abc_33898_n5654;
  wire REGFILE_SIM_reg_bank__abc_33898_n5655;
  wire REGFILE_SIM_reg_bank__abc_33898_n5657;
  wire REGFILE_SIM_reg_bank__abc_33898_n5658;
  wire REGFILE_SIM_reg_bank__abc_33898_n5659;
  wire REGFILE_SIM_reg_bank__abc_33898_n5660;
  wire REGFILE_SIM_reg_bank__abc_33898_n5661;
  wire REGFILE_SIM_reg_bank__abc_33898_n5662;
  wire REGFILE_SIM_reg_bank__abc_33898_n5663;
  wire REGFILE_SIM_reg_bank__abc_33898_n5664;
  wire REGFILE_SIM_reg_bank__abc_33898_n5665;
  wire REGFILE_SIM_reg_bank__abc_33898_n5666;
  wire REGFILE_SIM_reg_bank__abc_33898_n5667;
  wire REGFILE_SIM_reg_bank__abc_33898_n5668;
  wire REGFILE_SIM_reg_bank__abc_33898_n5669;
  wire REGFILE_SIM_reg_bank__abc_33898_n5670;
  wire REGFILE_SIM_reg_bank__abc_33898_n5671;
  wire REGFILE_SIM_reg_bank__abc_33898_n5672;
  wire REGFILE_SIM_reg_bank__abc_33898_n5673;
  wire REGFILE_SIM_reg_bank__abc_33898_n5674;
  wire REGFILE_SIM_reg_bank__abc_33898_n5675;
  wire REGFILE_SIM_reg_bank__abc_33898_n5676;
  wire REGFILE_SIM_reg_bank__abc_33898_n5677;
  wire REGFILE_SIM_reg_bank__abc_33898_n5678;
  wire REGFILE_SIM_reg_bank__abc_33898_n5679;
  wire REGFILE_SIM_reg_bank__abc_33898_n5680;
  wire REGFILE_SIM_reg_bank__abc_33898_n5681;
  wire REGFILE_SIM_reg_bank__abc_33898_n5682;
  wire REGFILE_SIM_reg_bank__abc_33898_n5683;
  wire REGFILE_SIM_reg_bank__abc_33898_n5684;
  wire REGFILE_SIM_reg_bank__abc_33898_n5685;
  wire REGFILE_SIM_reg_bank__abc_33898_n5686;
  wire REGFILE_SIM_reg_bank__abc_33898_n5687;
  wire REGFILE_SIM_reg_bank__abc_33898_n5688;
  wire REGFILE_SIM_reg_bank__abc_33898_n5689;
  wire REGFILE_SIM_reg_bank__abc_33898_n5690;
  wire REGFILE_SIM_reg_bank__abc_33898_n5691;
  wire REGFILE_SIM_reg_bank__abc_33898_n5692;
  wire REGFILE_SIM_reg_bank__abc_33898_n5693;
  wire REGFILE_SIM_reg_bank__abc_33898_n5694;
  wire REGFILE_SIM_reg_bank__abc_33898_n5695;
  wire REGFILE_SIM_reg_bank__abc_33898_n5696;
  wire REGFILE_SIM_reg_bank__abc_33898_n5697;
  wire REGFILE_SIM_reg_bank__abc_33898_n5698;
  wire REGFILE_SIM_reg_bank__abc_33898_n5699;
  wire REGFILE_SIM_reg_bank__abc_33898_n5700;
  wire REGFILE_SIM_reg_bank__abc_33898_n5701;
  wire REGFILE_SIM_reg_bank__abc_33898_n5702;
  wire REGFILE_SIM_reg_bank__abc_33898_n5703;
  wire REGFILE_SIM_reg_bank__abc_33898_n5704;
  wire REGFILE_SIM_reg_bank__abc_33898_n5705;
  wire REGFILE_SIM_reg_bank__abc_33898_n5706;
  wire REGFILE_SIM_reg_bank__abc_33898_n5707;
  wire REGFILE_SIM_reg_bank__abc_33898_n5708;
  wire REGFILE_SIM_reg_bank__abc_33898_n5709;
  wire REGFILE_SIM_reg_bank__abc_33898_n5710;
  wire REGFILE_SIM_reg_bank__abc_33898_n5711;
  wire REGFILE_SIM_reg_bank__abc_33898_n5712;
  wire REGFILE_SIM_reg_bank__abc_33898_n5713;
  wire REGFILE_SIM_reg_bank__abc_33898_n5714;
  wire REGFILE_SIM_reg_bank__abc_33898_n5715;
  wire REGFILE_SIM_reg_bank__abc_33898_n5716;
  wire REGFILE_SIM_reg_bank__abc_33898_n5718;
  wire REGFILE_SIM_reg_bank__abc_33898_n5719;
  wire REGFILE_SIM_reg_bank__abc_33898_n5720;
  wire REGFILE_SIM_reg_bank__abc_33898_n5721;
  wire REGFILE_SIM_reg_bank__abc_33898_n5722;
  wire REGFILE_SIM_reg_bank__abc_33898_n5723;
  wire REGFILE_SIM_reg_bank__abc_33898_n5724;
  wire REGFILE_SIM_reg_bank__abc_33898_n5725;
  wire REGFILE_SIM_reg_bank__abc_33898_n5726;
  wire REGFILE_SIM_reg_bank__abc_33898_n5727;
  wire REGFILE_SIM_reg_bank__abc_33898_n5728;
  wire REGFILE_SIM_reg_bank__abc_33898_n5729;
  wire REGFILE_SIM_reg_bank__abc_33898_n5730;
  wire REGFILE_SIM_reg_bank__abc_33898_n5731;
  wire REGFILE_SIM_reg_bank__abc_33898_n5732;
  wire REGFILE_SIM_reg_bank__abc_33898_n5733;
  wire REGFILE_SIM_reg_bank__abc_33898_n5734;
  wire REGFILE_SIM_reg_bank__abc_33898_n5735;
  wire REGFILE_SIM_reg_bank__abc_33898_n5736;
  wire REGFILE_SIM_reg_bank__abc_33898_n5737;
  wire REGFILE_SIM_reg_bank__abc_33898_n5738;
  wire REGFILE_SIM_reg_bank__abc_33898_n5739;
  wire REGFILE_SIM_reg_bank__abc_33898_n5740;
  wire REGFILE_SIM_reg_bank__abc_33898_n5741;
  wire REGFILE_SIM_reg_bank__abc_33898_n5742;
  wire REGFILE_SIM_reg_bank__abc_33898_n5743;
  wire REGFILE_SIM_reg_bank__abc_33898_n5744;
  wire REGFILE_SIM_reg_bank__abc_33898_n5745;
  wire REGFILE_SIM_reg_bank__abc_33898_n5746;
  wire REGFILE_SIM_reg_bank__abc_33898_n5747;
  wire REGFILE_SIM_reg_bank__abc_33898_n5748;
  wire REGFILE_SIM_reg_bank__abc_33898_n5749;
  wire REGFILE_SIM_reg_bank__abc_33898_n5750;
  wire REGFILE_SIM_reg_bank__abc_33898_n5751;
  wire REGFILE_SIM_reg_bank__abc_33898_n5752;
  wire REGFILE_SIM_reg_bank__abc_33898_n5753;
  wire REGFILE_SIM_reg_bank__abc_33898_n5754;
  wire REGFILE_SIM_reg_bank__abc_33898_n5755;
  wire REGFILE_SIM_reg_bank__abc_33898_n5756;
  wire REGFILE_SIM_reg_bank__abc_33898_n5757;
  wire REGFILE_SIM_reg_bank__abc_33898_n5758;
  wire REGFILE_SIM_reg_bank__abc_33898_n5759;
  wire REGFILE_SIM_reg_bank__abc_33898_n5760;
  wire REGFILE_SIM_reg_bank__abc_33898_n5761;
  wire REGFILE_SIM_reg_bank__abc_33898_n5762;
  wire REGFILE_SIM_reg_bank__abc_33898_n5763;
  wire REGFILE_SIM_reg_bank__abc_33898_n5764;
  wire REGFILE_SIM_reg_bank__abc_33898_n5765;
  wire REGFILE_SIM_reg_bank__abc_33898_n5766;
  wire REGFILE_SIM_reg_bank__abc_33898_n5767;
  wire REGFILE_SIM_reg_bank__abc_33898_n5768;
  wire REGFILE_SIM_reg_bank__abc_33898_n5769;
  wire REGFILE_SIM_reg_bank__abc_33898_n5770;
  wire REGFILE_SIM_reg_bank__abc_33898_n5771;
  wire REGFILE_SIM_reg_bank__abc_33898_n5772;
  wire REGFILE_SIM_reg_bank__abc_33898_n5773;
  wire REGFILE_SIM_reg_bank__abc_33898_n5774;
  wire REGFILE_SIM_reg_bank__abc_33898_n5775;
  wire REGFILE_SIM_reg_bank__abc_33898_n5776;
  wire REGFILE_SIM_reg_bank__abc_33898_n5777;
  wire REGFILE_SIM_reg_bank__abc_33898_n5779;
  wire REGFILE_SIM_reg_bank__abc_33898_n5780;
  wire REGFILE_SIM_reg_bank__abc_33898_n5781;
  wire REGFILE_SIM_reg_bank__abc_33898_n5782;
  wire REGFILE_SIM_reg_bank__abc_33898_n5783;
  wire REGFILE_SIM_reg_bank__abc_33898_n5784;
  wire REGFILE_SIM_reg_bank__abc_33898_n5785;
  wire REGFILE_SIM_reg_bank__abc_33898_n5786;
  wire REGFILE_SIM_reg_bank__abc_33898_n5787;
  wire REGFILE_SIM_reg_bank__abc_33898_n5788;
  wire REGFILE_SIM_reg_bank__abc_33898_n5789;
  wire REGFILE_SIM_reg_bank__abc_33898_n5790;
  wire REGFILE_SIM_reg_bank__abc_33898_n5791;
  wire REGFILE_SIM_reg_bank__abc_33898_n5792;
  wire REGFILE_SIM_reg_bank__abc_33898_n5793;
  wire REGFILE_SIM_reg_bank__abc_33898_n5794;
  wire REGFILE_SIM_reg_bank__abc_33898_n5795;
  wire REGFILE_SIM_reg_bank__abc_33898_n5796;
  wire REGFILE_SIM_reg_bank__abc_33898_n5797;
  wire REGFILE_SIM_reg_bank__abc_33898_n5798;
  wire REGFILE_SIM_reg_bank__abc_33898_n5799;
  wire REGFILE_SIM_reg_bank__abc_33898_n5800;
  wire REGFILE_SIM_reg_bank__abc_33898_n5801;
  wire REGFILE_SIM_reg_bank__abc_33898_n5802;
  wire REGFILE_SIM_reg_bank__abc_33898_n5803;
  wire REGFILE_SIM_reg_bank__abc_33898_n5804;
  wire REGFILE_SIM_reg_bank__abc_33898_n5805;
  wire REGFILE_SIM_reg_bank__abc_33898_n5806;
  wire REGFILE_SIM_reg_bank__abc_33898_n5807;
  wire REGFILE_SIM_reg_bank__abc_33898_n5808;
  wire REGFILE_SIM_reg_bank__abc_33898_n5809;
  wire REGFILE_SIM_reg_bank__abc_33898_n5810;
  wire REGFILE_SIM_reg_bank__abc_33898_n5811;
  wire REGFILE_SIM_reg_bank__abc_33898_n5812;
  wire REGFILE_SIM_reg_bank__abc_33898_n5813;
  wire REGFILE_SIM_reg_bank__abc_33898_n5814;
  wire REGFILE_SIM_reg_bank__abc_33898_n5815;
  wire REGFILE_SIM_reg_bank__abc_33898_n5816;
  wire REGFILE_SIM_reg_bank__abc_33898_n5817;
  wire REGFILE_SIM_reg_bank__abc_33898_n5818;
  wire REGFILE_SIM_reg_bank__abc_33898_n5819;
  wire REGFILE_SIM_reg_bank__abc_33898_n5820;
  wire REGFILE_SIM_reg_bank__abc_33898_n5821;
  wire REGFILE_SIM_reg_bank__abc_33898_n5822;
  wire REGFILE_SIM_reg_bank__abc_33898_n5823;
  wire REGFILE_SIM_reg_bank__abc_33898_n5824;
  wire REGFILE_SIM_reg_bank__abc_33898_n5825;
  wire REGFILE_SIM_reg_bank__abc_33898_n5826;
  wire REGFILE_SIM_reg_bank__abc_33898_n5827;
  wire REGFILE_SIM_reg_bank__abc_33898_n5828;
  wire REGFILE_SIM_reg_bank__abc_33898_n5829;
  wire REGFILE_SIM_reg_bank__abc_33898_n5830;
  wire REGFILE_SIM_reg_bank__abc_33898_n5831;
  wire REGFILE_SIM_reg_bank__abc_33898_n5832;
  wire REGFILE_SIM_reg_bank__abc_33898_n5833;
  wire REGFILE_SIM_reg_bank__abc_33898_n5834;
  wire REGFILE_SIM_reg_bank__abc_33898_n5835;
  wire REGFILE_SIM_reg_bank__abc_33898_n5836;
  wire REGFILE_SIM_reg_bank__abc_33898_n5837;
  wire REGFILE_SIM_reg_bank__abc_33898_n5838;
  wire REGFILE_SIM_reg_bank__abc_33898_n5840;
  wire REGFILE_SIM_reg_bank__abc_33898_n5841;
  wire REGFILE_SIM_reg_bank__abc_33898_n5842;
  wire REGFILE_SIM_reg_bank__abc_33898_n5843;
  wire REGFILE_SIM_reg_bank__abc_33898_n5844;
  wire REGFILE_SIM_reg_bank__abc_33898_n5845;
  wire REGFILE_SIM_reg_bank__abc_33898_n5846;
  wire REGFILE_SIM_reg_bank__abc_33898_n5847;
  wire REGFILE_SIM_reg_bank__abc_33898_n5848;
  wire REGFILE_SIM_reg_bank__abc_33898_n5849;
  wire REGFILE_SIM_reg_bank__abc_33898_n5850;
  wire REGFILE_SIM_reg_bank__abc_33898_n5851;
  wire REGFILE_SIM_reg_bank__abc_33898_n5852;
  wire REGFILE_SIM_reg_bank__abc_33898_n5853;
  wire REGFILE_SIM_reg_bank__abc_33898_n5854;
  wire REGFILE_SIM_reg_bank__abc_33898_n5855;
  wire REGFILE_SIM_reg_bank__abc_33898_n5856;
  wire REGFILE_SIM_reg_bank__abc_33898_n5857;
  wire REGFILE_SIM_reg_bank__abc_33898_n5858;
  wire REGFILE_SIM_reg_bank__abc_33898_n5859;
  wire REGFILE_SIM_reg_bank__abc_33898_n5860;
  wire REGFILE_SIM_reg_bank__abc_33898_n5861;
  wire REGFILE_SIM_reg_bank__abc_33898_n5862;
  wire REGFILE_SIM_reg_bank__abc_33898_n5863;
  wire REGFILE_SIM_reg_bank__abc_33898_n5864;
  wire REGFILE_SIM_reg_bank__abc_33898_n5865;
  wire REGFILE_SIM_reg_bank__abc_33898_n5866;
  wire REGFILE_SIM_reg_bank__abc_33898_n5867;
  wire REGFILE_SIM_reg_bank__abc_33898_n5868;
  wire REGFILE_SIM_reg_bank__abc_33898_n5869;
  wire REGFILE_SIM_reg_bank__abc_33898_n5870;
  wire REGFILE_SIM_reg_bank__abc_33898_n5871;
  wire REGFILE_SIM_reg_bank__abc_33898_n5872;
  wire REGFILE_SIM_reg_bank__abc_33898_n5873;
  wire REGFILE_SIM_reg_bank__abc_33898_n5874;
  wire REGFILE_SIM_reg_bank__abc_33898_n5875;
  wire REGFILE_SIM_reg_bank__abc_33898_n5876;
  wire REGFILE_SIM_reg_bank__abc_33898_n5877;
  wire REGFILE_SIM_reg_bank__abc_33898_n5878;
  wire REGFILE_SIM_reg_bank__abc_33898_n5879;
  wire REGFILE_SIM_reg_bank__abc_33898_n5880;
  wire REGFILE_SIM_reg_bank__abc_33898_n5881;
  wire REGFILE_SIM_reg_bank__abc_33898_n5882;
  wire REGFILE_SIM_reg_bank__abc_33898_n5883;
  wire REGFILE_SIM_reg_bank__abc_33898_n5884;
  wire REGFILE_SIM_reg_bank__abc_33898_n5885;
  wire REGFILE_SIM_reg_bank__abc_33898_n5886;
  wire REGFILE_SIM_reg_bank__abc_33898_n5887;
  wire REGFILE_SIM_reg_bank__abc_33898_n5888;
  wire REGFILE_SIM_reg_bank__abc_33898_n5889;
  wire REGFILE_SIM_reg_bank__abc_33898_n5890;
  wire REGFILE_SIM_reg_bank__abc_33898_n5891;
  wire REGFILE_SIM_reg_bank__abc_33898_n5892;
  wire REGFILE_SIM_reg_bank__abc_33898_n5893;
  wire REGFILE_SIM_reg_bank__abc_33898_n5894;
  wire REGFILE_SIM_reg_bank__abc_33898_n5895;
  wire REGFILE_SIM_reg_bank__abc_33898_n5896;
  wire REGFILE_SIM_reg_bank__abc_33898_n5897;
  wire REGFILE_SIM_reg_bank__abc_33898_n5898;
  wire REGFILE_SIM_reg_bank__abc_33898_n5899;
  wire REGFILE_SIM_reg_bank__abc_33898_n5901;
  wire REGFILE_SIM_reg_bank__abc_33898_n5902;
  wire REGFILE_SIM_reg_bank__abc_33898_n5903;
  wire REGFILE_SIM_reg_bank__abc_33898_n5904;
  wire REGFILE_SIM_reg_bank__abc_33898_n5905;
  wire REGFILE_SIM_reg_bank__abc_33898_n5906;
  wire REGFILE_SIM_reg_bank__abc_33898_n5907;
  wire REGFILE_SIM_reg_bank__abc_33898_n5908;
  wire REGFILE_SIM_reg_bank__abc_33898_n5909;
  wire REGFILE_SIM_reg_bank__abc_33898_n5910;
  wire REGFILE_SIM_reg_bank__abc_33898_n5911;
  wire REGFILE_SIM_reg_bank__abc_33898_n5912;
  wire REGFILE_SIM_reg_bank__abc_33898_n5913;
  wire REGFILE_SIM_reg_bank__abc_33898_n5914;
  wire REGFILE_SIM_reg_bank__abc_33898_n5915;
  wire REGFILE_SIM_reg_bank__abc_33898_n5916;
  wire REGFILE_SIM_reg_bank__abc_33898_n5917;
  wire REGFILE_SIM_reg_bank__abc_33898_n5918;
  wire REGFILE_SIM_reg_bank__abc_33898_n5919;
  wire REGFILE_SIM_reg_bank__abc_33898_n5920;
  wire REGFILE_SIM_reg_bank__abc_33898_n5921;
  wire REGFILE_SIM_reg_bank__abc_33898_n5922;
  wire REGFILE_SIM_reg_bank__abc_33898_n5923;
  wire REGFILE_SIM_reg_bank__abc_33898_n5924;
  wire REGFILE_SIM_reg_bank__abc_33898_n5925;
  wire REGFILE_SIM_reg_bank__abc_33898_n5926;
  wire REGFILE_SIM_reg_bank__abc_33898_n5927;
  wire REGFILE_SIM_reg_bank__abc_33898_n5928;
  wire REGFILE_SIM_reg_bank__abc_33898_n5929;
  wire REGFILE_SIM_reg_bank__abc_33898_n5930;
  wire REGFILE_SIM_reg_bank__abc_33898_n5931;
  wire REGFILE_SIM_reg_bank__abc_33898_n5932;
  wire REGFILE_SIM_reg_bank__abc_33898_n5933;
  wire REGFILE_SIM_reg_bank__abc_33898_n5934;
  wire REGFILE_SIM_reg_bank__abc_33898_n5935;
  wire REGFILE_SIM_reg_bank__abc_33898_n5936;
  wire REGFILE_SIM_reg_bank__abc_33898_n5937;
  wire REGFILE_SIM_reg_bank__abc_33898_n5938;
  wire REGFILE_SIM_reg_bank__abc_33898_n5939;
  wire REGFILE_SIM_reg_bank__abc_33898_n5940;
  wire REGFILE_SIM_reg_bank__abc_33898_n5941;
  wire REGFILE_SIM_reg_bank__abc_33898_n5942;
  wire REGFILE_SIM_reg_bank__abc_33898_n5943;
  wire REGFILE_SIM_reg_bank__abc_33898_n5944;
  wire REGFILE_SIM_reg_bank__abc_33898_n5945;
  wire REGFILE_SIM_reg_bank__abc_33898_n5946;
  wire REGFILE_SIM_reg_bank__abc_33898_n5947;
  wire REGFILE_SIM_reg_bank__abc_33898_n5948;
  wire REGFILE_SIM_reg_bank__abc_33898_n5949;
  wire REGFILE_SIM_reg_bank__abc_33898_n5950;
  wire REGFILE_SIM_reg_bank__abc_33898_n5951;
  wire REGFILE_SIM_reg_bank__abc_33898_n5952;
  wire REGFILE_SIM_reg_bank__abc_33898_n5953;
  wire REGFILE_SIM_reg_bank__abc_33898_n5954;
  wire REGFILE_SIM_reg_bank__abc_33898_n5955;
  wire REGFILE_SIM_reg_bank__abc_33898_n5956;
  wire REGFILE_SIM_reg_bank__abc_33898_n5957;
  wire REGFILE_SIM_reg_bank__abc_33898_n5958;
  wire REGFILE_SIM_reg_bank__abc_33898_n5959;
  wire REGFILE_SIM_reg_bank__abc_33898_n5960;
  wire REGFILE_SIM_reg_bank__abc_33898_n5962;
  wire REGFILE_SIM_reg_bank__abc_33898_n5963;
  wire REGFILE_SIM_reg_bank__abc_33898_n5964;
  wire REGFILE_SIM_reg_bank__abc_33898_n5965;
  wire REGFILE_SIM_reg_bank__abc_33898_n5966;
  wire REGFILE_SIM_reg_bank__abc_33898_n5967;
  wire REGFILE_SIM_reg_bank__abc_33898_n5968;
  wire REGFILE_SIM_reg_bank__abc_33898_n5969;
  wire REGFILE_SIM_reg_bank__abc_33898_n5970;
  wire REGFILE_SIM_reg_bank__abc_33898_n5971;
  wire REGFILE_SIM_reg_bank__abc_33898_n5972;
  wire REGFILE_SIM_reg_bank__abc_33898_n5973;
  wire REGFILE_SIM_reg_bank__abc_33898_n5974;
  wire REGFILE_SIM_reg_bank__abc_33898_n5975;
  wire REGFILE_SIM_reg_bank__abc_33898_n5976;
  wire REGFILE_SIM_reg_bank__abc_33898_n5977;
  wire REGFILE_SIM_reg_bank__abc_33898_n5978;
  wire REGFILE_SIM_reg_bank__abc_33898_n5979;
  wire REGFILE_SIM_reg_bank__abc_33898_n5980;
  wire REGFILE_SIM_reg_bank__abc_33898_n5981;
  wire REGFILE_SIM_reg_bank__abc_33898_n5982;
  wire REGFILE_SIM_reg_bank__abc_33898_n5983;
  wire REGFILE_SIM_reg_bank__abc_33898_n5984;
  wire REGFILE_SIM_reg_bank__abc_33898_n5985;
  wire REGFILE_SIM_reg_bank__abc_33898_n5986;
  wire REGFILE_SIM_reg_bank__abc_33898_n5987;
  wire REGFILE_SIM_reg_bank__abc_33898_n5988;
  wire REGFILE_SIM_reg_bank__abc_33898_n5989;
  wire REGFILE_SIM_reg_bank__abc_33898_n5990;
  wire REGFILE_SIM_reg_bank__abc_33898_n5991;
  wire REGFILE_SIM_reg_bank__abc_33898_n5992;
  wire REGFILE_SIM_reg_bank__abc_33898_n5993;
  wire REGFILE_SIM_reg_bank__abc_33898_n5994;
  wire REGFILE_SIM_reg_bank__abc_33898_n5995;
  wire REGFILE_SIM_reg_bank__abc_33898_n5996;
  wire REGFILE_SIM_reg_bank__abc_33898_n5997;
  wire REGFILE_SIM_reg_bank__abc_33898_n5998;
  wire REGFILE_SIM_reg_bank__abc_33898_n5999;
  wire REGFILE_SIM_reg_bank__abc_33898_n6000;
  wire REGFILE_SIM_reg_bank__abc_33898_n6001;
  wire REGFILE_SIM_reg_bank__abc_33898_n6002;
  wire REGFILE_SIM_reg_bank__abc_33898_n6003;
  wire REGFILE_SIM_reg_bank__abc_33898_n6004;
  wire REGFILE_SIM_reg_bank__abc_33898_n6005;
  wire REGFILE_SIM_reg_bank__abc_33898_n6006;
  wire REGFILE_SIM_reg_bank__abc_33898_n6007;
  wire REGFILE_SIM_reg_bank__abc_33898_n6008;
  wire REGFILE_SIM_reg_bank__abc_33898_n6009;
  wire REGFILE_SIM_reg_bank__abc_33898_n6010;
  wire REGFILE_SIM_reg_bank__abc_33898_n6011;
  wire REGFILE_SIM_reg_bank__abc_33898_n6012;
  wire REGFILE_SIM_reg_bank__abc_33898_n6013;
  wire REGFILE_SIM_reg_bank__abc_33898_n6014;
  wire REGFILE_SIM_reg_bank__abc_33898_n6015;
  wire REGFILE_SIM_reg_bank__abc_33898_n6016;
  wire REGFILE_SIM_reg_bank__abc_33898_n6017;
  wire REGFILE_SIM_reg_bank__abc_33898_n6018;
  wire REGFILE_SIM_reg_bank__abc_33898_n6019;
  wire REGFILE_SIM_reg_bank__abc_33898_n6020;
  wire REGFILE_SIM_reg_bank__abc_33898_n6021;
  wire REGFILE_SIM_reg_bank__abc_33898_n6023;
  wire REGFILE_SIM_reg_bank__abc_33898_n6024;
  wire REGFILE_SIM_reg_bank__abc_33898_n6025;
  wire REGFILE_SIM_reg_bank__abc_33898_n6026;
  wire REGFILE_SIM_reg_bank__abc_33898_n6027;
  wire REGFILE_SIM_reg_bank__abc_33898_n6028;
  wire REGFILE_SIM_reg_bank__abc_33898_n6029;
  wire REGFILE_SIM_reg_bank__abc_33898_n6030;
  wire REGFILE_SIM_reg_bank__abc_33898_n6031;
  wire REGFILE_SIM_reg_bank__abc_33898_n6032;
  wire REGFILE_SIM_reg_bank__abc_33898_n6033;
  wire REGFILE_SIM_reg_bank__abc_33898_n6034;
  wire REGFILE_SIM_reg_bank__abc_33898_n6035;
  wire REGFILE_SIM_reg_bank__abc_33898_n6036;
  wire REGFILE_SIM_reg_bank__abc_33898_n6037;
  wire REGFILE_SIM_reg_bank__abc_33898_n6038;
  wire REGFILE_SIM_reg_bank__abc_33898_n6039;
  wire REGFILE_SIM_reg_bank__abc_33898_n6040;
  wire REGFILE_SIM_reg_bank__abc_33898_n6041;
  wire REGFILE_SIM_reg_bank__abc_33898_n6042;
  wire REGFILE_SIM_reg_bank__abc_33898_n6043;
  wire REGFILE_SIM_reg_bank__abc_33898_n6044;
  wire REGFILE_SIM_reg_bank__abc_33898_n6045;
  wire REGFILE_SIM_reg_bank__abc_33898_n6046;
  wire REGFILE_SIM_reg_bank__abc_33898_n6047;
  wire REGFILE_SIM_reg_bank__abc_33898_n6048;
  wire REGFILE_SIM_reg_bank__abc_33898_n6049;
  wire REGFILE_SIM_reg_bank__abc_33898_n6050;
  wire REGFILE_SIM_reg_bank__abc_33898_n6051;
  wire REGFILE_SIM_reg_bank__abc_33898_n6052;
  wire REGFILE_SIM_reg_bank__abc_33898_n6053;
  wire REGFILE_SIM_reg_bank__abc_33898_n6054;
  wire REGFILE_SIM_reg_bank__abc_33898_n6055;
  wire REGFILE_SIM_reg_bank__abc_33898_n6056;
  wire REGFILE_SIM_reg_bank__abc_33898_n6057;
  wire REGFILE_SIM_reg_bank__abc_33898_n6058;
  wire REGFILE_SIM_reg_bank__abc_33898_n6059;
  wire REGFILE_SIM_reg_bank__abc_33898_n6060;
  wire REGFILE_SIM_reg_bank__abc_33898_n6061;
  wire REGFILE_SIM_reg_bank__abc_33898_n6062;
  wire REGFILE_SIM_reg_bank__abc_33898_n6063;
  wire REGFILE_SIM_reg_bank__abc_33898_n6064;
  wire REGFILE_SIM_reg_bank__abc_33898_n6065;
  wire REGFILE_SIM_reg_bank__abc_33898_n6066;
  wire REGFILE_SIM_reg_bank__abc_33898_n6067;
  wire REGFILE_SIM_reg_bank__abc_33898_n6068;
  wire REGFILE_SIM_reg_bank__abc_33898_n6069;
  wire REGFILE_SIM_reg_bank__abc_33898_n6070;
  wire REGFILE_SIM_reg_bank__abc_33898_n6071;
  wire REGFILE_SIM_reg_bank__abc_33898_n6072;
  wire REGFILE_SIM_reg_bank__abc_33898_n6073;
  wire REGFILE_SIM_reg_bank__abc_33898_n6074;
  wire REGFILE_SIM_reg_bank__abc_33898_n6075;
  wire REGFILE_SIM_reg_bank__abc_33898_n6076;
  wire REGFILE_SIM_reg_bank__abc_33898_n6077;
  wire REGFILE_SIM_reg_bank__abc_33898_n6078;
  wire REGFILE_SIM_reg_bank__abc_33898_n6079;
  wire REGFILE_SIM_reg_bank__abc_33898_n6080;
  wire REGFILE_SIM_reg_bank__abc_33898_n6081;
  wire REGFILE_SIM_reg_bank__abc_33898_n6082;
  wire REGFILE_SIM_reg_bank__abc_33898_n6084;
  wire REGFILE_SIM_reg_bank__abc_33898_n6085;
  wire REGFILE_SIM_reg_bank__abc_33898_n6086;
  wire REGFILE_SIM_reg_bank__abc_33898_n6087;
  wire REGFILE_SIM_reg_bank__abc_33898_n6088;
  wire REGFILE_SIM_reg_bank__abc_33898_n6089;
  wire REGFILE_SIM_reg_bank__abc_33898_n6090;
  wire REGFILE_SIM_reg_bank__abc_33898_n6091;
  wire REGFILE_SIM_reg_bank__abc_33898_n6092;
  wire REGFILE_SIM_reg_bank__abc_33898_n6093;
  wire REGFILE_SIM_reg_bank__abc_33898_n6094;
  wire REGFILE_SIM_reg_bank__abc_33898_n6095;
  wire REGFILE_SIM_reg_bank__abc_33898_n6096;
  wire REGFILE_SIM_reg_bank__abc_33898_n6097;
  wire REGFILE_SIM_reg_bank__abc_33898_n6098;
  wire REGFILE_SIM_reg_bank__abc_33898_n6099;
  wire REGFILE_SIM_reg_bank__abc_33898_n6100;
  wire REGFILE_SIM_reg_bank__abc_33898_n6101;
  wire REGFILE_SIM_reg_bank__abc_33898_n6102;
  wire REGFILE_SIM_reg_bank__abc_33898_n6103;
  wire REGFILE_SIM_reg_bank__abc_33898_n6104;
  wire REGFILE_SIM_reg_bank__abc_33898_n6105;
  wire REGFILE_SIM_reg_bank__abc_33898_n6106;
  wire REGFILE_SIM_reg_bank__abc_33898_n6107;
  wire REGFILE_SIM_reg_bank__abc_33898_n6108;
  wire REGFILE_SIM_reg_bank__abc_33898_n6109;
  wire REGFILE_SIM_reg_bank__abc_33898_n6110;
  wire REGFILE_SIM_reg_bank__abc_33898_n6111;
  wire REGFILE_SIM_reg_bank__abc_33898_n6112;
  wire REGFILE_SIM_reg_bank__abc_33898_n6113;
  wire REGFILE_SIM_reg_bank__abc_33898_n6114;
  wire REGFILE_SIM_reg_bank__abc_33898_n6115;
  wire REGFILE_SIM_reg_bank__abc_33898_n6116;
  wire REGFILE_SIM_reg_bank__abc_33898_n6117;
  wire REGFILE_SIM_reg_bank__abc_33898_n6118;
  wire REGFILE_SIM_reg_bank__abc_33898_n6119;
  wire REGFILE_SIM_reg_bank__abc_33898_n6120;
  wire REGFILE_SIM_reg_bank__abc_33898_n6121;
  wire REGFILE_SIM_reg_bank__abc_33898_n6122;
  wire REGFILE_SIM_reg_bank__abc_33898_n6123;
  wire REGFILE_SIM_reg_bank__abc_33898_n6124;
  wire REGFILE_SIM_reg_bank__abc_33898_n6125;
  wire REGFILE_SIM_reg_bank__abc_33898_n6126;
  wire REGFILE_SIM_reg_bank__abc_33898_n6127;
  wire REGFILE_SIM_reg_bank__abc_33898_n6128;
  wire REGFILE_SIM_reg_bank__abc_33898_n6129;
  wire REGFILE_SIM_reg_bank__abc_33898_n6130;
  wire REGFILE_SIM_reg_bank__abc_33898_n6131;
  wire REGFILE_SIM_reg_bank__abc_33898_n6132;
  wire REGFILE_SIM_reg_bank__abc_33898_n6133;
  wire REGFILE_SIM_reg_bank__abc_33898_n6134;
  wire REGFILE_SIM_reg_bank__abc_33898_n6135;
  wire REGFILE_SIM_reg_bank__abc_33898_n6136;
  wire REGFILE_SIM_reg_bank__abc_33898_n6137;
  wire REGFILE_SIM_reg_bank__abc_33898_n6138;
  wire REGFILE_SIM_reg_bank__abc_33898_n6139;
  wire REGFILE_SIM_reg_bank__abc_33898_n6140;
  wire REGFILE_SIM_reg_bank__abc_33898_n6141;
  wire REGFILE_SIM_reg_bank__abc_33898_n6142;
  wire REGFILE_SIM_reg_bank__abc_33898_n6143;
  wire REGFILE_SIM_reg_bank__abc_33898_n6145;
  wire REGFILE_SIM_reg_bank__abc_33898_n6146;
  wire REGFILE_SIM_reg_bank__abc_33898_n6147;
  wire REGFILE_SIM_reg_bank__abc_33898_n6148;
  wire REGFILE_SIM_reg_bank__abc_33898_n6149;
  wire REGFILE_SIM_reg_bank__abc_33898_n6150;
  wire REGFILE_SIM_reg_bank__abc_33898_n6151;
  wire REGFILE_SIM_reg_bank__abc_33898_n6152;
  wire REGFILE_SIM_reg_bank__abc_33898_n6153;
  wire REGFILE_SIM_reg_bank__abc_33898_n6154;
  wire REGFILE_SIM_reg_bank__abc_33898_n6155;
  wire REGFILE_SIM_reg_bank__abc_33898_n6156;
  wire REGFILE_SIM_reg_bank__abc_33898_n6157;
  wire REGFILE_SIM_reg_bank__abc_33898_n6158;
  wire REGFILE_SIM_reg_bank__abc_33898_n6159;
  wire REGFILE_SIM_reg_bank__abc_33898_n6160;
  wire REGFILE_SIM_reg_bank__abc_33898_n6161;
  wire REGFILE_SIM_reg_bank__abc_33898_n6162;
  wire REGFILE_SIM_reg_bank__abc_33898_n6163;
  wire REGFILE_SIM_reg_bank__abc_33898_n6164;
  wire REGFILE_SIM_reg_bank__abc_33898_n6165;
  wire REGFILE_SIM_reg_bank__abc_33898_n6166;
  wire REGFILE_SIM_reg_bank__abc_33898_n6167;
  wire REGFILE_SIM_reg_bank__abc_33898_n6168;
  wire REGFILE_SIM_reg_bank__abc_33898_n6169;
  wire REGFILE_SIM_reg_bank__abc_33898_n6170;
  wire REGFILE_SIM_reg_bank__abc_33898_n6171;
  wire REGFILE_SIM_reg_bank__abc_33898_n6172;
  wire REGFILE_SIM_reg_bank__abc_33898_n6173;
  wire REGFILE_SIM_reg_bank__abc_33898_n6174;
  wire REGFILE_SIM_reg_bank__abc_33898_n6175;
  wire REGFILE_SIM_reg_bank__abc_33898_n6176;
  wire REGFILE_SIM_reg_bank__abc_33898_n6177;
  wire REGFILE_SIM_reg_bank__abc_33898_n6178;
  wire REGFILE_SIM_reg_bank__abc_33898_n6179;
  wire REGFILE_SIM_reg_bank__abc_33898_n6180;
  wire REGFILE_SIM_reg_bank__abc_33898_n6181;
  wire REGFILE_SIM_reg_bank__abc_33898_n6182;
  wire REGFILE_SIM_reg_bank__abc_33898_n6183;
  wire REGFILE_SIM_reg_bank__abc_33898_n6184;
  wire REGFILE_SIM_reg_bank__abc_33898_n6185;
  wire REGFILE_SIM_reg_bank__abc_33898_n6186;
  wire REGFILE_SIM_reg_bank__abc_33898_n6187;
  wire REGFILE_SIM_reg_bank__abc_33898_n6188;
  wire REGFILE_SIM_reg_bank__abc_33898_n6189;
  wire REGFILE_SIM_reg_bank__abc_33898_n6190;
  wire REGFILE_SIM_reg_bank__abc_33898_n6191;
  wire REGFILE_SIM_reg_bank__abc_33898_n6192;
  wire REGFILE_SIM_reg_bank__abc_33898_n6193;
  wire REGFILE_SIM_reg_bank__abc_33898_n6194;
  wire REGFILE_SIM_reg_bank__abc_33898_n6195;
  wire REGFILE_SIM_reg_bank__abc_33898_n6196;
  wire REGFILE_SIM_reg_bank__abc_33898_n6197;
  wire REGFILE_SIM_reg_bank__abc_33898_n6198;
  wire REGFILE_SIM_reg_bank__abc_33898_n6199;
  wire REGFILE_SIM_reg_bank__abc_33898_n6200;
  wire REGFILE_SIM_reg_bank__abc_33898_n6201;
  wire REGFILE_SIM_reg_bank__abc_33898_n6202;
  wire REGFILE_SIM_reg_bank__abc_33898_n6203;
  wire REGFILE_SIM_reg_bank__abc_33898_n6204;
  wire REGFILE_SIM_reg_bank__abc_33898_n6206;
  wire REGFILE_SIM_reg_bank__abc_33898_n6207;
  wire REGFILE_SIM_reg_bank__abc_33898_n6208;
  wire REGFILE_SIM_reg_bank__abc_33898_n6209;
  wire REGFILE_SIM_reg_bank__abc_33898_n6210;
  wire REGFILE_SIM_reg_bank__abc_33898_n6211;
  wire REGFILE_SIM_reg_bank__abc_33898_n6212;
  wire REGFILE_SIM_reg_bank__abc_33898_n6213;
  wire REGFILE_SIM_reg_bank__abc_33898_n6214;
  wire REGFILE_SIM_reg_bank__abc_33898_n6215;
  wire REGFILE_SIM_reg_bank__abc_33898_n6216;
  wire REGFILE_SIM_reg_bank__abc_33898_n6217;
  wire REGFILE_SIM_reg_bank__abc_33898_n6218;
  wire REGFILE_SIM_reg_bank__abc_33898_n6219;
  wire REGFILE_SIM_reg_bank__abc_33898_n6220;
  wire REGFILE_SIM_reg_bank__abc_33898_n6221;
  wire REGFILE_SIM_reg_bank__abc_33898_n6222;
  wire REGFILE_SIM_reg_bank__abc_33898_n6223;
  wire REGFILE_SIM_reg_bank__abc_33898_n6224;
  wire REGFILE_SIM_reg_bank__abc_33898_n6225;
  wire REGFILE_SIM_reg_bank__abc_33898_n6226;
  wire REGFILE_SIM_reg_bank__abc_33898_n6227;
  wire REGFILE_SIM_reg_bank__abc_33898_n6228;
  wire REGFILE_SIM_reg_bank__abc_33898_n6229;
  wire REGFILE_SIM_reg_bank__abc_33898_n6230;
  wire REGFILE_SIM_reg_bank__abc_33898_n6231;
  wire REGFILE_SIM_reg_bank__abc_33898_n6232;
  wire REGFILE_SIM_reg_bank__abc_33898_n6233;
  wire REGFILE_SIM_reg_bank__abc_33898_n6234;
  wire REGFILE_SIM_reg_bank__abc_33898_n6235;
  wire REGFILE_SIM_reg_bank__abc_33898_n6236;
  wire REGFILE_SIM_reg_bank__abc_33898_n6237;
  wire REGFILE_SIM_reg_bank__abc_33898_n6238;
  wire REGFILE_SIM_reg_bank__abc_33898_n6239;
  wire REGFILE_SIM_reg_bank__abc_33898_n6240;
  wire REGFILE_SIM_reg_bank__abc_33898_n6241;
  wire REGFILE_SIM_reg_bank__abc_33898_n6242;
  wire REGFILE_SIM_reg_bank__abc_33898_n6243;
  wire REGFILE_SIM_reg_bank__abc_33898_n6244;
  wire REGFILE_SIM_reg_bank__abc_33898_n6245;
  wire REGFILE_SIM_reg_bank__abc_33898_n6246;
  wire REGFILE_SIM_reg_bank__abc_33898_n6247;
  wire REGFILE_SIM_reg_bank__abc_33898_n6248;
  wire REGFILE_SIM_reg_bank__abc_33898_n6249;
  wire REGFILE_SIM_reg_bank__abc_33898_n6250;
  wire REGFILE_SIM_reg_bank__abc_33898_n6251;
  wire REGFILE_SIM_reg_bank__abc_33898_n6252;
  wire REGFILE_SIM_reg_bank__abc_33898_n6253;
  wire REGFILE_SIM_reg_bank__abc_33898_n6254;
  wire REGFILE_SIM_reg_bank__abc_33898_n6255;
  wire REGFILE_SIM_reg_bank__abc_33898_n6256;
  wire REGFILE_SIM_reg_bank__abc_33898_n6257;
  wire REGFILE_SIM_reg_bank__abc_33898_n6258;
  wire REGFILE_SIM_reg_bank__abc_33898_n6259;
  wire REGFILE_SIM_reg_bank__abc_33898_n6260;
  wire REGFILE_SIM_reg_bank__abc_33898_n6261;
  wire REGFILE_SIM_reg_bank__abc_33898_n6262;
  wire REGFILE_SIM_reg_bank__abc_33898_n6263;
  wire REGFILE_SIM_reg_bank__abc_33898_n6264;
  wire REGFILE_SIM_reg_bank__abc_33898_n6265;
  wire REGFILE_SIM_reg_bank__abc_33898_n6267;
  wire REGFILE_SIM_reg_bank__abc_33898_n6268;
  wire REGFILE_SIM_reg_bank__abc_33898_n6269;
  wire REGFILE_SIM_reg_bank__abc_33898_n6270;
  wire REGFILE_SIM_reg_bank__abc_33898_n6271;
  wire REGFILE_SIM_reg_bank__abc_33898_n6272;
  wire REGFILE_SIM_reg_bank__abc_33898_n6273;
  wire REGFILE_SIM_reg_bank__abc_33898_n6274;
  wire REGFILE_SIM_reg_bank__abc_33898_n6275;
  wire REGFILE_SIM_reg_bank__abc_33898_n6276;
  wire REGFILE_SIM_reg_bank__abc_33898_n6277;
  wire REGFILE_SIM_reg_bank__abc_33898_n6278;
  wire REGFILE_SIM_reg_bank__abc_33898_n6279;
  wire REGFILE_SIM_reg_bank__abc_33898_n6280;
  wire REGFILE_SIM_reg_bank__abc_33898_n6281;
  wire REGFILE_SIM_reg_bank__abc_33898_n6282;
  wire REGFILE_SIM_reg_bank__abc_33898_n6283;
  wire REGFILE_SIM_reg_bank__abc_33898_n6284;
  wire REGFILE_SIM_reg_bank__abc_33898_n6285;
  wire REGFILE_SIM_reg_bank__abc_33898_n6286;
  wire REGFILE_SIM_reg_bank__abc_33898_n6287;
  wire REGFILE_SIM_reg_bank__abc_33898_n6288;
  wire REGFILE_SIM_reg_bank__abc_33898_n6289;
  wire REGFILE_SIM_reg_bank__abc_33898_n6290;
  wire REGFILE_SIM_reg_bank__abc_33898_n6291;
  wire REGFILE_SIM_reg_bank__abc_33898_n6292;
  wire REGFILE_SIM_reg_bank__abc_33898_n6293;
  wire REGFILE_SIM_reg_bank__abc_33898_n6294;
  wire REGFILE_SIM_reg_bank__abc_33898_n6295;
  wire REGFILE_SIM_reg_bank__abc_33898_n6296;
  wire REGFILE_SIM_reg_bank__abc_33898_n6297;
  wire REGFILE_SIM_reg_bank__abc_33898_n6298;
  wire REGFILE_SIM_reg_bank__abc_33898_n6299;
  wire REGFILE_SIM_reg_bank__abc_33898_n6300;
  wire REGFILE_SIM_reg_bank__abc_33898_n6301;
  wire REGFILE_SIM_reg_bank__abc_33898_n6302;
  wire REGFILE_SIM_reg_bank__abc_33898_n6303;
  wire REGFILE_SIM_reg_bank__abc_33898_n6304;
  wire REGFILE_SIM_reg_bank__abc_33898_n6305;
  wire REGFILE_SIM_reg_bank__abc_33898_n6306;
  wire REGFILE_SIM_reg_bank__abc_33898_n6307;
  wire REGFILE_SIM_reg_bank__abc_33898_n6308;
  wire REGFILE_SIM_reg_bank__abc_33898_n6309;
  wire REGFILE_SIM_reg_bank__abc_33898_n6310;
  wire REGFILE_SIM_reg_bank__abc_33898_n6311;
  wire REGFILE_SIM_reg_bank__abc_33898_n6312;
  wire REGFILE_SIM_reg_bank__abc_33898_n6313;
  wire REGFILE_SIM_reg_bank__abc_33898_n6314;
  wire REGFILE_SIM_reg_bank__abc_33898_n6315;
  wire REGFILE_SIM_reg_bank__abc_33898_n6316;
  wire REGFILE_SIM_reg_bank__abc_33898_n6317;
  wire REGFILE_SIM_reg_bank__abc_33898_n6318;
  wire REGFILE_SIM_reg_bank__abc_33898_n6319;
  wire REGFILE_SIM_reg_bank__abc_33898_n6320;
  wire REGFILE_SIM_reg_bank__abc_33898_n6321;
  wire REGFILE_SIM_reg_bank__abc_33898_n6322;
  wire REGFILE_SIM_reg_bank__abc_33898_n6323;
  wire REGFILE_SIM_reg_bank__abc_33898_n6324;
  wire REGFILE_SIM_reg_bank__abc_33898_n6325;
  wire REGFILE_SIM_reg_bank__abc_33898_n6326;
  wire REGFILE_SIM_reg_bank__abc_33898_n6328;
  wire REGFILE_SIM_reg_bank__abc_33898_n6329;
  wire REGFILE_SIM_reg_bank__abc_33898_n6330;
  wire REGFILE_SIM_reg_bank__abc_33898_n6331;
  wire REGFILE_SIM_reg_bank__abc_33898_n6332;
  wire REGFILE_SIM_reg_bank__abc_33898_n6333;
  wire REGFILE_SIM_reg_bank__abc_33898_n6334;
  wire REGFILE_SIM_reg_bank__abc_33898_n6335;
  wire REGFILE_SIM_reg_bank__abc_33898_n6336;
  wire REGFILE_SIM_reg_bank__abc_33898_n6337;
  wire REGFILE_SIM_reg_bank__abc_33898_n6338;
  wire REGFILE_SIM_reg_bank__abc_33898_n6339;
  wire REGFILE_SIM_reg_bank__abc_33898_n6340;
  wire REGFILE_SIM_reg_bank__abc_33898_n6341;
  wire REGFILE_SIM_reg_bank__abc_33898_n6342;
  wire REGFILE_SIM_reg_bank__abc_33898_n6343;
  wire REGFILE_SIM_reg_bank__abc_33898_n6344;
  wire REGFILE_SIM_reg_bank__abc_33898_n6345;
  wire REGFILE_SIM_reg_bank__abc_33898_n6346;
  wire REGFILE_SIM_reg_bank__abc_33898_n6347;
  wire REGFILE_SIM_reg_bank__abc_33898_n6348;
  wire REGFILE_SIM_reg_bank__abc_33898_n6349;
  wire REGFILE_SIM_reg_bank__abc_33898_n6350;
  wire REGFILE_SIM_reg_bank__abc_33898_n6351;
  wire REGFILE_SIM_reg_bank__abc_33898_n6352;
  wire REGFILE_SIM_reg_bank__abc_33898_n6353;
  wire REGFILE_SIM_reg_bank__abc_33898_n6354;
  wire REGFILE_SIM_reg_bank__abc_33898_n6355;
  wire REGFILE_SIM_reg_bank__abc_33898_n6356;
  wire REGFILE_SIM_reg_bank__abc_33898_n6357;
  wire REGFILE_SIM_reg_bank__abc_33898_n6358;
  wire REGFILE_SIM_reg_bank__abc_33898_n6359;
  wire REGFILE_SIM_reg_bank__abc_33898_n6360;
  wire REGFILE_SIM_reg_bank__abc_33898_n6361;
  wire REGFILE_SIM_reg_bank__abc_33898_n6362;
  wire REGFILE_SIM_reg_bank__abc_33898_n6363;
  wire REGFILE_SIM_reg_bank__abc_33898_n6364;
  wire REGFILE_SIM_reg_bank__abc_33898_n6365;
  wire REGFILE_SIM_reg_bank__abc_33898_n6366;
  wire REGFILE_SIM_reg_bank__abc_33898_n6367;
  wire REGFILE_SIM_reg_bank__abc_33898_n6368;
  wire REGFILE_SIM_reg_bank__abc_33898_n6369;
  wire REGFILE_SIM_reg_bank__abc_33898_n6370;
  wire REGFILE_SIM_reg_bank__abc_33898_n6371;
  wire REGFILE_SIM_reg_bank__abc_33898_n6372;
  wire REGFILE_SIM_reg_bank__abc_33898_n6373;
  wire REGFILE_SIM_reg_bank__abc_33898_n6374;
  wire REGFILE_SIM_reg_bank__abc_33898_n6375;
  wire REGFILE_SIM_reg_bank__abc_33898_n6376;
  wire REGFILE_SIM_reg_bank__abc_33898_n6377;
  wire REGFILE_SIM_reg_bank__abc_33898_n6378;
  wire REGFILE_SIM_reg_bank__abc_33898_n6379;
  wire REGFILE_SIM_reg_bank__abc_33898_n6380;
  wire REGFILE_SIM_reg_bank__abc_33898_n6381;
  wire REGFILE_SIM_reg_bank__abc_33898_n6382;
  wire REGFILE_SIM_reg_bank__abc_33898_n6383;
  wire REGFILE_SIM_reg_bank__abc_33898_n6384;
  wire REGFILE_SIM_reg_bank__abc_33898_n6385;
  wire REGFILE_SIM_reg_bank__abc_33898_n6386;
  wire REGFILE_SIM_reg_bank__abc_33898_n6387;
  wire REGFILE_SIM_reg_bank__abc_33898_n6389;
  wire REGFILE_SIM_reg_bank__abc_33898_n6390;
  wire REGFILE_SIM_reg_bank__abc_33898_n6391;
  wire REGFILE_SIM_reg_bank__abc_33898_n6392;
  wire REGFILE_SIM_reg_bank__abc_33898_n6393;
  wire REGFILE_SIM_reg_bank__abc_33898_n6394;
  wire REGFILE_SIM_reg_bank__abc_33898_n6395;
  wire REGFILE_SIM_reg_bank__abc_33898_n6396;
  wire REGFILE_SIM_reg_bank__abc_33898_n6397;
  wire REGFILE_SIM_reg_bank__abc_33898_n6398;
  wire REGFILE_SIM_reg_bank__abc_33898_n6399;
  wire REGFILE_SIM_reg_bank__abc_33898_n6400;
  wire REGFILE_SIM_reg_bank__abc_33898_n6401;
  wire REGFILE_SIM_reg_bank__abc_33898_n6402;
  wire REGFILE_SIM_reg_bank__abc_33898_n6403;
  wire REGFILE_SIM_reg_bank__abc_33898_n6404;
  wire REGFILE_SIM_reg_bank__abc_33898_n6405;
  wire REGFILE_SIM_reg_bank__abc_33898_n6406;
  wire REGFILE_SIM_reg_bank__abc_33898_n6407;
  wire REGFILE_SIM_reg_bank__abc_33898_n6408;
  wire REGFILE_SIM_reg_bank__abc_33898_n6409;
  wire REGFILE_SIM_reg_bank__abc_33898_n6410;
  wire REGFILE_SIM_reg_bank__abc_33898_n6411;
  wire REGFILE_SIM_reg_bank__abc_33898_n6412;
  wire REGFILE_SIM_reg_bank__abc_33898_n6413;
  wire REGFILE_SIM_reg_bank__abc_33898_n6414;
  wire REGFILE_SIM_reg_bank__abc_33898_n6415;
  wire REGFILE_SIM_reg_bank__abc_33898_n6416;
  wire REGFILE_SIM_reg_bank__abc_33898_n6417;
  wire REGFILE_SIM_reg_bank__abc_33898_n6418;
  wire REGFILE_SIM_reg_bank__abc_33898_n6419;
  wire REGFILE_SIM_reg_bank__abc_33898_n6420;
  wire REGFILE_SIM_reg_bank__abc_33898_n6421;
  wire REGFILE_SIM_reg_bank__abc_33898_n6422;
  wire REGFILE_SIM_reg_bank__abc_33898_n6423;
  wire REGFILE_SIM_reg_bank__abc_33898_n6424;
  wire REGFILE_SIM_reg_bank__abc_33898_n6425;
  wire REGFILE_SIM_reg_bank__abc_33898_n6426;
  wire REGFILE_SIM_reg_bank__abc_33898_n6427;
  wire REGFILE_SIM_reg_bank__abc_33898_n6428;
  wire REGFILE_SIM_reg_bank__abc_33898_n6429;
  wire REGFILE_SIM_reg_bank__abc_33898_n6430;
  wire REGFILE_SIM_reg_bank__abc_33898_n6431;
  wire REGFILE_SIM_reg_bank__abc_33898_n6432;
  wire REGFILE_SIM_reg_bank__abc_33898_n6433;
  wire REGFILE_SIM_reg_bank__abc_33898_n6434;
  wire REGFILE_SIM_reg_bank__abc_33898_n6435;
  wire REGFILE_SIM_reg_bank__abc_33898_n6436;
  wire REGFILE_SIM_reg_bank__abc_33898_n6437;
  wire REGFILE_SIM_reg_bank__abc_33898_n6438;
  wire REGFILE_SIM_reg_bank__abc_33898_n6439;
  wire REGFILE_SIM_reg_bank__abc_33898_n6440;
  wire REGFILE_SIM_reg_bank__abc_33898_n6441;
  wire REGFILE_SIM_reg_bank__abc_33898_n6442;
  wire REGFILE_SIM_reg_bank__abc_33898_n6443;
  wire REGFILE_SIM_reg_bank__abc_33898_n6444;
  wire REGFILE_SIM_reg_bank__abc_33898_n6445;
  wire REGFILE_SIM_reg_bank__abc_33898_n6446;
  wire REGFILE_SIM_reg_bank__abc_33898_n6447;
  wire REGFILE_SIM_reg_bank__abc_33898_n6448;
  wire REGFILE_SIM_reg_bank__abc_33898_n6450;
  wire REGFILE_SIM_reg_bank__abc_33898_n6451;
  wire REGFILE_SIM_reg_bank__abc_33898_n6452;
  wire REGFILE_SIM_reg_bank__abc_33898_n6453;
  wire REGFILE_SIM_reg_bank__abc_33898_n6454;
  wire REGFILE_SIM_reg_bank__abc_33898_n6455;
  wire REGFILE_SIM_reg_bank__abc_33898_n6456;
  wire REGFILE_SIM_reg_bank__abc_33898_n6457;
  wire REGFILE_SIM_reg_bank__abc_33898_n6458;
  wire REGFILE_SIM_reg_bank__abc_33898_n6459;
  wire REGFILE_SIM_reg_bank__abc_33898_n6460;
  wire REGFILE_SIM_reg_bank__abc_33898_n6461;
  wire REGFILE_SIM_reg_bank__abc_33898_n6462;
  wire REGFILE_SIM_reg_bank__abc_33898_n6463;
  wire REGFILE_SIM_reg_bank__abc_33898_n6464;
  wire REGFILE_SIM_reg_bank__abc_33898_n6465;
  wire REGFILE_SIM_reg_bank__abc_33898_n6466;
  wire REGFILE_SIM_reg_bank__abc_33898_n6467;
  wire REGFILE_SIM_reg_bank__abc_33898_n6468;
  wire REGFILE_SIM_reg_bank__abc_33898_n6469;
  wire REGFILE_SIM_reg_bank__abc_33898_n6470;
  wire REGFILE_SIM_reg_bank__abc_33898_n6471;
  wire REGFILE_SIM_reg_bank__abc_33898_n6472;
  wire REGFILE_SIM_reg_bank__abc_33898_n6473;
  wire REGFILE_SIM_reg_bank__abc_33898_n6474;
  wire REGFILE_SIM_reg_bank__abc_33898_n6475;
  wire REGFILE_SIM_reg_bank__abc_33898_n6476;
  wire REGFILE_SIM_reg_bank__abc_33898_n6477;
  wire REGFILE_SIM_reg_bank__abc_33898_n6478;
  wire REGFILE_SIM_reg_bank__abc_33898_n6479;
  wire REGFILE_SIM_reg_bank__abc_33898_n6480;
  wire REGFILE_SIM_reg_bank__abc_33898_n6481;
  wire REGFILE_SIM_reg_bank__abc_33898_n6482;
  wire REGFILE_SIM_reg_bank__abc_33898_n6483;
  wire REGFILE_SIM_reg_bank__abc_33898_n6484;
  wire REGFILE_SIM_reg_bank__abc_33898_n6485;
  wire REGFILE_SIM_reg_bank__abc_33898_n6486;
  wire REGFILE_SIM_reg_bank__abc_33898_n6487;
  wire REGFILE_SIM_reg_bank__abc_33898_n6488;
  wire REGFILE_SIM_reg_bank__abc_33898_n6489;
  wire REGFILE_SIM_reg_bank__abc_33898_n6490;
  wire REGFILE_SIM_reg_bank__abc_33898_n6491;
  wire REGFILE_SIM_reg_bank__abc_33898_n6492;
  wire REGFILE_SIM_reg_bank__abc_33898_n6493;
  wire REGFILE_SIM_reg_bank__abc_33898_n6494;
  wire REGFILE_SIM_reg_bank__abc_33898_n6495;
  wire REGFILE_SIM_reg_bank__abc_33898_n6496;
  wire REGFILE_SIM_reg_bank__abc_33898_n6497;
  wire REGFILE_SIM_reg_bank__abc_33898_n6498;
  wire REGFILE_SIM_reg_bank__abc_33898_n6499;
  wire REGFILE_SIM_reg_bank__abc_33898_n6500;
  wire REGFILE_SIM_reg_bank__abc_33898_n6501;
  wire REGFILE_SIM_reg_bank__abc_33898_n6502;
  wire REGFILE_SIM_reg_bank__abc_33898_n6503;
  wire REGFILE_SIM_reg_bank__abc_33898_n6504;
  wire REGFILE_SIM_reg_bank__abc_33898_n6505;
  wire REGFILE_SIM_reg_bank__abc_33898_n6506;
  wire REGFILE_SIM_reg_bank__abc_33898_n6507;
  wire REGFILE_SIM_reg_bank__abc_33898_n6508;
  wire REGFILE_SIM_reg_bank__abc_33898_n6509;
  wire REGFILE_SIM_reg_bank__abc_33898_n6511;
  wire REGFILE_SIM_reg_bank__abc_33898_n6512;
  wire REGFILE_SIM_reg_bank__abc_33898_n6513;
  wire REGFILE_SIM_reg_bank__abc_33898_n6514;
  wire REGFILE_SIM_reg_bank__abc_33898_n6515;
  wire REGFILE_SIM_reg_bank__abc_33898_n6516;
  wire REGFILE_SIM_reg_bank__abc_33898_n6517;
  wire REGFILE_SIM_reg_bank__abc_33898_n6518;
  wire REGFILE_SIM_reg_bank__abc_33898_n6519;
  wire REGFILE_SIM_reg_bank__abc_33898_n6520;
  wire REGFILE_SIM_reg_bank__abc_33898_n6521;
  wire REGFILE_SIM_reg_bank__abc_33898_n6522;
  wire REGFILE_SIM_reg_bank__abc_33898_n6523;
  wire REGFILE_SIM_reg_bank__abc_33898_n6524;
  wire REGFILE_SIM_reg_bank__abc_33898_n6525;
  wire REGFILE_SIM_reg_bank__abc_33898_n6526;
  wire REGFILE_SIM_reg_bank__abc_33898_n6527;
  wire REGFILE_SIM_reg_bank__abc_33898_n6528;
  wire REGFILE_SIM_reg_bank__abc_33898_n6529;
  wire REGFILE_SIM_reg_bank__abc_33898_n6530;
  wire REGFILE_SIM_reg_bank__abc_33898_n6531;
  wire REGFILE_SIM_reg_bank__abc_33898_n6532;
  wire REGFILE_SIM_reg_bank__abc_33898_n6533;
  wire REGFILE_SIM_reg_bank__abc_33898_n6534;
  wire REGFILE_SIM_reg_bank__abc_33898_n6535;
  wire REGFILE_SIM_reg_bank__abc_33898_n6536;
  wire REGFILE_SIM_reg_bank__abc_33898_n6537;
  wire REGFILE_SIM_reg_bank__abc_33898_n6538;
  wire REGFILE_SIM_reg_bank__abc_33898_n6539;
  wire REGFILE_SIM_reg_bank__abc_33898_n6540;
  wire REGFILE_SIM_reg_bank__abc_33898_n6541;
  wire REGFILE_SIM_reg_bank__abc_33898_n6542;
  wire REGFILE_SIM_reg_bank__abc_33898_n6543;
  wire REGFILE_SIM_reg_bank__abc_33898_n6544;
  wire REGFILE_SIM_reg_bank__abc_33898_n6545;
  wire REGFILE_SIM_reg_bank__abc_33898_n6546;
  wire REGFILE_SIM_reg_bank__abc_33898_n6547;
  wire REGFILE_SIM_reg_bank__abc_33898_n6548;
  wire REGFILE_SIM_reg_bank__abc_33898_n6549;
  wire REGFILE_SIM_reg_bank__abc_33898_n6550;
  wire REGFILE_SIM_reg_bank__abc_33898_n6551;
  wire REGFILE_SIM_reg_bank__abc_33898_n6552;
  wire REGFILE_SIM_reg_bank__abc_33898_n6553;
  wire REGFILE_SIM_reg_bank__abc_33898_n6554;
  wire REGFILE_SIM_reg_bank__abc_33898_n6555;
  wire REGFILE_SIM_reg_bank__abc_33898_n6556;
  wire REGFILE_SIM_reg_bank__abc_33898_n6557;
  wire REGFILE_SIM_reg_bank__abc_33898_n6558;
  wire REGFILE_SIM_reg_bank__abc_33898_n6559;
  wire REGFILE_SIM_reg_bank__abc_33898_n6560;
  wire REGFILE_SIM_reg_bank__abc_33898_n6561;
  wire REGFILE_SIM_reg_bank__abc_33898_n6562;
  wire REGFILE_SIM_reg_bank__abc_33898_n6563;
  wire REGFILE_SIM_reg_bank__abc_33898_n6564;
  wire REGFILE_SIM_reg_bank__abc_33898_n6565;
  wire REGFILE_SIM_reg_bank__abc_33898_n6566;
  wire REGFILE_SIM_reg_bank__abc_33898_n6567;
  wire REGFILE_SIM_reg_bank__abc_33898_n6568;
  wire REGFILE_SIM_reg_bank__abc_33898_n6569;
  wire REGFILE_SIM_reg_bank__abc_33898_n6570;
  wire REGFILE_SIM_reg_bank__abc_33898_n6572;
  wire REGFILE_SIM_reg_bank__abc_33898_n6573;
  wire REGFILE_SIM_reg_bank__abc_33898_n6574;
  wire REGFILE_SIM_reg_bank__abc_33898_n6575;
  wire REGFILE_SIM_reg_bank__abc_33898_n6576;
  wire REGFILE_SIM_reg_bank__abc_33898_n6577;
  wire REGFILE_SIM_reg_bank__abc_33898_n6578;
  wire REGFILE_SIM_reg_bank__abc_33898_n6579;
  wire REGFILE_SIM_reg_bank__abc_33898_n6580;
  wire REGFILE_SIM_reg_bank__abc_33898_n6581;
  wire REGFILE_SIM_reg_bank__abc_33898_n6582;
  wire REGFILE_SIM_reg_bank__abc_33898_n6583;
  wire REGFILE_SIM_reg_bank__abc_33898_n6584;
  wire REGFILE_SIM_reg_bank__abc_33898_n6585;
  wire REGFILE_SIM_reg_bank__abc_33898_n6586;
  wire REGFILE_SIM_reg_bank__abc_33898_n6587;
  wire REGFILE_SIM_reg_bank__abc_33898_n6588;
  wire REGFILE_SIM_reg_bank__abc_33898_n6589;
  wire REGFILE_SIM_reg_bank__abc_33898_n6590;
  wire REGFILE_SIM_reg_bank__abc_33898_n6591;
  wire REGFILE_SIM_reg_bank__abc_33898_n6592;
  wire REGFILE_SIM_reg_bank__abc_33898_n6593;
  wire REGFILE_SIM_reg_bank__abc_33898_n6594;
  wire REGFILE_SIM_reg_bank__abc_33898_n6595;
  wire REGFILE_SIM_reg_bank__abc_33898_n6596;
  wire REGFILE_SIM_reg_bank__abc_33898_n6597;
  wire REGFILE_SIM_reg_bank__abc_33898_n6598;
  wire REGFILE_SIM_reg_bank__abc_33898_n6599;
  wire REGFILE_SIM_reg_bank__abc_33898_n6600;
  wire REGFILE_SIM_reg_bank__abc_33898_n6601;
  wire REGFILE_SIM_reg_bank__abc_33898_n6602;
  wire REGFILE_SIM_reg_bank__abc_33898_n6603;
  wire REGFILE_SIM_reg_bank__abc_33898_n6604;
  wire REGFILE_SIM_reg_bank__abc_33898_n6605;
  wire REGFILE_SIM_reg_bank__abc_33898_n6606;
  wire REGFILE_SIM_reg_bank__abc_33898_n6607;
  wire REGFILE_SIM_reg_bank__abc_33898_n6608;
  wire REGFILE_SIM_reg_bank__abc_33898_n6609;
  wire REGFILE_SIM_reg_bank__abc_33898_n6610;
  wire REGFILE_SIM_reg_bank__abc_33898_n6611;
  wire REGFILE_SIM_reg_bank__abc_33898_n6612;
  wire REGFILE_SIM_reg_bank__abc_33898_n6613;
  wire REGFILE_SIM_reg_bank__abc_33898_n6614;
  wire REGFILE_SIM_reg_bank__abc_33898_n6615;
  wire REGFILE_SIM_reg_bank__abc_33898_n6616;
  wire REGFILE_SIM_reg_bank__abc_33898_n6617;
  wire REGFILE_SIM_reg_bank__abc_33898_n6618;
  wire REGFILE_SIM_reg_bank__abc_33898_n6619;
  wire REGFILE_SIM_reg_bank__abc_33898_n6620;
  wire REGFILE_SIM_reg_bank__abc_33898_n6621;
  wire REGFILE_SIM_reg_bank__abc_33898_n6622;
  wire REGFILE_SIM_reg_bank__abc_33898_n6623;
  wire REGFILE_SIM_reg_bank__abc_33898_n6624;
  wire REGFILE_SIM_reg_bank__abc_33898_n6625;
  wire REGFILE_SIM_reg_bank__abc_33898_n6626;
  wire REGFILE_SIM_reg_bank__abc_33898_n6627;
  wire REGFILE_SIM_reg_bank__abc_33898_n6628;
  wire REGFILE_SIM_reg_bank__abc_33898_n6629;
  wire REGFILE_SIM_reg_bank__abc_33898_n6630;
  wire REGFILE_SIM_reg_bank__abc_33898_n6631;
  wire REGFILE_SIM_reg_bank__abc_33898_n6633;
  wire REGFILE_SIM_reg_bank__abc_33898_n6634;
  wire REGFILE_SIM_reg_bank__abc_33898_n6635;
  wire REGFILE_SIM_reg_bank__abc_33898_n6636;
  wire REGFILE_SIM_reg_bank__abc_33898_n6637;
  wire REGFILE_SIM_reg_bank__abc_33898_n6638;
  wire REGFILE_SIM_reg_bank__abc_33898_n6639;
  wire REGFILE_SIM_reg_bank__abc_33898_n6640;
  wire REGFILE_SIM_reg_bank__abc_33898_n6641;
  wire REGFILE_SIM_reg_bank__abc_33898_n6642;
  wire REGFILE_SIM_reg_bank__abc_33898_n6643;
  wire REGFILE_SIM_reg_bank__abc_33898_n6644;
  wire REGFILE_SIM_reg_bank__abc_33898_n6645;
  wire REGFILE_SIM_reg_bank__abc_33898_n6646;
  wire REGFILE_SIM_reg_bank__abc_33898_n6647;
  wire REGFILE_SIM_reg_bank__abc_33898_n6648;
  wire REGFILE_SIM_reg_bank__abc_33898_n6649;
  wire REGFILE_SIM_reg_bank__abc_33898_n6650;
  wire REGFILE_SIM_reg_bank__abc_33898_n6651;
  wire REGFILE_SIM_reg_bank__abc_33898_n6652;
  wire REGFILE_SIM_reg_bank__abc_33898_n6653;
  wire REGFILE_SIM_reg_bank__abc_33898_n6654;
  wire REGFILE_SIM_reg_bank__abc_33898_n6655;
  wire REGFILE_SIM_reg_bank__abc_33898_n6656;
  wire REGFILE_SIM_reg_bank__abc_33898_n6657;
  wire REGFILE_SIM_reg_bank__abc_33898_n6658;
  wire REGFILE_SIM_reg_bank__abc_33898_n6659;
  wire REGFILE_SIM_reg_bank__abc_33898_n6660;
  wire REGFILE_SIM_reg_bank__abc_33898_n6661;
  wire REGFILE_SIM_reg_bank__abc_33898_n6662;
  wire REGFILE_SIM_reg_bank__abc_33898_n6663;
  wire REGFILE_SIM_reg_bank__abc_33898_n6664;
  wire REGFILE_SIM_reg_bank__abc_33898_n6665;
  wire REGFILE_SIM_reg_bank__abc_33898_n6666;
  wire REGFILE_SIM_reg_bank__abc_33898_n6667;
  wire REGFILE_SIM_reg_bank__abc_33898_n6668;
  wire REGFILE_SIM_reg_bank__abc_33898_n6669;
  wire REGFILE_SIM_reg_bank__abc_33898_n6670;
  wire REGFILE_SIM_reg_bank__abc_33898_n6671;
  wire REGFILE_SIM_reg_bank__abc_33898_n6672;
  wire REGFILE_SIM_reg_bank__abc_33898_n6673;
  wire REGFILE_SIM_reg_bank__abc_33898_n6674;
  wire REGFILE_SIM_reg_bank__abc_33898_n6675;
  wire REGFILE_SIM_reg_bank__abc_33898_n6676;
  wire REGFILE_SIM_reg_bank__abc_33898_n6677;
  wire REGFILE_SIM_reg_bank__abc_33898_n6678;
  wire REGFILE_SIM_reg_bank__abc_33898_n6679;
  wire REGFILE_SIM_reg_bank__abc_33898_n6680;
  wire REGFILE_SIM_reg_bank__abc_33898_n6681;
  wire REGFILE_SIM_reg_bank__abc_33898_n6682;
  wire REGFILE_SIM_reg_bank__abc_33898_n6683;
  wire REGFILE_SIM_reg_bank__abc_33898_n6684;
  wire REGFILE_SIM_reg_bank__abc_33898_n6685;
  wire REGFILE_SIM_reg_bank__abc_33898_n6686;
  wire REGFILE_SIM_reg_bank__abc_33898_n6687;
  wire REGFILE_SIM_reg_bank__abc_33898_n6688;
  wire REGFILE_SIM_reg_bank__abc_33898_n6689;
  wire REGFILE_SIM_reg_bank__abc_33898_n6690;
  wire REGFILE_SIM_reg_bank__abc_33898_n6691;
  wire REGFILE_SIM_reg_bank__abc_33898_n6692;
  wire REGFILE_SIM_reg_bank__abc_33898_n6694;
  wire REGFILE_SIM_reg_bank__abc_33898_n6695;
  wire REGFILE_SIM_reg_bank__abc_33898_n6696;
  wire REGFILE_SIM_reg_bank__abc_33898_n6697;
  wire REGFILE_SIM_reg_bank__abc_33898_n6698;
  wire REGFILE_SIM_reg_bank__abc_33898_n6699;
  wire REGFILE_SIM_reg_bank__abc_33898_n6700;
  wire REGFILE_SIM_reg_bank__abc_33898_n6701;
  wire REGFILE_SIM_reg_bank__abc_33898_n6702;
  wire REGFILE_SIM_reg_bank__abc_33898_n6703;
  wire REGFILE_SIM_reg_bank__abc_33898_n6704;
  wire REGFILE_SIM_reg_bank__abc_33898_n6705;
  wire REGFILE_SIM_reg_bank__abc_33898_n6706;
  wire REGFILE_SIM_reg_bank__abc_33898_n6707;
  wire REGFILE_SIM_reg_bank__abc_33898_n6708;
  wire REGFILE_SIM_reg_bank__abc_33898_n6709;
  wire REGFILE_SIM_reg_bank__abc_33898_n6710;
  wire REGFILE_SIM_reg_bank__abc_33898_n6711;
  wire REGFILE_SIM_reg_bank__abc_33898_n6712;
  wire REGFILE_SIM_reg_bank__abc_33898_n6713;
  wire REGFILE_SIM_reg_bank__abc_33898_n6714;
  wire REGFILE_SIM_reg_bank__abc_33898_n6715;
  wire REGFILE_SIM_reg_bank__abc_33898_n6716;
  wire REGFILE_SIM_reg_bank__abc_33898_n6717;
  wire REGFILE_SIM_reg_bank__abc_33898_n6718;
  wire REGFILE_SIM_reg_bank__abc_33898_n6719;
  wire REGFILE_SIM_reg_bank__abc_33898_n6720;
  wire REGFILE_SIM_reg_bank__abc_33898_n6721;
  wire REGFILE_SIM_reg_bank__abc_33898_n6722;
  wire REGFILE_SIM_reg_bank__abc_33898_n6723;
  wire REGFILE_SIM_reg_bank__abc_33898_n6724;
  wire REGFILE_SIM_reg_bank__abc_33898_n6725;
  wire REGFILE_SIM_reg_bank__abc_33898_n6726;
  wire REGFILE_SIM_reg_bank__abc_33898_n6727;
  wire REGFILE_SIM_reg_bank__abc_33898_n6728;
  wire REGFILE_SIM_reg_bank__abc_33898_n6729;
  wire REGFILE_SIM_reg_bank__abc_33898_n6730;
  wire REGFILE_SIM_reg_bank__abc_33898_n6731;
  wire REGFILE_SIM_reg_bank__abc_33898_n6732;
  wire REGFILE_SIM_reg_bank__abc_33898_n6733;
  wire REGFILE_SIM_reg_bank__abc_33898_n6734;
  wire REGFILE_SIM_reg_bank__abc_33898_n6735;
  wire REGFILE_SIM_reg_bank__abc_33898_n6736;
  wire REGFILE_SIM_reg_bank__abc_33898_n6737;
  wire REGFILE_SIM_reg_bank__abc_33898_n6738;
  wire REGFILE_SIM_reg_bank__abc_33898_n6739;
  wire REGFILE_SIM_reg_bank__abc_33898_n6740;
  wire REGFILE_SIM_reg_bank__abc_33898_n6741;
  wire REGFILE_SIM_reg_bank__abc_33898_n6742;
  wire REGFILE_SIM_reg_bank__abc_33898_n6743;
  wire REGFILE_SIM_reg_bank__abc_33898_n6744;
  wire REGFILE_SIM_reg_bank__abc_33898_n6745;
  wire REGFILE_SIM_reg_bank__abc_33898_n6746;
  wire REGFILE_SIM_reg_bank__abc_33898_n6747;
  wire REGFILE_SIM_reg_bank__abc_33898_n6748;
  wire REGFILE_SIM_reg_bank__abc_33898_n6749;
  wire REGFILE_SIM_reg_bank__abc_33898_n6750;
  wire REGFILE_SIM_reg_bank__abc_33898_n6751;
  wire REGFILE_SIM_reg_bank__abc_33898_n6752;
  wire REGFILE_SIM_reg_bank__abc_33898_n6753;
  wire REGFILE_SIM_reg_bank__abc_33898_n6755;
  wire REGFILE_SIM_reg_bank__abc_33898_n6756;
  wire REGFILE_SIM_reg_bank__abc_33898_n6757;
  wire REGFILE_SIM_reg_bank__abc_33898_n6758;
  wire REGFILE_SIM_reg_bank__abc_33898_n6759;
  wire REGFILE_SIM_reg_bank__abc_33898_n6760;
  wire REGFILE_SIM_reg_bank__abc_33898_n6761;
  wire REGFILE_SIM_reg_bank__abc_33898_n6762;
  wire REGFILE_SIM_reg_bank__abc_33898_n6763;
  wire REGFILE_SIM_reg_bank__abc_33898_n6764;
  wire REGFILE_SIM_reg_bank__abc_33898_n6765;
  wire REGFILE_SIM_reg_bank__abc_33898_n6766;
  wire REGFILE_SIM_reg_bank__abc_33898_n6767;
  wire REGFILE_SIM_reg_bank__abc_33898_n6768;
  wire REGFILE_SIM_reg_bank__abc_33898_n6769;
  wire REGFILE_SIM_reg_bank__abc_33898_n6770;
  wire REGFILE_SIM_reg_bank__abc_33898_n6771;
  wire REGFILE_SIM_reg_bank__abc_33898_n6772;
  wire REGFILE_SIM_reg_bank__abc_33898_n6773;
  wire REGFILE_SIM_reg_bank__abc_33898_n6774;
  wire REGFILE_SIM_reg_bank__abc_33898_n6775;
  wire REGFILE_SIM_reg_bank__abc_33898_n6776;
  wire REGFILE_SIM_reg_bank__abc_33898_n6777;
  wire REGFILE_SIM_reg_bank__abc_33898_n6778;
  wire REGFILE_SIM_reg_bank__abc_33898_n6779;
  wire REGFILE_SIM_reg_bank__abc_33898_n6780;
  wire REGFILE_SIM_reg_bank__abc_33898_n6781;
  wire REGFILE_SIM_reg_bank__abc_33898_n6782;
  wire REGFILE_SIM_reg_bank__abc_33898_n6783;
  wire REGFILE_SIM_reg_bank__abc_33898_n6784;
  wire REGFILE_SIM_reg_bank__abc_33898_n6785;
  wire REGFILE_SIM_reg_bank__abc_33898_n6786;
  wire REGFILE_SIM_reg_bank__abc_33898_n6787;
  wire REGFILE_SIM_reg_bank__abc_33898_n6788;
  wire REGFILE_SIM_reg_bank__abc_33898_n6789;
  wire REGFILE_SIM_reg_bank__abc_33898_n6790;
  wire REGFILE_SIM_reg_bank__abc_33898_n6791;
  wire REGFILE_SIM_reg_bank__abc_33898_n6792;
  wire REGFILE_SIM_reg_bank__abc_33898_n6793;
  wire REGFILE_SIM_reg_bank__abc_33898_n6794;
  wire REGFILE_SIM_reg_bank__abc_33898_n6795;
  wire REGFILE_SIM_reg_bank__abc_33898_n6796;
  wire REGFILE_SIM_reg_bank__abc_33898_n6797;
  wire REGFILE_SIM_reg_bank__abc_33898_n6798;
  wire REGFILE_SIM_reg_bank__abc_33898_n6799;
  wire REGFILE_SIM_reg_bank__abc_33898_n6800;
  wire REGFILE_SIM_reg_bank__abc_33898_n6801;
  wire REGFILE_SIM_reg_bank__abc_33898_n6802;
  wire REGFILE_SIM_reg_bank__abc_33898_n6803;
  wire REGFILE_SIM_reg_bank__abc_33898_n6804;
  wire REGFILE_SIM_reg_bank__abc_33898_n6805;
  wire REGFILE_SIM_reg_bank__abc_33898_n6806;
  wire REGFILE_SIM_reg_bank__abc_33898_n6807;
  wire REGFILE_SIM_reg_bank__abc_33898_n6808;
  wire REGFILE_SIM_reg_bank__abc_33898_n6809;
  wire REGFILE_SIM_reg_bank__abc_33898_n6810;
  wire REGFILE_SIM_reg_bank__abc_33898_n6811;
  wire REGFILE_SIM_reg_bank__abc_33898_n6812;
  wire REGFILE_SIM_reg_bank__abc_33898_n6813;
  wire REGFILE_SIM_reg_bank__abc_33898_n6814;
  wire REGFILE_SIM_reg_bank__abc_33898_n6816;
  wire REGFILE_SIM_reg_bank__abc_33898_n6817;
  wire REGFILE_SIM_reg_bank__abc_33898_n6818;
  wire REGFILE_SIM_reg_bank__abc_33898_n6819;
  wire REGFILE_SIM_reg_bank__abc_33898_n6820;
  wire REGFILE_SIM_reg_bank__abc_33898_n6821;
  wire REGFILE_SIM_reg_bank__abc_33898_n6822;
  wire REGFILE_SIM_reg_bank__abc_33898_n6823;
  wire REGFILE_SIM_reg_bank__abc_33898_n6824;
  wire REGFILE_SIM_reg_bank__abc_33898_n6825;
  wire REGFILE_SIM_reg_bank__abc_33898_n6826;
  wire REGFILE_SIM_reg_bank__abc_33898_n6827;
  wire REGFILE_SIM_reg_bank__abc_33898_n6828;
  wire REGFILE_SIM_reg_bank__abc_33898_n6829;
  wire REGFILE_SIM_reg_bank__abc_33898_n6830;
  wire REGFILE_SIM_reg_bank__abc_33898_n6831;
  wire REGFILE_SIM_reg_bank__abc_33898_n6832;
  wire REGFILE_SIM_reg_bank__abc_33898_n6833;
  wire REGFILE_SIM_reg_bank__abc_33898_n6834;
  wire REGFILE_SIM_reg_bank__abc_33898_n6835;
  wire REGFILE_SIM_reg_bank__abc_33898_n6836;
  wire REGFILE_SIM_reg_bank__abc_33898_n6837;
  wire REGFILE_SIM_reg_bank__abc_33898_n6838;
  wire REGFILE_SIM_reg_bank__abc_33898_n6839;
  wire REGFILE_SIM_reg_bank__abc_33898_n6840;
  wire REGFILE_SIM_reg_bank__abc_33898_n6841;
  wire REGFILE_SIM_reg_bank__abc_33898_n6842;
  wire REGFILE_SIM_reg_bank__abc_33898_n6843;
  wire REGFILE_SIM_reg_bank__abc_33898_n6844;
  wire REGFILE_SIM_reg_bank__abc_33898_n6845;
  wire REGFILE_SIM_reg_bank__abc_33898_n6846;
  wire REGFILE_SIM_reg_bank__abc_33898_n6847;
  wire REGFILE_SIM_reg_bank__abc_33898_n6848;
  wire REGFILE_SIM_reg_bank__abc_33898_n6849;
  wire REGFILE_SIM_reg_bank__abc_33898_n6850;
  wire REGFILE_SIM_reg_bank__abc_33898_n6851;
  wire REGFILE_SIM_reg_bank__abc_33898_n6852;
  wire REGFILE_SIM_reg_bank__abc_33898_n6853;
  wire REGFILE_SIM_reg_bank__abc_33898_n6854;
  wire REGFILE_SIM_reg_bank__abc_33898_n6855;
  wire REGFILE_SIM_reg_bank__abc_33898_n6856;
  wire REGFILE_SIM_reg_bank__abc_33898_n6857;
  wire REGFILE_SIM_reg_bank__abc_33898_n6858;
  wire REGFILE_SIM_reg_bank__abc_33898_n6859;
  wire REGFILE_SIM_reg_bank__abc_33898_n6860;
  wire REGFILE_SIM_reg_bank__abc_33898_n6861;
  wire REGFILE_SIM_reg_bank__abc_33898_n6862;
  wire REGFILE_SIM_reg_bank__abc_33898_n6863;
  wire REGFILE_SIM_reg_bank__abc_33898_n6864;
  wire REGFILE_SIM_reg_bank__abc_33898_n6865;
  wire REGFILE_SIM_reg_bank__abc_33898_n6866;
  wire REGFILE_SIM_reg_bank__abc_33898_n6867;
  wire REGFILE_SIM_reg_bank__abc_33898_n6868;
  wire REGFILE_SIM_reg_bank__abc_33898_n6869;
  wire REGFILE_SIM_reg_bank__abc_33898_n6870;
  wire REGFILE_SIM_reg_bank__abc_33898_n6871;
  wire REGFILE_SIM_reg_bank__abc_33898_n6872;
  wire REGFILE_SIM_reg_bank__abc_33898_n6873;
  wire REGFILE_SIM_reg_bank__abc_33898_n6874;
  wire REGFILE_SIM_reg_bank__abc_33898_n6875;
  wire REGFILE_SIM_reg_bank__abc_33898_n6877;
  wire REGFILE_SIM_reg_bank__abc_33898_n6878;
  wire REGFILE_SIM_reg_bank__abc_33898_n6879;
  wire REGFILE_SIM_reg_bank__abc_33898_n6880;
  wire REGFILE_SIM_reg_bank__abc_33898_n6881;
  wire REGFILE_SIM_reg_bank__abc_33898_n6882;
  wire REGFILE_SIM_reg_bank__abc_33898_n6883;
  wire REGFILE_SIM_reg_bank__abc_33898_n6884;
  wire REGFILE_SIM_reg_bank__abc_33898_n6885;
  wire REGFILE_SIM_reg_bank__abc_33898_n6886;
  wire REGFILE_SIM_reg_bank__abc_33898_n6887;
  wire REGFILE_SIM_reg_bank__abc_33898_n6888;
  wire REGFILE_SIM_reg_bank__abc_33898_n6889;
  wire REGFILE_SIM_reg_bank__abc_33898_n6890;
  wire REGFILE_SIM_reg_bank__abc_33898_n6891;
  wire REGFILE_SIM_reg_bank__abc_33898_n6892;
  wire REGFILE_SIM_reg_bank__abc_33898_n6893;
  wire REGFILE_SIM_reg_bank__abc_33898_n6894;
  wire REGFILE_SIM_reg_bank__abc_33898_n6895;
  wire REGFILE_SIM_reg_bank__abc_33898_n6896;
  wire REGFILE_SIM_reg_bank__abc_33898_n6897;
  wire REGFILE_SIM_reg_bank__abc_33898_n6898;
  wire REGFILE_SIM_reg_bank__abc_33898_n6899;
  wire REGFILE_SIM_reg_bank__abc_33898_n6900;
  wire REGFILE_SIM_reg_bank__abc_33898_n6901;
  wire REGFILE_SIM_reg_bank__abc_33898_n6902;
  wire REGFILE_SIM_reg_bank__abc_33898_n6903;
  wire REGFILE_SIM_reg_bank__abc_33898_n6904;
  wire REGFILE_SIM_reg_bank__abc_33898_n6905;
  wire REGFILE_SIM_reg_bank__abc_33898_n6906;
  wire REGFILE_SIM_reg_bank__abc_33898_n6907;
  wire REGFILE_SIM_reg_bank__abc_33898_n6908;
  wire REGFILE_SIM_reg_bank__abc_33898_n6909;
  wire REGFILE_SIM_reg_bank__abc_33898_n6910;
  wire REGFILE_SIM_reg_bank__abc_33898_n6911;
  wire REGFILE_SIM_reg_bank__abc_33898_n6912;
  wire REGFILE_SIM_reg_bank__abc_33898_n6913;
  wire REGFILE_SIM_reg_bank__abc_33898_n6914;
  wire REGFILE_SIM_reg_bank__abc_33898_n6915;
  wire REGFILE_SIM_reg_bank__abc_33898_n6916;
  wire REGFILE_SIM_reg_bank__abc_33898_n6917;
  wire REGFILE_SIM_reg_bank__abc_33898_n6918;
  wire REGFILE_SIM_reg_bank__abc_33898_n6919;
  wire REGFILE_SIM_reg_bank__abc_33898_n6920;
  wire REGFILE_SIM_reg_bank__abc_33898_n6921;
  wire REGFILE_SIM_reg_bank__abc_33898_n6922;
  wire REGFILE_SIM_reg_bank__abc_33898_n6923;
  wire REGFILE_SIM_reg_bank__abc_33898_n6924;
  wire REGFILE_SIM_reg_bank__abc_33898_n6925;
  wire REGFILE_SIM_reg_bank__abc_33898_n6926;
  wire REGFILE_SIM_reg_bank__abc_33898_n6927;
  wire REGFILE_SIM_reg_bank__abc_33898_n6928;
  wire REGFILE_SIM_reg_bank__abc_33898_n6929;
  wire REGFILE_SIM_reg_bank__abc_33898_n6930;
  wire REGFILE_SIM_reg_bank__abc_33898_n6931;
  wire REGFILE_SIM_reg_bank__abc_33898_n6932;
  wire REGFILE_SIM_reg_bank__abc_33898_n6933;
  wire REGFILE_SIM_reg_bank__abc_33898_n6934;
  wire REGFILE_SIM_reg_bank__abc_33898_n6935;
  wire REGFILE_SIM_reg_bank__abc_33898_n6936;
  wire REGFILE_SIM_reg_bank__abc_33898_n6938;
  wire REGFILE_SIM_reg_bank__abc_33898_n6939;
  wire REGFILE_SIM_reg_bank__abc_33898_n6940;
  wire REGFILE_SIM_reg_bank__abc_33898_n6941;
  wire REGFILE_SIM_reg_bank__abc_33898_n6942;
  wire REGFILE_SIM_reg_bank__abc_33898_n6943;
  wire REGFILE_SIM_reg_bank__abc_33898_n6944;
  wire REGFILE_SIM_reg_bank__abc_33898_n6945;
  wire REGFILE_SIM_reg_bank__abc_33898_n6946;
  wire REGFILE_SIM_reg_bank__abc_33898_n6947;
  wire REGFILE_SIM_reg_bank__abc_33898_n6948;
  wire REGFILE_SIM_reg_bank__abc_33898_n6949;
  wire REGFILE_SIM_reg_bank__abc_33898_n6950;
  wire REGFILE_SIM_reg_bank__abc_33898_n6951;
  wire REGFILE_SIM_reg_bank__abc_33898_n6952;
  wire REGFILE_SIM_reg_bank__abc_33898_n6953;
  wire REGFILE_SIM_reg_bank__abc_33898_n6954;
  wire REGFILE_SIM_reg_bank__abc_33898_n6955;
  wire REGFILE_SIM_reg_bank__abc_33898_n6956;
  wire REGFILE_SIM_reg_bank__abc_33898_n6957;
  wire REGFILE_SIM_reg_bank__abc_33898_n6958;
  wire REGFILE_SIM_reg_bank__abc_33898_n6959;
  wire REGFILE_SIM_reg_bank__abc_33898_n6960;
  wire REGFILE_SIM_reg_bank__abc_33898_n6961;
  wire REGFILE_SIM_reg_bank__abc_33898_n6962;
  wire REGFILE_SIM_reg_bank__abc_33898_n6963;
  wire REGFILE_SIM_reg_bank__abc_33898_n6964;
  wire REGFILE_SIM_reg_bank__abc_33898_n6965;
  wire REGFILE_SIM_reg_bank__abc_33898_n6966;
  wire REGFILE_SIM_reg_bank__abc_33898_n6967;
  wire REGFILE_SIM_reg_bank__abc_33898_n6968;
  wire REGFILE_SIM_reg_bank__abc_33898_n6969;
  wire REGFILE_SIM_reg_bank__abc_33898_n6970;
  wire REGFILE_SIM_reg_bank__abc_33898_n6971;
  wire REGFILE_SIM_reg_bank__abc_33898_n6972;
  wire REGFILE_SIM_reg_bank__abc_33898_n6973;
  wire REGFILE_SIM_reg_bank__abc_33898_n6974;
  wire REGFILE_SIM_reg_bank__abc_33898_n6975;
  wire REGFILE_SIM_reg_bank__abc_33898_n6976;
  wire REGFILE_SIM_reg_bank__abc_33898_n6977;
  wire REGFILE_SIM_reg_bank__abc_33898_n6978;
  wire REGFILE_SIM_reg_bank__abc_33898_n6979;
  wire REGFILE_SIM_reg_bank__abc_33898_n6980;
  wire REGFILE_SIM_reg_bank__abc_33898_n6981;
  wire REGFILE_SIM_reg_bank__abc_33898_n6982;
  wire REGFILE_SIM_reg_bank__abc_33898_n6983;
  wire REGFILE_SIM_reg_bank__abc_33898_n6984;
  wire REGFILE_SIM_reg_bank__abc_33898_n6985;
  wire REGFILE_SIM_reg_bank__abc_33898_n6986;
  wire REGFILE_SIM_reg_bank__abc_33898_n6987;
  wire REGFILE_SIM_reg_bank__abc_33898_n6988;
  wire REGFILE_SIM_reg_bank__abc_33898_n6989;
  wire REGFILE_SIM_reg_bank__abc_33898_n6990;
  wire REGFILE_SIM_reg_bank__abc_33898_n6991;
  wire REGFILE_SIM_reg_bank__abc_33898_n6992;
  wire REGFILE_SIM_reg_bank__abc_33898_n6993;
  wire REGFILE_SIM_reg_bank__abc_33898_n6994;
  wire REGFILE_SIM_reg_bank__abc_33898_n6995;
  wire REGFILE_SIM_reg_bank__abc_33898_n6996;
  wire REGFILE_SIM_reg_bank__abc_33898_n6997;
  wire REGFILE_SIM_reg_bank__abc_33898_n6999;
  wire REGFILE_SIM_reg_bank__abc_33898_n7000;
  wire REGFILE_SIM_reg_bank__abc_33898_n7001;
  wire REGFILE_SIM_reg_bank__abc_33898_n7002;
  wire REGFILE_SIM_reg_bank__abc_33898_n7003;
  wire REGFILE_SIM_reg_bank__abc_33898_n7004;
  wire REGFILE_SIM_reg_bank__abc_33898_n7005;
  wire REGFILE_SIM_reg_bank__abc_33898_n7006;
  wire REGFILE_SIM_reg_bank__abc_33898_n7007;
  wire REGFILE_SIM_reg_bank__abc_33898_n7008;
  wire REGFILE_SIM_reg_bank__abc_33898_n7009;
  wire REGFILE_SIM_reg_bank__abc_33898_n7010;
  wire REGFILE_SIM_reg_bank__abc_33898_n7011;
  wire REGFILE_SIM_reg_bank__abc_33898_n7012;
  wire REGFILE_SIM_reg_bank__abc_33898_n7013;
  wire REGFILE_SIM_reg_bank__abc_33898_n7014;
  wire REGFILE_SIM_reg_bank__abc_33898_n7015;
  wire REGFILE_SIM_reg_bank__abc_33898_n7016;
  wire REGFILE_SIM_reg_bank__abc_33898_n7017;
  wire REGFILE_SIM_reg_bank__abc_33898_n7018;
  wire REGFILE_SIM_reg_bank__abc_33898_n7019;
  wire REGFILE_SIM_reg_bank__abc_33898_n7020;
  wire REGFILE_SIM_reg_bank__abc_33898_n7021;
  wire REGFILE_SIM_reg_bank__abc_33898_n7022;
  wire REGFILE_SIM_reg_bank__abc_33898_n7023;
  wire REGFILE_SIM_reg_bank__abc_33898_n7024;
  wire REGFILE_SIM_reg_bank__abc_33898_n7025;
  wire REGFILE_SIM_reg_bank__abc_33898_n7026;
  wire REGFILE_SIM_reg_bank__abc_33898_n7027;
  wire REGFILE_SIM_reg_bank__abc_33898_n7028;
  wire REGFILE_SIM_reg_bank__abc_33898_n7029;
  wire REGFILE_SIM_reg_bank__abc_33898_n7030;
  wire REGFILE_SIM_reg_bank__abc_33898_n7031;
  wire REGFILE_SIM_reg_bank__abc_33898_n7032;
  wire REGFILE_SIM_reg_bank__abc_33898_n7033;
  wire REGFILE_SIM_reg_bank__abc_33898_n7034;
  wire REGFILE_SIM_reg_bank__abc_33898_n7035;
  wire REGFILE_SIM_reg_bank__abc_33898_n7036;
  wire REGFILE_SIM_reg_bank__abc_33898_n7037;
  wire REGFILE_SIM_reg_bank__abc_33898_n7038;
  wire REGFILE_SIM_reg_bank__abc_33898_n7039;
  wire REGFILE_SIM_reg_bank__abc_33898_n7040;
  wire REGFILE_SIM_reg_bank__abc_33898_n7041;
  wire REGFILE_SIM_reg_bank__abc_33898_n7042;
  wire REGFILE_SIM_reg_bank__abc_33898_n7043;
  wire REGFILE_SIM_reg_bank__abc_33898_n7044;
  wire REGFILE_SIM_reg_bank__abc_33898_n7045;
  wire REGFILE_SIM_reg_bank__abc_33898_n7046;
  wire REGFILE_SIM_reg_bank__abc_33898_n7047;
  wire REGFILE_SIM_reg_bank__abc_33898_n7048;
  wire REGFILE_SIM_reg_bank__abc_33898_n7049;
  wire REGFILE_SIM_reg_bank__abc_33898_n7050;
  wire REGFILE_SIM_reg_bank__abc_33898_n7051;
  wire REGFILE_SIM_reg_bank__abc_33898_n7052;
  wire REGFILE_SIM_reg_bank__abc_33898_n7053;
  wire REGFILE_SIM_reg_bank__abc_33898_n7054;
  wire REGFILE_SIM_reg_bank__abc_33898_n7055;
  wire REGFILE_SIM_reg_bank__abc_33898_n7056;
  wire REGFILE_SIM_reg_bank__abc_33898_n7057;
  wire REGFILE_SIM_reg_bank__abc_33898_n7058;
  wire REGFILE_SIM_reg_bank__abc_33898_n7060;
  wire REGFILE_SIM_reg_bank__abc_33898_n7061;
  wire REGFILE_SIM_reg_bank__abc_33898_n7062;
  wire REGFILE_SIM_reg_bank__abc_33898_n7063;
  wire REGFILE_SIM_reg_bank__abc_33898_n7064;
  wire REGFILE_SIM_reg_bank__abc_33898_n7065;
  wire REGFILE_SIM_reg_bank__abc_33898_n7066;
  wire REGFILE_SIM_reg_bank__abc_33898_n7067;
  wire REGFILE_SIM_reg_bank__abc_33898_n7068;
  wire REGFILE_SIM_reg_bank__abc_33898_n7069;
  wire REGFILE_SIM_reg_bank__abc_33898_n7070;
  wire REGFILE_SIM_reg_bank__abc_33898_n7071;
  wire REGFILE_SIM_reg_bank__abc_33898_n7072;
  wire REGFILE_SIM_reg_bank__abc_33898_n7073;
  wire REGFILE_SIM_reg_bank__abc_33898_n7074;
  wire REGFILE_SIM_reg_bank__abc_33898_n7075;
  wire REGFILE_SIM_reg_bank__abc_33898_n7076;
  wire REGFILE_SIM_reg_bank__abc_33898_n7077;
  wire REGFILE_SIM_reg_bank__abc_33898_n7078;
  wire REGFILE_SIM_reg_bank__abc_33898_n7079;
  wire REGFILE_SIM_reg_bank__abc_33898_n7080;
  wire REGFILE_SIM_reg_bank__abc_33898_n7081;
  wire REGFILE_SIM_reg_bank__abc_33898_n7082;
  wire REGFILE_SIM_reg_bank__abc_33898_n7083;
  wire REGFILE_SIM_reg_bank__abc_33898_n7084;
  wire REGFILE_SIM_reg_bank__abc_33898_n7085;
  wire REGFILE_SIM_reg_bank__abc_33898_n7086;
  wire REGFILE_SIM_reg_bank__abc_33898_n7087;
  wire REGFILE_SIM_reg_bank__abc_33898_n7088;
  wire REGFILE_SIM_reg_bank__abc_33898_n7089;
  wire REGFILE_SIM_reg_bank__abc_33898_n7090;
  wire REGFILE_SIM_reg_bank__abc_33898_n7091;
  wire REGFILE_SIM_reg_bank__abc_33898_n7092;
  wire REGFILE_SIM_reg_bank__abc_33898_n7093;
  wire REGFILE_SIM_reg_bank__abc_33898_n7094;
  wire REGFILE_SIM_reg_bank__abc_33898_n7095;
  wire REGFILE_SIM_reg_bank__abc_33898_n7096;
  wire REGFILE_SIM_reg_bank__abc_33898_n7097;
  wire REGFILE_SIM_reg_bank__abc_33898_n7098;
  wire REGFILE_SIM_reg_bank__abc_33898_n7099;
  wire REGFILE_SIM_reg_bank__abc_33898_n7100;
  wire REGFILE_SIM_reg_bank__abc_33898_n7101;
  wire REGFILE_SIM_reg_bank__abc_33898_n7102;
  wire REGFILE_SIM_reg_bank__abc_33898_n7103;
  wire REGFILE_SIM_reg_bank__abc_33898_n7104;
  wire REGFILE_SIM_reg_bank__abc_33898_n7105;
  wire REGFILE_SIM_reg_bank__abc_33898_n7106;
  wire REGFILE_SIM_reg_bank__abc_33898_n7107;
  wire REGFILE_SIM_reg_bank__abc_33898_n7108;
  wire REGFILE_SIM_reg_bank__abc_33898_n7109;
  wire REGFILE_SIM_reg_bank__abc_33898_n7110;
  wire REGFILE_SIM_reg_bank__abc_33898_n7111;
  wire REGFILE_SIM_reg_bank__abc_33898_n7112;
  wire REGFILE_SIM_reg_bank__abc_33898_n7113;
  wire REGFILE_SIM_reg_bank__abc_33898_n7114;
  wire REGFILE_SIM_reg_bank__abc_33898_n7115;
  wire REGFILE_SIM_reg_bank__abc_33898_n7116;
  wire REGFILE_SIM_reg_bank__abc_33898_n7117;
  wire REGFILE_SIM_reg_bank__abc_33898_n7118;
  wire REGFILE_SIM_reg_bank__abc_33898_n7119;
  wire REGFILE_SIM_reg_bank__abc_33898_n7121;
  wire REGFILE_SIM_reg_bank__abc_33898_n7122;
  wire REGFILE_SIM_reg_bank__abc_33898_n7123;
  wire REGFILE_SIM_reg_bank__abc_33898_n7124;
  wire REGFILE_SIM_reg_bank__abc_33898_n7125;
  wire REGFILE_SIM_reg_bank__abc_33898_n7126;
  wire REGFILE_SIM_reg_bank__abc_33898_n7127;
  wire REGFILE_SIM_reg_bank__abc_33898_n7128;
  wire REGFILE_SIM_reg_bank__abc_33898_n7129;
  wire REGFILE_SIM_reg_bank__abc_33898_n7130;
  wire REGFILE_SIM_reg_bank__abc_33898_n7131;
  wire REGFILE_SIM_reg_bank__abc_33898_n7132;
  wire REGFILE_SIM_reg_bank__abc_33898_n7133;
  wire REGFILE_SIM_reg_bank__abc_33898_n7134;
  wire REGFILE_SIM_reg_bank__abc_33898_n7135;
  wire REGFILE_SIM_reg_bank__abc_33898_n7136;
  wire REGFILE_SIM_reg_bank__abc_33898_n7137;
  wire REGFILE_SIM_reg_bank__abc_33898_n7138;
  wire REGFILE_SIM_reg_bank__abc_33898_n7139;
  wire REGFILE_SIM_reg_bank__abc_33898_n7140;
  wire REGFILE_SIM_reg_bank__abc_33898_n7141;
  wire REGFILE_SIM_reg_bank__abc_33898_n7142;
  wire REGFILE_SIM_reg_bank__abc_33898_n7143;
  wire REGFILE_SIM_reg_bank__abc_33898_n7144;
  wire REGFILE_SIM_reg_bank__abc_33898_n7145;
  wire REGFILE_SIM_reg_bank__abc_33898_n7146;
  wire REGFILE_SIM_reg_bank__abc_33898_n7147;
  wire REGFILE_SIM_reg_bank__abc_33898_n7148;
  wire REGFILE_SIM_reg_bank__abc_33898_n7149;
  wire REGFILE_SIM_reg_bank__abc_33898_n7150;
  wire REGFILE_SIM_reg_bank__abc_33898_n7151;
  wire REGFILE_SIM_reg_bank__abc_33898_n7152;
  wire REGFILE_SIM_reg_bank__abc_33898_n7153;
  wire REGFILE_SIM_reg_bank__abc_33898_n7154;
  wire REGFILE_SIM_reg_bank__abc_33898_n7155;
  wire REGFILE_SIM_reg_bank__abc_33898_n7156;
  wire REGFILE_SIM_reg_bank__abc_33898_n7157;
  wire REGFILE_SIM_reg_bank__abc_33898_n7158;
  wire REGFILE_SIM_reg_bank__abc_33898_n7159;
  wire REGFILE_SIM_reg_bank__abc_33898_n7160;
  wire REGFILE_SIM_reg_bank__abc_33898_n7161;
  wire REGFILE_SIM_reg_bank__abc_33898_n7162;
  wire REGFILE_SIM_reg_bank__abc_33898_n7163;
  wire REGFILE_SIM_reg_bank__abc_33898_n7164;
  wire REGFILE_SIM_reg_bank__abc_33898_n7165;
  wire REGFILE_SIM_reg_bank__abc_33898_n7166;
  wire REGFILE_SIM_reg_bank__abc_33898_n7167;
  wire REGFILE_SIM_reg_bank__abc_33898_n7168;
  wire REGFILE_SIM_reg_bank__abc_33898_n7169;
  wire REGFILE_SIM_reg_bank__abc_33898_n7170;
  wire REGFILE_SIM_reg_bank__abc_33898_n7171;
  wire REGFILE_SIM_reg_bank__abc_33898_n7172;
  wire REGFILE_SIM_reg_bank__abc_33898_n7173;
  wire REGFILE_SIM_reg_bank__abc_33898_n7174;
  wire REGFILE_SIM_reg_bank__abc_33898_n7175;
  wire REGFILE_SIM_reg_bank__abc_33898_n7176;
  wire REGFILE_SIM_reg_bank__abc_33898_n7177;
  wire REGFILE_SIM_reg_bank__abc_33898_n7178;
  wire REGFILE_SIM_reg_bank__abc_33898_n7179;
  wire REGFILE_SIM_reg_bank__abc_33898_n7180;
  wire REGFILE_SIM_reg_bank__abc_33898_n7182;
  wire REGFILE_SIM_reg_bank__abc_33898_n7183;
  wire REGFILE_SIM_reg_bank__abc_33898_n7184;
  wire REGFILE_SIM_reg_bank__abc_33898_n7185;
  wire REGFILE_SIM_reg_bank__abc_33898_n7186;
  wire REGFILE_SIM_reg_bank__abc_33898_n7187;
  wire REGFILE_SIM_reg_bank__abc_33898_n7188;
  wire REGFILE_SIM_reg_bank__abc_33898_n7189;
  wire REGFILE_SIM_reg_bank__abc_33898_n7190;
  wire REGFILE_SIM_reg_bank__abc_33898_n7191;
  wire REGFILE_SIM_reg_bank__abc_33898_n7192;
  wire REGFILE_SIM_reg_bank__abc_33898_n7193;
  wire REGFILE_SIM_reg_bank__abc_33898_n7194;
  wire REGFILE_SIM_reg_bank__abc_33898_n7195;
  wire REGFILE_SIM_reg_bank__abc_33898_n7196;
  wire REGFILE_SIM_reg_bank__abc_33898_n7197;
  wire REGFILE_SIM_reg_bank__abc_33898_n7198;
  wire REGFILE_SIM_reg_bank__abc_33898_n7199;
  wire REGFILE_SIM_reg_bank__abc_33898_n7200;
  wire REGFILE_SIM_reg_bank__abc_33898_n7201;
  wire REGFILE_SIM_reg_bank__abc_33898_n7202;
  wire REGFILE_SIM_reg_bank__abc_33898_n7203;
  wire REGFILE_SIM_reg_bank__abc_33898_n7204;
  wire REGFILE_SIM_reg_bank__abc_33898_n7205;
  wire REGFILE_SIM_reg_bank__abc_33898_n7206;
  wire REGFILE_SIM_reg_bank__abc_33898_n7207;
  wire REGFILE_SIM_reg_bank__abc_33898_n7208;
  wire REGFILE_SIM_reg_bank__abc_33898_n7209;
  wire REGFILE_SIM_reg_bank__abc_33898_n7210;
  wire REGFILE_SIM_reg_bank__abc_33898_n7211;
  wire REGFILE_SIM_reg_bank__abc_33898_n7212;
  wire REGFILE_SIM_reg_bank__abc_33898_n7213;
  wire REGFILE_SIM_reg_bank__abc_33898_n7214;
  wire REGFILE_SIM_reg_bank__abc_33898_n7215;
  wire REGFILE_SIM_reg_bank__abc_33898_n7216;
  wire REGFILE_SIM_reg_bank__abc_33898_n7217;
  wire REGFILE_SIM_reg_bank__abc_33898_n7218;
  wire REGFILE_SIM_reg_bank__abc_33898_n7219;
  wire REGFILE_SIM_reg_bank__abc_33898_n7220;
  wire REGFILE_SIM_reg_bank__abc_33898_n7221;
  wire REGFILE_SIM_reg_bank__abc_33898_n7222;
  wire REGFILE_SIM_reg_bank__abc_33898_n7223;
  wire REGFILE_SIM_reg_bank__abc_33898_n7224;
  wire REGFILE_SIM_reg_bank__abc_33898_n7225;
  wire REGFILE_SIM_reg_bank__abc_33898_n7226;
  wire REGFILE_SIM_reg_bank__abc_33898_n7227;
  wire REGFILE_SIM_reg_bank__abc_33898_n7228;
  wire REGFILE_SIM_reg_bank__abc_33898_n7229;
  wire REGFILE_SIM_reg_bank__abc_33898_n7230;
  wire REGFILE_SIM_reg_bank__abc_33898_n7231;
  wire REGFILE_SIM_reg_bank__abc_33898_n7232;
  wire REGFILE_SIM_reg_bank__abc_33898_n7233;
  wire REGFILE_SIM_reg_bank__abc_33898_n7234;
  wire REGFILE_SIM_reg_bank__abc_33898_n7235;
  wire REGFILE_SIM_reg_bank__abc_33898_n7236;
  wire REGFILE_SIM_reg_bank__abc_33898_n7237;
  wire REGFILE_SIM_reg_bank__abc_33898_n7238;
  wire REGFILE_SIM_reg_bank__abc_33898_n7239;
  wire REGFILE_SIM_reg_bank__abc_33898_n7240;
  wire REGFILE_SIM_reg_bank__abc_33898_n7241;
  wire REGFILE_SIM_reg_bank__abc_33898_n7243;
  wire REGFILE_SIM_reg_bank__abc_33898_n7244;
  wire REGFILE_SIM_reg_bank__abc_33898_n7245;
  wire REGFILE_SIM_reg_bank__abc_33898_n7246;
  wire REGFILE_SIM_reg_bank__abc_33898_n7247;
  wire REGFILE_SIM_reg_bank__abc_33898_n7248;
  wire REGFILE_SIM_reg_bank__abc_33898_n7249;
  wire REGFILE_SIM_reg_bank__abc_33898_n7250;
  wire REGFILE_SIM_reg_bank__abc_33898_n7251;
  wire REGFILE_SIM_reg_bank__abc_33898_n7252;
  wire REGFILE_SIM_reg_bank__abc_33898_n7253;
  wire REGFILE_SIM_reg_bank__abc_33898_n7254;
  wire REGFILE_SIM_reg_bank__abc_33898_n7255;
  wire REGFILE_SIM_reg_bank__abc_33898_n7256;
  wire REGFILE_SIM_reg_bank__abc_33898_n7257;
  wire REGFILE_SIM_reg_bank__abc_33898_n7258;
  wire REGFILE_SIM_reg_bank__abc_33898_n7259;
  wire REGFILE_SIM_reg_bank__abc_33898_n7260;
  wire REGFILE_SIM_reg_bank__abc_33898_n7261;
  wire REGFILE_SIM_reg_bank__abc_33898_n7262;
  wire REGFILE_SIM_reg_bank__abc_33898_n7263;
  wire REGFILE_SIM_reg_bank__abc_33898_n7264;
  wire REGFILE_SIM_reg_bank__abc_33898_n7265;
  wire REGFILE_SIM_reg_bank__abc_33898_n7266;
  wire REGFILE_SIM_reg_bank__abc_33898_n7267;
  wire REGFILE_SIM_reg_bank__abc_33898_n7268;
  wire REGFILE_SIM_reg_bank__abc_33898_n7269;
  wire REGFILE_SIM_reg_bank__abc_33898_n7270;
  wire REGFILE_SIM_reg_bank__abc_33898_n7271;
  wire REGFILE_SIM_reg_bank__abc_33898_n7272;
  wire REGFILE_SIM_reg_bank__abc_33898_n7273;
  wire REGFILE_SIM_reg_bank__abc_33898_n7274;
  wire REGFILE_SIM_reg_bank__abc_33898_n7275;
  wire REGFILE_SIM_reg_bank__abc_33898_n7276;
  wire REGFILE_SIM_reg_bank__abc_33898_n7277;
  wire REGFILE_SIM_reg_bank__abc_33898_n7278;
  wire REGFILE_SIM_reg_bank__abc_33898_n7279;
  wire REGFILE_SIM_reg_bank__abc_33898_n7280;
  wire REGFILE_SIM_reg_bank__abc_33898_n7281;
  wire REGFILE_SIM_reg_bank__abc_33898_n7282;
  wire REGFILE_SIM_reg_bank__abc_33898_n7283;
  wire REGFILE_SIM_reg_bank__abc_33898_n7284;
  wire REGFILE_SIM_reg_bank__abc_33898_n7285;
  wire REGFILE_SIM_reg_bank__abc_33898_n7286;
  wire REGFILE_SIM_reg_bank__abc_33898_n7287;
  wire REGFILE_SIM_reg_bank__abc_33898_n7288;
  wire REGFILE_SIM_reg_bank__abc_33898_n7289;
  wire REGFILE_SIM_reg_bank__abc_33898_n7290;
  wire REGFILE_SIM_reg_bank__abc_33898_n7291;
  wire REGFILE_SIM_reg_bank__abc_33898_n7292;
  wire REGFILE_SIM_reg_bank__abc_33898_n7293;
  wire REGFILE_SIM_reg_bank__abc_33898_n7294;
  wire REGFILE_SIM_reg_bank__abc_33898_n7295;
  wire REGFILE_SIM_reg_bank__abc_33898_n7296;
  wire REGFILE_SIM_reg_bank__abc_33898_n7297;
  wire REGFILE_SIM_reg_bank__abc_33898_n7298;
  wire REGFILE_SIM_reg_bank__abc_33898_n7299;
  wire REGFILE_SIM_reg_bank__abc_33898_n7300;
  wire REGFILE_SIM_reg_bank__abc_33898_n7301;
  wire REGFILE_SIM_reg_bank__abc_33898_n7302;
  wire REGFILE_SIM_reg_bank__abc_33898_n7304;
  wire REGFILE_SIM_reg_bank__abc_33898_n7305;
  wire REGFILE_SIM_reg_bank__abc_33898_n7306;
  wire REGFILE_SIM_reg_bank__abc_33898_n7307;
  wire REGFILE_SIM_reg_bank__abc_33898_n7308;
  wire REGFILE_SIM_reg_bank__abc_33898_n7309;
  wire REGFILE_SIM_reg_bank__abc_33898_n7310;
  wire REGFILE_SIM_reg_bank__abc_33898_n7311;
  wire REGFILE_SIM_reg_bank__abc_33898_n7312;
  wire REGFILE_SIM_reg_bank__abc_33898_n7313;
  wire REGFILE_SIM_reg_bank__abc_33898_n7314;
  wire REGFILE_SIM_reg_bank__abc_33898_n7315;
  wire REGFILE_SIM_reg_bank__abc_33898_n7316;
  wire REGFILE_SIM_reg_bank__abc_33898_n7317;
  wire REGFILE_SIM_reg_bank__abc_33898_n7318;
  wire REGFILE_SIM_reg_bank__abc_33898_n7319;
  wire REGFILE_SIM_reg_bank__abc_33898_n7320;
  wire REGFILE_SIM_reg_bank__abc_33898_n7321;
  wire REGFILE_SIM_reg_bank__abc_33898_n7322;
  wire REGFILE_SIM_reg_bank__abc_33898_n7323;
  wire REGFILE_SIM_reg_bank__abc_33898_n7324;
  wire REGFILE_SIM_reg_bank__abc_33898_n7325;
  wire REGFILE_SIM_reg_bank__abc_33898_n7326;
  wire REGFILE_SIM_reg_bank__abc_33898_n7327;
  wire REGFILE_SIM_reg_bank__abc_33898_n7328;
  wire REGFILE_SIM_reg_bank__abc_33898_n7329;
  wire REGFILE_SIM_reg_bank__abc_33898_n7330;
  wire REGFILE_SIM_reg_bank__abc_33898_n7331;
  wire REGFILE_SIM_reg_bank__abc_33898_n7332;
  wire REGFILE_SIM_reg_bank__abc_33898_n7333;
  wire REGFILE_SIM_reg_bank__abc_33898_n7334;
  wire REGFILE_SIM_reg_bank__abc_33898_n7335;
  wire REGFILE_SIM_reg_bank__abc_33898_n7336;
  wire REGFILE_SIM_reg_bank__abc_33898_n7337;
  wire REGFILE_SIM_reg_bank__abc_33898_n7338;
  wire REGFILE_SIM_reg_bank__abc_33898_n7339;
  wire REGFILE_SIM_reg_bank__abc_33898_n7340;
  wire REGFILE_SIM_reg_bank__abc_33898_n7341;
  wire REGFILE_SIM_reg_bank__abc_33898_n7342;
  wire REGFILE_SIM_reg_bank__abc_33898_n7343;
  wire REGFILE_SIM_reg_bank__abc_33898_n7344;
  wire REGFILE_SIM_reg_bank__abc_33898_n7345;
  wire REGFILE_SIM_reg_bank__abc_33898_n7346;
  wire REGFILE_SIM_reg_bank__abc_33898_n7347;
  wire REGFILE_SIM_reg_bank__abc_33898_n7348;
  wire REGFILE_SIM_reg_bank__abc_33898_n7349;
  wire REGFILE_SIM_reg_bank__abc_33898_n7350;
  wire REGFILE_SIM_reg_bank__abc_33898_n7351;
  wire REGFILE_SIM_reg_bank__abc_33898_n7352;
  wire REGFILE_SIM_reg_bank__abc_33898_n7353;
  wire REGFILE_SIM_reg_bank__abc_33898_n7354;
  wire REGFILE_SIM_reg_bank__abc_33898_n7355;
  wire REGFILE_SIM_reg_bank__abc_33898_n7356;
  wire REGFILE_SIM_reg_bank__abc_33898_n7357;
  wire REGFILE_SIM_reg_bank__abc_33898_n7358;
  wire REGFILE_SIM_reg_bank__abc_33898_n7359;
  wire REGFILE_SIM_reg_bank__abc_33898_n7360;
  wire REGFILE_SIM_reg_bank__abc_33898_n7361;
  wire REGFILE_SIM_reg_bank__abc_33898_n7362;
  wire REGFILE_SIM_reg_bank__abc_33898_n7363;
  wire REGFILE_SIM_reg_bank__abc_33898_n7365;
  wire REGFILE_SIM_reg_bank__abc_33898_n7366;
  wire REGFILE_SIM_reg_bank__abc_33898_n7367;
  wire REGFILE_SIM_reg_bank__abc_33898_n7368;
  wire REGFILE_SIM_reg_bank__abc_33898_n7369;
  wire REGFILE_SIM_reg_bank__abc_33898_n7370;
  wire REGFILE_SIM_reg_bank__abc_33898_n7371;
  wire REGFILE_SIM_reg_bank__abc_33898_n7372;
  wire REGFILE_SIM_reg_bank__abc_33898_n7373;
  wire REGFILE_SIM_reg_bank__abc_33898_n7374;
  wire REGFILE_SIM_reg_bank__abc_33898_n7375;
  wire REGFILE_SIM_reg_bank__abc_33898_n7376;
  wire REGFILE_SIM_reg_bank__abc_33898_n7377;
  wire REGFILE_SIM_reg_bank__abc_33898_n7378;
  wire REGFILE_SIM_reg_bank__abc_33898_n7379;
  wire REGFILE_SIM_reg_bank__abc_33898_n7380;
  wire REGFILE_SIM_reg_bank__abc_33898_n7381;
  wire REGFILE_SIM_reg_bank__abc_33898_n7382;
  wire REGFILE_SIM_reg_bank__abc_33898_n7383;
  wire REGFILE_SIM_reg_bank__abc_33898_n7384;
  wire REGFILE_SIM_reg_bank__abc_33898_n7385;
  wire REGFILE_SIM_reg_bank__abc_33898_n7386;
  wire REGFILE_SIM_reg_bank__abc_33898_n7387;
  wire REGFILE_SIM_reg_bank__abc_33898_n7388;
  wire REGFILE_SIM_reg_bank__abc_33898_n7389;
  wire REGFILE_SIM_reg_bank__abc_33898_n7390;
  wire REGFILE_SIM_reg_bank__abc_33898_n7391;
  wire REGFILE_SIM_reg_bank__abc_33898_n7392;
  wire REGFILE_SIM_reg_bank__abc_33898_n7393;
  wire REGFILE_SIM_reg_bank__abc_33898_n7394;
  wire REGFILE_SIM_reg_bank__abc_33898_n7395;
  wire REGFILE_SIM_reg_bank__abc_33898_n7396;
  wire REGFILE_SIM_reg_bank__abc_33898_n7397;
  wire REGFILE_SIM_reg_bank__abc_33898_n7398;
  wire REGFILE_SIM_reg_bank__abc_33898_n7399;
  wire REGFILE_SIM_reg_bank__abc_33898_n7400;
  wire REGFILE_SIM_reg_bank__abc_33898_n7401;
  wire REGFILE_SIM_reg_bank__abc_33898_n7402;
  wire REGFILE_SIM_reg_bank__abc_33898_n7403;
  wire REGFILE_SIM_reg_bank__abc_33898_n7404;
  wire REGFILE_SIM_reg_bank__abc_33898_n7405;
  wire REGFILE_SIM_reg_bank__abc_33898_n7406;
  wire REGFILE_SIM_reg_bank__abc_33898_n7407;
  wire REGFILE_SIM_reg_bank__abc_33898_n7408;
  wire REGFILE_SIM_reg_bank__abc_33898_n7409;
  wire REGFILE_SIM_reg_bank__abc_33898_n7410;
  wire REGFILE_SIM_reg_bank__abc_33898_n7411;
  wire REGFILE_SIM_reg_bank__abc_33898_n7412;
  wire REGFILE_SIM_reg_bank__abc_33898_n7413;
  wire REGFILE_SIM_reg_bank__abc_33898_n7414;
  wire REGFILE_SIM_reg_bank__abc_33898_n7415;
  wire REGFILE_SIM_reg_bank__abc_33898_n7416;
  wire REGFILE_SIM_reg_bank__abc_33898_n7417;
  wire REGFILE_SIM_reg_bank__abc_33898_n7418;
  wire REGFILE_SIM_reg_bank__abc_33898_n7419;
  wire REGFILE_SIM_reg_bank__abc_33898_n7420;
  wire REGFILE_SIM_reg_bank__abc_33898_n7421;
  wire REGFILE_SIM_reg_bank__abc_33898_n7422;
  wire REGFILE_SIM_reg_bank__abc_33898_n7423;
  wire REGFILE_SIM_reg_bank__abc_33898_n7424;
  wire REGFILE_SIM_reg_bank__abc_33898_n7426;
  wire REGFILE_SIM_reg_bank__abc_33898_n7427;
  wire REGFILE_SIM_reg_bank__abc_33898_n7428;
  wire REGFILE_SIM_reg_bank__abc_33898_n7429;
  wire REGFILE_SIM_reg_bank__abc_33898_n7430;
  wire REGFILE_SIM_reg_bank__abc_33898_n7431;
  wire REGFILE_SIM_reg_bank__abc_33898_n7432;
  wire REGFILE_SIM_reg_bank__abc_33898_n7433;
  wire REGFILE_SIM_reg_bank__abc_33898_n7434;
  wire REGFILE_SIM_reg_bank__abc_33898_n7435;
  wire REGFILE_SIM_reg_bank__abc_33898_n7436;
  wire REGFILE_SIM_reg_bank__abc_33898_n7437;
  wire REGFILE_SIM_reg_bank__abc_33898_n7438;
  wire REGFILE_SIM_reg_bank__abc_33898_n7439;
  wire REGFILE_SIM_reg_bank__abc_33898_n7440;
  wire REGFILE_SIM_reg_bank__abc_33898_n7441;
  wire REGFILE_SIM_reg_bank__abc_33898_n7442;
  wire REGFILE_SIM_reg_bank__abc_33898_n7443;
  wire REGFILE_SIM_reg_bank__abc_33898_n7444;
  wire REGFILE_SIM_reg_bank__abc_33898_n7445;
  wire REGFILE_SIM_reg_bank__abc_33898_n7446;
  wire REGFILE_SIM_reg_bank__abc_33898_n7447;
  wire REGFILE_SIM_reg_bank__abc_33898_n7448;
  wire REGFILE_SIM_reg_bank__abc_33898_n7449;
  wire REGFILE_SIM_reg_bank__abc_33898_n7450;
  wire REGFILE_SIM_reg_bank__abc_33898_n7451;
  wire REGFILE_SIM_reg_bank__abc_33898_n7452;
  wire REGFILE_SIM_reg_bank__abc_33898_n7453;
  wire REGFILE_SIM_reg_bank__abc_33898_n7454;
  wire REGFILE_SIM_reg_bank__abc_33898_n7455;
  wire REGFILE_SIM_reg_bank__abc_33898_n7456;
  wire REGFILE_SIM_reg_bank__abc_33898_n7457;
  wire REGFILE_SIM_reg_bank__abc_33898_n7458;
  wire REGFILE_SIM_reg_bank__abc_33898_n7459;
  wire REGFILE_SIM_reg_bank__abc_33898_n7460;
  wire REGFILE_SIM_reg_bank__abc_33898_n7461;
  wire REGFILE_SIM_reg_bank__abc_33898_n7462;
  wire REGFILE_SIM_reg_bank__abc_33898_n7463;
  wire REGFILE_SIM_reg_bank__abc_33898_n7464;
  wire REGFILE_SIM_reg_bank__abc_33898_n7465;
  wire REGFILE_SIM_reg_bank__abc_33898_n7466;
  wire REGFILE_SIM_reg_bank__abc_33898_n7467;
  wire REGFILE_SIM_reg_bank__abc_33898_n7468;
  wire REGFILE_SIM_reg_bank__abc_33898_n7469;
  wire REGFILE_SIM_reg_bank__abc_33898_n7470;
  wire REGFILE_SIM_reg_bank__abc_33898_n7471;
  wire REGFILE_SIM_reg_bank__abc_33898_n7472;
  wire REGFILE_SIM_reg_bank__abc_33898_n7473;
  wire REGFILE_SIM_reg_bank__abc_33898_n7474;
  wire REGFILE_SIM_reg_bank__abc_33898_n7475;
  wire REGFILE_SIM_reg_bank__abc_33898_n7476;
  wire REGFILE_SIM_reg_bank__abc_33898_n7477;
  wire REGFILE_SIM_reg_bank__abc_33898_n7478;
  wire REGFILE_SIM_reg_bank__abc_33898_n7479;
  wire REGFILE_SIM_reg_bank__abc_33898_n7480;
  wire REGFILE_SIM_reg_bank__abc_33898_n7481;
  wire REGFILE_SIM_reg_bank__abc_33898_n7482;
  wire REGFILE_SIM_reg_bank__abc_33898_n7483;
  wire REGFILE_SIM_reg_bank__abc_33898_n7484;
  wire REGFILE_SIM_reg_bank__abc_33898_n7485;
  wire REGFILE_SIM_reg_bank__abc_33898_n7487;
  wire REGFILE_SIM_reg_bank__abc_33898_n7488;
  wire REGFILE_SIM_reg_bank__abc_33898_n7489;
  wire REGFILE_SIM_reg_bank__abc_33898_n7490;
  wire REGFILE_SIM_reg_bank__abc_33898_n7491;
  wire REGFILE_SIM_reg_bank__abc_33898_n7492;
  wire REGFILE_SIM_reg_bank__abc_33898_n7493;
  wire REGFILE_SIM_reg_bank__abc_33898_n7494;
  wire REGFILE_SIM_reg_bank__abc_33898_n7495;
  wire REGFILE_SIM_reg_bank__abc_33898_n7496;
  wire REGFILE_SIM_reg_bank__abc_33898_n7497;
  wire REGFILE_SIM_reg_bank__abc_33898_n7498;
  wire REGFILE_SIM_reg_bank__abc_33898_n7499;
  wire REGFILE_SIM_reg_bank__abc_33898_n7500;
  wire REGFILE_SIM_reg_bank__abc_33898_n7501;
  wire REGFILE_SIM_reg_bank__abc_33898_n7502;
  wire REGFILE_SIM_reg_bank__abc_33898_n7503;
  wire REGFILE_SIM_reg_bank__abc_33898_n7504;
  wire REGFILE_SIM_reg_bank__abc_33898_n7505;
  wire REGFILE_SIM_reg_bank__abc_33898_n7506;
  wire REGFILE_SIM_reg_bank__abc_33898_n7507;
  wire REGFILE_SIM_reg_bank__abc_33898_n7508;
  wire REGFILE_SIM_reg_bank__abc_33898_n7509;
  wire REGFILE_SIM_reg_bank__abc_33898_n7510;
  wire REGFILE_SIM_reg_bank__abc_33898_n7511;
  wire REGFILE_SIM_reg_bank__abc_33898_n7512;
  wire REGFILE_SIM_reg_bank__abc_33898_n7513;
  wire REGFILE_SIM_reg_bank__abc_33898_n7514;
  wire REGFILE_SIM_reg_bank__abc_33898_n7515;
  wire REGFILE_SIM_reg_bank__abc_33898_n7516;
  wire REGFILE_SIM_reg_bank__abc_33898_n7517;
  wire REGFILE_SIM_reg_bank__abc_33898_n7518;
  wire REGFILE_SIM_reg_bank__abc_33898_n7519;
  wire REGFILE_SIM_reg_bank__abc_33898_n7520;
  wire REGFILE_SIM_reg_bank__abc_33898_n7521;
  wire REGFILE_SIM_reg_bank__abc_33898_n7522;
  wire REGFILE_SIM_reg_bank__abc_33898_n7523;
  wire REGFILE_SIM_reg_bank__abc_33898_n7524;
  wire REGFILE_SIM_reg_bank__abc_33898_n7525;
  wire REGFILE_SIM_reg_bank__abc_33898_n7526;
  wire REGFILE_SIM_reg_bank__abc_33898_n7527;
  wire REGFILE_SIM_reg_bank__abc_33898_n7528;
  wire REGFILE_SIM_reg_bank__abc_33898_n7529;
  wire REGFILE_SIM_reg_bank__abc_33898_n7530;
  wire REGFILE_SIM_reg_bank__abc_33898_n7531;
  wire REGFILE_SIM_reg_bank__abc_33898_n7532;
  wire REGFILE_SIM_reg_bank__abc_33898_n7533;
  wire REGFILE_SIM_reg_bank__abc_33898_n7534;
  wire REGFILE_SIM_reg_bank__abc_33898_n7535;
  wire REGFILE_SIM_reg_bank__abc_33898_n7536;
  wire REGFILE_SIM_reg_bank__abc_33898_n7537;
  wire REGFILE_SIM_reg_bank__abc_33898_n7538;
  wire REGFILE_SIM_reg_bank__abc_33898_n7539;
  wire REGFILE_SIM_reg_bank__abc_33898_n7540;
  wire REGFILE_SIM_reg_bank__abc_33898_n7541;
  wire REGFILE_SIM_reg_bank__abc_33898_n7542;
  wire REGFILE_SIM_reg_bank__abc_33898_n7543;
  wire REGFILE_SIM_reg_bank__abc_33898_n7544;
  wire REGFILE_SIM_reg_bank__abc_33898_n7545;
  wire REGFILE_SIM_reg_bank__abc_33898_n7546;
  wire REGFILE_SIM_reg_bank__abc_33898_n7548;
  wire REGFILE_SIM_reg_bank__abc_33898_n7549;
  wire REGFILE_SIM_reg_bank__abc_33898_n7550;
  wire REGFILE_SIM_reg_bank__abc_33898_n7551;
  wire REGFILE_SIM_reg_bank__abc_33898_n7552;
  wire REGFILE_SIM_reg_bank__abc_33898_n7553;
  wire REGFILE_SIM_reg_bank__abc_33898_n7554;
  wire REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7555;
  wire REGFILE_SIM_reg_bank__abc_33898_n7556;
  wire REGFILE_SIM_reg_bank__abc_33898_n7557;
  wire REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7558;
  wire REGFILE_SIM_reg_bank__abc_33898_n7559;
  wire REGFILE_SIM_reg_bank__abc_33898_n7560;
  wire REGFILE_SIM_reg_bank__abc_33898_n7561;
  wire REGFILE_SIM_reg_bank__abc_33898_n7562;
  wire REGFILE_SIM_reg_bank__abc_33898_n7563;
  wire REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7564;
  wire REGFILE_SIM_reg_bank__abc_33898_n7565;
  wire REGFILE_SIM_reg_bank__abc_33898_n7566;
  wire REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7567;
  wire REGFILE_SIM_reg_bank__abc_33898_n7568;
  wire REGFILE_SIM_reg_bank__abc_33898_n7569;
  wire REGFILE_SIM_reg_bank__abc_33898_n7570;
  wire REGFILE_SIM_reg_bank__abc_33898_n7571;
  wire REGFILE_SIM_reg_bank__abc_33898_n7572;
  wire REGFILE_SIM_reg_bank__abc_33898_n7573;
  wire REGFILE_SIM_reg_bank__abc_33898_n7574;
  wire REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7575;
  wire REGFILE_SIM_reg_bank__abc_33898_n7576;
  wire REGFILE_SIM_reg_bank__abc_33898_n7577;
  wire REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7578;
  wire REGFILE_SIM_reg_bank__abc_33898_n7579;
  wire REGFILE_SIM_reg_bank__abc_33898_n7580;
  wire REGFILE_SIM_reg_bank__abc_33898_n7581;
  wire REGFILE_SIM_reg_bank__abc_33898_n7582;
  wire REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7583;
  wire REGFILE_SIM_reg_bank__abc_33898_n7584;
  wire REGFILE_SIM_reg_bank__abc_33898_n7585;
  wire REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7586;
  wire REGFILE_SIM_reg_bank__abc_33898_n7587;
  wire REGFILE_SIM_reg_bank__abc_33898_n7588;
  wire REGFILE_SIM_reg_bank__abc_33898_n7589;
  wire REGFILE_SIM_reg_bank__abc_33898_n7590;
  wire REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7591;
  wire REGFILE_SIM_reg_bank__abc_33898_n7592;
  wire REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7593;
  wire REGFILE_SIM_reg_bank__abc_33898_n7594;
  wire REGFILE_SIM_reg_bank__abc_33898_n7595;
  wire REGFILE_SIM_reg_bank__abc_33898_n7596;
  wire REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7597;
  wire REGFILE_SIM_reg_bank__abc_33898_n7598;
  wire REGFILE_SIM_reg_bank__abc_33898_n7599;
  wire REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7600;
  wire REGFILE_SIM_reg_bank__abc_33898_n7601;
  wire REGFILE_SIM_reg_bank__abc_33898_n7602;
  wire REGFILE_SIM_reg_bank__abc_33898_n7603;
  wire REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7604;
  wire REGFILE_SIM_reg_bank__abc_33898_n7605;
  wire REGFILE_SIM_reg_bank__abc_33898_n7606;
  wire REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7607;
  wire REGFILE_SIM_reg_bank__abc_33898_n7608;
  wire REGFILE_SIM_reg_bank__abc_33898_n7609;
  wire REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7610;
  wire REGFILE_SIM_reg_bank__abc_33898_n7611;
  wire REGFILE_SIM_reg_bank__abc_33898_n7612;
  wire REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7613;
  wire REGFILE_SIM_reg_bank__abc_33898_n7614;
  wire REGFILE_SIM_reg_bank__abc_33898_n7615;
  wire REGFILE_SIM_reg_bank__abc_33898_n7616;
  wire REGFILE_SIM_reg_bank__abc_33898_n7617;
  wire REGFILE_SIM_reg_bank__abc_33898_n7618;
  wire REGFILE_SIM_reg_bank__abc_33898_n7619;
  wire REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7620;
  wire REGFILE_SIM_reg_bank__abc_33898_n7621;
  wire REGFILE_SIM_reg_bank__abc_33898_n7622;
  wire REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7623;
  wire REGFILE_SIM_reg_bank__abc_33898_n7624;
  wire REGFILE_SIM_reg_bank__abc_33898_n7625;
  wire REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7626;
  wire REGFILE_SIM_reg_bank__abc_33898_n7627;
  wire REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7628;
  wire REGFILE_SIM_reg_bank__abc_33898_n7629;
  wire REGFILE_SIM_reg_bank__abc_33898_n7630;
  wire REGFILE_SIM_reg_bank__abc_33898_n7631;
  wire REGFILE_SIM_reg_bank__abc_33898_n7632;
  wire REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7633;
  wire REGFILE_SIM_reg_bank__abc_33898_n7634;
  wire REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7635;
  wire REGFILE_SIM_reg_bank__abc_33898_n7636;
  wire REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7637;
  wire REGFILE_SIM_reg_bank__abc_33898_n7638;
  wire REGFILE_SIM_reg_bank__abc_33898_n7639;
  wire REGFILE_SIM_reg_bank__abc_33898_n7640;
  wire REGFILE_SIM_reg_bank__abc_33898_n7641;
  wire REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7642;
  wire REGFILE_SIM_reg_bank__abc_33898_n7643;
  wire REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7644;
  wire REGFILE_SIM_reg_bank__abc_33898_n7645;
  wire REGFILE_SIM_reg_bank__abc_33898_n7646;
  wire REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7647;
  wire REGFILE_SIM_reg_bank__abc_33898_n7648;
  wire REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7649;
  wire REGFILE_SIM_reg_bank__abc_33898_n7650;
  wire REGFILE_SIM_reg_bank__abc_33898_n7651;
  wire REGFILE_SIM_reg_bank__abc_33898_n7652;
  wire REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7653;
  wire REGFILE_SIM_reg_bank__abc_33898_n7654;
  wire REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7655;
  wire REGFILE_SIM_reg_bank__abc_33898_n7656;
  wire REGFILE_SIM_reg_bank__abc_33898_n7657;
  wire REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7658;
  wire REGFILE_SIM_reg_bank__abc_33898_n7659;
  wire REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf0;
  wire REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf1;
  wire REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf2;
  wire REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3;
  wire REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4;
  wire REGFILE_SIM_reg_bank__abc_33898_n7660;
  wire REGFILE_SIM_reg_bank__abc_33898_n7661;
  wire REGFILE_SIM_reg_bank__abc_33898_n7662;
  wire REGFILE_SIM_reg_bank__abc_33898_n7663;
  wire REGFILE_SIM_reg_bank__abc_33898_n7664;
  wire REGFILE_SIM_reg_bank__abc_33898_n7666;
  wire REGFILE_SIM_reg_bank__abc_33898_n7667;
  wire REGFILE_SIM_reg_bank__abc_33898_n7668;
  wire REGFILE_SIM_reg_bank__abc_33898_n7669;
  wire REGFILE_SIM_reg_bank__abc_33898_n7670;
  wire REGFILE_SIM_reg_bank__abc_33898_n7671;
  wire REGFILE_SIM_reg_bank__abc_33898_n7672;
  wire REGFILE_SIM_reg_bank__abc_33898_n7673;
  wire REGFILE_SIM_reg_bank__abc_33898_n7674;
  wire REGFILE_SIM_reg_bank__abc_33898_n7675;
  wire REGFILE_SIM_reg_bank__abc_33898_n7676;
  wire REGFILE_SIM_reg_bank__abc_33898_n7677;
  wire REGFILE_SIM_reg_bank__abc_33898_n7678;
  wire REGFILE_SIM_reg_bank__abc_33898_n7679;
  wire REGFILE_SIM_reg_bank__abc_33898_n7680;
  wire REGFILE_SIM_reg_bank__abc_33898_n7681;
  wire REGFILE_SIM_reg_bank__abc_33898_n7682;
  wire REGFILE_SIM_reg_bank__abc_33898_n7683;
  wire REGFILE_SIM_reg_bank__abc_33898_n7684;
  wire REGFILE_SIM_reg_bank__abc_33898_n7685;
  wire REGFILE_SIM_reg_bank__abc_33898_n7686;
  wire REGFILE_SIM_reg_bank__abc_33898_n7687;
  wire REGFILE_SIM_reg_bank__abc_33898_n7688;
  wire REGFILE_SIM_reg_bank__abc_33898_n7689;
  wire REGFILE_SIM_reg_bank__abc_33898_n7690;
  wire REGFILE_SIM_reg_bank__abc_33898_n7691;
  wire REGFILE_SIM_reg_bank__abc_33898_n7692;
  wire REGFILE_SIM_reg_bank__abc_33898_n7693;
  wire REGFILE_SIM_reg_bank__abc_33898_n7694;
  wire REGFILE_SIM_reg_bank__abc_33898_n7695;
  wire REGFILE_SIM_reg_bank__abc_33898_n7696;
  wire REGFILE_SIM_reg_bank__abc_33898_n7697;
  wire REGFILE_SIM_reg_bank__abc_33898_n7698;
  wire REGFILE_SIM_reg_bank__abc_33898_n7699;
  wire REGFILE_SIM_reg_bank__abc_33898_n7700;
  wire REGFILE_SIM_reg_bank__abc_33898_n7701;
  wire REGFILE_SIM_reg_bank__abc_33898_n7702;
  wire REGFILE_SIM_reg_bank__abc_33898_n7703;
  wire REGFILE_SIM_reg_bank__abc_33898_n7704;
  wire REGFILE_SIM_reg_bank__abc_33898_n7705;
  wire REGFILE_SIM_reg_bank__abc_33898_n7706;
  wire REGFILE_SIM_reg_bank__abc_33898_n7707;
  wire REGFILE_SIM_reg_bank__abc_33898_n7708;
  wire REGFILE_SIM_reg_bank__abc_33898_n7709;
  wire REGFILE_SIM_reg_bank__abc_33898_n7710;
  wire REGFILE_SIM_reg_bank__abc_33898_n7711;
  wire REGFILE_SIM_reg_bank__abc_33898_n7712;
  wire REGFILE_SIM_reg_bank__abc_33898_n7713;
  wire REGFILE_SIM_reg_bank__abc_33898_n7714;
  wire REGFILE_SIM_reg_bank__abc_33898_n7715;
  wire REGFILE_SIM_reg_bank__abc_33898_n7716;
  wire REGFILE_SIM_reg_bank__abc_33898_n7717;
  wire REGFILE_SIM_reg_bank__abc_33898_n7718;
  wire REGFILE_SIM_reg_bank__abc_33898_n7719;
  wire REGFILE_SIM_reg_bank__abc_33898_n7720;
  wire REGFILE_SIM_reg_bank__abc_33898_n7721;
  wire REGFILE_SIM_reg_bank__abc_33898_n7722;
  wire REGFILE_SIM_reg_bank__abc_33898_n7723;
  wire REGFILE_SIM_reg_bank__abc_33898_n7724;
  wire REGFILE_SIM_reg_bank__abc_33898_n7725;
  wire REGFILE_SIM_reg_bank__abc_33898_n7727;
  wire REGFILE_SIM_reg_bank__abc_33898_n7728;
  wire REGFILE_SIM_reg_bank__abc_33898_n7729;
  wire REGFILE_SIM_reg_bank__abc_33898_n7730;
  wire REGFILE_SIM_reg_bank__abc_33898_n7731;
  wire REGFILE_SIM_reg_bank__abc_33898_n7732;
  wire REGFILE_SIM_reg_bank__abc_33898_n7733;
  wire REGFILE_SIM_reg_bank__abc_33898_n7734;
  wire REGFILE_SIM_reg_bank__abc_33898_n7735;
  wire REGFILE_SIM_reg_bank__abc_33898_n7736;
  wire REGFILE_SIM_reg_bank__abc_33898_n7737;
  wire REGFILE_SIM_reg_bank__abc_33898_n7738;
  wire REGFILE_SIM_reg_bank__abc_33898_n7739;
  wire REGFILE_SIM_reg_bank__abc_33898_n7740;
  wire REGFILE_SIM_reg_bank__abc_33898_n7741;
  wire REGFILE_SIM_reg_bank__abc_33898_n7742;
  wire REGFILE_SIM_reg_bank__abc_33898_n7743;
  wire REGFILE_SIM_reg_bank__abc_33898_n7744;
  wire REGFILE_SIM_reg_bank__abc_33898_n7745;
  wire REGFILE_SIM_reg_bank__abc_33898_n7746;
  wire REGFILE_SIM_reg_bank__abc_33898_n7747;
  wire REGFILE_SIM_reg_bank__abc_33898_n7748;
  wire REGFILE_SIM_reg_bank__abc_33898_n7749;
  wire REGFILE_SIM_reg_bank__abc_33898_n7750;
  wire REGFILE_SIM_reg_bank__abc_33898_n7751;
  wire REGFILE_SIM_reg_bank__abc_33898_n7752;
  wire REGFILE_SIM_reg_bank__abc_33898_n7753;
  wire REGFILE_SIM_reg_bank__abc_33898_n7754;
  wire REGFILE_SIM_reg_bank__abc_33898_n7755;
  wire REGFILE_SIM_reg_bank__abc_33898_n7756;
  wire REGFILE_SIM_reg_bank__abc_33898_n7757;
  wire REGFILE_SIM_reg_bank__abc_33898_n7758;
  wire REGFILE_SIM_reg_bank__abc_33898_n7759;
  wire REGFILE_SIM_reg_bank__abc_33898_n7760;
  wire REGFILE_SIM_reg_bank__abc_33898_n7761;
  wire REGFILE_SIM_reg_bank__abc_33898_n7762;
  wire REGFILE_SIM_reg_bank__abc_33898_n7763;
  wire REGFILE_SIM_reg_bank__abc_33898_n7764;
  wire REGFILE_SIM_reg_bank__abc_33898_n7765;
  wire REGFILE_SIM_reg_bank__abc_33898_n7766;
  wire REGFILE_SIM_reg_bank__abc_33898_n7767;
  wire REGFILE_SIM_reg_bank__abc_33898_n7768;
  wire REGFILE_SIM_reg_bank__abc_33898_n7769;
  wire REGFILE_SIM_reg_bank__abc_33898_n7770;
  wire REGFILE_SIM_reg_bank__abc_33898_n7771;
  wire REGFILE_SIM_reg_bank__abc_33898_n7772;
  wire REGFILE_SIM_reg_bank__abc_33898_n7773;
  wire REGFILE_SIM_reg_bank__abc_33898_n7774;
  wire REGFILE_SIM_reg_bank__abc_33898_n7775;
  wire REGFILE_SIM_reg_bank__abc_33898_n7776;
  wire REGFILE_SIM_reg_bank__abc_33898_n7777;
  wire REGFILE_SIM_reg_bank__abc_33898_n7778;
  wire REGFILE_SIM_reg_bank__abc_33898_n7779;
  wire REGFILE_SIM_reg_bank__abc_33898_n7780;
  wire REGFILE_SIM_reg_bank__abc_33898_n7781;
  wire REGFILE_SIM_reg_bank__abc_33898_n7782;
  wire REGFILE_SIM_reg_bank__abc_33898_n7783;
  wire REGFILE_SIM_reg_bank__abc_33898_n7784;
  wire REGFILE_SIM_reg_bank__abc_33898_n7785;
  wire REGFILE_SIM_reg_bank__abc_33898_n7786;
  wire REGFILE_SIM_reg_bank__abc_33898_n7788;
  wire REGFILE_SIM_reg_bank__abc_33898_n7789;
  wire REGFILE_SIM_reg_bank__abc_33898_n7790;
  wire REGFILE_SIM_reg_bank__abc_33898_n7791;
  wire REGFILE_SIM_reg_bank__abc_33898_n7792;
  wire REGFILE_SIM_reg_bank__abc_33898_n7793;
  wire REGFILE_SIM_reg_bank__abc_33898_n7794;
  wire REGFILE_SIM_reg_bank__abc_33898_n7795;
  wire REGFILE_SIM_reg_bank__abc_33898_n7796;
  wire REGFILE_SIM_reg_bank__abc_33898_n7797;
  wire REGFILE_SIM_reg_bank__abc_33898_n7798;
  wire REGFILE_SIM_reg_bank__abc_33898_n7799;
  wire REGFILE_SIM_reg_bank__abc_33898_n7800;
  wire REGFILE_SIM_reg_bank__abc_33898_n7801;
  wire REGFILE_SIM_reg_bank__abc_33898_n7802;
  wire REGFILE_SIM_reg_bank__abc_33898_n7803;
  wire REGFILE_SIM_reg_bank__abc_33898_n7804;
  wire REGFILE_SIM_reg_bank__abc_33898_n7805;
  wire REGFILE_SIM_reg_bank__abc_33898_n7806;
  wire REGFILE_SIM_reg_bank__abc_33898_n7807;
  wire REGFILE_SIM_reg_bank__abc_33898_n7808;
  wire REGFILE_SIM_reg_bank__abc_33898_n7809;
  wire REGFILE_SIM_reg_bank__abc_33898_n7810;
  wire REGFILE_SIM_reg_bank__abc_33898_n7811;
  wire REGFILE_SIM_reg_bank__abc_33898_n7812;
  wire REGFILE_SIM_reg_bank__abc_33898_n7813;
  wire REGFILE_SIM_reg_bank__abc_33898_n7814;
  wire REGFILE_SIM_reg_bank__abc_33898_n7815;
  wire REGFILE_SIM_reg_bank__abc_33898_n7816;
  wire REGFILE_SIM_reg_bank__abc_33898_n7817;
  wire REGFILE_SIM_reg_bank__abc_33898_n7818;
  wire REGFILE_SIM_reg_bank__abc_33898_n7819;
  wire REGFILE_SIM_reg_bank__abc_33898_n7820;
  wire REGFILE_SIM_reg_bank__abc_33898_n7821;
  wire REGFILE_SIM_reg_bank__abc_33898_n7822;
  wire REGFILE_SIM_reg_bank__abc_33898_n7823;
  wire REGFILE_SIM_reg_bank__abc_33898_n7824;
  wire REGFILE_SIM_reg_bank__abc_33898_n7825;
  wire REGFILE_SIM_reg_bank__abc_33898_n7826;
  wire REGFILE_SIM_reg_bank__abc_33898_n7827;
  wire REGFILE_SIM_reg_bank__abc_33898_n7828;
  wire REGFILE_SIM_reg_bank__abc_33898_n7829;
  wire REGFILE_SIM_reg_bank__abc_33898_n7830;
  wire REGFILE_SIM_reg_bank__abc_33898_n7831;
  wire REGFILE_SIM_reg_bank__abc_33898_n7832;
  wire REGFILE_SIM_reg_bank__abc_33898_n7833;
  wire REGFILE_SIM_reg_bank__abc_33898_n7834;
  wire REGFILE_SIM_reg_bank__abc_33898_n7835;
  wire REGFILE_SIM_reg_bank__abc_33898_n7836;
  wire REGFILE_SIM_reg_bank__abc_33898_n7837;
  wire REGFILE_SIM_reg_bank__abc_33898_n7838;
  wire REGFILE_SIM_reg_bank__abc_33898_n7839;
  wire REGFILE_SIM_reg_bank__abc_33898_n7840;
  wire REGFILE_SIM_reg_bank__abc_33898_n7841;
  wire REGFILE_SIM_reg_bank__abc_33898_n7842;
  wire REGFILE_SIM_reg_bank__abc_33898_n7843;
  wire REGFILE_SIM_reg_bank__abc_33898_n7844;
  wire REGFILE_SIM_reg_bank__abc_33898_n7845;
  wire REGFILE_SIM_reg_bank__abc_33898_n7846;
  wire REGFILE_SIM_reg_bank__abc_33898_n7847;
  wire REGFILE_SIM_reg_bank__abc_33898_n7849;
  wire REGFILE_SIM_reg_bank__abc_33898_n7850;
  wire REGFILE_SIM_reg_bank__abc_33898_n7851;
  wire REGFILE_SIM_reg_bank__abc_33898_n7852;
  wire REGFILE_SIM_reg_bank__abc_33898_n7853;
  wire REGFILE_SIM_reg_bank__abc_33898_n7854;
  wire REGFILE_SIM_reg_bank__abc_33898_n7855;
  wire REGFILE_SIM_reg_bank__abc_33898_n7856;
  wire REGFILE_SIM_reg_bank__abc_33898_n7857;
  wire REGFILE_SIM_reg_bank__abc_33898_n7858;
  wire REGFILE_SIM_reg_bank__abc_33898_n7859;
  wire REGFILE_SIM_reg_bank__abc_33898_n7860;
  wire REGFILE_SIM_reg_bank__abc_33898_n7861;
  wire REGFILE_SIM_reg_bank__abc_33898_n7862;
  wire REGFILE_SIM_reg_bank__abc_33898_n7863;
  wire REGFILE_SIM_reg_bank__abc_33898_n7864;
  wire REGFILE_SIM_reg_bank__abc_33898_n7865;
  wire REGFILE_SIM_reg_bank__abc_33898_n7866;
  wire REGFILE_SIM_reg_bank__abc_33898_n7867;
  wire REGFILE_SIM_reg_bank__abc_33898_n7868;
  wire REGFILE_SIM_reg_bank__abc_33898_n7869;
  wire REGFILE_SIM_reg_bank__abc_33898_n7870;
  wire REGFILE_SIM_reg_bank__abc_33898_n7871;
  wire REGFILE_SIM_reg_bank__abc_33898_n7872;
  wire REGFILE_SIM_reg_bank__abc_33898_n7873;
  wire REGFILE_SIM_reg_bank__abc_33898_n7874;
  wire REGFILE_SIM_reg_bank__abc_33898_n7875;
  wire REGFILE_SIM_reg_bank__abc_33898_n7876;
  wire REGFILE_SIM_reg_bank__abc_33898_n7877;
  wire REGFILE_SIM_reg_bank__abc_33898_n7878;
  wire REGFILE_SIM_reg_bank__abc_33898_n7879;
  wire REGFILE_SIM_reg_bank__abc_33898_n7880;
  wire REGFILE_SIM_reg_bank__abc_33898_n7881;
  wire REGFILE_SIM_reg_bank__abc_33898_n7882;
  wire REGFILE_SIM_reg_bank__abc_33898_n7883;
  wire REGFILE_SIM_reg_bank__abc_33898_n7884;
  wire REGFILE_SIM_reg_bank__abc_33898_n7885;
  wire REGFILE_SIM_reg_bank__abc_33898_n7886;
  wire REGFILE_SIM_reg_bank__abc_33898_n7887;
  wire REGFILE_SIM_reg_bank__abc_33898_n7888;
  wire REGFILE_SIM_reg_bank__abc_33898_n7889;
  wire REGFILE_SIM_reg_bank__abc_33898_n7890;
  wire REGFILE_SIM_reg_bank__abc_33898_n7891;
  wire REGFILE_SIM_reg_bank__abc_33898_n7892;
  wire REGFILE_SIM_reg_bank__abc_33898_n7893;
  wire REGFILE_SIM_reg_bank__abc_33898_n7894;
  wire REGFILE_SIM_reg_bank__abc_33898_n7895;
  wire REGFILE_SIM_reg_bank__abc_33898_n7896;
  wire REGFILE_SIM_reg_bank__abc_33898_n7897;
  wire REGFILE_SIM_reg_bank__abc_33898_n7898;
  wire REGFILE_SIM_reg_bank__abc_33898_n7899;
  wire REGFILE_SIM_reg_bank__abc_33898_n7900;
  wire REGFILE_SIM_reg_bank__abc_33898_n7901;
  wire REGFILE_SIM_reg_bank__abc_33898_n7902;
  wire REGFILE_SIM_reg_bank__abc_33898_n7903;
  wire REGFILE_SIM_reg_bank__abc_33898_n7904;
  wire REGFILE_SIM_reg_bank__abc_33898_n7905;
  wire REGFILE_SIM_reg_bank__abc_33898_n7906;
  wire REGFILE_SIM_reg_bank__abc_33898_n7907;
  wire REGFILE_SIM_reg_bank__abc_33898_n7908;
  wire REGFILE_SIM_reg_bank__abc_33898_n7910;
  wire REGFILE_SIM_reg_bank__abc_33898_n7911;
  wire REGFILE_SIM_reg_bank__abc_33898_n7912;
  wire REGFILE_SIM_reg_bank__abc_33898_n7913;
  wire REGFILE_SIM_reg_bank__abc_33898_n7914;
  wire REGFILE_SIM_reg_bank__abc_33898_n7915;
  wire REGFILE_SIM_reg_bank__abc_33898_n7916;
  wire REGFILE_SIM_reg_bank__abc_33898_n7917;
  wire REGFILE_SIM_reg_bank__abc_33898_n7918;
  wire REGFILE_SIM_reg_bank__abc_33898_n7919;
  wire REGFILE_SIM_reg_bank__abc_33898_n7920;
  wire REGFILE_SIM_reg_bank__abc_33898_n7921;
  wire REGFILE_SIM_reg_bank__abc_33898_n7922;
  wire REGFILE_SIM_reg_bank__abc_33898_n7923;
  wire REGFILE_SIM_reg_bank__abc_33898_n7924;
  wire REGFILE_SIM_reg_bank__abc_33898_n7925;
  wire REGFILE_SIM_reg_bank__abc_33898_n7926;
  wire REGFILE_SIM_reg_bank__abc_33898_n7927;
  wire REGFILE_SIM_reg_bank__abc_33898_n7928;
  wire REGFILE_SIM_reg_bank__abc_33898_n7929;
  wire REGFILE_SIM_reg_bank__abc_33898_n7930;
  wire REGFILE_SIM_reg_bank__abc_33898_n7931;
  wire REGFILE_SIM_reg_bank__abc_33898_n7932;
  wire REGFILE_SIM_reg_bank__abc_33898_n7933;
  wire REGFILE_SIM_reg_bank__abc_33898_n7934;
  wire REGFILE_SIM_reg_bank__abc_33898_n7935;
  wire REGFILE_SIM_reg_bank__abc_33898_n7936;
  wire REGFILE_SIM_reg_bank__abc_33898_n7937;
  wire REGFILE_SIM_reg_bank__abc_33898_n7938;
  wire REGFILE_SIM_reg_bank__abc_33898_n7939;
  wire REGFILE_SIM_reg_bank__abc_33898_n7940;
  wire REGFILE_SIM_reg_bank__abc_33898_n7941;
  wire REGFILE_SIM_reg_bank__abc_33898_n7942;
  wire REGFILE_SIM_reg_bank__abc_33898_n7943;
  wire REGFILE_SIM_reg_bank__abc_33898_n7944;
  wire REGFILE_SIM_reg_bank__abc_33898_n7945;
  wire REGFILE_SIM_reg_bank__abc_33898_n7946;
  wire REGFILE_SIM_reg_bank__abc_33898_n7947;
  wire REGFILE_SIM_reg_bank__abc_33898_n7948;
  wire REGFILE_SIM_reg_bank__abc_33898_n7949;
  wire REGFILE_SIM_reg_bank__abc_33898_n7950;
  wire REGFILE_SIM_reg_bank__abc_33898_n7951;
  wire REGFILE_SIM_reg_bank__abc_33898_n7952;
  wire REGFILE_SIM_reg_bank__abc_33898_n7953;
  wire REGFILE_SIM_reg_bank__abc_33898_n7954;
  wire REGFILE_SIM_reg_bank__abc_33898_n7955;
  wire REGFILE_SIM_reg_bank__abc_33898_n7956;
  wire REGFILE_SIM_reg_bank__abc_33898_n7957;
  wire REGFILE_SIM_reg_bank__abc_33898_n7958;
  wire REGFILE_SIM_reg_bank__abc_33898_n7959;
  wire REGFILE_SIM_reg_bank__abc_33898_n7960;
  wire REGFILE_SIM_reg_bank__abc_33898_n7961;
  wire REGFILE_SIM_reg_bank__abc_33898_n7962;
  wire REGFILE_SIM_reg_bank__abc_33898_n7963;
  wire REGFILE_SIM_reg_bank__abc_33898_n7964;
  wire REGFILE_SIM_reg_bank__abc_33898_n7965;
  wire REGFILE_SIM_reg_bank__abc_33898_n7966;
  wire REGFILE_SIM_reg_bank__abc_33898_n7967;
  wire REGFILE_SIM_reg_bank__abc_33898_n7968;
  wire REGFILE_SIM_reg_bank__abc_33898_n7969;
  wire REGFILE_SIM_reg_bank__abc_33898_n7971;
  wire REGFILE_SIM_reg_bank__abc_33898_n7972;
  wire REGFILE_SIM_reg_bank__abc_33898_n7973;
  wire REGFILE_SIM_reg_bank__abc_33898_n7974;
  wire REGFILE_SIM_reg_bank__abc_33898_n7975;
  wire REGFILE_SIM_reg_bank__abc_33898_n7976;
  wire REGFILE_SIM_reg_bank__abc_33898_n7977;
  wire REGFILE_SIM_reg_bank__abc_33898_n7978;
  wire REGFILE_SIM_reg_bank__abc_33898_n7979;
  wire REGFILE_SIM_reg_bank__abc_33898_n7980;
  wire REGFILE_SIM_reg_bank__abc_33898_n7981;
  wire REGFILE_SIM_reg_bank__abc_33898_n7982;
  wire REGFILE_SIM_reg_bank__abc_33898_n7983;
  wire REGFILE_SIM_reg_bank__abc_33898_n7984;
  wire REGFILE_SIM_reg_bank__abc_33898_n7985;
  wire REGFILE_SIM_reg_bank__abc_33898_n7986;
  wire REGFILE_SIM_reg_bank__abc_33898_n7987;
  wire REGFILE_SIM_reg_bank__abc_33898_n7988;
  wire REGFILE_SIM_reg_bank__abc_33898_n7989;
  wire REGFILE_SIM_reg_bank__abc_33898_n7990;
  wire REGFILE_SIM_reg_bank__abc_33898_n7991;
  wire REGFILE_SIM_reg_bank__abc_33898_n7992;
  wire REGFILE_SIM_reg_bank__abc_33898_n7993;
  wire REGFILE_SIM_reg_bank__abc_33898_n7994;
  wire REGFILE_SIM_reg_bank__abc_33898_n7995;
  wire REGFILE_SIM_reg_bank__abc_33898_n7996;
  wire REGFILE_SIM_reg_bank__abc_33898_n7997;
  wire REGFILE_SIM_reg_bank__abc_33898_n7998;
  wire REGFILE_SIM_reg_bank__abc_33898_n7999;
  wire REGFILE_SIM_reg_bank__abc_33898_n8000;
  wire REGFILE_SIM_reg_bank__abc_33898_n8001;
  wire REGFILE_SIM_reg_bank__abc_33898_n8002;
  wire REGFILE_SIM_reg_bank__abc_33898_n8003;
  wire REGFILE_SIM_reg_bank__abc_33898_n8004;
  wire REGFILE_SIM_reg_bank__abc_33898_n8005;
  wire REGFILE_SIM_reg_bank__abc_33898_n8006;
  wire REGFILE_SIM_reg_bank__abc_33898_n8007;
  wire REGFILE_SIM_reg_bank__abc_33898_n8008;
  wire REGFILE_SIM_reg_bank__abc_33898_n8009;
  wire REGFILE_SIM_reg_bank__abc_33898_n8010;
  wire REGFILE_SIM_reg_bank__abc_33898_n8011;
  wire REGFILE_SIM_reg_bank__abc_33898_n8012;
  wire REGFILE_SIM_reg_bank__abc_33898_n8013;
  wire REGFILE_SIM_reg_bank__abc_33898_n8014;
  wire REGFILE_SIM_reg_bank__abc_33898_n8015;
  wire REGFILE_SIM_reg_bank__abc_33898_n8016;
  wire REGFILE_SIM_reg_bank__abc_33898_n8017;
  wire REGFILE_SIM_reg_bank__abc_33898_n8018;
  wire REGFILE_SIM_reg_bank__abc_33898_n8019;
  wire REGFILE_SIM_reg_bank__abc_33898_n8020;
  wire REGFILE_SIM_reg_bank__abc_33898_n8021;
  wire REGFILE_SIM_reg_bank__abc_33898_n8022;
  wire REGFILE_SIM_reg_bank__abc_33898_n8023;
  wire REGFILE_SIM_reg_bank__abc_33898_n8024;
  wire REGFILE_SIM_reg_bank__abc_33898_n8025;
  wire REGFILE_SIM_reg_bank__abc_33898_n8026;
  wire REGFILE_SIM_reg_bank__abc_33898_n8027;
  wire REGFILE_SIM_reg_bank__abc_33898_n8028;
  wire REGFILE_SIM_reg_bank__abc_33898_n8029;
  wire REGFILE_SIM_reg_bank__abc_33898_n8030;
  wire REGFILE_SIM_reg_bank__abc_33898_n8032;
  wire REGFILE_SIM_reg_bank__abc_33898_n8033;
  wire REGFILE_SIM_reg_bank__abc_33898_n8034;
  wire REGFILE_SIM_reg_bank__abc_33898_n8035;
  wire REGFILE_SIM_reg_bank__abc_33898_n8036;
  wire REGFILE_SIM_reg_bank__abc_33898_n8037;
  wire REGFILE_SIM_reg_bank__abc_33898_n8038;
  wire REGFILE_SIM_reg_bank__abc_33898_n8039;
  wire REGFILE_SIM_reg_bank__abc_33898_n8040;
  wire REGFILE_SIM_reg_bank__abc_33898_n8041;
  wire REGFILE_SIM_reg_bank__abc_33898_n8042;
  wire REGFILE_SIM_reg_bank__abc_33898_n8043;
  wire REGFILE_SIM_reg_bank__abc_33898_n8044;
  wire REGFILE_SIM_reg_bank__abc_33898_n8045;
  wire REGFILE_SIM_reg_bank__abc_33898_n8046;
  wire REGFILE_SIM_reg_bank__abc_33898_n8047;
  wire REGFILE_SIM_reg_bank__abc_33898_n8048;
  wire REGFILE_SIM_reg_bank__abc_33898_n8049;
  wire REGFILE_SIM_reg_bank__abc_33898_n8050;
  wire REGFILE_SIM_reg_bank__abc_33898_n8051;
  wire REGFILE_SIM_reg_bank__abc_33898_n8052;
  wire REGFILE_SIM_reg_bank__abc_33898_n8053;
  wire REGFILE_SIM_reg_bank__abc_33898_n8054;
  wire REGFILE_SIM_reg_bank__abc_33898_n8055;
  wire REGFILE_SIM_reg_bank__abc_33898_n8056;
  wire REGFILE_SIM_reg_bank__abc_33898_n8057;
  wire REGFILE_SIM_reg_bank__abc_33898_n8058;
  wire REGFILE_SIM_reg_bank__abc_33898_n8059;
  wire REGFILE_SIM_reg_bank__abc_33898_n8060;
  wire REGFILE_SIM_reg_bank__abc_33898_n8061;
  wire REGFILE_SIM_reg_bank__abc_33898_n8062;
  wire REGFILE_SIM_reg_bank__abc_33898_n8063;
  wire REGFILE_SIM_reg_bank__abc_33898_n8064;
  wire REGFILE_SIM_reg_bank__abc_33898_n8065;
  wire REGFILE_SIM_reg_bank__abc_33898_n8066;
  wire REGFILE_SIM_reg_bank__abc_33898_n8067;
  wire REGFILE_SIM_reg_bank__abc_33898_n8068;
  wire REGFILE_SIM_reg_bank__abc_33898_n8069;
  wire REGFILE_SIM_reg_bank__abc_33898_n8070;
  wire REGFILE_SIM_reg_bank__abc_33898_n8071;
  wire REGFILE_SIM_reg_bank__abc_33898_n8072;
  wire REGFILE_SIM_reg_bank__abc_33898_n8073;
  wire REGFILE_SIM_reg_bank__abc_33898_n8074;
  wire REGFILE_SIM_reg_bank__abc_33898_n8075;
  wire REGFILE_SIM_reg_bank__abc_33898_n8076;
  wire REGFILE_SIM_reg_bank__abc_33898_n8077;
  wire REGFILE_SIM_reg_bank__abc_33898_n8078;
  wire REGFILE_SIM_reg_bank__abc_33898_n8079;
  wire REGFILE_SIM_reg_bank__abc_33898_n8080;
  wire REGFILE_SIM_reg_bank__abc_33898_n8081;
  wire REGFILE_SIM_reg_bank__abc_33898_n8082;
  wire REGFILE_SIM_reg_bank__abc_33898_n8083;
  wire REGFILE_SIM_reg_bank__abc_33898_n8084;
  wire REGFILE_SIM_reg_bank__abc_33898_n8085;
  wire REGFILE_SIM_reg_bank__abc_33898_n8086;
  wire REGFILE_SIM_reg_bank__abc_33898_n8087;
  wire REGFILE_SIM_reg_bank__abc_33898_n8088;
  wire REGFILE_SIM_reg_bank__abc_33898_n8089;
  wire REGFILE_SIM_reg_bank__abc_33898_n8090;
  wire REGFILE_SIM_reg_bank__abc_33898_n8091;
  wire REGFILE_SIM_reg_bank__abc_33898_n8093;
  wire REGFILE_SIM_reg_bank__abc_33898_n8094;
  wire REGFILE_SIM_reg_bank__abc_33898_n8095;
  wire REGFILE_SIM_reg_bank__abc_33898_n8096;
  wire REGFILE_SIM_reg_bank__abc_33898_n8097;
  wire REGFILE_SIM_reg_bank__abc_33898_n8098;
  wire REGFILE_SIM_reg_bank__abc_33898_n8099;
  wire REGFILE_SIM_reg_bank__abc_33898_n8100;
  wire REGFILE_SIM_reg_bank__abc_33898_n8101;
  wire REGFILE_SIM_reg_bank__abc_33898_n8102;
  wire REGFILE_SIM_reg_bank__abc_33898_n8103;
  wire REGFILE_SIM_reg_bank__abc_33898_n8104;
  wire REGFILE_SIM_reg_bank__abc_33898_n8105;
  wire REGFILE_SIM_reg_bank__abc_33898_n8106;
  wire REGFILE_SIM_reg_bank__abc_33898_n8107;
  wire REGFILE_SIM_reg_bank__abc_33898_n8108;
  wire REGFILE_SIM_reg_bank__abc_33898_n8109;
  wire REGFILE_SIM_reg_bank__abc_33898_n8110;
  wire REGFILE_SIM_reg_bank__abc_33898_n8111;
  wire REGFILE_SIM_reg_bank__abc_33898_n8112;
  wire REGFILE_SIM_reg_bank__abc_33898_n8113;
  wire REGFILE_SIM_reg_bank__abc_33898_n8114;
  wire REGFILE_SIM_reg_bank__abc_33898_n8115;
  wire REGFILE_SIM_reg_bank__abc_33898_n8116;
  wire REGFILE_SIM_reg_bank__abc_33898_n8117;
  wire REGFILE_SIM_reg_bank__abc_33898_n8118;
  wire REGFILE_SIM_reg_bank__abc_33898_n8119;
  wire REGFILE_SIM_reg_bank__abc_33898_n8120;
  wire REGFILE_SIM_reg_bank__abc_33898_n8121;
  wire REGFILE_SIM_reg_bank__abc_33898_n8122;
  wire REGFILE_SIM_reg_bank__abc_33898_n8123;
  wire REGFILE_SIM_reg_bank__abc_33898_n8124;
  wire REGFILE_SIM_reg_bank__abc_33898_n8125;
  wire REGFILE_SIM_reg_bank__abc_33898_n8126;
  wire REGFILE_SIM_reg_bank__abc_33898_n8127;
  wire REGFILE_SIM_reg_bank__abc_33898_n8128;
  wire REGFILE_SIM_reg_bank__abc_33898_n8129;
  wire REGFILE_SIM_reg_bank__abc_33898_n8130;
  wire REGFILE_SIM_reg_bank__abc_33898_n8131;
  wire REGFILE_SIM_reg_bank__abc_33898_n8132;
  wire REGFILE_SIM_reg_bank__abc_33898_n8133;
  wire REGFILE_SIM_reg_bank__abc_33898_n8134;
  wire REGFILE_SIM_reg_bank__abc_33898_n8135;
  wire REGFILE_SIM_reg_bank__abc_33898_n8136;
  wire REGFILE_SIM_reg_bank__abc_33898_n8137;
  wire REGFILE_SIM_reg_bank__abc_33898_n8138;
  wire REGFILE_SIM_reg_bank__abc_33898_n8139;
  wire REGFILE_SIM_reg_bank__abc_33898_n8140;
  wire REGFILE_SIM_reg_bank__abc_33898_n8141;
  wire REGFILE_SIM_reg_bank__abc_33898_n8142;
  wire REGFILE_SIM_reg_bank__abc_33898_n8143;
  wire REGFILE_SIM_reg_bank__abc_33898_n8144;
  wire REGFILE_SIM_reg_bank__abc_33898_n8145;
  wire REGFILE_SIM_reg_bank__abc_33898_n8146;
  wire REGFILE_SIM_reg_bank__abc_33898_n8147;
  wire REGFILE_SIM_reg_bank__abc_33898_n8148;
  wire REGFILE_SIM_reg_bank__abc_33898_n8149;
  wire REGFILE_SIM_reg_bank__abc_33898_n8150;
  wire REGFILE_SIM_reg_bank__abc_33898_n8151;
  wire REGFILE_SIM_reg_bank__abc_33898_n8152;
  wire REGFILE_SIM_reg_bank__abc_33898_n8154;
  wire REGFILE_SIM_reg_bank__abc_33898_n8155;
  wire REGFILE_SIM_reg_bank__abc_33898_n8156;
  wire REGFILE_SIM_reg_bank__abc_33898_n8157;
  wire REGFILE_SIM_reg_bank__abc_33898_n8158;
  wire REGFILE_SIM_reg_bank__abc_33898_n8159;
  wire REGFILE_SIM_reg_bank__abc_33898_n8160;
  wire REGFILE_SIM_reg_bank__abc_33898_n8161;
  wire REGFILE_SIM_reg_bank__abc_33898_n8162;
  wire REGFILE_SIM_reg_bank__abc_33898_n8163;
  wire REGFILE_SIM_reg_bank__abc_33898_n8164;
  wire REGFILE_SIM_reg_bank__abc_33898_n8165;
  wire REGFILE_SIM_reg_bank__abc_33898_n8166;
  wire REGFILE_SIM_reg_bank__abc_33898_n8167;
  wire REGFILE_SIM_reg_bank__abc_33898_n8168;
  wire REGFILE_SIM_reg_bank__abc_33898_n8169;
  wire REGFILE_SIM_reg_bank__abc_33898_n8170;
  wire REGFILE_SIM_reg_bank__abc_33898_n8171;
  wire REGFILE_SIM_reg_bank__abc_33898_n8172;
  wire REGFILE_SIM_reg_bank__abc_33898_n8173;
  wire REGFILE_SIM_reg_bank__abc_33898_n8174;
  wire REGFILE_SIM_reg_bank__abc_33898_n8175;
  wire REGFILE_SIM_reg_bank__abc_33898_n8176;
  wire REGFILE_SIM_reg_bank__abc_33898_n8177;
  wire REGFILE_SIM_reg_bank__abc_33898_n8178;
  wire REGFILE_SIM_reg_bank__abc_33898_n8179;
  wire REGFILE_SIM_reg_bank__abc_33898_n8180;
  wire REGFILE_SIM_reg_bank__abc_33898_n8181;
  wire REGFILE_SIM_reg_bank__abc_33898_n8182;
  wire REGFILE_SIM_reg_bank__abc_33898_n8183;
  wire REGFILE_SIM_reg_bank__abc_33898_n8184;
  wire REGFILE_SIM_reg_bank__abc_33898_n8185;
  wire REGFILE_SIM_reg_bank__abc_33898_n8186;
  wire REGFILE_SIM_reg_bank__abc_33898_n8187;
  wire REGFILE_SIM_reg_bank__abc_33898_n8188;
  wire REGFILE_SIM_reg_bank__abc_33898_n8189;
  wire REGFILE_SIM_reg_bank__abc_33898_n8190;
  wire REGFILE_SIM_reg_bank__abc_33898_n8191;
  wire REGFILE_SIM_reg_bank__abc_33898_n8192;
  wire REGFILE_SIM_reg_bank__abc_33898_n8193;
  wire REGFILE_SIM_reg_bank__abc_33898_n8194;
  wire REGFILE_SIM_reg_bank__abc_33898_n8195;
  wire REGFILE_SIM_reg_bank__abc_33898_n8196;
  wire REGFILE_SIM_reg_bank__abc_33898_n8197;
  wire REGFILE_SIM_reg_bank__abc_33898_n8198;
  wire REGFILE_SIM_reg_bank__abc_33898_n8199;
  wire REGFILE_SIM_reg_bank__abc_33898_n8200;
  wire REGFILE_SIM_reg_bank__abc_33898_n8201;
  wire REGFILE_SIM_reg_bank__abc_33898_n8202;
  wire REGFILE_SIM_reg_bank__abc_33898_n8203;
  wire REGFILE_SIM_reg_bank__abc_33898_n8204;
  wire REGFILE_SIM_reg_bank__abc_33898_n8205;
  wire REGFILE_SIM_reg_bank__abc_33898_n8206;
  wire REGFILE_SIM_reg_bank__abc_33898_n8207;
  wire REGFILE_SIM_reg_bank__abc_33898_n8208;
  wire REGFILE_SIM_reg_bank__abc_33898_n8209;
  wire REGFILE_SIM_reg_bank__abc_33898_n8210;
  wire REGFILE_SIM_reg_bank__abc_33898_n8211;
  wire REGFILE_SIM_reg_bank__abc_33898_n8212;
  wire REGFILE_SIM_reg_bank__abc_33898_n8213;
  wire REGFILE_SIM_reg_bank__abc_33898_n8215;
  wire REGFILE_SIM_reg_bank__abc_33898_n8216;
  wire REGFILE_SIM_reg_bank__abc_33898_n8217;
  wire REGFILE_SIM_reg_bank__abc_33898_n8218;
  wire REGFILE_SIM_reg_bank__abc_33898_n8219;
  wire REGFILE_SIM_reg_bank__abc_33898_n8220;
  wire REGFILE_SIM_reg_bank__abc_33898_n8221;
  wire REGFILE_SIM_reg_bank__abc_33898_n8222;
  wire REGFILE_SIM_reg_bank__abc_33898_n8223;
  wire REGFILE_SIM_reg_bank__abc_33898_n8224;
  wire REGFILE_SIM_reg_bank__abc_33898_n8225;
  wire REGFILE_SIM_reg_bank__abc_33898_n8226;
  wire REGFILE_SIM_reg_bank__abc_33898_n8227;
  wire REGFILE_SIM_reg_bank__abc_33898_n8228;
  wire REGFILE_SIM_reg_bank__abc_33898_n8229;
  wire REGFILE_SIM_reg_bank__abc_33898_n8230;
  wire REGFILE_SIM_reg_bank__abc_33898_n8231;
  wire REGFILE_SIM_reg_bank__abc_33898_n8232;
  wire REGFILE_SIM_reg_bank__abc_33898_n8233;
  wire REGFILE_SIM_reg_bank__abc_33898_n8234;
  wire REGFILE_SIM_reg_bank__abc_33898_n8235;
  wire REGFILE_SIM_reg_bank__abc_33898_n8236;
  wire REGFILE_SIM_reg_bank__abc_33898_n8237;
  wire REGFILE_SIM_reg_bank__abc_33898_n8238;
  wire REGFILE_SIM_reg_bank__abc_33898_n8239;
  wire REGFILE_SIM_reg_bank__abc_33898_n8240;
  wire REGFILE_SIM_reg_bank__abc_33898_n8241;
  wire REGFILE_SIM_reg_bank__abc_33898_n8242;
  wire REGFILE_SIM_reg_bank__abc_33898_n8243;
  wire REGFILE_SIM_reg_bank__abc_33898_n8244;
  wire REGFILE_SIM_reg_bank__abc_33898_n8245;
  wire REGFILE_SIM_reg_bank__abc_33898_n8246;
  wire REGFILE_SIM_reg_bank__abc_33898_n8247;
  wire REGFILE_SIM_reg_bank__abc_33898_n8248;
  wire REGFILE_SIM_reg_bank__abc_33898_n8249;
  wire REGFILE_SIM_reg_bank__abc_33898_n8250;
  wire REGFILE_SIM_reg_bank__abc_33898_n8251;
  wire REGFILE_SIM_reg_bank__abc_33898_n8252;
  wire REGFILE_SIM_reg_bank__abc_33898_n8253;
  wire REGFILE_SIM_reg_bank__abc_33898_n8254;
  wire REGFILE_SIM_reg_bank__abc_33898_n8255;
  wire REGFILE_SIM_reg_bank__abc_33898_n8256;
  wire REGFILE_SIM_reg_bank__abc_33898_n8257;
  wire REGFILE_SIM_reg_bank__abc_33898_n8258;
  wire REGFILE_SIM_reg_bank__abc_33898_n8259;
  wire REGFILE_SIM_reg_bank__abc_33898_n8260;
  wire REGFILE_SIM_reg_bank__abc_33898_n8261;
  wire REGFILE_SIM_reg_bank__abc_33898_n8262;
  wire REGFILE_SIM_reg_bank__abc_33898_n8263;
  wire REGFILE_SIM_reg_bank__abc_33898_n8264;
  wire REGFILE_SIM_reg_bank__abc_33898_n8265;
  wire REGFILE_SIM_reg_bank__abc_33898_n8266;
  wire REGFILE_SIM_reg_bank__abc_33898_n8267;
  wire REGFILE_SIM_reg_bank__abc_33898_n8268;
  wire REGFILE_SIM_reg_bank__abc_33898_n8269;
  wire REGFILE_SIM_reg_bank__abc_33898_n8270;
  wire REGFILE_SIM_reg_bank__abc_33898_n8271;
  wire REGFILE_SIM_reg_bank__abc_33898_n8272;
  wire REGFILE_SIM_reg_bank__abc_33898_n8273;
  wire REGFILE_SIM_reg_bank__abc_33898_n8274;
  wire REGFILE_SIM_reg_bank__abc_33898_n8276;
  wire REGFILE_SIM_reg_bank__abc_33898_n8277;
  wire REGFILE_SIM_reg_bank__abc_33898_n8278;
  wire REGFILE_SIM_reg_bank__abc_33898_n8279;
  wire REGFILE_SIM_reg_bank__abc_33898_n8280;
  wire REGFILE_SIM_reg_bank__abc_33898_n8281;
  wire REGFILE_SIM_reg_bank__abc_33898_n8282;
  wire REGFILE_SIM_reg_bank__abc_33898_n8283;
  wire REGFILE_SIM_reg_bank__abc_33898_n8284;
  wire REGFILE_SIM_reg_bank__abc_33898_n8285;
  wire REGFILE_SIM_reg_bank__abc_33898_n8286;
  wire REGFILE_SIM_reg_bank__abc_33898_n8287;
  wire REGFILE_SIM_reg_bank__abc_33898_n8288;
  wire REGFILE_SIM_reg_bank__abc_33898_n8289;
  wire REGFILE_SIM_reg_bank__abc_33898_n8290;
  wire REGFILE_SIM_reg_bank__abc_33898_n8291;
  wire REGFILE_SIM_reg_bank__abc_33898_n8292;
  wire REGFILE_SIM_reg_bank__abc_33898_n8293;
  wire REGFILE_SIM_reg_bank__abc_33898_n8294;
  wire REGFILE_SIM_reg_bank__abc_33898_n8295;
  wire REGFILE_SIM_reg_bank__abc_33898_n8296;
  wire REGFILE_SIM_reg_bank__abc_33898_n8297;
  wire REGFILE_SIM_reg_bank__abc_33898_n8298;
  wire REGFILE_SIM_reg_bank__abc_33898_n8299;
  wire REGFILE_SIM_reg_bank__abc_33898_n8300;
  wire REGFILE_SIM_reg_bank__abc_33898_n8301;
  wire REGFILE_SIM_reg_bank__abc_33898_n8302;
  wire REGFILE_SIM_reg_bank__abc_33898_n8303;
  wire REGFILE_SIM_reg_bank__abc_33898_n8304;
  wire REGFILE_SIM_reg_bank__abc_33898_n8305;
  wire REGFILE_SIM_reg_bank__abc_33898_n8306;
  wire REGFILE_SIM_reg_bank__abc_33898_n8307;
  wire REGFILE_SIM_reg_bank__abc_33898_n8308;
  wire REGFILE_SIM_reg_bank__abc_33898_n8309;
  wire REGFILE_SIM_reg_bank__abc_33898_n8310;
  wire REGFILE_SIM_reg_bank__abc_33898_n8311;
  wire REGFILE_SIM_reg_bank__abc_33898_n8312;
  wire REGFILE_SIM_reg_bank__abc_33898_n8313;
  wire REGFILE_SIM_reg_bank__abc_33898_n8314;
  wire REGFILE_SIM_reg_bank__abc_33898_n8315;
  wire REGFILE_SIM_reg_bank__abc_33898_n8316;
  wire REGFILE_SIM_reg_bank__abc_33898_n8317;
  wire REGFILE_SIM_reg_bank__abc_33898_n8318;
  wire REGFILE_SIM_reg_bank__abc_33898_n8319;
  wire REGFILE_SIM_reg_bank__abc_33898_n8320;
  wire REGFILE_SIM_reg_bank__abc_33898_n8321;
  wire REGFILE_SIM_reg_bank__abc_33898_n8322;
  wire REGFILE_SIM_reg_bank__abc_33898_n8323;
  wire REGFILE_SIM_reg_bank__abc_33898_n8324;
  wire REGFILE_SIM_reg_bank__abc_33898_n8325;
  wire REGFILE_SIM_reg_bank__abc_33898_n8326;
  wire REGFILE_SIM_reg_bank__abc_33898_n8327;
  wire REGFILE_SIM_reg_bank__abc_33898_n8328;
  wire REGFILE_SIM_reg_bank__abc_33898_n8329;
  wire REGFILE_SIM_reg_bank__abc_33898_n8330;
  wire REGFILE_SIM_reg_bank__abc_33898_n8331;
  wire REGFILE_SIM_reg_bank__abc_33898_n8332;
  wire REGFILE_SIM_reg_bank__abc_33898_n8333;
  wire REGFILE_SIM_reg_bank__abc_33898_n8334;
  wire REGFILE_SIM_reg_bank__abc_33898_n8335;
  wire REGFILE_SIM_reg_bank__abc_33898_n8337;
  wire REGFILE_SIM_reg_bank__abc_33898_n8338;
  wire REGFILE_SIM_reg_bank__abc_33898_n8339;
  wire REGFILE_SIM_reg_bank__abc_33898_n8340;
  wire REGFILE_SIM_reg_bank__abc_33898_n8341;
  wire REGFILE_SIM_reg_bank__abc_33898_n8342;
  wire REGFILE_SIM_reg_bank__abc_33898_n8343;
  wire REGFILE_SIM_reg_bank__abc_33898_n8344;
  wire REGFILE_SIM_reg_bank__abc_33898_n8345;
  wire REGFILE_SIM_reg_bank__abc_33898_n8346;
  wire REGFILE_SIM_reg_bank__abc_33898_n8347;
  wire REGFILE_SIM_reg_bank__abc_33898_n8348;
  wire REGFILE_SIM_reg_bank__abc_33898_n8349;
  wire REGFILE_SIM_reg_bank__abc_33898_n8350;
  wire REGFILE_SIM_reg_bank__abc_33898_n8351;
  wire REGFILE_SIM_reg_bank__abc_33898_n8352;
  wire REGFILE_SIM_reg_bank__abc_33898_n8353;
  wire REGFILE_SIM_reg_bank__abc_33898_n8354;
  wire REGFILE_SIM_reg_bank__abc_33898_n8355;
  wire REGFILE_SIM_reg_bank__abc_33898_n8356;
  wire REGFILE_SIM_reg_bank__abc_33898_n8357;
  wire REGFILE_SIM_reg_bank__abc_33898_n8358;
  wire REGFILE_SIM_reg_bank__abc_33898_n8359;
  wire REGFILE_SIM_reg_bank__abc_33898_n8360;
  wire REGFILE_SIM_reg_bank__abc_33898_n8361;
  wire REGFILE_SIM_reg_bank__abc_33898_n8362;
  wire REGFILE_SIM_reg_bank__abc_33898_n8363;
  wire REGFILE_SIM_reg_bank__abc_33898_n8364;
  wire REGFILE_SIM_reg_bank__abc_33898_n8365;
  wire REGFILE_SIM_reg_bank__abc_33898_n8366;
  wire REGFILE_SIM_reg_bank__abc_33898_n8367;
  wire REGFILE_SIM_reg_bank__abc_33898_n8368;
  wire REGFILE_SIM_reg_bank__abc_33898_n8369;
  wire REGFILE_SIM_reg_bank__abc_33898_n8370;
  wire REGFILE_SIM_reg_bank__abc_33898_n8371;
  wire REGFILE_SIM_reg_bank__abc_33898_n8372;
  wire REGFILE_SIM_reg_bank__abc_33898_n8373;
  wire REGFILE_SIM_reg_bank__abc_33898_n8374;
  wire REGFILE_SIM_reg_bank__abc_33898_n8375;
  wire REGFILE_SIM_reg_bank__abc_33898_n8376;
  wire REGFILE_SIM_reg_bank__abc_33898_n8377;
  wire REGFILE_SIM_reg_bank__abc_33898_n8378;
  wire REGFILE_SIM_reg_bank__abc_33898_n8379;
  wire REGFILE_SIM_reg_bank__abc_33898_n8380;
  wire REGFILE_SIM_reg_bank__abc_33898_n8381;
  wire REGFILE_SIM_reg_bank__abc_33898_n8382;
  wire REGFILE_SIM_reg_bank__abc_33898_n8383;
  wire REGFILE_SIM_reg_bank__abc_33898_n8384;
  wire REGFILE_SIM_reg_bank__abc_33898_n8385;
  wire REGFILE_SIM_reg_bank__abc_33898_n8386;
  wire REGFILE_SIM_reg_bank__abc_33898_n8387;
  wire REGFILE_SIM_reg_bank__abc_33898_n8388;
  wire REGFILE_SIM_reg_bank__abc_33898_n8389;
  wire REGFILE_SIM_reg_bank__abc_33898_n8390;
  wire REGFILE_SIM_reg_bank__abc_33898_n8391;
  wire REGFILE_SIM_reg_bank__abc_33898_n8392;
  wire REGFILE_SIM_reg_bank__abc_33898_n8393;
  wire REGFILE_SIM_reg_bank__abc_33898_n8394;
  wire REGFILE_SIM_reg_bank__abc_33898_n8395;
  wire REGFILE_SIM_reg_bank__abc_33898_n8396;
  wire REGFILE_SIM_reg_bank__abc_33898_n8398;
  wire REGFILE_SIM_reg_bank__abc_33898_n8399;
  wire REGFILE_SIM_reg_bank__abc_33898_n8400;
  wire REGFILE_SIM_reg_bank__abc_33898_n8401;
  wire REGFILE_SIM_reg_bank__abc_33898_n8402;
  wire REGFILE_SIM_reg_bank__abc_33898_n8403;
  wire REGFILE_SIM_reg_bank__abc_33898_n8404;
  wire REGFILE_SIM_reg_bank__abc_33898_n8405;
  wire REGFILE_SIM_reg_bank__abc_33898_n8406;
  wire REGFILE_SIM_reg_bank__abc_33898_n8407;
  wire REGFILE_SIM_reg_bank__abc_33898_n8408;
  wire REGFILE_SIM_reg_bank__abc_33898_n8409;
  wire REGFILE_SIM_reg_bank__abc_33898_n8410;
  wire REGFILE_SIM_reg_bank__abc_33898_n8411;
  wire REGFILE_SIM_reg_bank__abc_33898_n8412;
  wire REGFILE_SIM_reg_bank__abc_33898_n8413;
  wire REGFILE_SIM_reg_bank__abc_33898_n8414;
  wire REGFILE_SIM_reg_bank__abc_33898_n8415;
  wire REGFILE_SIM_reg_bank__abc_33898_n8416;
  wire REGFILE_SIM_reg_bank__abc_33898_n8417;
  wire REGFILE_SIM_reg_bank__abc_33898_n8418;
  wire REGFILE_SIM_reg_bank__abc_33898_n8419;
  wire REGFILE_SIM_reg_bank__abc_33898_n8420;
  wire REGFILE_SIM_reg_bank__abc_33898_n8421;
  wire REGFILE_SIM_reg_bank__abc_33898_n8422;
  wire REGFILE_SIM_reg_bank__abc_33898_n8423;
  wire REGFILE_SIM_reg_bank__abc_33898_n8424;
  wire REGFILE_SIM_reg_bank__abc_33898_n8425;
  wire REGFILE_SIM_reg_bank__abc_33898_n8426;
  wire REGFILE_SIM_reg_bank__abc_33898_n8427;
  wire REGFILE_SIM_reg_bank__abc_33898_n8428;
  wire REGFILE_SIM_reg_bank__abc_33898_n8429;
  wire REGFILE_SIM_reg_bank__abc_33898_n8430;
  wire REGFILE_SIM_reg_bank__abc_33898_n8431;
  wire REGFILE_SIM_reg_bank__abc_33898_n8432;
  wire REGFILE_SIM_reg_bank__abc_33898_n8433;
  wire REGFILE_SIM_reg_bank__abc_33898_n8434;
  wire REGFILE_SIM_reg_bank__abc_33898_n8435;
  wire REGFILE_SIM_reg_bank__abc_33898_n8436;
  wire REGFILE_SIM_reg_bank__abc_33898_n8437;
  wire REGFILE_SIM_reg_bank__abc_33898_n8438;
  wire REGFILE_SIM_reg_bank__abc_33898_n8439;
  wire REGFILE_SIM_reg_bank__abc_33898_n8440;
  wire REGFILE_SIM_reg_bank__abc_33898_n8441;
  wire REGFILE_SIM_reg_bank__abc_33898_n8442;
  wire REGFILE_SIM_reg_bank__abc_33898_n8443;
  wire REGFILE_SIM_reg_bank__abc_33898_n8444;
  wire REGFILE_SIM_reg_bank__abc_33898_n8445;
  wire REGFILE_SIM_reg_bank__abc_33898_n8446;
  wire REGFILE_SIM_reg_bank__abc_33898_n8447;
  wire REGFILE_SIM_reg_bank__abc_33898_n8448;
  wire REGFILE_SIM_reg_bank__abc_33898_n8449;
  wire REGFILE_SIM_reg_bank__abc_33898_n8450;
  wire REGFILE_SIM_reg_bank__abc_33898_n8451;
  wire REGFILE_SIM_reg_bank__abc_33898_n8452;
  wire REGFILE_SIM_reg_bank__abc_33898_n8453;
  wire REGFILE_SIM_reg_bank__abc_33898_n8454;
  wire REGFILE_SIM_reg_bank__abc_33898_n8455;
  wire REGFILE_SIM_reg_bank__abc_33898_n8456;
  wire REGFILE_SIM_reg_bank__abc_33898_n8457;
  wire REGFILE_SIM_reg_bank__abc_33898_n8459;
  wire REGFILE_SIM_reg_bank__abc_33898_n8460;
  wire REGFILE_SIM_reg_bank__abc_33898_n8461;
  wire REGFILE_SIM_reg_bank__abc_33898_n8462;
  wire REGFILE_SIM_reg_bank__abc_33898_n8463;
  wire REGFILE_SIM_reg_bank__abc_33898_n8464;
  wire REGFILE_SIM_reg_bank__abc_33898_n8465;
  wire REGFILE_SIM_reg_bank__abc_33898_n8466;
  wire REGFILE_SIM_reg_bank__abc_33898_n8467;
  wire REGFILE_SIM_reg_bank__abc_33898_n8468;
  wire REGFILE_SIM_reg_bank__abc_33898_n8469;
  wire REGFILE_SIM_reg_bank__abc_33898_n8470;
  wire REGFILE_SIM_reg_bank__abc_33898_n8471;
  wire REGFILE_SIM_reg_bank__abc_33898_n8472;
  wire REGFILE_SIM_reg_bank__abc_33898_n8473;
  wire REGFILE_SIM_reg_bank__abc_33898_n8474;
  wire REGFILE_SIM_reg_bank__abc_33898_n8475;
  wire REGFILE_SIM_reg_bank__abc_33898_n8476;
  wire REGFILE_SIM_reg_bank__abc_33898_n8477;
  wire REGFILE_SIM_reg_bank__abc_33898_n8478;
  wire REGFILE_SIM_reg_bank__abc_33898_n8479;
  wire REGFILE_SIM_reg_bank__abc_33898_n8480;
  wire REGFILE_SIM_reg_bank__abc_33898_n8481;
  wire REGFILE_SIM_reg_bank__abc_33898_n8482;
  wire REGFILE_SIM_reg_bank__abc_33898_n8483;
  wire REGFILE_SIM_reg_bank__abc_33898_n8484;
  wire REGFILE_SIM_reg_bank__abc_33898_n8485;
  wire REGFILE_SIM_reg_bank__abc_33898_n8486;
  wire REGFILE_SIM_reg_bank__abc_33898_n8487;
  wire REGFILE_SIM_reg_bank__abc_33898_n8488;
  wire REGFILE_SIM_reg_bank__abc_33898_n8489;
  wire REGFILE_SIM_reg_bank__abc_33898_n8490;
  wire REGFILE_SIM_reg_bank__abc_33898_n8491;
  wire REGFILE_SIM_reg_bank__abc_33898_n8492;
  wire REGFILE_SIM_reg_bank__abc_33898_n8493;
  wire REGFILE_SIM_reg_bank__abc_33898_n8494;
  wire REGFILE_SIM_reg_bank__abc_33898_n8495;
  wire REGFILE_SIM_reg_bank__abc_33898_n8496;
  wire REGFILE_SIM_reg_bank__abc_33898_n8497;
  wire REGFILE_SIM_reg_bank__abc_33898_n8498;
  wire REGFILE_SIM_reg_bank__abc_33898_n8499;
  wire REGFILE_SIM_reg_bank__abc_33898_n8500;
  wire REGFILE_SIM_reg_bank__abc_33898_n8501;
  wire REGFILE_SIM_reg_bank__abc_33898_n8502;
  wire REGFILE_SIM_reg_bank__abc_33898_n8503;
  wire REGFILE_SIM_reg_bank__abc_33898_n8504;
  wire REGFILE_SIM_reg_bank__abc_33898_n8505;
  wire REGFILE_SIM_reg_bank__abc_33898_n8506;
  wire REGFILE_SIM_reg_bank__abc_33898_n8507;
  wire REGFILE_SIM_reg_bank__abc_33898_n8508;
  wire REGFILE_SIM_reg_bank__abc_33898_n8509;
  wire REGFILE_SIM_reg_bank__abc_33898_n8510;
  wire REGFILE_SIM_reg_bank__abc_33898_n8511;
  wire REGFILE_SIM_reg_bank__abc_33898_n8512;
  wire REGFILE_SIM_reg_bank__abc_33898_n8513;
  wire REGFILE_SIM_reg_bank__abc_33898_n8514;
  wire REGFILE_SIM_reg_bank__abc_33898_n8515;
  wire REGFILE_SIM_reg_bank__abc_33898_n8516;
  wire REGFILE_SIM_reg_bank__abc_33898_n8517;
  wire REGFILE_SIM_reg_bank__abc_33898_n8518;
  wire REGFILE_SIM_reg_bank__abc_33898_n8520;
  wire REGFILE_SIM_reg_bank__abc_33898_n8521;
  wire REGFILE_SIM_reg_bank__abc_33898_n8522;
  wire REGFILE_SIM_reg_bank__abc_33898_n8523;
  wire REGFILE_SIM_reg_bank__abc_33898_n8524;
  wire REGFILE_SIM_reg_bank__abc_33898_n8525;
  wire REGFILE_SIM_reg_bank__abc_33898_n8526;
  wire REGFILE_SIM_reg_bank__abc_33898_n8527;
  wire REGFILE_SIM_reg_bank__abc_33898_n8528;
  wire REGFILE_SIM_reg_bank__abc_33898_n8529;
  wire REGFILE_SIM_reg_bank__abc_33898_n8530;
  wire REGFILE_SIM_reg_bank__abc_33898_n8531;
  wire REGFILE_SIM_reg_bank__abc_33898_n8532;
  wire REGFILE_SIM_reg_bank__abc_33898_n8533;
  wire REGFILE_SIM_reg_bank__abc_33898_n8534;
  wire REGFILE_SIM_reg_bank__abc_33898_n8535;
  wire REGFILE_SIM_reg_bank__abc_33898_n8536;
  wire REGFILE_SIM_reg_bank__abc_33898_n8537;
  wire REGFILE_SIM_reg_bank__abc_33898_n8538;
  wire REGFILE_SIM_reg_bank__abc_33898_n8539;
  wire REGFILE_SIM_reg_bank__abc_33898_n8540;
  wire REGFILE_SIM_reg_bank__abc_33898_n8541;
  wire REGFILE_SIM_reg_bank__abc_33898_n8542;
  wire REGFILE_SIM_reg_bank__abc_33898_n8543;
  wire REGFILE_SIM_reg_bank__abc_33898_n8544;
  wire REGFILE_SIM_reg_bank__abc_33898_n8545;
  wire REGFILE_SIM_reg_bank__abc_33898_n8546;
  wire REGFILE_SIM_reg_bank__abc_33898_n8547;
  wire REGFILE_SIM_reg_bank__abc_33898_n8548;
  wire REGFILE_SIM_reg_bank__abc_33898_n8549;
  wire REGFILE_SIM_reg_bank__abc_33898_n8550;
  wire REGFILE_SIM_reg_bank__abc_33898_n8551;
  wire REGFILE_SIM_reg_bank__abc_33898_n8552;
  wire REGFILE_SIM_reg_bank__abc_33898_n8553;
  wire REGFILE_SIM_reg_bank__abc_33898_n8554;
  wire REGFILE_SIM_reg_bank__abc_33898_n8555;
  wire REGFILE_SIM_reg_bank__abc_33898_n8556;
  wire REGFILE_SIM_reg_bank__abc_33898_n8557;
  wire REGFILE_SIM_reg_bank__abc_33898_n8558;
  wire REGFILE_SIM_reg_bank__abc_33898_n8559;
  wire REGFILE_SIM_reg_bank__abc_33898_n8560;
  wire REGFILE_SIM_reg_bank__abc_33898_n8561;
  wire REGFILE_SIM_reg_bank__abc_33898_n8562;
  wire REGFILE_SIM_reg_bank__abc_33898_n8563;
  wire REGFILE_SIM_reg_bank__abc_33898_n8564;
  wire REGFILE_SIM_reg_bank__abc_33898_n8565;
  wire REGFILE_SIM_reg_bank__abc_33898_n8566;
  wire REGFILE_SIM_reg_bank__abc_33898_n8567;
  wire REGFILE_SIM_reg_bank__abc_33898_n8568;
  wire REGFILE_SIM_reg_bank__abc_33898_n8569;
  wire REGFILE_SIM_reg_bank__abc_33898_n8570;
  wire REGFILE_SIM_reg_bank__abc_33898_n8571;
  wire REGFILE_SIM_reg_bank__abc_33898_n8572;
  wire REGFILE_SIM_reg_bank__abc_33898_n8573;
  wire REGFILE_SIM_reg_bank__abc_33898_n8574;
  wire REGFILE_SIM_reg_bank__abc_33898_n8575;
  wire REGFILE_SIM_reg_bank__abc_33898_n8576;
  wire REGFILE_SIM_reg_bank__abc_33898_n8577;
  wire REGFILE_SIM_reg_bank__abc_33898_n8578;
  wire REGFILE_SIM_reg_bank__abc_33898_n8579;
  wire REGFILE_SIM_reg_bank__abc_33898_n8581;
  wire REGFILE_SIM_reg_bank__abc_33898_n8582;
  wire REGFILE_SIM_reg_bank__abc_33898_n8583;
  wire REGFILE_SIM_reg_bank__abc_33898_n8584;
  wire REGFILE_SIM_reg_bank__abc_33898_n8585;
  wire REGFILE_SIM_reg_bank__abc_33898_n8586;
  wire REGFILE_SIM_reg_bank__abc_33898_n8587;
  wire REGFILE_SIM_reg_bank__abc_33898_n8588;
  wire REGFILE_SIM_reg_bank__abc_33898_n8589;
  wire REGFILE_SIM_reg_bank__abc_33898_n8590;
  wire REGFILE_SIM_reg_bank__abc_33898_n8591;
  wire REGFILE_SIM_reg_bank__abc_33898_n8592;
  wire REGFILE_SIM_reg_bank__abc_33898_n8593;
  wire REGFILE_SIM_reg_bank__abc_33898_n8594;
  wire REGFILE_SIM_reg_bank__abc_33898_n8595;
  wire REGFILE_SIM_reg_bank__abc_33898_n8596;
  wire REGFILE_SIM_reg_bank__abc_33898_n8597;
  wire REGFILE_SIM_reg_bank__abc_33898_n8598;
  wire REGFILE_SIM_reg_bank__abc_33898_n8599;
  wire REGFILE_SIM_reg_bank__abc_33898_n8600;
  wire REGFILE_SIM_reg_bank__abc_33898_n8601;
  wire REGFILE_SIM_reg_bank__abc_33898_n8602;
  wire REGFILE_SIM_reg_bank__abc_33898_n8603;
  wire REGFILE_SIM_reg_bank__abc_33898_n8604;
  wire REGFILE_SIM_reg_bank__abc_33898_n8605;
  wire REGFILE_SIM_reg_bank__abc_33898_n8606;
  wire REGFILE_SIM_reg_bank__abc_33898_n8607;
  wire REGFILE_SIM_reg_bank__abc_33898_n8608;
  wire REGFILE_SIM_reg_bank__abc_33898_n8609;
  wire REGFILE_SIM_reg_bank__abc_33898_n8610;
  wire REGFILE_SIM_reg_bank__abc_33898_n8611;
  wire REGFILE_SIM_reg_bank__abc_33898_n8612;
  wire REGFILE_SIM_reg_bank__abc_33898_n8613;
  wire REGFILE_SIM_reg_bank__abc_33898_n8614;
  wire REGFILE_SIM_reg_bank__abc_33898_n8615;
  wire REGFILE_SIM_reg_bank__abc_33898_n8616;
  wire REGFILE_SIM_reg_bank__abc_33898_n8617;
  wire REGFILE_SIM_reg_bank__abc_33898_n8618;
  wire REGFILE_SIM_reg_bank__abc_33898_n8619;
  wire REGFILE_SIM_reg_bank__abc_33898_n8620;
  wire REGFILE_SIM_reg_bank__abc_33898_n8621;
  wire REGFILE_SIM_reg_bank__abc_33898_n8622;
  wire REGFILE_SIM_reg_bank__abc_33898_n8623;
  wire REGFILE_SIM_reg_bank__abc_33898_n8624;
  wire REGFILE_SIM_reg_bank__abc_33898_n8625;
  wire REGFILE_SIM_reg_bank__abc_33898_n8626;
  wire REGFILE_SIM_reg_bank__abc_33898_n8627;
  wire REGFILE_SIM_reg_bank__abc_33898_n8628;
  wire REGFILE_SIM_reg_bank__abc_33898_n8629;
  wire REGFILE_SIM_reg_bank__abc_33898_n8630;
  wire REGFILE_SIM_reg_bank__abc_33898_n8631;
  wire REGFILE_SIM_reg_bank__abc_33898_n8632;
  wire REGFILE_SIM_reg_bank__abc_33898_n8633;
  wire REGFILE_SIM_reg_bank__abc_33898_n8634;
  wire REGFILE_SIM_reg_bank__abc_33898_n8635;
  wire REGFILE_SIM_reg_bank__abc_33898_n8636;
  wire REGFILE_SIM_reg_bank__abc_33898_n8637;
  wire REGFILE_SIM_reg_bank__abc_33898_n8638;
  wire REGFILE_SIM_reg_bank__abc_33898_n8639;
  wire REGFILE_SIM_reg_bank__abc_33898_n8640;
  wire REGFILE_SIM_reg_bank__abc_33898_n8642;
  wire REGFILE_SIM_reg_bank__abc_33898_n8643;
  wire REGFILE_SIM_reg_bank__abc_33898_n8644;
  wire REGFILE_SIM_reg_bank__abc_33898_n8645;
  wire REGFILE_SIM_reg_bank__abc_33898_n8646;
  wire REGFILE_SIM_reg_bank__abc_33898_n8647;
  wire REGFILE_SIM_reg_bank__abc_33898_n8648;
  wire REGFILE_SIM_reg_bank__abc_33898_n8649;
  wire REGFILE_SIM_reg_bank__abc_33898_n8650;
  wire REGFILE_SIM_reg_bank__abc_33898_n8651;
  wire REGFILE_SIM_reg_bank__abc_33898_n8652;
  wire REGFILE_SIM_reg_bank__abc_33898_n8653;
  wire REGFILE_SIM_reg_bank__abc_33898_n8654;
  wire REGFILE_SIM_reg_bank__abc_33898_n8655;
  wire REGFILE_SIM_reg_bank__abc_33898_n8656;
  wire REGFILE_SIM_reg_bank__abc_33898_n8657;
  wire REGFILE_SIM_reg_bank__abc_33898_n8658;
  wire REGFILE_SIM_reg_bank__abc_33898_n8659;
  wire REGFILE_SIM_reg_bank__abc_33898_n8660;
  wire REGFILE_SIM_reg_bank__abc_33898_n8661;
  wire REGFILE_SIM_reg_bank__abc_33898_n8662;
  wire REGFILE_SIM_reg_bank__abc_33898_n8663;
  wire REGFILE_SIM_reg_bank__abc_33898_n8664;
  wire REGFILE_SIM_reg_bank__abc_33898_n8665;
  wire REGFILE_SIM_reg_bank__abc_33898_n8666;
  wire REGFILE_SIM_reg_bank__abc_33898_n8667;
  wire REGFILE_SIM_reg_bank__abc_33898_n8668;
  wire REGFILE_SIM_reg_bank__abc_33898_n8669;
  wire REGFILE_SIM_reg_bank__abc_33898_n8670;
  wire REGFILE_SIM_reg_bank__abc_33898_n8671;
  wire REGFILE_SIM_reg_bank__abc_33898_n8672;
  wire REGFILE_SIM_reg_bank__abc_33898_n8673;
  wire REGFILE_SIM_reg_bank__abc_33898_n8674;
  wire REGFILE_SIM_reg_bank__abc_33898_n8675;
  wire REGFILE_SIM_reg_bank__abc_33898_n8676;
  wire REGFILE_SIM_reg_bank__abc_33898_n8677;
  wire REGFILE_SIM_reg_bank__abc_33898_n8678;
  wire REGFILE_SIM_reg_bank__abc_33898_n8679;
  wire REGFILE_SIM_reg_bank__abc_33898_n8680;
  wire REGFILE_SIM_reg_bank__abc_33898_n8681;
  wire REGFILE_SIM_reg_bank__abc_33898_n8682;
  wire REGFILE_SIM_reg_bank__abc_33898_n8683;
  wire REGFILE_SIM_reg_bank__abc_33898_n8684;
  wire REGFILE_SIM_reg_bank__abc_33898_n8685;
  wire REGFILE_SIM_reg_bank__abc_33898_n8686;
  wire REGFILE_SIM_reg_bank__abc_33898_n8687;
  wire REGFILE_SIM_reg_bank__abc_33898_n8688;
  wire REGFILE_SIM_reg_bank__abc_33898_n8689;
  wire REGFILE_SIM_reg_bank__abc_33898_n8690;
  wire REGFILE_SIM_reg_bank__abc_33898_n8691;
  wire REGFILE_SIM_reg_bank__abc_33898_n8692;
  wire REGFILE_SIM_reg_bank__abc_33898_n8693;
  wire REGFILE_SIM_reg_bank__abc_33898_n8694;
  wire REGFILE_SIM_reg_bank__abc_33898_n8695;
  wire REGFILE_SIM_reg_bank__abc_33898_n8696;
  wire REGFILE_SIM_reg_bank__abc_33898_n8697;
  wire REGFILE_SIM_reg_bank__abc_33898_n8698;
  wire REGFILE_SIM_reg_bank__abc_33898_n8699;
  wire REGFILE_SIM_reg_bank__abc_33898_n8700;
  wire REGFILE_SIM_reg_bank__abc_33898_n8701;
  wire REGFILE_SIM_reg_bank__abc_33898_n8703;
  wire REGFILE_SIM_reg_bank__abc_33898_n8704;
  wire REGFILE_SIM_reg_bank__abc_33898_n8705;
  wire REGFILE_SIM_reg_bank__abc_33898_n8706;
  wire REGFILE_SIM_reg_bank__abc_33898_n8707;
  wire REGFILE_SIM_reg_bank__abc_33898_n8708;
  wire REGFILE_SIM_reg_bank__abc_33898_n8709;
  wire REGFILE_SIM_reg_bank__abc_33898_n8710;
  wire REGFILE_SIM_reg_bank__abc_33898_n8711;
  wire REGFILE_SIM_reg_bank__abc_33898_n8712;
  wire REGFILE_SIM_reg_bank__abc_33898_n8713;
  wire REGFILE_SIM_reg_bank__abc_33898_n8714;
  wire REGFILE_SIM_reg_bank__abc_33898_n8715;
  wire REGFILE_SIM_reg_bank__abc_33898_n8716;
  wire REGFILE_SIM_reg_bank__abc_33898_n8717;
  wire REGFILE_SIM_reg_bank__abc_33898_n8718;
  wire REGFILE_SIM_reg_bank__abc_33898_n8719;
  wire REGFILE_SIM_reg_bank__abc_33898_n8720;
  wire REGFILE_SIM_reg_bank__abc_33898_n8721;
  wire REGFILE_SIM_reg_bank__abc_33898_n8722;
  wire REGFILE_SIM_reg_bank__abc_33898_n8723;
  wire REGFILE_SIM_reg_bank__abc_33898_n8724;
  wire REGFILE_SIM_reg_bank__abc_33898_n8725;
  wire REGFILE_SIM_reg_bank__abc_33898_n8726;
  wire REGFILE_SIM_reg_bank__abc_33898_n8727;
  wire REGFILE_SIM_reg_bank__abc_33898_n8728;
  wire REGFILE_SIM_reg_bank__abc_33898_n8729;
  wire REGFILE_SIM_reg_bank__abc_33898_n8730;
  wire REGFILE_SIM_reg_bank__abc_33898_n8731;
  wire REGFILE_SIM_reg_bank__abc_33898_n8732;
  wire REGFILE_SIM_reg_bank__abc_33898_n8733;
  wire REGFILE_SIM_reg_bank__abc_33898_n8734;
  wire REGFILE_SIM_reg_bank__abc_33898_n8735;
  wire REGFILE_SIM_reg_bank__abc_33898_n8736;
  wire REGFILE_SIM_reg_bank__abc_33898_n8737;
  wire REGFILE_SIM_reg_bank__abc_33898_n8738;
  wire REGFILE_SIM_reg_bank__abc_33898_n8739;
  wire REGFILE_SIM_reg_bank__abc_33898_n8740;
  wire REGFILE_SIM_reg_bank__abc_33898_n8741;
  wire REGFILE_SIM_reg_bank__abc_33898_n8742;
  wire REGFILE_SIM_reg_bank__abc_33898_n8743;
  wire REGFILE_SIM_reg_bank__abc_33898_n8744;
  wire REGFILE_SIM_reg_bank__abc_33898_n8745;
  wire REGFILE_SIM_reg_bank__abc_33898_n8746;
  wire REGFILE_SIM_reg_bank__abc_33898_n8747;
  wire REGFILE_SIM_reg_bank__abc_33898_n8748;
  wire REGFILE_SIM_reg_bank__abc_33898_n8749;
  wire REGFILE_SIM_reg_bank__abc_33898_n8750;
  wire REGFILE_SIM_reg_bank__abc_33898_n8751;
  wire REGFILE_SIM_reg_bank__abc_33898_n8752;
  wire REGFILE_SIM_reg_bank__abc_33898_n8753;
  wire REGFILE_SIM_reg_bank__abc_33898_n8754;
  wire REGFILE_SIM_reg_bank__abc_33898_n8755;
  wire REGFILE_SIM_reg_bank__abc_33898_n8756;
  wire REGFILE_SIM_reg_bank__abc_33898_n8757;
  wire REGFILE_SIM_reg_bank__abc_33898_n8758;
  wire REGFILE_SIM_reg_bank__abc_33898_n8759;
  wire REGFILE_SIM_reg_bank__abc_33898_n8760;
  wire REGFILE_SIM_reg_bank__abc_33898_n8761;
  wire REGFILE_SIM_reg_bank__abc_33898_n8762;
  wire REGFILE_SIM_reg_bank__abc_33898_n8764;
  wire REGFILE_SIM_reg_bank__abc_33898_n8765;
  wire REGFILE_SIM_reg_bank__abc_33898_n8766;
  wire REGFILE_SIM_reg_bank__abc_33898_n8767;
  wire REGFILE_SIM_reg_bank__abc_33898_n8768;
  wire REGFILE_SIM_reg_bank__abc_33898_n8769;
  wire REGFILE_SIM_reg_bank__abc_33898_n8770;
  wire REGFILE_SIM_reg_bank__abc_33898_n8771;
  wire REGFILE_SIM_reg_bank__abc_33898_n8772;
  wire REGFILE_SIM_reg_bank__abc_33898_n8773;
  wire REGFILE_SIM_reg_bank__abc_33898_n8774;
  wire REGFILE_SIM_reg_bank__abc_33898_n8775;
  wire REGFILE_SIM_reg_bank__abc_33898_n8776;
  wire REGFILE_SIM_reg_bank__abc_33898_n8777;
  wire REGFILE_SIM_reg_bank__abc_33898_n8778;
  wire REGFILE_SIM_reg_bank__abc_33898_n8779;
  wire REGFILE_SIM_reg_bank__abc_33898_n8780;
  wire REGFILE_SIM_reg_bank__abc_33898_n8781;
  wire REGFILE_SIM_reg_bank__abc_33898_n8782;
  wire REGFILE_SIM_reg_bank__abc_33898_n8783;
  wire REGFILE_SIM_reg_bank__abc_33898_n8784;
  wire REGFILE_SIM_reg_bank__abc_33898_n8785;
  wire REGFILE_SIM_reg_bank__abc_33898_n8786;
  wire REGFILE_SIM_reg_bank__abc_33898_n8787;
  wire REGFILE_SIM_reg_bank__abc_33898_n8788;
  wire REGFILE_SIM_reg_bank__abc_33898_n8789;
  wire REGFILE_SIM_reg_bank__abc_33898_n8790;
  wire REGFILE_SIM_reg_bank__abc_33898_n8791;
  wire REGFILE_SIM_reg_bank__abc_33898_n8792;
  wire REGFILE_SIM_reg_bank__abc_33898_n8793;
  wire REGFILE_SIM_reg_bank__abc_33898_n8794;
  wire REGFILE_SIM_reg_bank__abc_33898_n8795;
  wire REGFILE_SIM_reg_bank__abc_33898_n8796;
  wire REGFILE_SIM_reg_bank__abc_33898_n8797;
  wire REGFILE_SIM_reg_bank__abc_33898_n8798;
  wire REGFILE_SIM_reg_bank__abc_33898_n8799;
  wire REGFILE_SIM_reg_bank__abc_33898_n8800;
  wire REGFILE_SIM_reg_bank__abc_33898_n8801;
  wire REGFILE_SIM_reg_bank__abc_33898_n8802;
  wire REGFILE_SIM_reg_bank__abc_33898_n8803;
  wire REGFILE_SIM_reg_bank__abc_33898_n8804;
  wire REGFILE_SIM_reg_bank__abc_33898_n8805;
  wire REGFILE_SIM_reg_bank__abc_33898_n8806;
  wire REGFILE_SIM_reg_bank__abc_33898_n8807;
  wire REGFILE_SIM_reg_bank__abc_33898_n8808;
  wire REGFILE_SIM_reg_bank__abc_33898_n8809;
  wire REGFILE_SIM_reg_bank__abc_33898_n8810;
  wire REGFILE_SIM_reg_bank__abc_33898_n8811;
  wire REGFILE_SIM_reg_bank__abc_33898_n8812;
  wire REGFILE_SIM_reg_bank__abc_33898_n8813;
  wire REGFILE_SIM_reg_bank__abc_33898_n8814;
  wire REGFILE_SIM_reg_bank__abc_33898_n8815;
  wire REGFILE_SIM_reg_bank__abc_33898_n8816;
  wire REGFILE_SIM_reg_bank__abc_33898_n8817;
  wire REGFILE_SIM_reg_bank__abc_33898_n8818;
  wire REGFILE_SIM_reg_bank__abc_33898_n8819;
  wire REGFILE_SIM_reg_bank__abc_33898_n8820;
  wire REGFILE_SIM_reg_bank__abc_33898_n8821;
  wire REGFILE_SIM_reg_bank__abc_33898_n8822;
  wire REGFILE_SIM_reg_bank__abc_33898_n8823;
  wire REGFILE_SIM_reg_bank__abc_33898_n8825;
  wire REGFILE_SIM_reg_bank__abc_33898_n8826;
  wire REGFILE_SIM_reg_bank__abc_33898_n8827;
  wire REGFILE_SIM_reg_bank__abc_33898_n8828;
  wire REGFILE_SIM_reg_bank__abc_33898_n8829;
  wire REGFILE_SIM_reg_bank__abc_33898_n8830;
  wire REGFILE_SIM_reg_bank__abc_33898_n8831;
  wire REGFILE_SIM_reg_bank__abc_33898_n8832;
  wire REGFILE_SIM_reg_bank__abc_33898_n8833;
  wire REGFILE_SIM_reg_bank__abc_33898_n8834;
  wire REGFILE_SIM_reg_bank__abc_33898_n8835;
  wire REGFILE_SIM_reg_bank__abc_33898_n8836;
  wire REGFILE_SIM_reg_bank__abc_33898_n8837;
  wire REGFILE_SIM_reg_bank__abc_33898_n8838;
  wire REGFILE_SIM_reg_bank__abc_33898_n8839;
  wire REGFILE_SIM_reg_bank__abc_33898_n8840;
  wire REGFILE_SIM_reg_bank__abc_33898_n8841;
  wire REGFILE_SIM_reg_bank__abc_33898_n8842;
  wire REGFILE_SIM_reg_bank__abc_33898_n8843;
  wire REGFILE_SIM_reg_bank__abc_33898_n8844;
  wire REGFILE_SIM_reg_bank__abc_33898_n8845;
  wire REGFILE_SIM_reg_bank__abc_33898_n8846;
  wire REGFILE_SIM_reg_bank__abc_33898_n8847;
  wire REGFILE_SIM_reg_bank__abc_33898_n8848;
  wire REGFILE_SIM_reg_bank__abc_33898_n8849;
  wire REGFILE_SIM_reg_bank__abc_33898_n8850;
  wire REGFILE_SIM_reg_bank__abc_33898_n8851;
  wire REGFILE_SIM_reg_bank__abc_33898_n8852;
  wire REGFILE_SIM_reg_bank__abc_33898_n8853;
  wire REGFILE_SIM_reg_bank__abc_33898_n8854;
  wire REGFILE_SIM_reg_bank__abc_33898_n8855;
  wire REGFILE_SIM_reg_bank__abc_33898_n8856;
  wire REGFILE_SIM_reg_bank__abc_33898_n8857;
  wire REGFILE_SIM_reg_bank__abc_33898_n8858;
  wire REGFILE_SIM_reg_bank__abc_33898_n8859;
  wire REGFILE_SIM_reg_bank__abc_33898_n8860;
  wire REGFILE_SIM_reg_bank__abc_33898_n8861;
  wire REGFILE_SIM_reg_bank__abc_33898_n8862;
  wire REGFILE_SIM_reg_bank__abc_33898_n8863;
  wire REGFILE_SIM_reg_bank__abc_33898_n8864;
  wire REGFILE_SIM_reg_bank__abc_33898_n8865;
  wire REGFILE_SIM_reg_bank__abc_33898_n8866;
  wire REGFILE_SIM_reg_bank__abc_33898_n8867;
  wire REGFILE_SIM_reg_bank__abc_33898_n8868;
  wire REGFILE_SIM_reg_bank__abc_33898_n8869;
  wire REGFILE_SIM_reg_bank__abc_33898_n8870;
  wire REGFILE_SIM_reg_bank__abc_33898_n8871;
  wire REGFILE_SIM_reg_bank__abc_33898_n8872;
  wire REGFILE_SIM_reg_bank__abc_33898_n8873;
  wire REGFILE_SIM_reg_bank__abc_33898_n8874;
  wire REGFILE_SIM_reg_bank__abc_33898_n8875;
  wire REGFILE_SIM_reg_bank__abc_33898_n8876;
  wire REGFILE_SIM_reg_bank__abc_33898_n8877;
  wire REGFILE_SIM_reg_bank__abc_33898_n8878;
  wire REGFILE_SIM_reg_bank__abc_33898_n8879;
  wire REGFILE_SIM_reg_bank__abc_33898_n8880;
  wire REGFILE_SIM_reg_bank__abc_33898_n8881;
  wire REGFILE_SIM_reg_bank__abc_33898_n8882;
  wire REGFILE_SIM_reg_bank__abc_33898_n8883;
  wire REGFILE_SIM_reg_bank__abc_33898_n8884;
  wire REGFILE_SIM_reg_bank__abc_33898_n8886;
  wire REGFILE_SIM_reg_bank__abc_33898_n8887;
  wire REGFILE_SIM_reg_bank__abc_33898_n8888;
  wire REGFILE_SIM_reg_bank__abc_33898_n8889;
  wire REGFILE_SIM_reg_bank__abc_33898_n8890;
  wire REGFILE_SIM_reg_bank__abc_33898_n8891;
  wire REGFILE_SIM_reg_bank__abc_33898_n8892;
  wire REGFILE_SIM_reg_bank__abc_33898_n8893;
  wire REGFILE_SIM_reg_bank__abc_33898_n8894;
  wire REGFILE_SIM_reg_bank__abc_33898_n8895;
  wire REGFILE_SIM_reg_bank__abc_33898_n8896;
  wire REGFILE_SIM_reg_bank__abc_33898_n8897;
  wire REGFILE_SIM_reg_bank__abc_33898_n8898;
  wire REGFILE_SIM_reg_bank__abc_33898_n8899;
  wire REGFILE_SIM_reg_bank__abc_33898_n8900;
  wire REGFILE_SIM_reg_bank__abc_33898_n8901;
  wire REGFILE_SIM_reg_bank__abc_33898_n8902;
  wire REGFILE_SIM_reg_bank__abc_33898_n8903;
  wire REGFILE_SIM_reg_bank__abc_33898_n8904;
  wire REGFILE_SIM_reg_bank__abc_33898_n8905;
  wire REGFILE_SIM_reg_bank__abc_33898_n8906;
  wire REGFILE_SIM_reg_bank__abc_33898_n8907;
  wire REGFILE_SIM_reg_bank__abc_33898_n8908;
  wire REGFILE_SIM_reg_bank__abc_33898_n8909;
  wire REGFILE_SIM_reg_bank__abc_33898_n8910;
  wire REGFILE_SIM_reg_bank__abc_33898_n8911;
  wire REGFILE_SIM_reg_bank__abc_33898_n8912;
  wire REGFILE_SIM_reg_bank__abc_33898_n8913;
  wire REGFILE_SIM_reg_bank__abc_33898_n8914;
  wire REGFILE_SIM_reg_bank__abc_33898_n8915;
  wire REGFILE_SIM_reg_bank__abc_33898_n8916;
  wire REGFILE_SIM_reg_bank__abc_33898_n8917;
  wire REGFILE_SIM_reg_bank__abc_33898_n8918;
  wire REGFILE_SIM_reg_bank__abc_33898_n8919;
  wire REGFILE_SIM_reg_bank__abc_33898_n8920;
  wire REGFILE_SIM_reg_bank__abc_33898_n8921;
  wire REGFILE_SIM_reg_bank__abc_33898_n8922;
  wire REGFILE_SIM_reg_bank__abc_33898_n8923;
  wire REGFILE_SIM_reg_bank__abc_33898_n8924;
  wire REGFILE_SIM_reg_bank__abc_33898_n8925;
  wire REGFILE_SIM_reg_bank__abc_33898_n8926;
  wire REGFILE_SIM_reg_bank__abc_33898_n8927;
  wire REGFILE_SIM_reg_bank__abc_33898_n8928;
  wire REGFILE_SIM_reg_bank__abc_33898_n8929;
  wire REGFILE_SIM_reg_bank__abc_33898_n8930;
  wire REGFILE_SIM_reg_bank__abc_33898_n8931;
  wire REGFILE_SIM_reg_bank__abc_33898_n8932;
  wire REGFILE_SIM_reg_bank__abc_33898_n8933;
  wire REGFILE_SIM_reg_bank__abc_33898_n8934;
  wire REGFILE_SIM_reg_bank__abc_33898_n8935;
  wire REGFILE_SIM_reg_bank__abc_33898_n8936;
  wire REGFILE_SIM_reg_bank__abc_33898_n8937;
  wire REGFILE_SIM_reg_bank__abc_33898_n8938;
  wire REGFILE_SIM_reg_bank__abc_33898_n8939;
  wire REGFILE_SIM_reg_bank__abc_33898_n8940;
  wire REGFILE_SIM_reg_bank__abc_33898_n8941;
  wire REGFILE_SIM_reg_bank__abc_33898_n8942;
  wire REGFILE_SIM_reg_bank__abc_33898_n8943;
  wire REGFILE_SIM_reg_bank__abc_33898_n8944;
  wire REGFILE_SIM_reg_bank__abc_33898_n8945;
  wire REGFILE_SIM_reg_bank__abc_33898_n8947;
  wire REGFILE_SIM_reg_bank__abc_33898_n8948;
  wire REGFILE_SIM_reg_bank__abc_33898_n8949;
  wire REGFILE_SIM_reg_bank__abc_33898_n8950;
  wire REGFILE_SIM_reg_bank__abc_33898_n8951;
  wire REGFILE_SIM_reg_bank__abc_33898_n8952;
  wire REGFILE_SIM_reg_bank__abc_33898_n8953;
  wire REGFILE_SIM_reg_bank__abc_33898_n8954;
  wire REGFILE_SIM_reg_bank__abc_33898_n8955;
  wire REGFILE_SIM_reg_bank__abc_33898_n8956;
  wire REGFILE_SIM_reg_bank__abc_33898_n8957;
  wire REGFILE_SIM_reg_bank__abc_33898_n8958;
  wire REGFILE_SIM_reg_bank__abc_33898_n8959;
  wire REGFILE_SIM_reg_bank__abc_33898_n8960;
  wire REGFILE_SIM_reg_bank__abc_33898_n8961;
  wire REGFILE_SIM_reg_bank__abc_33898_n8962;
  wire REGFILE_SIM_reg_bank__abc_33898_n8963;
  wire REGFILE_SIM_reg_bank__abc_33898_n8964;
  wire REGFILE_SIM_reg_bank__abc_33898_n8965;
  wire REGFILE_SIM_reg_bank__abc_33898_n8966;
  wire REGFILE_SIM_reg_bank__abc_33898_n8967;
  wire REGFILE_SIM_reg_bank__abc_33898_n8968;
  wire REGFILE_SIM_reg_bank__abc_33898_n8969;
  wire REGFILE_SIM_reg_bank__abc_33898_n8970;
  wire REGFILE_SIM_reg_bank__abc_33898_n8971;
  wire REGFILE_SIM_reg_bank__abc_33898_n8972;
  wire REGFILE_SIM_reg_bank__abc_33898_n8973;
  wire REGFILE_SIM_reg_bank__abc_33898_n8974;
  wire REGFILE_SIM_reg_bank__abc_33898_n8975;
  wire REGFILE_SIM_reg_bank__abc_33898_n8976;
  wire REGFILE_SIM_reg_bank__abc_33898_n8977;
  wire REGFILE_SIM_reg_bank__abc_33898_n8978;
  wire REGFILE_SIM_reg_bank__abc_33898_n8979;
  wire REGFILE_SIM_reg_bank__abc_33898_n8980;
  wire REGFILE_SIM_reg_bank__abc_33898_n8981;
  wire REGFILE_SIM_reg_bank__abc_33898_n8982;
  wire REGFILE_SIM_reg_bank__abc_33898_n8983;
  wire REGFILE_SIM_reg_bank__abc_33898_n8984;
  wire REGFILE_SIM_reg_bank__abc_33898_n8985;
  wire REGFILE_SIM_reg_bank__abc_33898_n8986;
  wire REGFILE_SIM_reg_bank__abc_33898_n8987;
  wire REGFILE_SIM_reg_bank__abc_33898_n8988;
  wire REGFILE_SIM_reg_bank__abc_33898_n8989;
  wire REGFILE_SIM_reg_bank__abc_33898_n8990;
  wire REGFILE_SIM_reg_bank__abc_33898_n8991;
  wire REGFILE_SIM_reg_bank__abc_33898_n8992;
  wire REGFILE_SIM_reg_bank__abc_33898_n8993;
  wire REGFILE_SIM_reg_bank__abc_33898_n8994;
  wire REGFILE_SIM_reg_bank__abc_33898_n8995;
  wire REGFILE_SIM_reg_bank__abc_33898_n8996;
  wire REGFILE_SIM_reg_bank__abc_33898_n8997;
  wire REGFILE_SIM_reg_bank__abc_33898_n8998;
  wire REGFILE_SIM_reg_bank__abc_33898_n8999;
  wire REGFILE_SIM_reg_bank__abc_33898_n9000;
  wire REGFILE_SIM_reg_bank__abc_33898_n9001;
  wire REGFILE_SIM_reg_bank__abc_33898_n9002;
  wire REGFILE_SIM_reg_bank__abc_33898_n9003;
  wire REGFILE_SIM_reg_bank__abc_33898_n9004;
  wire REGFILE_SIM_reg_bank__abc_33898_n9005;
  wire REGFILE_SIM_reg_bank__abc_33898_n9006;
  wire REGFILE_SIM_reg_bank__abc_33898_n9008;
  wire REGFILE_SIM_reg_bank__abc_33898_n9009;
  wire REGFILE_SIM_reg_bank__abc_33898_n9010;
  wire REGFILE_SIM_reg_bank__abc_33898_n9011;
  wire REGFILE_SIM_reg_bank__abc_33898_n9012;
  wire REGFILE_SIM_reg_bank__abc_33898_n9013;
  wire REGFILE_SIM_reg_bank__abc_33898_n9014;
  wire REGFILE_SIM_reg_bank__abc_33898_n9015;
  wire REGFILE_SIM_reg_bank__abc_33898_n9016;
  wire REGFILE_SIM_reg_bank__abc_33898_n9017;
  wire REGFILE_SIM_reg_bank__abc_33898_n9018;
  wire REGFILE_SIM_reg_bank__abc_33898_n9019;
  wire REGFILE_SIM_reg_bank__abc_33898_n9020;
  wire REGFILE_SIM_reg_bank__abc_33898_n9021;
  wire REGFILE_SIM_reg_bank__abc_33898_n9022;
  wire REGFILE_SIM_reg_bank__abc_33898_n9023;
  wire REGFILE_SIM_reg_bank__abc_33898_n9024;
  wire REGFILE_SIM_reg_bank__abc_33898_n9025;
  wire REGFILE_SIM_reg_bank__abc_33898_n9026;
  wire REGFILE_SIM_reg_bank__abc_33898_n9027;
  wire REGFILE_SIM_reg_bank__abc_33898_n9028;
  wire REGFILE_SIM_reg_bank__abc_33898_n9029;
  wire REGFILE_SIM_reg_bank__abc_33898_n9030;
  wire REGFILE_SIM_reg_bank__abc_33898_n9031;
  wire REGFILE_SIM_reg_bank__abc_33898_n9032;
  wire REGFILE_SIM_reg_bank__abc_33898_n9033;
  wire REGFILE_SIM_reg_bank__abc_33898_n9034;
  wire REGFILE_SIM_reg_bank__abc_33898_n9035;
  wire REGFILE_SIM_reg_bank__abc_33898_n9036;
  wire REGFILE_SIM_reg_bank__abc_33898_n9037;
  wire REGFILE_SIM_reg_bank__abc_33898_n9038;
  wire REGFILE_SIM_reg_bank__abc_33898_n9039;
  wire REGFILE_SIM_reg_bank__abc_33898_n9040;
  wire REGFILE_SIM_reg_bank__abc_33898_n9041;
  wire REGFILE_SIM_reg_bank__abc_33898_n9042;
  wire REGFILE_SIM_reg_bank__abc_33898_n9043;
  wire REGFILE_SIM_reg_bank__abc_33898_n9044;
  wire REGFILE_SIM_reg_bank__abc_33898_n9045;
  wire REGFILE_SIM_reg_bank__abc_33898_n9046;
  wire REGFILE_SIM_reg_bank__abc_33898_n9047;
  wire REGFILE_SIM_reg_bank__abc_33898_n9048;
  wire REGFILE_SIM_reg_bank__abc_33898_n9049;
  wire REGFILE_SIM_reg_bank__abc_33898_n9050;
  wire REGFILE_SIM_reg_bank__abc_33898_n9051;
  wire REGFILE_SIM_reg_bank__abc_33898_n9052;
  wire REGFILE_SIM_reg_bank__abc_33898_n9053;
  wire REGFILE_SIM_reg_bank__abc_33898_n9054;
  wire REGFILE_SIM_reg_bank__abc_33898_n9055;
  wire REGFILE_SIM_reg_bank__abc_33898_n9056;
  wire REGFILE_SIM_reg_bank__abc_33898_n9057;
  wire REGFILE_SIM_reg_bank__abc_33898_n9058;
  wire REGFILE_SIM_reg_bank__abc_33898_n9059;
  wire REGFILE_SIM_reg_bank__abc_33898_n9060;
  wire REGFILE_SIM_reg_bank__abc_33898_n9061;
  wire REGFILE_SIM_reg_bank__abc_33898_n9062;
  wire REGFILE_SIM_reg_bank__abc_33898_n9063;
  wire REGFILE_SIM_reg_bank__abc_33898_n9064;
  wire REGFILE_SIM_reg_bank__abc_33898_n9065;
  wire REGFILE_SIM_reg_bank__abc_33898_n9066;
  wire REGFILE_SIM_reg_bank__abc_33898_n9067;
  wire REGFILE_SIM_reg_bank__abc_33898_n9069;
  wire REGFILE_SIM_reg_bank__abc_33898_n9070;
  wire REGFILE_SIM_reg_bank__abc_33898_n9071;
  wire REGFILE_SIM_reg_bank__abc_33898_n9072;
  wire REGFILE_SIM_reg_bank__abc_33898_n9073;
  wire REGFILE_SIM_reg_bank__abc_33898_n9074;
  wire REGFILE_SIM_reg_bank__abc_33898_n9075;
  wire REGFILE_SIM_reg_bank__abc_33898_n9076;
  wire REGFILE_SIM_reg_bank__abc_33898_n9077;
  wire REGFILE_SIM_reg_bank__abc_33898_n9078;
  wire REGFILE_SIM_reg_bank__abc_33898_n9079;
  wire REGFILE_SIM_reg_bank__abc_33898_n9080;
  wire REGFILE_SIM_reg_bank__abc_33898_n9081;
  wire REGFILE_SIM_reg_bank__abc_33898_n9082;
  wire REGFILE_SIM_reg_bank__abc_33898_n9083;
  wire REGFILE_SIM_reg_bank__abc_33898_n9084;
  wire REGFILE_SIM_reg_bank__abc_33898_n9085;
  wire REGFILE_SIM_reg_bank__abc_33898_n9086;
  wire REGFILE_SIM_reg_bank__abc_33898_n9087;
  wire REGFILE_SIM_reg_bank__abc_33898_n9088;
  wire REGFILE_SIM_reg_bank__abc_33898_n9089;
  wire REGFILE_SIM_reg_bank__abc_33898_n9090;
  wire REGFILE_SIM_reg_bank__abc_33898_n9091;
  wire REGFILE_SIM_reg_bank__abc_33898_n9092;
  wire REGFILE_SIM_reg_bank__abc_33898_n9093;
  wire REGFILE_SIM_reg_bank__abc_33898_n9094;
  wire REGFILE_SIM_reg_bank__abc_33898_n9095;
  wire REGFILE_SIM_reg_bank__abc_33898_n9096;
  wire REGFILE_SIM_reg_bank__abc_33898_n9097;
  wire REGFILE_SIM_reg_bank__abc_33898_n9098;
  wire REGFILE_SIM_reg_bank__abc_33898_n9099;
  wire REGFILE_SIM_reg_bank__abc_33898_n9100;
  wire REGFILE_SIM_reg_bank__abc_33898_n9101;
  wire REGFILE_SIM_reg_bank__abc_33898_n9102;
  wire REGFILE_SIM_reg_bank__abc_33898_n9103;
  wire REGFILE_SIM_reg_bank__abc_33898_n9104;
  wire REGFILE_SIM_reg_bank__abc_33898_n9105;
  wire REGFILE_SIM_reg_bank__abc_33898_n9106;
  wire REGFILE_SIM_reg_bank__abc_33898_n9107;
  wire REGFILE_SIM_reg_bank__abc_33898_n9108;
  wire REGFILE_SIM_reg_bank__abc_33898_n9109;
  wire REGFILE_SIM_reg_bank__abc_33898_n9110;
  wire REGFILE_SIM_reg_bank__abc_33898_n9111;
  wire REGFILE_SIM_reg_bank__abc_33898_n9112;
  wire REGFILE_SIM_reg_bank__abc_33898_n9113;
  wire REGFILE_SIM_reg_bank__abc_33898_n9114;
  wire REGFILE_SIM_reg_bank__abc_33898_n9115;
  wire REGFILE_SIM_reg_bank__abc_33898_n9116;
  wire REGFILE_SIM_reg_bank__abc_33898_n9117;
  wire REGFILE_SIM_reg_bank__abc_33898_n9118;
  wire REGFILE_SIM_reg_bank__abc_33898_n9119;
  wire REGFILE_SIM_reg_bank__abc_33898_n9120;
  wire REGFILE_SIM_reg_bank__abc_33898_n9121;
  wire REGFILE_SIM_reg_bank__abc_33898_n9122;
  wire REGFILE_SIM_reg_bank__abc_33898_n9123;
  wire REGFILE_SIM_reg_bank__abc_33898_n9124;
  wire REGFILE_SIM_reg_bank__abc_33898_n9125;
  wire REGFILE_SIM_reg_bank__abc_33898_n9126;
  wire REGFILE_SIM_reg_bank__abc_33898_n9127;
  wire REGFILE_SIM_reg_bank__abc_33898_n9128;
  wire REGFILE_SIM_reg_bank__abc_33898_n9130;
  wire REGFILE_SIM_reg_bank__abc_33898_n9131;
  wire REGFILE_SIM_reg_bank__abc_33898_n9132;
  wire REGFILE_SIM_reg_bank__abc_33898_n9133;
  wire REGFILE_SIM_reg_bank__abc_33898_n9134;
  wire REGFILE_SIM_reg_bank__abc_33898_n9135;
  wire REGFILE_SIM_reg_bank__abc_33898_n9136;
  wire REGFILE_SIM_reg_bank__abc_33898_n9137;
  wire REGFILE_SIM_reg_bank__abc_33898_n9138;
  wire REGFILE_SIM_reg_bank__abc_33898_n9139;
  wire REGFILE_SIM_reg_bank__abc_33898_n9140;
  wire REGFILE_SIM_reg_bank__abc_33898_n9141;
  wire REGFILE_SIM_reg_bank__abc_33898_n9142;
  wire REGFILE_SIM_reg_bank__abc_33898_n9143;
  wire REGFILE_SIM_reg_bank__abc_33898_n9144;
  wire REGFILE_SIM_reg_bank__abc_33898_n9145;
  wire REGFILE_SIM_reg_bank__abc_33898_n9146;
  wire REGFILE_SIM_reg_bank__abc_33898_n9147;
  wire REGFILE_SIM_reg_bank__abc_33898_n9148;
  wire REGFILE_SIM_reg_bank__abc_33898_n9149;
  wire REGFILE_SIM_reg_bank__abc_33898_n9150;
  wire REGFILE_SIM_reg_bank__abc_33898_n9151;
  wire REGFILE_SIM_reg_bank__abc_33898_n9152;
  wire REGFILE_SIM_reg_bank__abc_33898_n9153;
  wire REGFILE_SIM_reg_bank__abc_33898_n9154;
  wire REGFILE_SIM_reg_bank__abc_33898_n9155;
  wire REGFILE_SIM_reg_bank__abc_33898_n9156;
  wire REGFILE_SIM_reg_bank__abc_33898_n9157;
  wire REGFILE_SIM_reg_bank__abc_33898_n9158;
  wire REGFILE_SIM_reg_bank__abc_33898_n9159;
  wire REGFILE_SIM_reg_bank__abc_33898_n9160;
  wire REGFILE_SIM_reg_bank__abc_33898_n9161;
  wire REGFILE_SIM_reg_bank__abc_33898_n9162;
  wire REGFILE_SIM_reg_bank__abc_33898_n9163;
  wire REGFILE_SIM_reg_bank__abc_33898_n9164;
  wire REGFILE_SIM_reg_bank__abc_33898_n9165;
  wire REGFILE_SIM_reg_bank__abc_33898_n9166;
  wire REGFILE_SIM_reg_bank__abc_33898_n9167;
  wire REGFILE_SIM_reg_bank__abc_33898_n9168;
  wire REGFILE_SIM_reg_bank__abc_33898_n9169;
  wire REGFILE_SIM_reg_bank__abc_33898_n9170;
  wire REGFILE_SIM_reg_bank__abc_33898_n9171;
  wire REGFILE_SIM_reg_bank__abc_33898_n9172;
  wire REGFILE_SIM_reg_bank__abc_33898_n9173;
  wire REGFILE_SIM_reg_bank__abc_33898_n9174;
  wire REGFILE_SIM_reg_bank__abc_33898_n9175;
  wire REGFILE_SIM_reg_bank__abc_33898_n9176;
  wire REGFILE_SIM_reg_bank__abc_33898_n9177;
  wire REGFILE_SIM_reg_bank__abc_33898_n9178;
  wire REGFILE_SIM_reg_bank__abc_33898_n9179;
  wire REGFILE_SIM_reg_bank__abc_33898_n9180;
  wire REGFILE_SIM_reg_bank__abc_33898_n9181;
  wire REGFILE_SIM_reg_bank__abc_33898_n9182;
  wire REGFILE_SIM_reg_bank__abc_33898_n9183;
  wire REGFILE_SIM_reg_bank__abc_33898_n9184;
  wire REGFILE_SIM_reg_bank__abc_33898_n9185;
  wire REGFILE_SIM_reg_bank__abc_33898_n9186;
  wire REGFILE_SIM_reg_bank__abc_33898_n9187;
  wire REGFILE_SIM_reg_bank__abc_33898_n9188;
  wire REGFILE_SIM_reg_bank__abc_33898_n9189;
  wire REGFILE_SIM_reg_bank__abc_33898_n9191;
  wire REGFILE_SIM_reg_bank__abc_33898_n9192;
  wire REGFILE_SIM_reg_bank__abc_33898_n9193;
  wire REGFILE_SIM_reg_bank__abc_33898_n9194;
  wire REGFILE_SIM_reg_bank__abc_33898_n9195;
  wire REGFILE_SIM_reg_bank__abc_33898_n9196;
  wire REGFILE_SIM_reg_bank__abc_33898_n9197;
  wire REGFILE_SIM_reg_bank__abc_33898_n9198;
  wire REGFILE_SIM_reg_bank__abc_33898_n9199;
  wire REGFILE_SIM_reg_bank__abc_33898_n9200;
  wire REGFILE_SIM_reg_bank__abc_33898_n9201;
  wire REGFILE_SIM_reg_bank__abc_33898_n9202;
  wire REGFILE_SIM_reg_bank__abc_33898_n9203;
  wire REGFILE_SIM_reg_bank__abc_33898_n9204;
  wire REGFILE_SIM_reg_bank__abc_33898_n9205;
  wire REGFILE_SIM_reg_bank__abc_33898_n9206;
  wire REGFILE_SIM_reg_bank__abc_33898_n9207;
  wire REGFILE_SIM_reg_bank__abc_33898_n9208;
  wire REGFILE_SIM_reg_bank__abc_33898_n9209;
  wire REGFILE_SIM_reg_bank__abc_33898_n9210;
  wire REGFILE_SIM_reg_bank__abc_33898_n9211;
  wire REGFILE_SIM_reg_bank__abc_33898_n9212;
  wire REGFILE_SIM_reg_bank__abc_33898_n9213;
  wire REGFILE_SIM_reg_bank__abc_33898_n9214;
  wire REGFILE_SIM_reg_bank__abc_33898_n9215;
  wire REGFILE_SIM_reg_bank__abc_33898_n9216;
  wire REGFILE_SIM_reg_bank__abc_33898_n9217;
  wire REGFILE_SIM_reg_bank__abc_33898_n9218;
  wire REGFILE_SIM_reg_bank__abc_33898_n9219;
  wire REGFILE_SIM_reg_bank__abc_33898_n9220;
  wire REGFILE_SIM_reg_bank__abc_33898_n9221;
  wire REGFILE_SIM_reg_bank__abc_33898_n9222;
  wire REGFILE_SIM_reg_bank__abc_33898_n9223;
  wire REGFILE_SIM_reg_bank__abc_33898_n9224;
  wire REGFILE_SIM_reg_bank__abc_33898_n9225;
  wire REGFILE_SIM_reg_bank__abc_33898_n9226;
  wire REGFILE_SIM_reg_bank__abc_33898_n9227;
  wire REGFILE_SIM_reg_bank__abc_33898_n9228;
  wire REGFILE_SIM_reg_bank__abc_33898_n9229;
  wire REGFILE_SIM_reg_bank__abc_33898_n9230;
  wire REGFILE_SIM_reg_bank__abc_33898_n9231;
  wire REGFILE_SIM_reg_bank__abc_33898_n9232;
  wire REGFILE_SIM_reg_bank__abc_33898_n9233;
  wire REGFILE_SIM_reg_bank__abc_33898_n9234;
  wire REGFILE_SIM_reg_bank__abc_33898_n9235;
  wire REGFILE_SIM_reg_bank__abc_33898_n9236;
  wire REGFILE_SIM_reg_bank__abc_33898_n9237;
  wire REGFILE_SIM_reg_bank__abc_33898_n9238;
  wire REGFILE_SIM_reg_bank__abc_33898_n9239;
  wire REGFILE_SIM_reg_bank__abc_33898_n9240;
  wire REGFILE_SIM_reg_bank__abc_33898_n9241;
  wire REGFILE_SIM_reg_bank__abc_33898_n9242;
  wire REGFILE_SIM_reg_bank__abc_33898_n9243;
  wire REGFILE_SIM_reg_bank__abc_33898_n9244;
  wire REGFILE_SIM_reg_bank__abc_33898_n9245;
  wire REGFILE_SIM_reg_bank__abc_33898_n9246;
  wire REGFILE_SIM_reg_bank__abc_33898_n9247;
  wire REGFILE_SIM_reg_bank__abc_33898_n9248;
  wire REGFILE_SIM_reg_bank__abc_33898_n9249;
  wire REGFILE_SIM_reg_bank__abc_33898_n9250;
  wire REGFILE_SIM_reg_bank__abc_33898_n9252;
  wire REGFILE_SIM_reg_bank__abc_33898_n9253;
  wire REGFILE_SIM_reg_bank__abc_33898_n9254;
  wire REGFILE_SIM_reg_bank__abc_33898_n9255;
  wire REGFILE_SIM_reg_bank__abc_33898_n9256;
  wire REGFILE_SIM_reg_bank__abc_33898_n9257;
  wire REGFILE_SIM_reg_bank__abc_33898_n9258;
  wire REGFILE_SIM_reg_bank__abc_33898_n9259;
  wire REGFILE_SIM_reg_bank__abc_33898_n9260;
  wire REGFILE_SIM_reg_bank__abc_33898_n9261;
  wire REGFILE_SIM_reg_bank__abc_33898_n9262;
  wire REGFILE_SIM_reg_bank__abc_33898_n9263;
  wire REGFILE_SIM_reg_bank__abc_33898_n9264;
  wire REGFILE_SIM_reg_bank__abc_33898_n9265;
  wire REGFILE_SIM_reg_bank__abc_33898_n9266;
  wire REGFILE_SIM_reg_bank__abc_33898_n9267;
  wire REGFILE_SIM_reg_bank__abc_33898_n9268;
  wire REGFILE_SIM_reg_bank__abc_33898_n9269;
  wire REGFILE_SIM_reg_bank__abc_33898_n9270;
  wire REGFILE_SIM_reg_bank__abc_33898_n9271;
  wire REGFILE_SIM_reg_bank__abc_33898_n9272;
  wire REGFILE_SIM_reg_bank__abc_33898_n9273;
  wire REGFILE_SIM_reg_bank__abc_33898_n9274;
  wire REGFILE_SIM_reg_bank__abc_33898_n9275;
  wire REGFILE_SIM_reg_bank__abc_33898_n9276;
  wire REGFILE_SIM_reg_bank__abc_33898_n9277;
  wire REGFILE_SIM_reg_bank__abc_33898_n9278;
  wire REGFILE_SIM_reg_bank__abc_33898_n9279;
  wire REGFILE_SIM_reg_bank__abc_33898_n9280;
  wire REGFILE_SIM_reg_bank__abc_33898_n9281;
  wire REGFILE_SIM_reg_bank__abc_33898_n9282;
  wire REGFILE_SIM_reg_bank__abc_33898_n9283;
  wire REGFILE_SIM_reg_bank__abc_33898_n9284;
  wire REGFILE_SIM_reg_bank__abc_33898_n9285;
  wire REGFILE_SIM_reg_bank__abc_33898_n9286;
  wire REGFILE_SIM_reg_bank__abc_33898_n9287;
  wire REGFILE_SIM_reg_bank__abc_33898_n9288;
  wire REGFILE_SIM_reg_bank__abc_33898_n9289;
  wire REGFILE_SIM_reg_bank__abc_33898_n9290;
  wire REGFILE_SIM_reg_bank__abc_33898_n9291;
  wire REGFILE_SIM_reg_bank__abc_33898_n9292;
  wire REGFILE_SIM_reg_bank__abc_33898_n9293;
  wire REGFILE_SIM_reg_bank__abc_33898_n9294;
  wire REGFILE_SIM_reg_bank__abc_33898_n9295;
  wire REGFILE_SIM_reg_bank__abc_33898_n9296;
  wire REGFILE_SIM_reg_bank__abc_33898_n9297;
  wire REGFILE_SIM_reg_bank__abc_33898_n9298;
  wire REGFILE_SIM_reg_bank__abc_33898_n9299;
  wire REGFILE_SIM_reg_bank__abc_33898_n9300;
  wire REGFILE_SIM_reg_bank__abc_33898_n9301;
  wire REGFILE_SIM_reg_bank__abc_33898_n9302;
  wire REGFILE_SIM_reg_bank__abc_33898_n9303;
  wire REGFILE_SIM_reg_bank__abc_33898_n9304;
  wire REGFILE_SIM_reg_bank__abc_33898_n9305;
  wire REGFILE_SIM_reg_bank__abc_33898_n9306;
  wire REGFILE_SIM_reg_bank__abc_33898_n9307;
  wire REGFILE_SIM_reg_bank__abc_33898_n9308;
  wire REGFILE_SIM_reg_bank__abc_33898_n9309;
  wire REGFILE_SIM_reg_bank__abc_33898_n9310;
  wire REGFILE_SIM_reg_bank__abc_33898_n9311;
  wire REGFILE_SIM_reg_bank__abc_33898_n9313;
  wire REGFILE_SIM_reg_bank__abc_33898_n9314;
  wire REGFILE_SIM_reg_bank__abc_33898_n9315;
  wire REGFILE_SIM_reg_bank__abc_33898_n9316;
  wire REGFILE_SIM_reg_bank__abc_33898_n9317;
  wire REGFILE_SIM_reg_bank__abc_33898_n9318;
  wire REGFILE_SIM_reg_bank__abc_33898_n9319;
  wire REGFILE_SIM_reg_bank__abc_33898_n9320;
  wire REGFILE_SIM_reg_bank__abc_33898_n9321;
  wire REGFILE_SIM_reg_bank__abc_33898_n9322;
  wire REGFILE_SIM_reg_bank__abc_33898_n9323;
  wire REGFILE_SIM_reg_bank__abc_33898_n9324;
  wire REGFILE_SIM_reg_bank__abc_33898_n9325;
  wire REGFILE_SIM_reg_bank__abc_33898_n9326;
  wire REGFILE_SIM_reg_bank__abc_33898_n9327;
  wire REGFILE_SIM_reg_bank__abc_33898_n9328;
  wire REGFILE_SIM_reg_bank__abc_33898_n9329;
  wire REGFILE_SIM_reg_bank__abc_33898_n9330;
  wire REGFILE_SIM_reg_bank__abc_33898_n9331;
  wire REGFILE_SIM_reg_bank__abc_33898_n9332;
  wire REGFILE_SIM_reg_bank__abc_33898_n9333;
  wire REGFILE_SIM_reg_bank__abc_33898_n9334;
  wire REGFILE_SIM_reg_bank__abc_33898_n9335;
  wire REGFILE_SIM_reg_bank__abc_33898_n9336;
  wire REGFILE_SIM_reg_bank__abc_33898_n9337;
  wire REGFILE_SIM_reg_bank__abc_33898_n9338;
  wire REGFILE_SIM_reg_bank__abc_33898_n9339;
  wire REGFILE_SIM_reg_bank__abc_33898_n9340;
  wire REGFILE_SIM_reg_bank__abc_33898_n9341;
  wire REGFILE_SIM_reg_bank__abc_33898_n9342;
  wire REGFILE_SIM_reg_bank__abc_33898_n9343;
  wire REGFILE_SIM_reg_bank__abc_33898_n9344;
  wire REGFILE_SIM_reg_bank__abc_33898_n9345;
  wire REGFILE_SIM_reg_bank__abc_33898_n9346;
  wire REGFILE_SIM_reg_bank__abc_33898_n9347;
  wire REGFILE_SIM_reg_bank__abc_33898_n9348;
  wire REGFILE_SIM_reg_bank__abc_33898_n9349;
  wire REGFILE_SIM_reg_bank__abc_33898_n9350;
  wire REGFILE_SIM_reg_bank__abc_33898_n9351;
  wire REGFILE_SIM_reg_bank__abc_33898_n9352;
  wire REGFILE_SIM_reg_bank__abc_33898_n9353;
  wire REGFILE_SIM_reg_bank__abc_33898_n9354;
  wire REGFILE_SIM_reg_bank__abc_33898_n9355;
  wire REGFILE_SIM_reg_bank__abc_33898_n9356;
  wire REGFILE_SIM_reg_bank__abc_33898_n9357;
  wire REGFILE_SIM_reg_bank__abc_33898_n9358;
  wire REGFILE_SIM_reg_bank__abc_33898_n9359;
  wire REGFILE_SIM_reg_bank__abc_33898_n9360;
  wire REGFILE_SIM_reg_bank__abc_33898_n9361;
  wire REGFILE_SIM_reg_bank__abc_33898_n9362;
  wire REGFILE_SIM_reg_bank__abc_33898_n9363;
  wire REGFILE_SIM_reg_bank__abc_33898_n9364;
  wire REGFILE_SIM_reg_bank__abc_33898_n9365;
  wire REGFILE_SIM_reg_bank__abc_33898_n9366;
  wire REGFILE_SIM_reg_bank__abc_33898_n9367;
  wire REGFILE_SIM_reg_bank__abc_33898_n9368;
  wire REGFILE_SIM_reg_bank__abc_33898_n9369;
  wire REGFILE_SIM_reg_bank__abc_33898_n9370;
  wire REGFILE_SIM_reg_bank__abc_33898_n9371;
  wire REGFILE_SIM_reg_bank__abc_33898_n9372;
  wire REGFILE_SIM_reg_bank__abc_33898_n9374;
  wire REGFILE_SIM_reg_bank__abc_33898_n9375;
  wire REGFILE_SIM_reg_bank__abc_33898_n9376;
  wire REGFILE_SIM_reg_bank__abc_33898_n9377;
  wire REGFILE_SIM_reg_bank__abc_33898_n9378;
  wire REGFILE_SIM_reg_bank__abc_33898_n9379;
  wire REGFILE_SIM_reg_bank__abc_33898_n9380;
  wire REGFILE_SIM_reg_bank__abc_33898_n9381;
  wire REGFILE_SIM_reg_bank__abc_33898_n9382;
  wire REGFILE_SIM_reg_bank__abc_33898_n9383;
  wire REGFILE_SIM_reg_bank__abc_33898_n9384;
  wire REGFILE_SIM_reg_bank__abc_33898_n9385;
  wire REGFILE_SIM_reg_bank__abc_33898_n9386;
  wire REGFILE_SIM_reg_bank__abc_33898_n9387;
  wire REGFILE_SIM_reg_bank__abc_33898_n9388;
  wire REGFILE_SIM_reg_bank__abc_33898_n9389;
  wire REGFILE_SIM_reg_bank__abc_33898_n9390;
  wire REGFILE_SIM_reg_bank__abc_33898_n9391;
  wire REGFILE_SIM_reg_bank__abc_33898_n9392;
  wire REGFILE_SIM_reg_bank__abc_33898_n9393;
  wire REGFILE_SIM_reg_bank__abc_33898_n9394;
  wire REGFILE_SIM_reg_bank__abc_33898_n9395;
  wire REGFILE_SIM_reg_bank__abc_33898_n9396;
  wire REGFILE_SIM_reg_bank__abc_33898_n9397;
  wire REGFILE_SIM_reg_bank__abc_33898_n9398;
  wire REGFILE_SIM_reg_bank__abc_33898_n9399;
  wire REGFILE_SIM_reg_bank__abc_33898_n9400;
  wire REGFILE_SIM_reg_bank__abc_33898_n9401;
  wire REGFILE_SIM_reg_bank__abc_33898_n9402;
  wire REGFILE_SIM_reg_bank__abc_33898_n9403;
  wire REGFILE_SIM_reg_bank__abc_33898_n9404;
  wire REGFILE_SIM_reg_bank__abc_33898_n9405;
  wire REGFILE_SIM_reg_bank__abc_33898_n9406;
  wire REGFILE_SIM_reg_bank__abc_33898_n9407;
  wire REGFILE_SIM_reg_bank__abc_33898_n9408;
  wire REGFILE_SIM_reg_bank__abc_33898_n9409;
  wire REGFILE_SIM_reg_bank__abc_33898_n9410;
  wire REGFILE_SIM_reg_bank__abc_33898_n9411;
  wire REGFILE_SIM_reg_bank__abc_33898_n9412;
  wire REGFILE_SIM_reg_bank__abc_33898_n9413;
  wire REGFILE_SIM_reg_bank__abc_33898_n9414;
  wire REGFILE_SIM_reg_bank__abc_33898_n9415;
  wire REGFILE_SIM_reg_bank__abc_33898_n9416;
  wire REGFILE_SIM_reg_bank__abc_33898_n9417;
  wire REGFILE_SIM_reg_bank__abc_33898_n9418;
  wire REGFILE_SIM_reg_bank__abc_33898_n9419;
  wire REGFILE_SIM_reg_bank__abc_33898_n9420;
  wire REGFILE_SIM_reg_bank__abc_33898_n9421;
  wire REGFILE_SIM_reg_bank__abc_33898_n9422;
  wire REGFILE_SIM_reg_bank__abc_33898_n9423;
  wire REGFILE_SIM_reg_bank__abc_33898_n9424;
  wire REGFILE_SIM_reg_bank__abc_33898_n9425;
  wire REGFILE_SIM_reg_bank__abc_33898_n9426;
  wire REGFILE_SIM_reg_bank__abc_33898_n9427;
  wire REGFILE_SIM_reg_bank__abc_33898_n9428;
  wire REGFILE_SIM_reg_bank__abc_33898_n9429;
  wire REGFILE_SIM_reg_bank__abc_33898_n9430;
  wire REGFILE_SIM_reg_bank__abc_33898_n9431;
  wire REGFILE_SIM_reg_bank__abc_33898_n9432;
  wire REGFILE_SIM_reg_bank__abc_33898_n9433;
  wire REGFILE_SIM_reg_bank__abc_33898_n9435;
  wire REGFILE_SIM_reg_bank__abc_33898_n9436;
  wire REGFILE_SIM_reg_bank__abc_33898_n9437;
  wire REGFILE_SIM_reg_bank__abc_33898_n9438;
  wire REGFILE_SIM_reg_bank__abc_33898_n9439;
  wire REGFILE_SIM_reg_bank__abc_33898_n9440;
  wire REGFILE_SIM_reg_bank__abc_33898_n9441;
  wire REGFILE_SIM_reg_bank__abc_33898_n9442;
  wire REGFILE_SIM_reg_bank__abc_33898_n9443;
  wire REGFILE_SIM_reg_bank__abc_33898_n9444;
  wire REGFILE_SIM_reg_bank__abc_33898_n9445;
  wire REGFILE_SIM_reg_bank__abc_33898_n9446;
  wire REGFILE_SIM_reg_bank__abc_33898_n9447;
  wire REGFILE_SIM_reg_bank__abc_33898_n9448;
  wire REGFILE_SIM_reg_bank__abc_33898_n9449;
  wire REGFILE_SIM_reg_bank__abc_33898_n9450;
  wire REGFILE_SIM_reg_bank__abc_33898_n9451;
  wire REGFILE_SIM_reg_bank__abc_33898_n9452;
  wire REGFILE_SIM_reg_bank__abc_33898_n9453;
  wire REGFILE_SIM_reg_bank__abc_33898_n9454;
  wire REGFILE_SIM_reg_bank__abc_33898_n9455;
  wire REGFILE_SIM_reg_bank__abc_33898_n9456;
  wire REGFILE_SIM_reg_bank__abc_33898_n9457;
  wire REGFILE_SIM_reg_bank__abc_33898_n9458;
  wire REGFILE_SIM_reg_bank__abc_33898_n9459;
  wire REGFILE_SIM_reg_bank__abc_33898_n9460;
  wire REGFILE_SIM_reg_bank__abc_33898_n9461;
  wire REGFILE_SIM_reg_bank__abc_33898_n9462;
  wire REGFILE_SIM_reg_bank__abc_33898_n9463;
  wire REGFILE_SIM_reg_bank__abc_33898_n9464;
  wire REGFILE_SIM_reg_bank__abc_33898_n9465;
  wire REGFILE_SIM_reg_bank__abc_33898_n9466;
  wire REGFILE_SIM_reg_bank__abc_33898_n9467;
  wire REGFILE_SIM_reg_bank__abc_33898_n9468;
  wire REGFILE_SIM_reg_bank__abc_33898_n9469;
  wire REGFILE_SIM_reg_bank__abc_33898_n9470;
  wire REGFILE_SIM_reg_bank__abc_33898_n9471;
  wire REGFILE_SIM_reg_bank__abc_33898_n9472;
  wire REGFILE_SIM_reg_bank__abc_33898_n9473;
  wire REGFILE_SIM_reg_bank__abc_33898_n9474;
  wire REGFILE_SIM_reg_bank__abc_33898_n9475;
  wire REGFILE_SIM_reg_bank__abc_33898_n9476;
  wire REGFILE_SIM_reg_bank__abc_33898_n9477;
  wire REGFILE_SIM_reg_bank__abc_33898_n9478;
  wire REGFILE_SIM_reg_bank__abc_33898_n9479;
  wire REGFILE_SIM_reg_bank__abc_33898_n9480;
  wire REGFILE_SIM_reg_bank__abc_33898_n9481;
  wire REGFILE_SIM_reg_bank__abc_33898_n9482;
  wire REGFILE_SIM_reg_bank__abc_33898_n9483;
  wire REGFILE_SIM_reg_bank__abc_33898_n9484;
  wire REGFILE_SIM_reg_bank__abc_33898_n9485;
  wire REGFILE_SIM_reg_bank__abc_33898_n9486;
  wire REGFILE_SIM_reg_bank__abc_33898_n9487;
  wire REGFILE_SIM_reg_bank__abc_33898_n9488;
  wire REGFILE_SIM_reg_bank__abc_33898_n9489;
  wire REGFILE_SIM_reg_bank__abc_33898_n9490;
  wire REGFILE_SIM_reg_bank__abc_33898_n9491;
  wire REGFILE_SIM_reg_bank__abc_33898_n9492;
  wire REGFILE_SIM_reg_bank__abc_33898_n9493;
  wire REGFILE_SIM_reg_bank__abc_33898_n9494;
  wire REGFILE_SIM_reg_bank__abc_33898_n9496;
  wire REGFILE_SIM_reg_bank__abc_33898_n9497;
  wire REGFILE_SIM_reg_bank__abc_33898_n9498;
  wire REGFILE_SIM_reg_bank__abc_33898_n9499;
  wire REGFILE_SIM_reg_bank__abc_33898_n9500;
  wire REGFILE_SIM_reg_bank__abc_33898_n9501;
  wire REGFILE_SIM_reg_bank__abc_33898_n9502;
  wire REGFILE_SIM_reg_bank__abc_33898_n9503;
  wire REGFILE_SIM_reg_bank__abc_33898_n9504;
  wire REGFILE_SIM_reg_bank__abc_33898_n9505;
  wire REGFILE_SIM_reg_bank__abc_33898_n9506;
  wire REGFILE_SIM_reg_bank__abc_33898_n9507;
  wire REGFILE_SIM_reg_bank__abc_33898_n9508;
  wire REGFILE_SIM_reg_bank__abc_33898_n9509;
  wire REGFILE_SIM_reg_bank__abc_33898_n9510;
  wire REGFILE_SIM_reg_bank__abc_33898_n9511;
  wire REGFILE_SIM_reg_bank__abc_33898_n9512;
  wire REGFILE_SIM_reg_bank__abc_33898_n9513;
  wire REGFILE_SIM_reg_bank__abc_33898_n9514;
  wire REGFILE_SIM_reg_bank__abc_33898_n9515;
  wire REGFILE_SIM_reg_bank__abc_33898_n9516;
  wire REGFILE_SIM_reg_bank__abc_33898_n9517;
  wire REGFILE_SIM_reg_bank__abc_33898_n9518;
  wire REGFILE_SIM_reg_bank__abc_33898_n9519;
  wire REGFILE_SIM_reg_bank__abc_33898_n9520;
  wire REGFILE_SIM_reg_bank__abc_33898_n9521;
  wire REGFILE_SIM_reg_bank__abc_33898_n9522;
  wire REGFILE_SIM_reg_bank__abc_33898_n9523;
  wire REGFILE_SIM_reg_bank__abc_33898_n9524;
  wire REGFILE_SIM_reg_bank__abc_33898_n9525;
  wire REGFILE_SIM_reg_bank__abc_33898_n9526;
  wire REGFILE_SIM_reg_bank__abc_33898_n9527;
  wire REGFILE_SIM_reg_bank__abc_33898_n9528;
  wire REGFILE_SIM_reg_bank__abc_33898_n9529;
  wire REGFILE_SIM_reg_bank__abc_33898_n9530;
  wire REGFILE_SIM_reg_bank__abc_33898_n9531;
  wire REGFILE_SIM_reg_bank__abc_33898_n9532;
  wire REGFILE_SIM_reg_bank__abc_33898_n9533;
  wire REGFILE_SIM_reg_bank__abc_33898_n9534;
  wire REGFILE_SIM_reg_bank__abc_33898_n9535;
  wire REGFILE_SIM_reg_bank__abc_33898_n9536;
  wire REGFILE_SIM_reg_bank__abc_33898_n9537;
  wire REGFILE_SIM_reg_bank__abc_33898_n9538;
  wire REGFILE_SIM_reg_bank__abc_33898_n9539;
  wire REGFILE_SIM_reg_bank__abc_33898_n9540;
  wire REGFILE_SIM_reg_bank__abc_33898_n9541;
  wire REGFILE_SIM_reg_bank__abc_33898_n9542;
  wire REGFILE_SIM_reg_bank__abc_33898_n9543;
  wire REGFILE_SIM_reg_bank__abc_33898_n9544;
  wire REGFILE_SIM_reg_bank__abc_33898_n9545;
  wire REGFILE_SIM_reg_bank__abc_33898_n9546;
  wire REGFILE_SIM_reg_bank__abc_33898_n9547;
  wire REGFILE_SIM_reg_bank__abc_33898_n9548;
  wire REGFILE_SIM_reg_bank__abc_33898_n9549;
  wire REGFILE_SIM_reg_bank__abc_33898_n9550;
  wire REGFILE_SIM_reg_bank__abc_33898_n9551;
  wire REGFILE_SIM_reg_bank__abc_33898_n9552;
  wire REGFILE_SIM_reg_bank__abc_33898_n9553;
  wire REGFILE_SIM_reg_bank__abc_33898_n9554;
  wire REGFILE_SIM_reg_bank__abc_33898_n9555;
  wire REGFILE_SIM_reg_bank_ra_i_0_;
  wire REGFILE_SIM_reg_bank_ra_i_1_;
  wire REGFILE_SIM_reg_bank_ra_i_2_;
  wire REGFILE_SIM_reg_bank_ra_i_3_;
  wire REGFILE_SIM_reg_bank_ra_i_4_;
  wire REGFILE_SIM_reg_bank_rb_i_0_;
  wire REGFILE_SIM_reg_bank_rb_i_1_;
  wire REGFILE_SIM_reg_bank_rb_i_2_;
  wire REGFILE_SIM_reg_bank_rb_i_3_;
  wire REGFILE_SIM_reg_bank_rb_i_4_;
  wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf0;
  wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf1;
  wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf2;
  wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf3;
  wire REGFILE_SIM_reg_bank_rd_i_0_;
  wire REGFILE_SIM_reg_bank_rd_i_1_;
  wire REGFILE_SIM_reg_bank_rd_i_2_;
  wire REGFILE_SIM_reg_bank_rd_i_3_;
  wire REGFILE_SIM_reg_bank_rd_i_4_;
  wire REGFILE_SIM_reg_bank_reg_r10_0_;
  wire REGFILE_SIM_reg_bank_reg_r10_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_10_;
  wire REGFILE_SIM_reg_bank_reg_r10_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_11_;
  wire REGFILE_SIM_reg_bank_reg_r10_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_12_;
  wire REGFILE_SIM_reg_bank_reg_r10_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_13_;
  wire REGFILE_SIM_reg_bank_reg_r10_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_14_;
  wire REGFILE_SIM_reg_bank_reg_r10_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_15_;
  wire REGFILE_SIM_reg_bank_reg_r10_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_16_;
  wire REGFILE_SIM_reg_bank_reg_r10_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_17_;
  wire REGFILE_SIM_reg_bank_reg_r10_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_18_;
  wire REGFILE_SIM_reg_bank_reg_r10_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_19_;
  wire REGFILE_SIM_reg_bank_reg_r10_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_1_;
  wire REGFILE_SIM_reg_bank_reg_r10_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_20_;
  wire REGFILE_SIM_reg_bank_reg_r10_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_21_;
  wire REGFILE_SIM_reg_bank_reg_r10_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_22_;
  wire REGFILE_SIM_reg_bank_reg_r10_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_23_;
  wire REGFILE_SIM_reg_bank_reg_r10_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_24_;
  wire REGFILE_SIM_reg_bank_reg_r10_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_25_;
  wire REGFILE_SIM_reg_bank_reg_r10_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_26_;
  wire REGFILE_SIM_reg_bank_reg_r10_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_27_;
  wire REGFILE_SIM_reg_bank_reg_r10_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_28_;
  wire REGFILE_SIM_reg_bank_reg_r10_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_29_;
  wire REGFILE_SIM_reg_bank_reg_r10_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_2_;
  wire REGFILE_SIM_reg_bank_reg_r10_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_30_;
  wire REGFILE_SIM_reg_bank_reg_r10_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_31_;
  wire REGFILE_SIM_reg_bank_reg_r10_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_3_;
  wire REGFILE_SIM_reg_bank_reg_r10_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_4_;
  wire REGFILE_SIM_reg_bank_reg_r10_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_5_;
  wire REGFILE_SIM_reg_bank_reg_r10_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_6_;
  wire REGFILE_SIM_reg_bank_reg_r10_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_7_;
  wire REGFILE_SIM_reg_bank_reg_r10_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_8_;
  wire REGFILE_SIM_reg_bank_reg_r10_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r10_9_;
  wire REGFILE_SIM_reg_bank_reg_r10_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_0_;
  wire REGFILE_SIM_reg_bank_reg_r11_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_10_;
  wire REGFILE_SIM_reg_bank_reg_r11_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_11_;
  wire REGFILE_SIM_reg_bank_reg_r11_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_12_;
  wire REGFILE_SIM_reg_bank_reg_r11_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_13_;
  wire REGFILE_SIM_reg_bank_reg_r11_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_14_;
  wire REGFILE_SIM_reg_bank_reg_r11_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_15_;
  wire REGFILE_SIM_reg_bank_reg_r11_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_16_;
  wire REGFILE_SIM_reg_bank_reg_r11_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_17_;
  wire REGFILE_SIM_reg_bank_reg_r11_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_18_;
  wire REGFILE_SIM_reg_bank_reg_r11_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_19_;
  wire REGFILE_SIM_reg_bank_reg_r11_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_1_;
  wire REGFILE_SIM_reg_bank_reg_r11_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_20_;
  wire REGFILE_SIM_reg_bank_reg_r11_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_21_;
  wire REGFILE_SIM_reg_bank_reg_r11_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_22_;
  wire REGFILE_SIM_reg_bank_reg_r11_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_23_;
  wire REGFILE_SIM_reg_bank_reg_r11_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_24_;
  wire REGFILE_SIM_reg_bank_reg_r11_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_25_;
  wire REGFILE_SIM_reg_bank_reg_r11_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_26_;
  wire REGFILE_SIM_reg_bank_reg_r11_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_27_;
  wire REGFILE_SIM_reg_bank_reg_r11_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_28_;
  wire REGFILE_SIM_reg_bank_reg_r11_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_29_;
  wire REGFILE_SIM_reg_bank_reg_r11_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_2_;
  wire REGFILE_SIM_reg_bank_reg_r11_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_30_;
  wire REGFILE_SIM_reg_bank_reg_r11_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_31_;
  wire REGFILE_SIM_reg_bank_reg_r11_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_3_;
  wire REGFILE_SIM_reg_bank_reg_r11_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_4_;
  wire REGFILE_SIM_reg_bank_reg_r11_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_5_;
  wire REGFILE_SIM_reg_bank_reg_r11_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_6_;
  wire REGFILE_SIM_reg_bank_reg_r11_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_7_;
  wire REGFILE_SIM_reg_bank_reg_r11_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_8_;
  wire REGFILE_SIM_reg_bank_reg_r11_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r11_9_;
  wire REGFILE_SIM_reg_bank_reg_r11_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_0_;
  wire REGFILE_SIM_reg_bank_reg_r12_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_10_;
  wire REGFILE_SIM_reg_bank_reg_r12_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_11_;
  wire REGFILE_SIM_reg_bank_reg_r12_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_12_;
  wire REGFILE_SIM_reg_bank_reg_r12_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_13_;
  wire REGFILE_SIM_reg_bank_reg_r12_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_14_;
  wire REGFILE_SIM_reg_bank_reg_r12_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_15_;
  wire REGFILE_SIM_reg_bank_reg_r12_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_16_;
  wire REGFILE_SIM_reg_bank_reg_r12_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_17_;
  wire REGFILE_SIM_reg_bank_reg_r12_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_18_;
  wire REGFILE_SIM_reg_bank_reg_r12_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_19_;
  wire REGFILE_SIM_reg_bank_reg_r12_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_1_;
  wire REGFILE_SIM_reg_bank_reg_r12_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_20_;
  wire REGFILE_SIM_reg_bank_reg_r12_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_21_;
  wire REGFILE_SIM_reg_bank_reg_r12_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_22_;
  wire REGFILE_SIM_reg_bank_reg_r12_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_23_;
  wire REGFILE_SIM_reg_bank_reg_r12_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_24_;
  wire REGFILE_SIM_reg_bank_reg_r12_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_25_;
  wire REGFILE_SIM_reg_bank_reg_r12_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_26_;
  wire REGFILE_SIM_reg_bank_reg_r12_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_27_;
  wire REGFILE_SIM_reg_bank_reg_r12_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_28_;
  wire REGFILE_SIM_reg_bank_reg_r12_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_29_;
  wire REGFILE_SIM_reg_bank_reg_r12_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_2_;
  wire REGFILE_SIM_reg_bank_reg_r12_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_30_;
  wire REGFILE_SIM_reg_bank_reg_r12_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_31_;
  wire REGFILE_SIM_reg_bank_reg_r12_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_3_;
  wire REGFILE_SIM_reg_bank_reg_r12_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_4_;
  wire REGFILE_SIM_reg_bank_reg_r12_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_5_;
  wire REGFILE_SIM_reg_bank_reg_r12_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_6_;
  wire REGFILE_SIM_reg_bank_reg_r12_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_7_;
  wire REGFILE_SIM_reg_bank_reg_r12_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_8_;
  wire REGFILE_SIM_reg_bank_reg_r12_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r12_9_;
  wire REGFILE_SIM_reg_bank_reg_r12_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_0_;
  wire REGFILE_SIM_reg_bank_reg_r13_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_10_;
  wire REGFILE_SIM_reg_bank_reg_r13_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_11_;
  wire REGFILE_SIM_reg_bank_reg_r13_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_12_;
  wire REGFILE_SIM_reg_bank_reg_r13_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_13_;
  wire REGFILE_SIM_reg_bank_reg_r13_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_14_;
  wire REGFILE_SIM_reg_bank_reg_r13_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_15_;
  wire REGFILE_SIM_reg_bank_reg_r13_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_16_;
  wire REGFILE_SIM_reg_bank_reg_r13_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_17_;
  wire REGFILE_SIM_reg_bank_reg_r13_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_18_;
  wire REGFILE_SIM_reg_bank_reg_r13_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_19_;
  wire REGFILE_SIM_reg_bank_reg_r13_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_1_;
  wire REGFILE_SIM_reg_bank_reg_r13_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_20_;
  wire REGFILE_SIM_reg_bank_reg_r13_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_21_;
  wire REGFILE_SIM_reg_bank_reg_r13_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_22_;
  wire REGFILE_SIM_reg_bank_reg_r13_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_23_;
  wire REGFILE_SIM_reg_bank_reg_r13_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_24_;
  wire REGFILE_SIM_reg_bank_reg_r13_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_25_;
  wire REGFILE_SIM_reg_bank_reg_r13_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_26_;
  wire REGFILE_SIM_reg_bank_reg_r13_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_27_;
  wire REGFILE_SIM_reg_bank_reg_r13_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_28_;
  wire REGFILE_SIM_reg_bank_reg_r13_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_29_;
  wire REGFILE_SIM_reg_bank_reg_r13_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_2_;
  wire REGFILE_SIM_reg_bank_reg_r13_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_30_;
  wire REGFILE_SIM_reg_bank_reg_r13_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_31_;
  wire REGFILE_SIM_reg_bank_reg_r13_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_3_;
  wire REGFILE_SIM_reg_bank_reg_r13_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_4_;
  wire REGFILE_SIM_reg_bank_reg_r13_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_5_;
  wire REGFILE_SIM_reg_bank_reg_r13_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_6_;
  wire REGFILE_SIM_reg_bank_reg_r13_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_7_;
  wire REGFILE_SIM_reg_bank_reg_r13_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_8_;
  wire REGFILE_SIM_reg_bank_reg_r13_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r13_9_;
  wire REGFILE_SIM_reg_bank_reg_r13_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_0_;
  wire REGFILE_SIM_reg_bank_reg_r14_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_10_;
  wire REGFILE_SIM_reg_bank_reg_r14_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_11_;
  wire REGFILE_SIM_reg_bank_reg_r14_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_12_;
  wire REGFILE_SIM_reg_bank_reg_r14_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_13_;
  wire REGFILE_SIM_reg_bank_reg_r14_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_14_;
  wire REGFILE_SIM_reg_bank_reg_r14_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_15_;
  wire REGFILE_SIM_reg_bank_reg_r14_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_16_;
  wire REGFILE_SIM_reg_bank_reg_r14_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_17_;
  wire REGFILE_SIM_reg_bank_reg_r14_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_18_;
  wire REGFILE_SIM_reg_bank_reg_r14_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_19_;
  wire REGFILE_SIM_reg_bank_reg_r14_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_1_;
  wire REGFILE_SIM_reg_bank_reg_r14_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_20_;
  wire REGFILE_SIM_reg_bank_reg_r14_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_21_;
  wire REGFILE_SIM_reg_bank_reg_r14_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_22_;
  wire REGFILE_SIM_reg_bank_reg_r14_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_23_;
  wire REGFILE_SIM_reg_bank_reg_r14_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_24_;
  wire REGFILE_SIM_reg_bank_reg_r14_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_25_;
  wire REGFILE_SIM_reg_bank_reg_r14_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_26_;
  wire REGFILE_SIM_reg_bank_reg_r14_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_27_;
  wire REGFILE_SIM_reg_bank_reg_r14_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_28_;
  wire REGFILE_SIM_reg_bank_reg_r14_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_29_;
  wire REGFILE_SIM_reg_bank_reg_r14_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_2_;
  wire REGFILE_SIM_reg_bank_reg_r14_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_30_;
  wire REGFILE_SIM_reg_bank_reg_r14_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_31_;
  wire REGFILE_SIM_reg_bank_reg_r14_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_3_;
  wire REGFILE_SIM_reg_bank_reg_r14_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_4_;
  wire REGFILE_SIM_reg_bank_reg_r14_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_5_;
  wire REGFILE_SIM_reg_bank_reg_r14_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_6_;
  wire REGFILE_SIM_reg_bank_reg_r14_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_7_;
  wire REGFILE_SIM_reg_bank_reg_r14_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_8_;
  wire REGFILE_SIM_reg_bank_reg_r14_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r14_9_;
  wire REGFILE_SIM_reg_bank_reg_r14_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_0_;
  wire REGFILE_SIM_reg_bank_reg_r15_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_10_;
  wire REGFILE_SIM_reg_bank_reg_r15_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_11_;
  wire REGFILE_SIM_reg_bank_reg_r15_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_12_;
  wire REGFILE_SIM_reg_bank_reg_r15_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_13_;
  wire REGFILE_SIM_reg_bank_reg_r15_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_14_;
  wire REGFILE_SIM_reg_bank_reg_r15_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_15_;
  wire REGFILE_SIM_reg_bank_reg_r15_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_16_;
  wire REGFILE_SIM_reg_bank_reg_r15_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_17_;
  wire REGFILE_SIM_reg_bank_reg_r15_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_18_;
  wire REGFILE_SIM_reg_bank_reg_r15_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_19_;
  wire REGFILE_SIM_reg_bank_reg_r15_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_1_;
  wire REGFILE_SIM_reg_bank_reg_r15_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_20_;
  wire REGFILE_SIM_reg_bank_reg_r15_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_21_;
  wire REGFILE_SIM_reg_bank_reg_r15_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_22_;
  wire REGFILE_SIM_reg_bank_reg_r15_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_23_;
  wire REGFILE_SIM_reg_bank_reg_r15_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_24_;
  wire REGFILE_SIM_reg_bank_reg_r15_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_25_;
  wire REGFILE_SIM_reg_bank_reg_r15_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_26_;
  wire REGFILE_SIM_reg_bank_reg_r15_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_27_;
  wire REGFILE_SIM_reg_bank_reg_r15_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_28_;
  wire REGFILE_SIM_reg_bank_reg_r15_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_29_;
  wire REGFILE_SIM_reg_bank_reg_r15_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_2_;
  wire REGFILE_SIM_reg_bank_reg_r15_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_30_;
  wire REGFILE_SIM_reg_bank_reg_r15_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_31_;
  wire REGFILE_SIM_reg_bank_reg_r15_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_3_;
  wire REGFILE_SIM_reg_bank_reg_r15_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_4_;
  wire REGFILE_SIM_reg_bank_reg_r15_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_5_;
  wire REGFILE_SIM_reg_bank_reg_r15_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_6_;
  wire REGFILE_SIM_reg_bank_reg_r15_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_7_;
  wire REGFILE_SIM_reg_bank_reg_r15_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_8_;
  wire REGFILE_SIM_reg_bank_reg_r15_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r15_9_;
  wire REGFILE_SIM_reg_bank_reg_r15_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_0_;
  wire REGFILE_SIM_reg_bank_reg_r16_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_10_;
  wire REGFILE_SIM_reg_bank_reg_r16_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_11_;
  wire REGFILE_SIM_reg_bank_reg_r16_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_12_;
  wire REGFILE_SIM_reg_bank_reg_r16_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_13_;
  wire REGFILE_SIM_reg_bank_reg_r16_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_14_;
  wire REGFILE_SIM_reg_bank_reg_r16_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_15_;
  wire REGFILE_SIM_reg_bank_reg_r16_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_16_;
  wire REGFILE_SIM_reg_bank_reg_r16_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_17_;
  wire REGFILE_SIM_reg_bank_reg_r16_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_18_;
  wire REGFILE_SIM_reg_bank_reg_r16_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_19_;
  wire REGFILE_SIM_reg_bank_reg_r16_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_1_;
  wire REGFILE_SIM_reg_bank_reg_r16_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_20_;
  wire REGFILE_SIM_reg_bank_reg_r16_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_21_;
  wire REGFILE_SIM_reg_bank_reg_r16_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_22_;
  wire REGFILE_SIM_reg_bank_reg_r16_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_23_;
  wire REGFILE_SIM_reg_bank_reg_r16_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_24_;
  wire REGFILE_SIM_reg_bank_reg_r16_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_25_;
  wire REGFILE_SIM_reg_bank_reg_r16_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_26_;
  wire REGFILE_SIM_reg_bank_reg_r16_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_27_;
  wire REGFILE_SIM_reg_bank_reg_r16_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_28_;
  wire REGFILE_SIM_reg_bank_reg_r16_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_29_;
  wire REGFILE_SIM_reg_bank_reg_r16_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_2_;
  wire REGFILE_SIM_reg_bank_reg_r16_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_30_;
  wire REGFILE_SIM_reg_bank_reg_r16_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_31_;
  wire REGFILE_SIM_reg_bank_reg_r16_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_3_;
  wire REGFILE_SIM_reg_bank_reg_r16_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_4_;
  wire REGFILE_SIM_reg_bank_reg_r16_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_5_;
  wire REGFILE_SIM_reg_bank_reg_r16_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_6_;
  wire REGFILE_SIM_reg_bank_reg_r16_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_7_;
  wire REGFILE_SIM_reg_bank_reg_r16_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_8_;
  wire REGFILE_SIM_reg_bank_reg_r16_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r16_9_;
  wire REGFILE_SIM_reg_bank_reg_r16_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_0_;
  wire REGFILE_SIM_reg_bank_reg_r17_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_10_;
  wire REGFILE_SIM_reg_bank_reg_r17_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_11_;
  wire REGFILE_SIM_reg_bank_reg_r17_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_12_;
  wire REGFILE_SIM_reg_bank_reg_r17_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_13_;
  wire REGFILE_SIM_reg_bank_reg_r17_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_14_;
  wire REGFILE_SIM_reg_bank_reg_r17_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_15_;
  wire REGFILE_SIM_reg_bank_reg_r17_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_16_;
  wire REGFILE_SIM_reg_bank_reg_r17_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_17_;
  wire REGFILE_SIM_reg_bank_reg_r17_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_18_;
  wire REGFILE_SIM_reg_bank_reg_r17_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_19_;
  wire REGFILE_SIM_reg_bank_reg_r17_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_1_;
  wire REGFILE_SIM_reg_bank_reg_r17_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_20_;
  wire REGFILE_SIM_reg_bank_reg_r17_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_21_;
  wire REGFILE_SIM_reg_bank_reg_r17_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_22_;
  wire REGFILE_SIM_reg_bank_reg_r17_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_23_;
  wire REGFILE_SIM_reg_bank_reg_r17_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_24_;
  wire REGFILE_SIM_reg_bank_reg_r17_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_25_;
  wire REGFILE_SIM_reg_bank_reg_r17_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_26_;
  wire REGFILE_SIM_reg_bank_reg_r17_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_27_;
  wire REGFILE_SIM_reg_bank_reg_r17_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_28_;
  wire REGFILE_SIM_reg_bank_reg_r17_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_29_;
  wire REGFILE_SIM_reg_bank_reg_r17_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_2_;
  wire REGFILE_SIM_reg_bank_reg_r17_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_30_;
  wire REGFILE_SIM_reg_bank_reg_r17_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_31_;
  wire REGFILE_SIM_reg_bank_reg_r17_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_3_;
  wire REGFILE_SIM_reg_bank_reg_r17_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_4_;
  wire REGFILE_SIM_reg_bank_reg_r17_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_5_;
  wire REGFILE_SIM_reg_bank_reg_r17_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_6_;
  wire REGFILE_SIM_reg_bank_reg_r17_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_7_;
  wire REGFILE_SIM_reg_bank_reg_r17_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_8_;
  wire REGFILE_SIM_reg_bank_reg_r17_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r17_9_;
  wire REGFILE_SIM_reg_bank_reg_r17_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_0_;
  wire REGFILE_SIM_reg_bank_reg_r18_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_10_;
  wire REGFILE_SIM_reg_bank_reg_r18_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_11_;
  wire REGFILE_SIM_reg_bank_reg_r18_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_12_;
  wire REGFILE_SIM_reg_bank_reg_r18_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_13_;
  wire REGFILE_SIM_reg_bank_reg_r18_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_14_;
  wire REGFILE_SIM_reg_bank_reg_r18_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_15_;
  wire REGFILE_SIM_reg_bank_reg_r18_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_16_;
  wire REGFILE_SIM_reg_bank_reg_r18_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_17_;
  wire REGFILE_SIM_reg_bank_reg_r18_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_18_;
  wire REGFILE_SIM_reg_bank_reg_r18_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_19_;
  wire REGFILE_SIM_reg_bank_reg_r18_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_1_;
  wire REGFILE_SIM_reg_bank_reg_r18_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_20_;
  wire REGFILE_SIM_reg_bank_reg_r18_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_21_;
  wire REGFILE_SIM_reg_bank_reg_r18_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_22_;
  wire REGFILE_SIM_reg_bank_reg_r18_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_23_;
  wire REGFILE_SIM_reg_bank_reg_r18_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_24_;
  wire REGFILE_SIM_reg_bank_reg_r18_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_25_;
  wire REGFILE_SIM_reg_bank_reg_r18_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_26_;
  wire REGFILE_SIM_reg_bank_reg_r18_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_27_;
  wire REGFILE_SIM_reg_bank_reg_r18_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_28_;
  wire REGFILE_SIM_reg_bank_reg_r18_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_29_;
  wire REGFILE_SIM_reg_bank_reg_r18_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_2_;
  wire REGFILE_SIM_reg_bank_reg_r18_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_30_;
  wire REGFILE_SIM_reg_bank_reg_r18_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_31_;
  wire REGFILE_SIM_reg_bank_reg_r18_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_3_;
  wire REGFILE_SIM_reg_bank_reg_r18_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_4_;
  wire REGFILE_SIM_reg_bank_reg_r18_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_5_;
  wire REGFILE_SIM_reg_bank_reg_r18_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_6_;
  wire REGFILE_SIM_reg_bank_reg_r18_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_7_;
  wire REGFILE_SIM_reg_bank_reg_r18_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_8_;
  wire REGFILE_SIM_reg_bank_reg_r18_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r18_9_;
  wire REGFILE_SIM_reg_bank_reg_r18_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_0_;
  wire REGFILE_SIM_reg_bank_reg_r19_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_10_;
  wire REGFILE_SIM_reg_bank_reg_r19_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_11_;
  wire REGFILE_SIM_reg_bank_reg_r19_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_12_;
  wire REGFILE_SIM_reg_bank_reg_r19_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_13_;
  wire REGFILE_SIM_reg_bank_reg_r19_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_14_;
  wire REGFILE_SIM_reg_bank_reg_r19_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_15_;
  wire REGFILE_SIM_reg_bank_reg_r19_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_16_;
  wire REGFILE_SIM_reg_bank_reg_r19_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_17_;
  wire REGFILE_SIM_reg_bank_reg_r19_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_18_;
  wire REGFILE_SIM_reg_bank_reg_r19_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_19_;
  wire REGFILE_SIM_reg_bank_reg_r19_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_1_;
  wire REGFILE_SIM_reg_bank_reg_r19_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_20_;
  wire REGFILE_SIM_reg_bank_reg_r19_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_21_;
  wire REGFILE_SIM_reg_bank_reg_r19_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_22_;
  wire REGFILE_SIM_reg_bank_reg_r19_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_23_;
  wire REGFILE_SIM_reg_bank_reg_r19_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_24_;
  wire REGFILE_SIM_reg_bank_reg_r19_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_25_;
  wire REGFILE_SIM_reg_bank_reg_r19_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_26_;
  wire REGFILE_SIM_reg_bank_reg_r19_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_27_;
  wire REGFILE_SIM_reg_bank_reg_r19_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_28_;
  wire REGFILE_SIM_reg_bank_reg_r19_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_29_;
  wire REGFILE_SIM_reg_bank_reg_r19_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_2_;
  wire REGFILE_SIM_reg_bank_reg_r19_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_30_;
  wire REGFILE_SIM_reg_bank_reg_r19_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_31_;
  wire REGFILE_SIM_reg_bank_reg_r19_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_3_;
  wire REGFILE_SIM_reg_bank_reg_r19_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_4_;
  wire REGFILE_SIM_reg_bank_reg_r19_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_5_;
  wire REGFILE_SIM_reg_bank_reg_r19_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_6_;
  wire REGFILE_SIM_reg_bank_reg_r19_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_7_;
  wire REGFILE_SIM_reg_bank_reg_r19_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_8_;
  wire REGFILE_SIM_reg_bank_reg_r19_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r19_9_;
  wire REGFILE_SIM_reg_bank_reg_r19_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_0_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_10_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_11_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_12_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_13_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_14_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_15_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_16_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_17_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_18_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_19_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_1_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_20_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_21_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_22_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_23_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_24_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_25_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_26_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_27_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_28_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_29_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_2_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_30_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_31_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_3_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_4_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_5_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_6_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_7_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_8_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_9_;
  wire REGFILE_SIM_reg_bank_reg_r1_sp_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_0_;
  wire REGFILE_SIM_reg_bank_reg_r20_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_10_;
  wire REGFILE_SIM_reg_bank_reg_r20_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_11_;
  wire REGFILE_SIM_reg_bank_reg_r20_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_12_;
  wire REGFILE_SIM_reg_bank_reg_r20_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_13_;
  wire REGFILE_SIM_reg_bank_reg_r20_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_14_;
  wire REGFILE_SIM_reg_bank_reg_r20_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_15_;
  wire REGFILE_SIM_reg_bank_reg_r20_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_16_;
  wire REGFILE_SIM_reg_bank_reg_r20_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_17_;
  wire REGFILE_SIM_reg_bank_reg_r20_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_18_;
  wire REGFILE_SIM_reg_bank_reg_r20_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_19_;
  wire REGFILE_SIM_reg_bank_reg_r20_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_1_;
  wire REGFILE_SIM_reg_bank_reg_r20_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_20_;
  wire REGFILE_SIM_reg_bank_reg_r20_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_21_;
  wire REGFILE_SIM_reg_bank_reg_r20_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_22_;
  wire REGFILE_SIM_reg_bank_reg_r20_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_23_;
  wire REGFILE_SIM_reg_bank_reg_r20_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_24_;
  wire REGFILE_SIM_reg_bank_reg_r20_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_25_;
  wire REGFILE_SIM_reg_bank_reg_r20_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_26_;
  wire REGFILE_SIM_reg_bank_reg_r20_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_27_;
  wire REGFILE_SIM_reg_bank_reg_r20_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_28_;
  wire REGFILE_SIM_reg_bank_reg_r20_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_29_;
  wire REGFILE_SIM_reg_bank_reg_r20_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_2_;
  wire REGFILE_SIM_reg_bank_reg_r20_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_30_;
  wire REGFILE_SIM_reg_bank_reg_r20_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_31_;
  wire REGFILE_SIM_reg_bank_reg_r20_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_3_;
  wire REGFILE_SIM_reg_bank_reg_r20_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_4_;
  wire REGFILE_SIM_reg_bank_reg_r20_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_5_;
  wire REGFILE_SIM_reg_bank_reg_r20_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_6_;
  wire REGFILE_SIM_reg_bank_reg_r20_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_7_;
  wire REGFILE_SIM_reg_bank_reg_r20_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_8_;
  wire REGFILE_SIM_reg_bank_reg_r20_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r20_9_;
  wire REGFILE_SIM_reg_bank_reg_r20_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_0_;
  wire REGFILE_SIM_reg_bank_reg_r21_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_10_;
  wire REGFILE_SIM_reg_bank_reg_r21_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_11_;
  wire REGFILE_SIM_reg_bank_reg_r21_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_12_;
  wire REGFILE_SIM_reg_bank_reg_r21_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_13_;
  wire REGFILE_SIM_reg_bank_reg_r21_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_14_;
  wire REGFILE_SIM_reg_bank_reg_r21_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_15_;
  wire REGFILE_SIM_reg_bank_reg_r21_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_16_;
  wire REGFILE_SIM_reg_bank_reg_r21_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_17_;
  wire REGFILE_SIM_reg_bank_reg_r21_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_18_;
  wire REGFILE_SIM_reg_bank_reg_r21_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_19_;
  wire REGFILE_SIM_reg_bank_reg_r21_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_1_;
  wire REGFILE_SIM_reg_bank_reg_r21_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_20_;
  wire REGFILE_SIM_reg_bank_reg_r21_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_21_;
  wire REGFILE_SIM_reg_bank_reg_r21_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_22_;
  wire REGFILE_SIM_reg_bank_reg_r21_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_23_;
  wire REGFILE_SIM_reg_bank_reg_r21_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_24_;
  wire REGFILE_SIM_reg_bank_reg_r21_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_25_;
  wire REGFILE_SIM_reg_bank_reg_r21_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_26_;
  wire REGFILE_SIM_reg_bank_reg_r21_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_27_;
  wire REGFILE_SIM_reg_bank_reg_r21_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_28_;
  wire REGFILE_SIM_reg_bank_reg_r21_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_29_;
  wire REGFILE_SIM_reg_bank_reg_r21_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_2_;
  wire REGFILE_SIM_reg_bank_reg_r21_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_30_;
  wire REGFILE_SIM_reg_bank_reg_r21_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_31_;
  wire REGFILE_SIM_reg_bank_reg_r21_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_3_;
  wire REGFILE_SIM_reg_bank_reg_r21_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_4_;
  wire REGFILE_SIM_reg_bank_reg_r21_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_5_;
  wire REGFILE_SIM_reg_bank_reg_r21_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_6_;
  wire REGFILE_SIM_reg_bank_reg_r21_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_7_;
  wire REGFILE_SIM_reg_bank_reg_r21_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_8_;
  wire REGFILE_SIM_reg_bank_reg_r21_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r21_9_;
  wire REGFILE_SIM_reg_bank_reg_r21_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_0_;
  wire REGFILE_SIM_reg_bank_reg_r22_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_10_;
  wire REGFILE_SIM_reg_bank_reg_r22_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_11_;
  wire REGFILE_SIM_reg_bank_reg_r22_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_12_;
  wire REGFILE_SIM_reg_bank_reg_r22_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_13_;
  wire REGFILE_SIM_reg_bank_reg_r22_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_14_;
  wire REGFILE_SIM_reg_bank_reg_r22_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_15_;
  wire REGFILE_SIM_reg_bank_reg_r22_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_16_;
  wire REGFILE_SIM_reg_bank_reg_r22_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_17_;
  wire REGFILE_SIM_reg_bank_reg_r22_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_18_;
  wire REGFILE_SIM_reg_bank_reg_r22_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_19_;
  wire REGFILE_SIM_reg_bank_reg_r22_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_1_;
  wire REGFILE_SIM_reg_bank_reg_r22_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_20_;
  wire REGFILE_SIM_reg_bank_reg_r22_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_21_;
  wire REGFILE_SIM_reg_bank_reg_r22_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_22_;
  wire REGFILE_SIM_reg_bank_reg_r22_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_23_;
  wire REGFILE_SIM_reg_bank_reg_r22_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_24_;
  wire REGFILE_SIM_reg_bank_reg_r22_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_25_;
  wire REGFILE_SIM_reg_bank_reg_r22_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_26_;
  wire REGFILE_SIM_reg_bank_reg_r22_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_27_;
  wire REGFILE_SIM_reg_bank_reg_r22_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_28_;
  wire REGFILE_SIM_reg_bank_reg_r22_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_29_;
  wire REGFILE_SIM_reg_bank_reg_r22_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_2_;
  wire REGFILE_SIM_reg_bank_reg_r22_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_30_;
  wire REGFILE_SIM_reg_bank_reg_r22_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_31_;
  wire REGFILE_SIM_reg_bank_reg_r22_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_3_;
  wire REGFILE_SIM_reg_bank_reg_r22_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_4_;
  wire REGFILE_SIM_reg_bank_reg_r22_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_5_;
  wire REGFILE_SIM_reg_bank_reg_r22_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_6_;
  wire REGFILE_SIM_reg_bank_reg_r22_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_7_;
  wire REGFILE_SIM_reg_bank_reg_r22_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_8_;
  wire REGFILE_SIM_reg_bank_reg_r22_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r22_9_;
  wire REGFILE_SIM_reg_bank_reg_r22_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_0_;
  wire REGFILE_SIM_reg_bank_reg_r23_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_10_;
  wire REGFILE_SIM_reg_bank_reg_r23_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_11_;
  wire REGFILE_SIM_reg_bank_reg_r23_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_12_;
  wire REGFILE_SIM_reg_bank_reg_r23_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_13_;
  wire REGFILE_SIM_reg_bank_reg_r23_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_14_;
  wire REGFILE_SIM_reg_bank_reg_r23_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_15_;
  wire REGFILE_SIM_reg_bank_reg_r23_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_16_;
  wire REGFILE_SIM_reg_bank_reg_r23_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_17_;
  wire REGFILE_SIM_reg_bank_reg_r23_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_18_;
  wire REGFILE_SIM_reg_bank_reg_r23_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_19_;
  wire REGFILE_SIM_reg_bank_reg_r23_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_1_;
  wire REGFILE_SIM_reg_bank_reg_r23_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_20_;
  wire REGFILE_SIM_reg_bank_reg_r23_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_21_;
  wire REGFILE_SIM_reg_bank_reg_r23_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_22_;
  wire REGFILE_SIM_reg_bank_reg_r23_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_23_;
  wire REGFILE_SIM_reg_bank_reg_r23_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_24_;
  wire REGFILE_SIM_reg_bank_reg_r23_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_25_;
  wire REGFILE_SIM_reg_bank_reg_r23_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_26_;
  wire REGFILE_SIM_reg_bank_reg_r23_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_27_;
  wire REGFILE_SIM_reg_bank_reg_r23_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_28_;
  wire REGFILE_SIM_reg_bank_reg_r23_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_29_;
  wire REGFILE_SIM_reg_bank_reg_r23_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_2_;
  wire REGFILE_SIM_reg_bank_reg_r23_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_30_;
  wire REGFILE_SIM_reg_bank_reg_r23_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_31_;
  wire REGFILE_SIM_reg_bank_reg_r23_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_3_;
  wire REGFILE_SIM_reg_bank_reg_r23_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_4_;
  wire REGFILE_SIM_reg_bank_reg_r23_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_5_;
  wire REGFILE_SIM_reg_bank_reg_r23_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_6_;
  wire REGFILE_SIM_reg_bank_reg_r23_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_7_;
  wire REGFILE_SIM_reg_bank_reg_r23_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_8_;
  wire REGFILE_SIM_reg_bank_reg_r23_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r23_9_;
  wire REGFILE_SIM_reg_bank_reg_r23_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_0_;
  wire REGFILE_SIM_reg_bank_reg_r24_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_10_;
  wire REGFILE_SIM_reg_bank_reg_r24_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_11_;
  wire REGFILE_SIM_reg_bank_reg_r24_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_12_;
  wire REGFILE_SIM_reg_bank_reg_r24_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_13_;
  wire REGFILE_SIM_reg_bank_reg_r24_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_14_;
  wire REGFILE_SIM_reg_bank_reg_r24_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_15_;
  wire REGFILE_SIM_reg_bank_reg_r24_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_16_;
  wire REGFILE_SIM_reg_bank_reg_r24_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_17_;
  wire REGFILE_SIM_reg_bank_reg_r24_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_18_;
  wire REGFILE_SIM_reg_bank_reg_r24_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_19_;
  wire REGFILE_SIM_reg_bank_reg_r24_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_1_;
  wire REGFILE_SIM_reg_bank_reg_r24_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_20_;
  wire REGFILE_SIM_reg_bank_reg_r24_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_21_;
  wire REGFILE_SIM_reg_bank_reg_r24_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_22_;
  wire REGFILE_SIM_reg_bank_reg_r24_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_23_;
  wire REGFILE_SIM_reg_bank_reg_r24_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_24_;
  wire REGFILE_SIM_reg_bank_reg_r24_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_25_;
  wire REGFILE_SIM_reg_bank_reg_r24_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_26_;
  wire REGFILE_SIM_reg_bank_reg_r24_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_27_;
  wire REGFILE_SIM_reg_bank_reg_r24_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_28_;
  wire REGFILE_SIM_reg_bank_reg_r24_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_29_;
  wire REGFILE_SIM_reg_bank_reg_r24_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_2_;
  wire REGFILE_SIM_reg_bank_reg_r24_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_30_;
  wire REGFILE_SIM_reg_bank_reg_r24_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_31_;
  wire REGFILE_SIM_reg_bank_reg_r24_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_3_;
  wire REGFILE_SIM_reg_bank_reg_r24_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_4_;
  wire REGFILE_SIM_reg_bank_reg_r24_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_5_;
  wire REGFILE_SIM_reg_bank_reg_r24_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_6_;
  wire REGFILE_SIM_reg_bank_reg_r24_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_7_;
  wire REGFILE_SIM_reg_bank_reg_r24_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_8_;
  wire REGFILE_SIM_reg_bank_reg_r24_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r24_9_;
  wire REGFILE_SIM_reg_bank_reg_r24_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_0_;
  wire REGFILE_SIM_reg_bank_reg_r25_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_10_;
  wire REGFILE_SIM_reg_bank_reg_r25_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_11_;
  wire REGFILE_SIM_reg_bank_reg_r25_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_12_;
  wire REGFILE_SIM_reg_bank_reg_r25_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_13_;
  wire REGFILE_SIM_reg_bank_reg_r25_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_14_;
  wire REGFILE_SIM_reg_bank_reg_r25_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_15_;
  wire REGFILE_SIM_reg_bank_reg_r25_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_16_;
  wire REGFILE_SIM_reg_bank_reg_r25_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_17_;
  wire REGFILE_SIM_reg_bank_reg_r25_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_18_;
  wire REGFILE_SIM_reg_bank_reg_r25_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_19_;
  wire REGFILE_SIM_reg_bank_reg_r25_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_1_;
  wire REGFILE_SIM_reg_bank_reg_r25_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_20_;
  wire REGFILE_SIM_reg_bank_reg_r25_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_21_;
  wire REGFILE_SIM_reg_bank_reg_r25_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_22_;
  wire REGFILE_SIM_reg_bank_reg_r25_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_23_;
  wire REGFILE_SIM_reg_bank_reg_r25_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_24_;
  wire REGFILE_SIM_reg_bank_reg_r25_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_25_;
  wire REGFILE_SIM_reg_bank_reg_r25_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_26_;
  wire REGFILE_SIM_reg_bank_reg_r25_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_27_;
  wire REGFILE_SIM_reg_bank_reg_r25_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_28_;
  wire REGFILE_SIM_reg_bank_reg_r25_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_29_;
  wire REGFILE_SIM_reg_bank_reg_r25_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_2_;
  wire REGFILE_SIM_reg_bank_reg_r25_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_30_;
  wire REGFILE_SIM_reg_bank_reg_r25_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_31_;
  wire REGFILE_SIM_reg_bank_reg_r25_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_3_;
  wire REGFILE_SIM_reg_bank_reg_r25_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_4_;
  wire REGFILE_SIM_reg_bank_reg_r25_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_5_;
  wire REGFILE_SIM_reg_bank_reg_r25_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_6_;
  wire REGFILE_SIM_reg_bank_reg_r25_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_7_;
  wire REGFILE_SIM_reg_bank_reg_r25_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_8_;
  wire REGFILE_SIM_reg_bank_reg_r25_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r25_9_;
  wire REGFILE_SIM_reg_bank_reg_r25_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_0_;
  wire REGFILE_SIM_reg_bank_reg_r26_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_10_;
  wire REGFILE_SIM_reg_bank_reg_r26_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_11_;
  wire REGFILE_SIM_reg_bank_reg_r26_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_12_;
  wire REGFILE_SIM_reg_bank_reg_r26_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_13_;
  wire REGFILE_SIM_reg_bank_reg_r26_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_14_;
  wire REGFILE_SIM_reg_bank_reg_r26_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_15_;
  wire REGFILE_SIM_reg_bank_reg_r26_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_16_;
  wire REGFILE_SIM_reg_bank_reg_r26_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_17_;
  wire REGFILE_SIM_reg_bank_reg_r26_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_18_;
  wire REGFILE_SIM_reg_bank_reg_r26_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_19_;
  wire REGFILE_SIM_reg_bank_reg_r26_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_1_;
  wire REGFILE_SIM_reg_bank_reg_r26_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_20_;
  wire REGFILE_SIM_reg_bank_reg_r26_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_21_;
  wire REGFILE_SIM_reg_bank_reg_r26_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_22_;
  wire REGFILE_SIM_reg_bank_reg_r26_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_23_;
  wire REGFILE_SIM_reg_bank_reg_r26_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_24_;
  wire REGFILE_SIM_reg_bank_reg_r26_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_25_;
  wire REGFILE_SIM_reg_bank_reg_r26_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_26_;
  wire REGFILE_SIM_reg_bank_reg_r26_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_27_;
  wire REGFILE_SIM_reg_bank_reg_r26_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_28_;
  wire REGFILE_SIM_reg_bank_reg_r26_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_29_;
  wire REGFILE_SIM_reg_bank_reg_r26_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_2_;
  wire REGFILE_SIM_reg_bank_reg_r26_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_30_;
  wire REGFILE_SIM_reg_bank_reg_r26_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_31_;
  wire REGFILE_SIM_reg_bank_reg_r26_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_3_;
  wire REGFILE_SIM_reg_bank_reg_r26_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_4_;
  wire REGFILE_SIM_reg_bank_reg_r26_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_5_;
  wire REGFILE_SIM_reg_bank_reg_r26_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_6_;
  wire REGFILE_SIM_reg_bank_reg_r26_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_7_;
  wire REGFILE_SIM_reg_bank_reg_r26_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_8_;
  wire REGFILE_SIM_reg_bank_reg_r26_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r26_9_;
  wire REGFILE_SIM_reg_bank_reg_r26_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_0_;
  wire REGFILE_SIM_reg_bank_reg_r27_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_10_;
  wire REGFILE_SIM_reg_bank_reg_r27_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_11_;
  wire REGFILE_SIM_reg_bank_reg_r27_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_12_;
  wire REGFILE_SIM_reg_bank_reg_r27_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_13_;
  wire REGFILE_SIM_reg_bank_reg_r27_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_14_;
  wire REGFILE_SIM_reg_bank_reg_r27_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_15_;
  wire REGFILE_SIM_reg_bank_reg_r27_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_16_;
  wire REGFILE_SIM_reg_bank_reg_r27_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_17_;
  wire REGFILE_SIM_reg_bank_reg_r27_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_18_;
  wire REGFILE_SIM_reg_bank_reg_r27_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_19_;
  wire REGFILE_SIM_reg_bank_reg_r27_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_1_;
  wire REGFILE_SIM_reg_bank_reg_r27_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_20_;
  wire REGFILE_SIM_reg_bank_reg_r27_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_21_;
  wire REGFILE_SIM_reg_bank_reg_r27_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_22_;
  wire REGFILE_SIM_reg_bank_reg_r27_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_23_;
  wire REGFILE_SIM_reg_bank_reg_r27_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_24_;
  wire REGFILE_SIM_reg_bank_reg_r27_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_25_;
  wire REGFILE_SIM_reg_bank_reg_r27_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_26_;
  wire REGFILE_SIM_reg_bank_reg_r27_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_27_;
  wire REGFILE_SIM_reg_bank_reg_r27_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_28_;
  wire REGFILE_SIM_reg_bank_reg_r27_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_29_;
  wire REGFILE_SIM_reg_bank_reg_r27_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_2_;
  wire REGFILE_SIM_reg_bank_reg_r27_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_30_;
  wire REGFILE_SIM_reg_bank_reg_r27_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_31_;
  wire REGFILE_SIM_reg_bank_reg_r27_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_3_;
  wire REGFILE_SIM_reg_bank_reg_r27_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_4_;
  wire REGFILE_SIM_reg_bank_reg_r27_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_5_;
  wire REGFILE_SIM_reg_bank_reg_r27_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_6_;
  wire REGFILE_SIM_reg_bank_reg_r27_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_7_;
  wire REGFILE_SIM_reg_bank_reg_r27_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_8_;
  wire REGFILE_SIM_reg_bank_reg_r27_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r27_9_;
  wire REGFILE_SIM_reg_bank_reg_r27_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_0_;
  wire REGFILE_SIM_reg_bank_reg_r28_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_10_;
  wire REGFILE_SIM_reg_bank_reg_r28_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_11_;
  wire REGFILE_SIM_reg_bank_reg_r28_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_12_;
  wire REGFILE_SIM_reg_bank_reg_r28_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_13_;
  wire REGFILE_SIM_reg_bank_reg_r28_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_14_;
  wire REGFILE_SIM_reg_bank_reg_r28_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_15_;
  wire REGFILE_SIM_reg_bank_reg_r28_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_16_;
  wire REGFILE_SIM_reg_bank_reg_r28_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_17_;
  wire REGFILE_SIM_reg_bank_reg_r28_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_18_;
  wire REGFILE_SIM_reg_bank_reg_r28_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_19_;
  wire REGFILE_SIM_reg_bank_reg_r28_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_1_;
  wire REGFILE_SIM_reg_bank_reg_r28_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_20_;
  wire REGFILE_SIM_reg_bank_reg_r28_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_21_;
  wire REGFILE_SIM_reg_bank_reg_r28_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_22_;
  wire REGFILE_SIM_reg_bank_reg_r28_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_23_;
  wire REGFILE_SIM_reg_bank_reg_r28_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_24_;
  wire REGFILE_SIM_reg_bank_reg_r28_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_25_;
  wire REGFILE_SIM_reg_bank_reg_r28_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_26_;
  wire REGFILE_SIM_reg_bank_reg_r28_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_27_;
  wire REGFILE_SIM_reg_bank_reg_r28_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_28_;
  wire REGFILE_SIM_reg_bank_reg_r28_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_29_;
  wire REGFILE_SIM_reg_bank_reg_r28_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_2_;
  wire REGFILE_SIM_reg_bank_reg_r28_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_30_;
  wire REGFILE_SIM_reg_bank_reg_r28_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_31_;
  wire REGFILE_SIM_reg_bank_reg_r28_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_3_;
  wire REGFILE_SIM_reg_bank_reg_r28_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_4_;
  wire REGFILE_SIM_reg_bank_reg_r28_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_5_;
  wire REGFILE_SIM_reg_bank_reg_r28_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_6_;
  wire REGFILE_SIM_reg_bank_reg_r28_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_7_;
  wire REGFILE_SIM_reg_bank_reg_r28_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_8_;
  wire REGFILE_SIM_reg_bank_reg_r28_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r28_9_;
  wire REGFILE_SIM_reg_bank_reg_r28_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_0_;
  wire REGFILE_SIM_reg_bank_reg_r29_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_10_;
  wire REGFILE_SIM_reg_bank_reg_r29_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_11_;
  wire REGFILE_SIM_reg_bank_reg_r29_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_12_;
  wire REGFILE_SIM_reg_bank_reg_r29_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_13_;
  wire REGFILE_SIM_reg_bank_reg_r29_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_14_;
  wire REGFILE_SIM_reg_bank_reg_r29_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_15_;
  wire REGFILE_SIM_reg_bank_reg_r29_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_16_;
  wire REGFILE_SIM_reg_bank_reg_r29_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_17_;
  wire REGFILE_SIM_reg_bank_reg_r29_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_18_;
  wire REGFILE_SIM_reg_bank_reg_r29_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_19_;
  wire REGFILE_SIM_reg_bank_reg_r29_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_1_;
  wire REGFILE_SIM_reg_bank_reg_r29_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_20_;
  wire REGFILE_SIM_reg_bank_reg_r29_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_21_;
  wire REGFILE_SIM_reg_bank_reg_r29_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_22_;
  wire REGFILE_SIM_reg_bank_reg_r29_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_23_;
  wire REGFILE_SIM_reg_bank_reg_r29_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_24_;
  wire REGFILE_SIM_reg_bank_reg_r29_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_25_;
  wire REGFILE_SIM_reg_bank_reg_r29_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_26_;
  wire REGFILE_SIM_reg_bank_reg_r29_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_27_;
  wire REGFILE_SIM_reg_bank_reg_r29_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_28_;
  wire REGFILE_SIM_reg_bank_reg_r29_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_29_;
  wire REGFILE_SIM_reg_bank_reg_r29_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_2_;
  wire REGFILE_SIM_reg_bank_reg_r29_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_30_;
  wire REGFILE_SIM_reg_bank_reg_r29_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_31_;
  wire REGFILE_SIM_reg_bank_reg_r29_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_3_;
  wire REGFILE_SIM_reg_bank_reg_r29_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_4_;
  wire REGFILE_SIM_reg_bank_reg_r29_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_5_;
  wire REGFILE_SIM_reg_bank_reg_r29_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_6_;
  wire REGFILE_SIM_reg_bank_reg_r29_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_7_;
  wire REGFILE_SIM_reg_bank_reg_r29_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_8_;
  wire REGFILE_SIM_reg_bank_reg_r29_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r29_9_;
  wire REGFILE_SIM_reg_bank_reg_r29_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_0_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_10_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_11_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_12_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_13_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_14_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_15_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_16_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_17_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_18_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_19_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_1_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_20_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_21_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_22_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_23_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_24_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_25_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_26_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_27_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_28_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_29_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_2_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_30_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_31_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_3_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_4_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_5_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_6_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_7_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_8_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_9_;
  wire REGFILE_SIM_reg_bank_reg_r2_fp_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_0_;
  wire REGFILE_SIM_reg_bank_reg_r30_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_10_;
  wire REGFILE_SIM_reg_bank_reg_r30_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_11_;
  wire REGFILE_SIM_reg_bank_reg_r30_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_12_;
  wire REGFILE_SIM_reg_bank_reg_r30_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_13_;
  wire REGFILE_SIM_reg_bank_reg_r30_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_14_;
  wire REGFILE_SIM_reg_bank_reg_r30_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_15_;
  wire REGFILE_SIM_reg_bank_reg_r30_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_16_;
  wire REGFILE_SIM_reg_bank_reg_r30_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_17_;
  wire REGFILE_SIM_reg_bank_reg_r30_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_18_;
  wire REGFILE_SIM_reg_bank_reg_r30_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_19_;
  wire REGFILE_SIM_reg_bank_reg_r30_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_1_;
  wire REGFILE_SIM_reg_bank_reg_r30_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_20_;
  wire REGFILE_SIM_reg_bank_reg_r30_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_21_;
  wire REGFILE_SIM_reg_bank_reg_r30_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_22_;
  wire REGFILE_SIM_reg_bank_reg_r30_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_23_;
  wire REGFILE_SIM_reg_bank_reg_r30_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_24_;
  wire REGFILE_SIM_reg_bank_reg_r30_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_25_;
  wire REGFILE_SIM_reg_bank_reg_r30_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_26_;
  wire REGFILE_SIM_reg_bank_reg_r30_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_27_;
  wire REGFILE_SIM_reg_bank_reg_r30_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_28_;
  wire REGFILE_SIM_reg_bank_reg_r30_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_29_;
  wire REGFILE_SIM_reg_bank_reg_r30_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_2_;
  wire REGFILE_SIM_reg_bank_reg_r30_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_30_;
  wire REGFILE_SIM_reg_bank_reg_r30_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_31_;
  wire REGFILE_SIM_reg_bank_reg_r30_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_3_;
  wire REGFILE_SIM_reg_bank_reg_r30_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_4_;
  wire REGFILE_SIM_reg_bank_reg_r30_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_5_;
  wire REGFILE_SIM_reg_bank_reg_r30_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_6_;
  wire REGFILE_SIM_reg_bank_reg_r30_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_7_;
  wire REGFILE_SIM_reg_bank_reg_r30_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_8_;
  wire REGFILE_SIM_reg_bank_reg_r30_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r30_9_;
  wire REGFILE_SIM_reg_bank_reg_r30_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_0_;
  wire REGFILE_SIM_reg_bank_reg_r31_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_10_;
  wire REGFILE_SIM_reg_bank_reg_r31_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_11_;
  wire REGFILE_SIM_reg_bank_reg_r31_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_12_;
  wire REGFILE_SIM_reg_bank_reg_r31_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_13_;
  wire REGFILE_SIM_reg_bank_reg_r31_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_14_;
  wire REGFILE_SIM_reg_bank_reg_r31_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_15_;
  wire REGFILE_SIM_reg_bank_reg_r31_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_16_;
  wire REGFILE_SIM_reg_bank_reg_r31_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_17_;
  wire REGFILE_SIM_reg_bank_reg_r31_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_18_;
  wire REGFILE_SIM_reg_bank_reg_r31_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_19_;
  wire REGFILE_SIM_reg_bank_reg_r31_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_1_;
  wire REGFILE_SIM_reg_bank_reg_r31_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_20_;
  wire REGFILE_SIM_reg_bank_reg_r31_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_21_;
  wire REGFILE_SIM_reg_bank_reg_r31_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_22_;
  wire REGFILE_SIM_reg_bank_reg_r31_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_23_;
  wire REGFILE_SIM_reg_bank_reg_r31_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_24_;
  wire REGFILE_SIM_reg_bank_reg_r31_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_25_;
  wire REGFILE_SIM_reg_bank_reg_r31_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_26_;
  wire REGFILE_SIM_reg_bank_reg_r31_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_27_;
  wire REGFILE_SIM_reg_bank_reg_r31_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_28_;
  wire REGFILE_SIM_reg_bank_reg_r31_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_29_;
  wire REGFILE_SIM_reg_bank_reg_r31_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_2_;
  wire REGFILE_SIM_reg_bank_reg_r31_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_30_;
  wire REGFILE_SIM_reg_bank_reg_r31_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_31_;
  wire REGFILE_SIM_reg_bank_reg_r31_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_3_;
  wire REGFILE_SIM_reg_bank_reg_r31_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_4_;
  wire REGFILE_SIM_reg_bank_reg_r31_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_5_;
  wire REGFILE_SIM_reg_bank_reg_r31_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_6_;
  wire REGFILE_SIM_reg_bank_reg_r31_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_7_;
  wire REGFILE_SIM_reg_bank_reg_r31_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_8_;
  wire REGFILE_SIM_reg_bank_reg_r31_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r31_9_;
  wire REGFILE_SIM_reg_bank_reg_r31_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_0_;
  wire REGFILE_SIM_reg_bank_reg_r3_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_10_;
  wire REGFILE_SIM_reg_bank_reg_r3_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_11_;
  wire REGFILE_SIM_reg_bank_reg_r3_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_12_;
  wire REGFILE_SIM_reg_bank_reg_r3_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_13_;
  wire REGFILE_SIM_reg_bank_reg_r3_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_14_;
  wire REGFILE_SIM_reg_bank_reg_r3_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_15_;
  wire REGFILE_SIM_reg_bank_reg_r3_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_16_;
  wire REGFILE_SIM_reg_bank_reg_r3_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_17_;
  wire REGFILE_SIM_reg_bank_reg_r3_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_18_;
  wire REGFILE_SIM_reg_bank_reg_r3_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_19_;
  wire REGFILE_SIM_reg_bank_reg_r3_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_1_;
  wire REGFILE_SIM_reg_bank_reg_r3_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_20_;
  wire REGFILE_SIM_reg_bank_reg_r3_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_21_;
  wire REGFILE_SIM_reg_bank_reg_r3_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_22_;
  wire REGFILE_SIM_reg_bank_reg_r3_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_23_;
  wire REGFILE_SIM_reg_bank_reg_r3_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_24_;
  wire REGFILE_SIM_reg_bank_reg_r3_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_25_;
  wire REGFILE_SIM_reg_bank_reg_r3_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_26_;
  wire REGFILE_SIM_reg_bank_reg_r3_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_27_;
  wire REGFILE_SIM_reg_bank_reg_r3_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_28_;
  wire REGFILE_SIM_reg_bank_reg_r3_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_29_;
  wire REGFILE_SIM_reg_bank_reg_r3_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_2_;
  wire REGFILE_SIM_reg_bank_reg_r3_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_30_;
  wire REGFILE_SIM_reg_bank_reg_r3_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_31_;
  wire REGFILE_SIM_reg_bank_reg_r3_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_3_;
  wire REGFILE_SIM_reg_bank_reg_r3_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_4_;
  wire REGFILE_SIM_reg_bank_reg_r3_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_5_;
  wire REGFILE_SIM_reg_bank_reg_r3_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_6_;
  wire REGFILE_SIM_reg_bank_reg_r3_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_7_;
  wire REGFILE_SIM_reg_bank_reg_r3_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_8_;
  wire REGFILE_SIM_reg_bank_reg_r3_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r3_9_;
  wire REGFILE_SIM_reg_bank_reg_r3_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_0_;
  wire REGFILE_SIM_reg_bank_reg_r4_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_10_;
  wire REGFILE_SIM_reg_bank_reg_r4_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_11_;
  wire REGFILE_SIM_reg_bank_reg_r4_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_12_;
  wire REGFILE_SIM_reg_bank_reg_r4_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_13_;
  wire REGFILE_SIM_reg_bank_reg_r4_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_14_;
  wire REGFILE_SIM_reg_bank_reg_r4_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_15_;
  wire REGFILE_SIM_reg_bank_reg_r4_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_16_;
  wire REGFILE_SIM_reg_bank_reg_r4_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_17_;
  wire REGFILE_SIM_reg_bank_reg_r4_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_18_;
  wire REGFILE_SIM_reg_bank_reg_r4_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_19_;
  wire REGFILE_SIM_reg_bank_reg_r4_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_1_;
  wire REGFILE_SIM_reg_bank_reg_r4_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_20_;
  wire REGFILE_SIM_reg_bank_reg_r4_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_21_;
  wire REGFILE_SIM_reg_bank_reg_r4_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_22_;
  wire REGFILE_SIM_reg_bank_reg_r4_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_23_;
  wire REGFILE_SIM_reg_bank_reg_r4_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_24_;
  wire REGFILE_SIM_reg_bank_reg_r4_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_25_;
  wire REGFILE_SIM_reg_bank_reg_r4_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_26_;
  wire REGFILE_SIM_reg_bank_reg_r4_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_27_;
  wire REGFILE_SIM_reg_bank_reg_r4_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_28_;
  wire REGFILE_SIM_reg_bank_reg_r4_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_29_;
  wire REGFILE_SIM_reg_bank_reg_r4_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_2_;
  wire REGFILE_SIM_reg_bank_reg_r4_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_30_;
  wire REGFILE_SIM_reg_bank_reg_r4_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_31_;
  wire REGFILE_SIM_reg_bank_reg_r4_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_3_;
  wire REGFILE_SIM_reg_bank_reg_r4_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_4_;
  wire REGFILE_SIM_reg_bank_reg_r4_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_5_;
  wire REGFILE_SIM_reg_bank_reg_r4_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_6_;
  wire REGFILE_SIM_reg_bank_reg_r4_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_7_;
  wire REGFILE_SIM_reg_bank_reg_r4_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_8_;
  wire REGFILE_SIM_reg_bank_reg_r4_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r4_9_;
  wire REGFILE_SIM_reg_bank_reg_r4_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_0_;
  wire REGFILE_SIM_reg_bank_reg_r5_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_10_;
  wire REGFILE_SIM_reg_bank_reg_r5_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_11_;
  wire REGFILE_SIM_reg_bank_reg_r5_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_12_;
  wire REGFILE_SIM_reg_bank_reg_r5_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_13_;
  wire REGFILE_SIM_reg_bank_reg_r5_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_14_;
  wire REGFILE_SIM_reg_bank_reg_r5_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_15_;
  wire REGFILE_SIM_reg_bank_reg_r5_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_16_;
  wire REGFILE_SIM_reg_bank_reg_r5_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_17_;
  wire REGFILE_SIM_reg_bank_reg_r5_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_18_;
  wire REGFILE_SIM_reg_bank_reg_r5_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_19_;
  wire REGFILE_SIM_reg_bank_reg_r5_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_1_;
  wire REGFILE_SIM_reg_bank_reg_r5_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_20_;
  wire REGFILE_SIM_reg_bank_reg_r5_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_21_;
  wire REGFILE_SIM_reg_bank_reg_r5_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_22_;
  wire REGFILE_SIM_reg_bank_reg_r5_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_23_;
  wire REGFILE_SIM_reg_bank_reg_r5_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_24_;
  wire REGFILE_SIM_reg_bank_reg_r5_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_25_;
  wire REGFILE_SIM_reg_bank_reg_r5_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_26_;
  wire REGFILE_SIM_reg_bank_reg_r5_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_27_;
  wire REGFILE_SIM_reg_bank_reg_r5_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_28_;
  wire REGFILE_SIM_reg_bank_reg_r5_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_29_;
  wire REGFILE_SIM_reg_bank_reg_r5_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_2_;
  wire REGFILE_SIM_reg_bank_reg_r5_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_30_;
  wire REGFILE_SIM_reg_bank_reg_r5_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_31_;
  wire REGFILE_SIM_reg_bank_reg_r5_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_3_;
  wire REGFILE_SIM_reg_bank_reg_r5_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_4_;
  wire REGFILE_SIM_reg_bank_reg_r5_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_5_;
  wire REGFILE_SIM_reg_bank_reg_r5_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_6_;
  wire REGFILE_SIM_reg_bank_reg_r5_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_7_;
  wire REGFILE_SIM_reg_bank_reg_r5_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_8_;
  wire REGFILE_SIM_reg_bank_reg_r5_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r5_9_;
  wire REGFILE_SIM_reg_bank_reg_r5_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_0_;
  wire REGFILE_SIM_reg_bank_reg_r6_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_10_;
  wire REGFILE_SIM_reg_bank_reg_r6_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_11_;
  wire REGFILE_SIM_reg_bank_reg_r6_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_12_;
  wire REGFILE_SIM_reg_bank_reg_r6_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_13_;
  wire REGFILE_SIM_reg_bank_reg_r6_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_14_;
  wire REGFILE_SIM_reg_bank_reg_r6_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_15_;
  wire REGFILE_SIM_reg_bank_reg_r6_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_16_;
  wire REGFILE_SIM_reg_bank_reg_r6_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_17_;
  wire REGFILE_SIM_reg_bank_reg_r6_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_18_;
  wire REGFILE_SIM_reg_bank_reg_r6_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_19_;
  wire REGFILE_SIM_reg_bank_reg_r6_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_1_;
  wire REGFILE_SIM_reg_bank_reg_r6_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_20_;
  wire REGFILE_SIM_reg_bank_reg_r6_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_21_;
  wire REGFILE_SIM_reg_bank_reg_r6_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_22_;
  wire REGFILE_SIM_reg_bank_reg_r6_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_23_;
  wire REGFILE_SIM_reg_bank_reg_r6_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_24_;
  wire REGFILE_SIM_reg_bank_reg_r6_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_25_;
  wire REGFILE_SIM_reg_bank_reg_r6_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_26_;
  wire REGFILE_SIM_reg_bank_reg_r6_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_27_;
  wire REGFILE_SIM_reg_bank_reg_r6_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_28_;
  wire REGFILE_SIM_reg_bank_reg_r6_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_29_;
  wire REGFILE_SIM_reg_bank_reg_r6_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_2_;
  wire REGFILE_SIM_reg_bank_reg_r6_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_30_;
  wire REGFILE_SIM_reg_bank_reg_r6_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_31_;
  wire REGFILE_SIM_reg_bank_reg_r6_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_3_;
  wire REGFILE_SIM_reg_bank_reg_r6_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_4_;
  wire REGFILE_SIM_reg_bank_reg_r6_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_5_;
  wire REGFILE_SIM_reg_bank_reg_r6_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_6_;
  wire REGFILE_SIM_reg_bank_reg_r6_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_7_;
  wire REGFILE_SIM_reg_bank_reg_r6_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_8_;
  wire REGFILE_SIM_reg_bank_reg_r6_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r6_9_;
  wire REGFILE_SIM_reg_bank_reg_r6_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_0_;
  wire REGFILE_SIM_reg_bank_reg_r7_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_10_;
  wire REGFILE_SIM_reg_bank_reg_r7_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_11_;
  wire REGFILE_SIM_reg_bank_reg_r7_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_12_;
  wire REGFILE_SIM_reg_bank_reg_r7_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_13_;
  wire REGFILE_SIM_reg_bank_reg_r7_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_14_;
  wire REGFILE_SIM_reg_bank_reg_r7_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_15_;
  wire REGFILE_SIM_reg_bank_reg_r7_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_16_;
  wire REGFILE_SIM_reg_bank_reg_r7_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_17_;
  wire REGFILE_SIM_reg_bank_reg_r7_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_18_;
  wire REGFILE_SIM_reg_bank_reg_r7_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_19_;
  wire REGFILE_SIM_reg_bank_reg_r7_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_1_;
  wire REGFILE_SIM_reg_bank_reg_r7_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_20_;
  wire REGFILE_SIM_reg_bank_reg_r7_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_21_;
  wire REGFILE_SIM_reg_bank_reg_r7_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_22_;
  wire REGFILE_SIM_reg_bank_reg_r7_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_23_;
  wire REGFILE_SIM_reg_bank_reg_r7_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_24_;
  wire REGFILE_SIM_reg_bank_reg_r7_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_25_;
  wire REGFILE_SIM_reg_bank_reg_r7_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_26_;
  wire REGFILE_SIM_reg_bank_reg_r7_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_27_;
  wire REGFILE_SIM_reg_bank_reg_r7_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_28_;
  wire REGFILE_SIM_reg_bank_reg_r7_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_29_;
  wire REGFILE_SIM_reg_bank_reg_r7_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_2_;
  wire REGFILE_SIM_reg_bank_reg_r7_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_30_;
  wire REGFILE_SIM_reg_bank_reg_r7_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_31_;
  wire REGFILE_SIM_reg_bank_reg_r7_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_3_;
  wire REGFILE_SIM_reg_bank_reg_r7_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_4_;
  wire REGFILE_SIM_reg_bank_reg_r7_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_5_;
  wire REGFILE_SIM_reg_bank_reg_r7_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_6_;
  wire REGFILE_SIM_reg_bank_reg_r7_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_7_;
  wire REGFILE_SIM_reg_bank_reg_r7_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_8_;
  wire REGFILE_SIM_reg_bank_reg_r7_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r7_9_;
  wire REGFILE_SIM_reg_bank_reg_r7_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_0_;
  wire REGFILE_SIM_reg_bank_reg_r8_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_10_;
  wire REGFILE_SIM_reg_bank_reg_r8_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_11_;
  wire REGFILE_SIM_reg_bank_reg_r8_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_12_;
  wire REGFILE_SIM_reg_bank_reg_r8_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_13_;
  wire REGFILE_SIM_reg_bank_reg_r8_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_14_;
  wire REGFILE_SIM_reg_bank_reg_r8_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_15_;
  wire REGFILE_SIM_reg_bank_reg_r8_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_16_;
  wire REGFILE_SIM_reg_bank_reg_r8_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_17_;
  wire REGFILE_SIM_reg_bank_reg_r8_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_18_;
  wire REGFILE_SIM_reg_bank_reg_r8_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_19_;
  wire REGFILE_SIM_reg_bank_reg_r8_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_1_;
  wire REGFILE_SIM_reg_bank_reg_r8_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_20_;
  wire REGFILE_SIM_reg_bank_reg_r8_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_21_;
  wire REGFILE_SIM_reg_bank_reg_r8_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_22_;
  wire REGFILE_SIM_reg_bank_reg_r8_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_23_;
  wire REGFILE_SIM_reg_bank_reg_r8_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_24_;
  wire REGFILE_SIM_reg_bank_reg_r8_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_25_;
  wire REGFILE_SIM_reg_bank_reg_r8_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_26_;
  wire REGFILE_SIM_reg_bank_reg_r8_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_27_;
  wire REGFILE_SIM_reg_bank_reg_r8_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_28_;
  wire REGFILE_SIM_reg_bank_reg_r8_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_29_;
  wire REGFILE_SIM_reg_bank_reg_r8_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_2_;
  wire REGFILE_SIM_reg_bank_reg_r8_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_30_;
  wire REGFILE_SIM_reg_bank_reg_r8_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_31_;
  wire REGFILE_SIM_reg_bank_reg_r8_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_3_;
  wire REGFILE_SIM_reg_bank_reg_r8_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_4_;
  wire REGFILE_SIM_reg_bank_reg_r8_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_5_;
  wire REGFILE_SIM_reg_bank_reg_r8_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_6_;
  wire REGFILE_SIM_reg_bank_reg_r8_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_7_;
  wire REGFILE_SIM_reg_bank_reg_r8_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_8_;
  wire REGFILE_SIM_reg_bank_reg_r8_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r8_9_;
  wire REGFILE_SIM_reg_bank_reg_r8_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_0_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_0__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_10_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_10__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_11_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_11__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_12_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_12__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_13_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_13__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_14_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_14__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_15_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_15__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_16_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_16__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_17_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_17__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_18_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_18__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_19_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_19__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_1_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_1__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_20_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_20__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_21_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_21__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_22_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_22__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_23_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_23__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_24_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_24__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_25_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_25__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_26_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_26__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_27_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_27__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_28_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_28__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_29_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_29__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_2_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_2__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_30_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_30__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_31_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_31__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_3_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_3__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_4_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_4__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_5_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_5__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_6_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_6__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_7_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_7__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_8_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_8__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_9_;
  wire REGFILE_SIM_reg_bank_reg_r9_lr_9__FF_INPUT;
  wire REGFILE_SIM_reg_bank_reg_ra_o_0_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_10_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_11_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_12_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_13_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_14_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_15_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_16_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_17_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_18_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_19_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_1_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_20_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_21_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_22_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_23_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_24_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_25_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_26_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_27_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_28_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_29_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_2_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_30_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_31_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_3_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_4_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_5_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_6_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_7_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_8_;
  wire REGFILE_SIM_reg_bank_reg_ra_o_9_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_0_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_10_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_11_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_12_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_13_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_14_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_15_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_16_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_17_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_18_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_19_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_1_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_20_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_21_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_22_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_23_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_24_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_25_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_26_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_27_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_28_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_29_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_2_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_30_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_31_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_3_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_4_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_5_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_6_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_7_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_8_;
  wire REGFILE_SIM_reg_bank_reg_rb_o_9_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_0_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_10_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_11_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_12_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_13_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_14_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_15_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_16_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_17_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_18_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_19_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_1_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_20_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_21_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_22_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_23_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_24_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_25_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_26_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_27_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_28_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_29_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_2_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_30_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_31_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_3_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_4_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_5_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_6_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_7_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_8_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3;
  wire REGFILE_SIM_reg_bank_reg_rd_i_9_;
  wire REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0;
  wire REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1;
  wire REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2;
  wire REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3;
  wire REGFILE_SIM_reg_bank_wr_i;
  wire REGFILE_SIM_reg_bank_wr_i_bF_buf0;
  wire REGFILE_SIM_reg_bank_wr_i_bF_buf1;
  wire REGFILE_SIM_reg_bank_wr_i_bF_buf2;
  wire REGFILE_SIM_reg_bank_wr_i_bF_buf3;
  wire REGFILE_SIM_reg_bank_wr_i_bF_buf4;
  wire REGFILE_SIM_reg_bank_wr_i_bF_buf5;
  wire _abc_27555_n185;
  wire _abc_27555_n288;
  wire _abc_27555_n343;
  wire _abc_27555_n353;
  wire _abc_27555_n4360;
  wire _abc_27555_n4367;
  wire _abc_27555_n4367_bF_buf0;
  wire _abc_27555_n4367_bF_buf1;
  wire _abc_27555_n4367_bF_buf2;
  wire _abc_27555_n4367_bF_buf3;
  wire _abc_27555_n4367_bF_buf4;
  wire _abc_27555_n4367_bF_buf5;
  wire _abc_27555_n4367_bF_buf6;
  wire _abc_27555_n4367_bF_buf7;
  wire _abc_43815_n1000;
  wire _abc_43815_n1001;
  wire _abc_43815_n1002;
  wire _abc_43815_n1003;
  wire _abc_43815_n1004;
  wire _abc_43815_n1005;
  wire _abc_43815_n1006;
  wire _abc_43815_n1007;
  wire _abc_43815_n1008;
  wire _abc_43815_n1009_1;
  wire _abc_43815_n1010;
  wire _abc_43815_n1011;
  wire _abc_43815_n1012;
  wire _abc_43815_n1013;
  wire _abc_43815_n1014;
  wire _abc_43815_n1015;
  wire _abc_43815_n1016;
  wire _abc_43815_n1017;
  wire _abc_43815_n1018;
  wire _abc_43815_n1019;
  wire _abc_43815_n1020;
  wire _abc_43815_n1021;
  wire _abc_43815_n1022;
  wire _abc_43815_n1023;
  wire _abc_43815_n1024;
  wire _abc_43815_n1025;
  wire _abc_43815_n1026;
  wire _abc_43815_n1027;
  wire _abc_43815_n1028;
  wire _abc_43815_n1029;
  wire _abc_43815_n1030;
  wire _abc_43815_n1031_1;
  wire _abc_43815_n1032_1;
  wire _abc_43815_n1033;
  wire _abc_43815_n1034;
  wire _abc_43815_n1035;
  wire _abc_43815_n1036;
  wire _abc_43815_n1037;
  wire _abc_43815_n1038;
  wire _abc_43815_n1039;
  wire _abc_43815_n1040;
  wire _abc_43815_n1041;
  wire _abc_43815_n1042;
  wire _abc_43815_n1043_1;
  wire _abc_43815_n1044;
  wire _abc_43815_n1045;
  wire _abc_43815_n1046_1;
  wire _abc_43815_n1047;
  wire _abc_43815_n1048;
  wire _abc_43815_n1049;
  wire _abc_43815_n1050;
  wire _abc_43815_n1051;
  wire _abc_43815_n1052;
  wire _abc_43815_n1053;
  wire _abc_43815_n1054;
  wire _abc_43815_n1055;
  wire _abc_43815_n1056;
  wire _abc_43815_n1057;
  wire _abc_43815_n1058;
  wire _abc_43815_n1059;
  wire _abc_43815_n1060;
  wire _abc_43815_n1060_bF_buf0;
  wire _abc_43815_n1060_bF_buf1;
  wire _abc_43815_n1060_bF_buf2;
  wire _abc_43815_n1060_bF_buf3;
  wire _abc_43815_n1061;
  wire _abc_43815_n1062;
  wire _abc_43815_n1063;
  wire _abc_43815_n1064_1;
  wire _abc_43815_n1065_1;
  wire _abc_43815_n1065_1_bF_buf0;
  wire _abc_43815_n1065_1_bF_buf1;
  wire _abc_43815_n1065_1_bF_buf2;
  wire _abc_43815_n1065_1_bF_buf3;
  wire _abc_43815_n1065_1_bF_buf4;
  wire _abc_43815_n1066;
  wire _abc_43815_n1067;
  wire _abc_43815_n1068;
  wire _abc_43815_n1069;
  wire _abc_43815_n1070;
  wire _abc_43815_n1071;
  wire _abc_43815_n1072;
  wire _abc_43815_n1073;
  wire _abc_43815_n1074;
  wire _abc_43815_n1075;
  wire _abc_43815_n1076;
  wire _abc_43815_n1077;
  wire _abc_43815_n1078;
  wire _abc_43815_n1079;
  wire _abc_43815_n1080;
  wire _abc_43815_n1081;
  wire _abc_43815_n1082;
  wire _abc_43815_n1083_1;
  wire _abc_43815_n1084;
  wire _abc_43815_n1085;
  wire _abc_43815_n1086_1;
  wire _abc_43815_n1087;
  wire _abc_43815_n1088;
  wire _abc_43815_n1089;
  wire _abc_43815_n1090;
  wire _abc_43815_n1091;
  wire _abc_43815_n1092;
  wire _abc_43815_n1093;
  wire _abc_43815_n1094;
  wire _abc_43815_n1095;
  wire _abc_43815_n1096;
  wire _abc_43815_n1097;
  wire _abc_43815_n1098;
  wire _abc_43815_n1099;
  wire _abc_43815_n1100;
  wire _abc_43815_n1101;
  wire _abc_43815_n1102_1;
  wire _abc_43815_n1103_1;
  wire _abc_43815_n1104;
  wire _abc_43815_n1105;
  wire _abc_43815_n1106;
  wire _abc_43815_n1107;
  wire _abc_43815_n1108_1;
  wire _abc_43815_n1109;
  wire _abc_43815_n1110;
  wire _abc_43815_n1111;
  wire _abc_43815_n1112;
  wire _abc_43815_n1113;
  wire _abc_43815_n1114;
  wire _abc_43815_n1115;
  wire _abc_43815_n1116_1;
  wire _abc_43815_n1117;
  wire _abc_43815_n1118;
  wire _abc_43815_n1119_1;
  wire _abc_43815_n1120;
  wire _abc_43815_n1121;
  wire _abc_43815_n1122;
  wire _abc_43815_n1123;
  wire _abc_43815_n1124;
  wire _abc_43815_n1125;
  wire _abc_43815_n1126;
  wire _abc_43815_n1127;
  wire _abc_43815_n1128;
  wire _abc_43815_n1129;
  wire _abc_43815_n1130;
  wire _abc_43815_n1131;
  wire _abc_43815_n1132;
  wire _abc_43815_n1133;
  wire _abc_43815_n1134;
  wire _abc_43815_n1135_1;
  wire _abc_43815_n1136_1;
  wire _abc_43815_n1137;
  wire _abc_43815_n1138;
  wire _abc_43815_n1139;
  wire _abc_43815_n1140;
  wire _abc_43815_n1141;
  wire _abc_43815_n1142_1;
  wire _abc_43815_n1143;
  wire _abc_43815_n1144;
  wire _abc_43815_n1145;
  wire _abc_43815_n1146;
  wire _abc_43815_n1147;
  wire _abc_43815_n1148;
  wire _abc_43815_n1149;
  wire _abc_43815_n1150;
  wire _abc_43815_n1151;
  wire _abc_43815_n1152;
  wire _abc_43815_n1153_1;
  wire _abc_43815_n1154;
  wire _abc_43815_n1155;
  wire _abc_43815_n1156_1;
  wire _abc_43815_n1157;
  wire _abc_43815_n1158;
  wire _abc_43815_n1159;
  wire _abc_43815_n1160;
  wire _abc_43815_n1161;
  wire _abc_43815_n1162;
  wire _abc_43815_n1163;
  wire _abc_43815_n1164;
  wire _abc_43815_n1165;
  wire _abc_43815_n1166;
  wire _abc_43815_n1167;
  wire _abc_43815_n1168;
  wire _abc_43815_n1169;
  wire _abc_43815_n1170;
  wire _abc_43815_n1171;
  wire _abc_43815_n1171_bF_buf0;
  wire _abc_43815_n1171_bF_buf1;
  wire _abc_43815_n1171_bF_buf2;
  wire _abc_43815_n1171_bF_buf3;
  wire _abc_43815_n1171_bF_buf4;
  wire _abc_43815_n1171_bF_buf5;
  wire _abc_43815_n1172_1;
  wire _abc_43815_n1172_1_bF_buf0;
  wire _abc_43815_n1172_1_bF_buf1;
  wire _abc_43815_n1172_1_bF_buf2;
  wire _abc_43815_n1172_1_bF_buf3;
  wire _abc_43815_n1172_1_bF_buf4;
  wire _abc_43815_n1173_1;
  wire _abc_43815_n1174;
  wire _abc_43815_n1175;
  wire _abc_43815_n1176;
  wire _abc_43815_n1177;
  wire _abc_43815_n1178_1;
  wire _abc_43815_n1179;
  wire _abc_43815_n1180;
  wire _abc_43815_n1181;
  wire _abc_43815_n1182;
  wire _abc_43815_n1183;
  wire _abc_43815_n1184;
  wire _abc_43815_n1185;
  wire _abc_43815_n1186_1;
  wire _abc_43815_n1187;
  wire _abc_43815_n1188;
  wire _abc_43815_n1189_1;
  wire _abc_43815_n1190;
  wire _abc_43815_n1191;
  wire _abc_43815_n1192;
  wire _abc_43815_n1193;
  wire _abc_43815_n1194;
  wire _abc_43815_n1195;
  wire _abc_43815_n1196;
  wire _abc_43815_n1197;
  wire _abc_43815_n1198;
  wire _abc_43815_n1199;
  wire _abc_43815_n1200;
  wire _abc_43815_n1201;
  wire _abc_43815_n1202;
  wire _abc_43815_n1203;
  wire _abc_43815_n1204;
  wire _abc_43815_n1205_1;
  wire _abc_43815_n1206_1;
  wire _abc_43815_n1207;
  wire _abc_43815_n1208;
  wire _abc_43815_n1209;
  wire _abc_43815_n1210;
  wire _abc_43815_n1211;
  wire _abc_43815_n1212;
  wire _abc_43815_n1213;
  wire _abc_43815_n1214_1;
  wire _abc_43815_n1215;
  wire _abc_43815_n1216;
  wire _abc_43815_n1217;
  wire _abc_43815_n1218;
  wire _abc_43815_n1219;
  wire _abc_43815_n1220;
  wire _abc_43815_n1221;
  wire _abc_43815_n1222;
  wire _abc_43815_n1223;
  wire _abc_43815_n1224;
  wire _abc_43815_n1225;
  wire _abc_43815_n1226;
  wire _abc_43815_n1227;
  wire _abc_43815_n1228;
  wire _abc_43815_n1229;
  wire _abc_43815_n1230_1;
  wire _abc_43815_n1231;
  wire _abc_43815_n1232;
  wire _abc_43815_n1233_1;
  wire _abc_43815_n1234;
  wire _abc_43815_n1235;
  wire _abc_43815_n1236;
  wire _abc_43815_n1237;
  wire _abc_43815_n1238;
  wire _abc_43815_n1239;
  wire _abc_43815_n1240;
  wire _abc_43815_n1241;
  wire _abc_43815_n1242;
  wire _abc_43815_n1243;
  wire _abc_43815_n1244;
  wire _abc_43815_n1245;
  wire _abc_43815_n1246;
  wire _abc_43815_n1247;
  wire _abc_43815_n1248;
  wire _abc_43815_n1249_1;
  wire _abc_43815_n1250_1;
  wire _abc_43815_n1251;
  wire _abc_43815_n1252;
  wire _abc_43815_n1253;
  wire _abc_43815_n1254;
  wire _abc_43815_n1255_1;
  wire _abc_43815_n1256;
  wire _abc_43815_n1257;
  wire _abc_43815_n1258;
  wire _abc_43815_n1259;
  wire _abc_43815_n1260;
  wire _abc_43815_n1261;
  wire _abc_43815_n1262;
  wire _abc_43815_n1263_1;
  wire _abc_43815_n1264;
  wire _abc_43815_n1265;
  wire _abc_43815_n1266_1;
  wire _abc_43815_n1267;
  wire _abc_43815_n1268;
  wire _abc_43815_n1269;
  wire _abc_43815_n1270;
  wire _abc_43815_n1271;
  wire _abc_43815_n1272;
  wire _abc_43815_n1273;
  wire _abc_43815_n1274;
  wire _abc_43815_n1275;
  wire _abc_43815_n1276;
  wire _abc_43815_n1277;
  wire _abc_43815_n1278;
  wire _abc_43815_n1278_bF_buf0;
  wire _abc_43815_n1278_bF_buf1;
  wire _abc_43815_n1278_bF_buf2;
  wire _abc_43815_n1278_bF_buf3;
  wire _abc_43815_n1278_bF_buf4;
  wire _abc_43815_n1278_bF_buf5;
  wire _abc_43815_n1278_bF_buf6;
  wire _abc_43815_n1278_bF_buf7;
  wire _abc_43815_n1279;
  wire _abc_43815_n1280;
  wire _abc_43815_n1281;
  wire _abc_43815_n1282_1;
  wire _abc_43815_n1283_1;
  wire _abc_43815_n1285;
  wire _abc_43815_n1286;
  wire _abc_43815_n1287;
  wire _abc_43815_n1288;
  wire _abc_43815_n1289_1;
  wire _abc_43815_n1290;
  wire _abc_43815_n1291;
  wire _abc_43815_n1292;
  wire _abc_43815_n1293;
  wire _abc_43815_n1294;
  wire _abc_43815_n1295;
  wire _abc_43815_n1296;
  wire _abc_43815_n1297;
  wire _abc_43815_n1298;
  wire _abc_43815_n1299;
  wire _abc_43815_n1300_1;
  wire _abc_43815_n1301;
  wire _abc_43815_n1302;
  wire _abc_43815_n1303_1;
  wire _abc_43815_n1304;
  wire _abc_43815_n1305;
  wire _abc_43815_n1306;
  wire _abc_43815_n1307;
  wire _abc_43815_n1308;
  wire _abc_43815_n1309;
  wire _abc_43815_n1310;
  wire _abc_43815_n1311;
  wire _abc_43815_n1312;
  wire _abc_43815_n1313;
  wire _abc_43815_n1314;
  wire _abc_43815_n1315;
  wire _abc_43815_n1316;
  wire _abc_43815_n1317;
  wire _abc_43815_n1318;
  wire _abc_43815_n1319_1;
  wire _abc_43815_n1320_1;
  wire _abc_43815_n1321;
  wire _abc_43815_n1322;
  wire _abc_43815_n1323;
  wire _abc_43815_n1324;
  wire _abc_43815_n1325_1;
  wire _abc_43815_n1326;
  wire _abc_43815_n1327;
  wire _abc_43815_n1328;
  wire _abc_43815_n1329;
  wire _abc_43815_n1330;
  wire _abc_43815_n1331;
  wire _abc_43815_n1332;
  wire _abc_43815_n1333_1;
  wire _abc_43815_n1334;
  wire _abc_43815_n1335;
  wire _abc_43815_n1336_1;
  wire _abc_43815_n1337;
  wire _abc_43815_n1338;
  wire _abc_43815_n1339;
  wire _abc_43815_n1340;
  wire _abc_43815_n1341;
  wire _abc_43815_n1342;
  wire _abc_43815_n1343;
  wire _abc_43815_n1344;
  wire _abc_43815_n1345;
  wire _abc_43815_n1346;
  wire _abc_43815_n1347;
  wire _abc_43815_n1348;
  wire _abc_43815_n1349;
  wire _abc_43815_n1350;
  wire _abc_43815_n1350_bF_buf0;
  wire _abc_43815_n1350_bF_buf1;
  wire _abc_43815_n1350_bF_buf2;
  wire _abc_43815_n1350_bF_buf3;
  wire _abc_43815_n1350_bF_buf4;
  wire _abc_43815_n1351;
  wire _abc_43815_n1351_bF_buf0;
  wire _abc_43815_n1351_bF_buf1;
  wire _abc_43815_n1351_bF_buf2;
  wire _abc_43815_n1351_bF_buf3;
  wire _abc_43815_n1351_bF_buf4;
  wire _abc_43815_n1352_1;
  wire _abc_43815_n1353_1;
  wire _abc_43815_n1354;
  wire _abc_43815_n1355;
  wire _abc_43815_n1356;
  wire _abc_43815_n1357;
  wire _abc_43815_n1358;
  wire _abc_43815_n1359;
  wire _abc_43815_n1360_1;
  wire _abc_43815_n1361;
  wire _abc_43815_n1362;
  wire _abc_43815_n1363;
  wire _abc_43815_n1364;
  wire _abc_43815_n1366;
  wire _abc_43815_n1367;
  wire _abc_43815_n1368;
  wire _abc_43815_n1369;
  wire _abc_43815_n1370;
  wire _abc_43815_n1371;
  wire _abc_43815_n1372_1;
  wire _abc_43815_n1373;
  wire _abc_43815_n1374;
  wire _abc_43815_n1375_1;
  wire _abc_43815_n1376;
  wire _abc_43815_n1377;
  wire _abc_43815_n1378;
  wire _abc_43815_n1379;
  wire _abc_43815_n1380;
  wire _abc_43815_n1381;
  wire _abc_43815_n1382;
  wire _abc_43815_n1383;
  wire _abc_43815_n1384;
  wire _abc_43815_n1385;
  wire _abc_43815_n1386;
  wire _abc_43815_n1387;
  wire _abc_43815_n1388;
  wire _abc_43815_n1389;
  wire _abc_43815_n1390;
  wire _abc_43815_n1391_1;
  wire _abc_43815_n1392_1;
  wire _abc_43815_n1393;
  wire _abc_43815_n1394;
  wire _abc_43815_n1395;
  wire _abc_43815_n1396;
  wire _abc_43815_n1398;
  wire _abc_43815_n1399;
  wire _abc_43815_n1399_bF_buf0;
  wire _abc_43815_n1399_bF_buf1;
  wire _abc_43815_n1399_bF_buf2;
  wire _abc_43815_n1399_bF_buf3;
  wire _abc_43815_n1399_bF_buf4;
  wire _abc_43815_n1400;
  wire _abc_43815_n1401;
  wire _abc_43815_n1402;
  wire _abc_43815_n1404;
  wire _abc_43815_n1405_1;
  wire _abc_43815_n1406;
  wire _abc_43815_n1408_1;
  wire _abc_43815_n1409;
  wire _abc_43815_n1410;
  wire _abc_43815_n1412;
  wire _abc_43815_n1413;
  wire _abc_43815_n1413_bF_buf0;
  wire _abc_43815_n1413_bF_buf1;
  wire _abc_43815_n1413_bF_buf2;
  wire _abc_43815_n1413_bF_buf3;
  wire _abc_43815_n1413_bF_buf4;
  wire _abc_43815_n1414;
  wire _abc_43815_n1415;
  wire _abc_43815_n1416;
  wire _abc_43815_n1417;
  wire _abc_43815_n1418;
  wire _abc_43815_n1418_bF_buf0;
  wire _abc_43815_n1418_bF_buf1;
  wire _abc_43815_n1418_bF_buf2;
  wire _abc_43815_n1418_bF_buf3;
  wire _abc_43815_n1418_bF_buf4;
  wire _abc_43815_n1418_bF_buf5;
  wire _abc_43815_n1419;
  wire _abc_43815_n1420;
  wire _abc_43815_n1421;
  wire _abc_43815_n1422;
  wire _abc_43815_n1423;
  wire _abc_43815_n1424_1;
  wire _abc_43815_n1425_1;
  wire _abc_43815_n1425_1_bF_buf0;
  wire _abc_43815_n1425_1_bF_buf1;
  wire _abc_43815_n1425_1_bF_buf2;
  wire _abc_43815_n1425_1_bF_buf3;
  wire _abc_43815_n1425_1_bF_buf4;
  wire _abc_43815_n1426;
  wire _abc_43815_n1427;
  wire _abc_43815_n1428;
  wire _abc_43815_n1428_bF_buf0;
  wire _abc_43815_n1428_bF_buf1;
  wire _abc_43815_n1428_bF_buf2;
  wire _abc_43815_n1428_bF_buf3;
  wire _abc_43815_n1428_bF_buf4;
  wire _abc_43815_n1429;
  wire _abc_43815_n1430;
  wire _abc_43815_n1431_1;
  wire _abc_43815_n1431_1_bF_buf0;
  wire _abc_43815_n1431_1_bF_buf1;
  wire _abc_43815_n1431_1_bF_buf2;
  wire _abc_43815_n1431_1_bF_buf3;
  wire _abc_43815_n1431_1_bF_buf4;
  wire _abc_43815_n1432;
  wire _abc_43815_n1433;
  wire _abc_43815_n1434;
  wire _abc_43815_n1435;
  wire _abc_43815_n1436;
  wire _abc_43815_n1437;
  wire _abc_43815_n1438;
  wire _abc_43815_n1439;
  wire _abc_43815_n1441;
  wire _abc_43815_n1442;
  wire _abc_43815_n1443_1;
  wire _abc_43815_n1444;
  wire _abc_43815_n1445;
  wire _abc_43815_n1446;
  wire _abc_43815_n1447;
  wire _abc_43815_n1448;
  wire _abc_43815_n1449;
  wire _abc_43815_n1450;
  wire _abc_43815_n1451;
  wire _abc_43815_n1452;
  wire _abc_43815_n1453;
  wire _abc_43815_n1454;
  wire _abc_43815_n1455;
  wire _abc_43815_n1456;
  wire _abc_43815_n1457;
  wire _abc_43815_n1458;
  wire _abc_43815_n1459_1;
  wire _abc_43815_n1461;
  wire _abc_43815_n1461_bF_buf0;
  wire _abc_43815_n1461_bF_buf1;
  wire _abc_43815_n1461_bF_buf2;
  wire _abc_43815_n1461_bF_buf3;
  wire _abc_43815_n1462;
  wire _abc_43815_n1463;
  wire _abc_43815_n1464;
  wire _abc_43815_n1465;
  wire _abc_43815_n1466;
  wire _abc_43815_n1467;
  wire _abc_43815_n1468;
  wire _abc_43815_n1469;
  wire _abc_43815_n1470;
  wire _abc_43815_n1471;
  wire _abc_43815_n1472_1;
  wire _abc_43815_n1472_1_bF_buf0;
  wire _abc_43815_n1472_1_bF_buf1;
  wire _abc_43815_n1472_1_bF_buf2;
  wire _abc_43815_n1472_1_bF_buf3;
  wire _abc_43815_n1472_1_bF_buf4;
  wire _abc_43815_n1473;
  wire _abc_43815_n1473_bF_buf0;
  wire _abc_43815_n1473_bF_buf1;
  wire _abc_43815_n1473_bF_buf2;
  wire _abc_43815_n1473_bF_buf3;
  wire _abc_43815_n1473_bF_buf4;
  wire _abc_43815_n1474;
  wire _abc_43815_n1475_1;
  wire _abc_43815_n1476;
  wire _abc_43815_n1477;
  wire _abc_43815_n1478;
  wire _abc_43815_n1479;
  wire _abc_43815_n1480;
  wire _abc_43815_n1481;
  wire _abc_43815_n1482;
  wire _abc_43815_n1483;
  wire _abc_43815_n1484;
  wire _abc_43815_n1485;
  wire _abc_43815_n1486;
  wire _abc_43815_n1487;
  wire _abc_43815_n1488;
  wire _abc_43815_n1489;
  wire _abc_43815_n1489_bF_buf0;
  wire _abc_43815_n1489_bF_buf1;
  wire _abc_43815_n1489_bF_buf2;
  wire _abc_43815_n1489_bF_buf3;
  wire _abc_43815_n1489_bF_buf4;
  wire _abc_43815_n1490;
  wire _abc_43815_n1491_1;
  wire _abc_43815_n1492_1;
  wire _abc_43815_n1493;
  wire _abc_43815_n1494;
  wire _abc_43815_n1495;
  wire _abc_43815_n1496;
  wire _abc_43815_n1497;
  wire _abc_43815_n1498;
  wire _abc_43815_n1499;
  wire _abc_43815_n1500;
  wire _abc_43815_n1502;
  wire _abc_43815_n1503;
  wire _abc_43815_n1504;
  wire _abc_43815_n1505;
  wire _abc_43815_n1506;
  wire _abc_43815_n1507;
  wire _abc_43815_n1508;
  wire _abc_43815_n1509;
  wire _abc_43815_n1510;
  wire _abc_43815_n1511;
  wire _abc_43815_n1512;
  wire _abc_43815_n1513;
  wire _abc_43815_n1514;
  wire _abc_43815_n1515_1;
  wire _abc_43815_n1516;
  wire _abc_43815_n1517;
  wire _abc_43815_n1518_1;
  wire _abc_43815_n1519;
  wire _abc_43815_n1520;
  wire _abc_43815_n1521;
  wire _abc_43815_n1522;
  wire _abc_43815_n1523;
  wire _abc_43815_n1524;
  wire _abc_43815_n1525;
  wire _abc_43815_n1526;
  wire _abc_43815_n1527;
  wire _abc_43815_n1528;
  wire _abc_43815_n1529;
  wire _abc_43815_n1530;
  wire _abc_43815_n1531;
  wire _abc_43815_n1532;
  wire _abc_43815_n1533;
  wire _abc_43815_n1534_1;
  wire _abc_43815_n1535_1;
  wire _abc_43815_n1536;
  wire _abc_43815_n1538;
  wire _abc_43815_n1539;
  wire _abc_43815_n1540;
  wire _abc_43815_n1541;
  wire _abc_43815_n1542;
  wire _abc_43815_n1543;
  wire _abc_43815_n1544;
  wire _abc_43815_n1545;
  wire _abc_43815_n1546;
  wire _abc_43815_n1547_1;
  wire _abc_43815_n1548;
  wire _abc_43815_n1549;
  wire _abc_43815_n1550_1;
  wire _abc_43815_n1551;
  wire _abc_43815_n1552;
  wire _abc_43815_n1553;
  wire _abc_43815_n1554;
  wire _abc_43815_n1555;
  wire _abc_43815_n1556;
  wire _abc_43815_n1557;
  wire _abc_43815_n1558;
  wire _abc_43815_n1559;
  wire _abc_43815_n1560;
  wire _abc_43815_n1561;
  wire _abc_43815_n1562;
  wire _abc_43815_n1563;
  wire _abc_43815_n1564;
  wire _abc_43815_n1565;
  wire _abc_43815_n1566_1;
  wire _abc_43815_n1567_1;
  wire _abc_43815_n1568;
  wire _abc_43815_n1569;
  wire _abc_43815_n1570;
  wire _abc_43815_n1571;
  wire _abc_43815_n1572;
  wire _abc_43815_n1573;
  wire _abc_43815_n1575;
  wire _abc_43815_n1576;
  wire _abc_43815_n1577;
  wire _abc_43815_n1578;
  wire _abc_43815_n1579;
  wire _abc_43815_n1580;
  wire _abc_43815_n1581;
  wire _abc_43815_n1582;
  wire _abc_43815_n1583_1;
  wire _abc_43815_n1584;
  wire _abc_43815_n1585;
  wire _abc_43815_n1586_1;
  wire _abc_43815_n1587;
  wire _abc_43815_n1588;
  wire _abc_43815_n1589;
  wire _abc_43815_n1590;
  wire _abc_43815_n1591;
  wire _abc_43815_n1592;
  wire _abc_43815_n1593;
  wire _abc_43815_n1594;
  wire _abc_43815_n1595;
  wire _abc_43815_n1596;
  wire _abc_43815_n1597;
  wire _abc_43815_n1598;
  wire _abc_43815_n1599;
  wire _abc_43815_n1600;
  wire _abc_43815_n1601;
  wire _abc_43815_n1602_1;
  wire _abc_43815_n1603_1;
  wire _abc_43815_n1604;
  wire _abc_43815_n1605;
  wire _abc_43815_n1606;
  wire _abc_43815_n1607;
  wire _abc_43815_n1608;
  wire _abc_43815_n1609;
  wire _abc_43815_n1610;
  wire _abc_43815_n1611;
  wire _abc_43815_n1612;
  wire _abc_43815_n1613;
  wire _abc_43815_n1615_1;
  wire _abc_43815_n1616;
  wire _abc_43815_n1617;
  wire _abc_43815_n1618_1;
  wire _abc_43815_n1619;
  wire _abc_43815_n1620;
  wire _abc_43815_n1621;
  wire _abc_43815_n1622;
  wire _abc_43815_n1623;
  wire _abc_43815_n1624;
  wire _abc_43815_n1625;
  wire _abc_43815_n1626;
  wire _abc_43815_n1627;
  wire _abc_43815_n1628;
  wire _abc_43815_n1629;
  wire _abc_43815_n1630;
  wire _abc_43815_n1631;
  wire _abc_43815_n1632;
  wire _abc_43815_n1633;
  wire _abc_43815_n1634_1;
  wire _abc_43815_n1635_1;
  wire _abc_43815_n1636;
  wire _abc_43815_n1637;
  wire _abc_43815_n1638;
  wire _abc_43815_n1639;
  wire _abc_43815_n1640;
  wire _abc_43815_n1641;
  wire _abc_43815_n1642;
  wire _abc_43815_n1643;
  wire _abc_43815_n1644;
  wire _abc_43815_n1645;
  wire _abc_43815_n1646;
  wire _abc_43815_n1647;
  wire _abc_43815_n1648;
  wire _abc_43815_n1649;
  wire _abc_43815_n1651;
  wire _abc_43815_n1652;
  wire _abc_43815_n1653;
  wire _abc_43815_n1654;
  wire _abc_43815_n1655_1;
  wire _abc_43815_n1656;
  wire _abc_43815_n1657;
  wire _abc_43815_n1658_1;
  wire _abc_43815_n1659;
  wire _abc_43815_n1660;
  wire _abc_43815_n1661;
  wire _abc_43815_n1662;
  wire _abc_43815_n1663;
  wire _abc_43815_n1664;
  wire _abc_43815_n1665;
  wire _abc_43815_n1666;
  wire _abc_43815_n1667;
  wire _abc_43815_n1668;
  wire _abc_43815_n1669;
  wire _abc_43815_n1670;
  wire _abc_43815_n1671;
  wire _abc_43815_n1672;
  wire _abc_43815_n1673;
  wire _abc_43815_n1674_1;
  wire _abc_43815_n1675_1;
  wire _abc_43815_n1676;
  wire _abc_43815_n1677;
  wire _abc_43815_n1678;
  wire _abc_43815_n1679;
  wire _abc_43815_n1680;
  wire _abc_43815_n1681;
  wire _abc_43815_n1682;
  wire _abc_43815_n1683;
  wire _abc_43815_n1684;
  wire _abc_43815_n1685;
  wire _abc_43815_n1686_1;
  wire _abc_43815_n1687;
  wire _abc_43815_n1688;
  wire _abc_43815_n1689_1;
  wire _abc_43815_n1690;
  wire _abc_43815_n1692;
  wire _abc_43815_n1693;
  wire _abc_43815_n1694;
  wire _abc_43815_n1695;
  wire _abc_43815_n1696;
  wire _abc_43815_n1697;
  wire _abc_43815_n1698;
  wire _abc_43815_n1699;
  wire _abc_43815_n1700;
  wire _abc_43815_n1701;
  wire _abc_43815_n1702;
  wire _abc_43815_n1703;
  wire _abc_43815_n1704;
  wire _abc_43815_n1705_1;
  wire _abc_43815_n1706_1;
  wire _abc_43815_n1707;
  wire _abc_43815_n1708;
  wire _abc_43815_n1709;
  wire _abc_43815_n1710;
  wire _abc_43815_n1711;
  wire _abc_43815_n1712;
  wire _abc_43815_n1713;
  wire _abc_43815_n1714;
  wire _abc_43815_n1715;
  wire _abc_43815_n1716;
  wire _abc_43815_n1717;
  wire _abc_43815_n1718;
  wire _abc_43815_n1719_1;
  wire _abc_43815_n1720;
  wire _abc_43815_n1721;
  wire _abc_43815_n1722_1;
  wire _abc_43815_n1723;
  wire _abc_43815_n1724;
  wire _abc_43815_n1725;
  wire _abc_43815_n1726;
  wire _abc_43815_n1727;
  wire _abc_43815_n1728;
  wire _abc_43815_n1730;
  wire _abc_43815_n1731;
  wire _abc_43815_n1732;
  wire _abc_43815_n1733;
  wire _abc_43815_n1734;
  wire _abc_43815_n1735;
  wire _abc_43815_n1736;
  wire _abc_43815_n1737;
  wire _abc_43815_n1738_1;
  wire _abc_43815_n1739_1;
  wire _abc_43815_n1740;
  wire _abc_43815_n1741;
  wire _abc_43815_n1742;
  wire _abc_43815_n1743;
  wire _abc_43815_n1744;
  wire _abc_43815_n1745;
  wire _abc_43815_n1746;
  wire _abc_43815_n1747;
  wire _abc_43815_n1748;
  wire _abc_43815_n1749;
  wire _abc_43815_n1750_1;
  wire _abc_43815_n1751;
  wire _abc_43815_n1752;
  wire _abc_43815_n1753_1;
  wire _abc_43815_n1754;
  wire _abc_43815_n1755;
  wire _abc_43815_n1756;
  wire _abc_43815_n1757;
  wire _abc_43815_n1758;
  wire _abc_43815_n1759;
  wire _abc_43815_n1760;
  wire _abc_43815_n1761;
  wire _abc_43815_n1762;
  wire _abc_43815_n1763;
  wire _abc_43815_n1764;
  wire _abc_43815_n1765;
  wire _abc_43815_n1766;
  wire _abc_43815_n1767;
  wire _abc_43815_n1769_1;
  wire _abc_43815_n1770;
  wire _abc_43815_n1771;
  wire _abc_43815_n1772;
  wire _abc_43815_n1773;
  wire _abc_43815_n1774;
  wire _abc_43815_n1775_1;
  wire _abc_43815_n1776;
  wire _abc_43815_n1777;
  wire _abc_43815_n1778_1;
  wire _abc_43815_n1779;
  wire _abc_43815_n1780;
  wire _abc_43815_n1781_1;
  wire _abc_43815_n1782;
  wire _abc_43815_n1783;
  wire _abc_43815_n1784;
  wire _abc_43815_n1785_1;
  wire _abc_43815_n1786;
  wire _abc_43815_n1787;
  wire _abc_43815_n1788_1;
  wire _abc_43815_n1789;
  wire _abc_43815_n1790;
  wire _abc_43815_n1791_1;
  wire _abc_43815_n1792;
  wire _abc_43815_n1793;
  wire _abc_43815_n1794_1;
  wire _abc_43815_n1795;
  wire _abc_43815_n1796;
  wire _abc_43815_n1797_1;
  wire _abc_43815_n1798;
  wire _abc_43815_n1799;
  wire _abc_43815_n1800;
  wire _abc_43815_n1801;
  wire _abc_43815_n1802_1;
  wire _abc_43815_n1803;
  wire _abc_43815_n1804;
  wire _abc_43815_n1805;
  wire _abc_43815_n1806;
  wire _abc_43815_n1807;
  wire _abc_43815_n1808;
  wire _abc_43815_n1810_1;
  wire _abc_43815_n1811;
  wire _abc_43815_n1812;
  wire _abc_43815_n1813;
  wire _abc_43815_n1814;
  wire _abc_43815_n1815_1;
  wire _abc_43815_n1816;
  wire _abc_43815_n1817;
  wire _abc_43815_n1818;
  wire _abc_43815_n1819;
  wire _abc_43815_n1820_1;
  wire _abc_43815_n1821;
  wire _abc_43815_n1822;
  wire _abc_43815_n1823_1;
  wire _abc_43815_n1824;
  wire _abc_43815_n1825;
  wire _abc_43815_n1826_1;
  wire _abc_43815_n1827;
  wire _abc_43815_n1828;
  wire _abc_43815_n1829_1;
  wire _abc_43815_n1830;
  wire _abc_43815_n1831;
  wire _abc_43815_n1832_1;
  wire _abc_43815_n1833;
  wire _abc_43815_n1834;
  wire _abc_43815_n1835_1;
  wire _abc_43815_n1836;
  wire _abc_43815_n1837;
  wire _abc_43815_n1838_1;
  wire _abc_43815_n1839;
  wire _abc_43815_n1840;
  wire _abc_43815_n1841_1;
  wire _abc_43815_n1842;
  wire _abc_43815_n1843;
  wire _abc_43815_n1844_1;
  wire _abc_43815_n1846;
  wire _abc_43815_n1847_1;
  wire _abc_43815_n1848;
  wire _abc_43815_n1849;
  wire _abc_43815_n1850_1;
  wire _abc_43815_n1851;
  wire _abc_43815_n1852;
  wire _abc_43815_n1853_1;
  wire _abc_43815_n1854;
  wire _abc_43815_n1855;
  wire _abc_43815_n1856_1;
  wire _abc_43815_n1857;
  wire _abc_43815_n1858;
  wire _abc_43815_n1859_1;
  wire _abc_43815_n1860;
  wire _abc_43815_n1861;
  wire _abc_43815_n1862_1;
  wire _abc_43815_n1863;
  wire _abc_43815_n1864;
  wire _abc_43815_n1865_1;
  wire _abc_43815_n1866;
  wire _abc_43815_n1867;
  wire _abc_43815_n1868_1;
  wire _abc_43815_n1869;
  wire _abc_43815_n1870;
  wire _abc_43815_n1871_1;
  wire _abc_43815_n1872;
  wire _abc_43815_n1873;
  wire _abc_43815_n1874_1;
  wire _abc_43815_n1875;
  wire _abc_43815_n1876;
  wire _abc_43815_n1877_1;
  wire _abc_43815_n1878;
  wire _abc_43815_n1879;
  wire _abc_43815_n1880_1;
  wire _abc_43815_n1881;
  wire _abc_43815_n1882;
  wire _abc_43815_n1883;
  wire _abc_43815_n1884;
  wire _abc_43815_n1885;
  wire _abc_43815_n1886;
  wire _abc_43815_n1887;
  wire _abc_43815_n1888;
  wire _abc_43815_n1890;
  wire _abc_43815_n1891;
  wire _abc_43815_n1892;
  wire _abc_43815_n1893;
  wire _abc_43815_n1894;
  wire _abc_43815_n1895;
  wire _abc_43815_n1896;
  wire _abc_43815_n1897;
  wire _abc_43815_n1898;
  wire _abc_43815_n1899;
  wire _abc_43815_n1900;
  wire _abc_43815_n1901;
  wire _abc_43815_n1902;
  wire _abc_43815_n1903;
  wire _abc_43815_n1904;
  wire _abc_43815_n1905;
  wire _abc_43815_n1906;
  wire _abc_43815_n1907;
  wire _abc_43815_n1908;
  wire _abc_43815_n1909;
  wire _abc_43815_n1910;
  wire _abc_43815_n1911;
  wire _abc_43815_n1912;
  wire _abc_43815_n1913;
  wire _abc_43815_n1914;
  wire _abc_43815_n1915;
  wire _abc_43815_n1916;
  wire _abc_43815_n1917;
  wire _abc_43815_n1918_1;
  wire _abc_43815_n1919;
  wire _abc_43815_n1920_1;
  wire _abc_43815_n1921;
  wire _abc_43815_n1922_1;
  wire _abc_43815_n1923_1;
  wire _abc_43815_n1924;
  wire _abc_43815_n1925_1;
  wire _abc_43815_n1926;
  wire _abc_43815_n1927;
  wire _abc_43815_n1929;
  wire _abc_43815_n1930;
  wire _abc_43815_n1931;
  wire _abc_43815_n1932;
  wire _abc_43815_n1933;
  wire _abc_43815_n1934;
  wire _abc_43815_n1935;
  wire _abc_43815_n1936;
  wire _abc_43815_n1937;
  wire _abc_43815_n1938;
  wire _abc_43815_n1939;
  wire _abc_43815_n1940;
  wire _abc_43815_n1941;
  wire _abc_43815_n1942;
  wire _abc_43815_n1943;
  wire _abc_43815_n1944;
  wire _abc_43815_n1945;
  wire _abc_43815_n1946;
  wire _abc_43815_n1947;
  wire _abc_43815_n1948;
  wire _abc_43815_n1949;
  wire _abc_43815_n1950;
  wire _abc_43815_n1951;
  wire _abc_43815_n1952;
  wire _abc_43815_n1953;
  wire _abc_43815_n1954_1;
  wire _abc_43815_n1955;
  wire _abc_43815_n1956;
  wire _abc_43815_n1957;
  wire _abc_43815_n1958;
  wire _abc_43815_n1959;
  wire _abc_43815_n1960;
  wire _abc_43815_n1961;
  wire _abc_43815_n1962;
  wire _abc_43815_n1963;
  wire _abc_43815_n1964;
  wire _abc_43815_n1966;
  wire _abc_43815_n1967;
  wire _abc_43815_n1968;
  wire _abc_43815_n1969;
  wire _abc_43815_n1970;
  wire _abc_43815_n1971;
  wire _abc_43815_n1972;
  wire _abc_43815_n1973;
  wire _abc_43815_n1974_1;
  wire _abc_43815_n1975;
  wire _abc_43815_n1976;
  wire _abc_43815_n1977;
  wire _abc_43815_n1978;
  wire _abc_43815_n1979;
  wire _abc_43815_n1980;
  wire _abc_43815_n1981;
  wire _abc_43815_n1982;
  wire _abc_43815_n1983;
  wire _abc_43815_n1984;
  wire _abc_43815_n1985;
  wire _abc_43815_n1986;
  wire _abc_43815_n1987;
  wire _abc_43815_n1988;
  wire _abc_43815_n1989;
  wire _abc_43815_n1990;
  wire _abc_43815_n1991;
  wire _abc_43815_n1992;
  wire _abc_43815_n1993_1;
  wire _abc_43815_n1994;
  wire _abc_43815_n1995;
  wire _abc_43815_n1996;
  wire _abc_43815_n1997;
  wire _abc_43815_n1998;
  wire _abc_43815_n1999;
  wire _abc_43815_n2000;
  wire _abc_43815_n2002;
  wire _abc_43815_n2003;
  wire _abc_43815_n2004;
  wire _abc_43815_n2005;
  wire _abc_43815_n2006;
  wire _abc_43815_n2007;
  wire _abc_43815_n2008;
  wire _abc_43815_n2009;
  wire _abc_43815_n2010;
  wire _abc_43815_n2011;
  wire _abc_43815_n2012;
  wire _abc_43815_n2013_1;
  wire _abc_43815_n2014;
  wire _abc_43815_n2015;
  wire _abc_43815_n2016;
  wire _abc_43815_n2017;
  wire _abc_43815_n2018;
  wire _abc_43815_n2019;
  wire _abc_43815_n2020;
  wire _abc_43815_n2021;
  wire _abc_43815_n2022;
  wire _abc_43815_n2023;
  wire _abc_43815_n2024;
  wire _abc_43815_n2025;
  wire _abc_43815_n2026;
  wire _abc_43815_n2027;
  wire _abc_43815_n2028;
  wire _abc_43815_n2029;
  wire _abc_43815_n2030;
  wire _abc_43815_n2031;
  wire _abc_43815_n2032;
  wire _abc_43815_n2033;
  wire _abc_43815_n2034_1;
  wire _abc_43815_n2035;
  wire _abc_43815_n2036;
  wire _abc_43815_n2037;
  wire _abc_43815_n2038;
  wire _abc_43815_n2039;
  wire _abc_43815_n2040;
  wire _abc_43815_n2041;
  wire _abc_43815_n2042;
  wire _abc_43815_n2043;
  wire _abc_43815_n2044;
  wire _abc_43815_n2045;
  wire _abc_43815_n2047;
  wire _abc_43815_n2048;
  wire _abc_43815_n2049;
  wire _abc_43815_n2050;
  wire _abc_43815_n2051;
  wire _abc_43815_n2052;
  wire _abc_43815_n2053;
  wire _abc_43815_n2054;
  wire _abc_43815_n2055_1;
  wire _abc_43815_n2056;
  wire _abc_43815_n2057;
  wire _abc_43815_n2058;
  wire _abc_43815_n2059;
  wire _abc_43815_n2060;
  wire _abc_43815_n2061;
  wire _abc_43815_n2062;
  wire _abc_43815_n2063;
  wire _abc_43815_n2064;
  wire _abc_43815_n2065;
  wire _abc_43815_n2066;
  wire _abc_43815_n2067;
  wire _abc_43815_n2068;
  wire _abc_43815_n2069;
  wire _abc_43815_n2070;
  wire _abc_43815_n2071;
  wire _abc_43815_n2072;
  wire _abc_43815_n2073_1;
  wire _abc_43815_n2074;
  wire _abc_43815_n2075;
  wire _abc_43815_n2076;
  wire _abc_43815_n2077;
  wire _abc_43815_n2078;
  wire _abc_43815_n2079;
  wire _abc_43815_n2080;
  wire _abc_43815_n2081;
  wire _abc_43815_n2082;
  wire _abc_43815_n2083;
  wire _abc_43815_n2084;
  wire _abc_43815_n2086;
  wire _abc_43815_n2087_1;
  wire _abc_43815_n2088;
  wire _abc_43815_n2089;
  wire _abc_43815_n2090;
  wire _abc_43815_n2091;
  wire _abc_43815_n2092;
  wire _abc_43815_n2093;
  wire _abc_43815_n2094;
  wire _abc_43815_n2095;
  wire _abc_43815_n2096;
  wire _abc_43815_n2097;
  wire _abc_43815_n2098;
  wire _abc_43815_n2099;
  wire _abc_43815_n2100;
  wire _abc_43815_n2101_1;
  wire _abc_43815_n2102;
  wire _abc_43815_n2103;
  wire _abc_43815_n2104;
  wire _abc_43815_n2105;
  wire _abc_43815_n2106;
  wire _abc_43815_n2107;
  wire _abc_43815_n2108;
  wire _abc_43815_n2109;
  wire _abc_43815_n2110;
  wire _abc_43815_n2111;
  wire _abc_43815_n2112;
  wire _abc_43815_n2113;
  wire _abc_43815_n2114;
  wire _abc_43815_n2115_1;
  wire _abc_43815_n2116;
  wire _abc_43815_n2117;
  wire _abc_43815_n2118;
  wire _abc_43815_n2119;
  wire _abc_43815_n2120;
  wire _abc_43815_n2121;
  wire _abc_43815_n2123;
  wire _abc_43815_n2124;
  wire _abc_43815_n2125;
  wire _abc_43815_n2126;
  wire _abc_43815_n2127;
  wire _abc_43815_n2128;
  wire _abc_43815_n2129_1;
  wire _abc_43815_n2130;
  wire _abc_43815_n2131;
  wire _abc_43815_n2132;
  wire _abc_43815_n2133;
  wire _abc_43815_n2134;
  wire _abc_43815_n2135;
  wire _abc_43815_n2136;
  wire _abc_43815_n2137;
  wire _abc_43815_n2138;
  wire _abc_43815_n2139;
  wire _abc_43815_n2140;
  wire _abc_43815_n2141;
  wire _abc_43815_n2142;
  wire _abc_43815_n2143_1;
  wire _abc_43815_n2144;
  wire _abc_43815_n2145;
  wire _abc_43815_n2146;
  wire _abc_43815_n2147;
  wire _abc_43815_n2148;
  wire _abc_43815_n2149;
  wire _abc_43815_n2150;
  wire _abc_43815_n2151;
  wire _abc_43815_n2152;
  wire _abc_43815_n2153;
  wire _abc_43815_n2154;
  wire _abc_43815_n2155;
  wire _abc_43815_n2156;
  wire _abc_43815_n2157;
  wire _abc_43815_n2159;
  wire _abc_43815_n2160;
  wire _abc_43815_n2161;
  wire _abc_43815_n2162;
  wire _abc_43815_n2163;
  wire _abc_43815_n2164;
  wire _abc_43815_n2165;
  wire _abc_43815_n2166;
  wire _abc_43815_n2167;
  wire _abc_43815_n2168;
  wire _abc_43815_n2169;
  wire _abc_43815_n2170;
  wire _abc_43815_n2171;
  wire _abc_43815_n2172;
  wire _abc_43815_n2173_1;
  wire _abc_43815_n2174;
  wire _abc_43815_n2175;
  wire _abc_43815_n2176;
  wire _abc_43815_n2177;
  wire _abc_43815_n2178;
  wire _abc_43815_n2179;
  wire _abc_43815_n2180;
  wire _abc_43815_n2181;
  wire _abc_43815_n2182;
  wire _abc_43815_n2183;
  wire _abc_43815_n2184;
  wire _abc_43815_n2185;
  wire _abc_43815_n2186;
  wire _abc_43815_n2187;
  wire _abc_43815_n2188_1;
  wire _abc_43815_n2189;
  wire _abc_43815_n2190;
  wire _abc_43815_n2191;
  wire _abc_43815_n2192;
  wire _abc_43815_n2193;
  wire _abc_43815_n2194;
  wire _abc_43815_n2195;
  wire _abc_43815_n2196;
  wire _abc_43815_n2197;
  wire _abc_43815_n2198;
  wire _abc_43815_n2199;
  wire _abc_43815_n2200;
  wire _abc_43815_n2202;
  wire _abc_43815_n2203_1;
  wire _abc_43815_n2204;
  wire _abc_43815_n2205;
  wire _abc_43815_n2206;
  wire _abc_43815_n2207;
  wire _abc_43815_n2208;
  wire _abc_43815_n2209;
  wire _abc_43815_n2210;
  wire _abc_43815_n2211;
  wire _abc_43815_n2212;
  wire _abc_43815_n2213;
  wire _abc_43815_n2214;
  wire _abc_43815_n2215;
  wire _abc_43815_n2216;
  wire _abc_43815_n2217;
  wire _abc_43815_n2218;
  wire _abc_43815_n2219;
  wire _abc_43815_n2220;
  wire _abc_43815_n2221;
  wire _abc_43815_n2222_1;
  wire _abc_43815_n2223;
  wire _abc_43815_n2224;
  wire _abc_43815_n2225;
  wire _abc_43815_n2226;
  wire _abc_43815_n2227;
  wire _abc_43815_n2228;
  wire _abc_43815_n2229;
  wire _abc_43815_n2230;
  wire _abc_43815_n2231;
  wire _abc_43815_n2232_1;
  wire _abc_43815_n2233;
  wire _abc_43815_n2234;
  wire _abc_43815_n2235;
  wire _abc_43815_n2236;
  wire _abc_43815_n2237;
  wire _abc_43815_n2238;
  wire _abc_43815_n2240;
  wire _abc_43815_n2241;
  wire _abc_43815_n2242_1;
  wire _abc_43815_n2243;
  wire _abc_43815_n2244;
  wire _abc_43815_n2245;
  wire _abc_43815_n2246;
  wire _abc_43815_n2247;
  wire _abc_43815_n2248;
  wire _abc_43815_n2249;
  wire _abc_43815_n2250;
  wire _abc_43815_n2251;
  wire _abc_43815_n2252_1;
  wire _abc_43815_n2253;
  wire _abc_43815_n2254;
  wire _abc_43815_n2255;
  wire _abc_43815_n2256;
  wire _abc_43815_n2257;
  wire _abc_43815_n2258;
  wire _abc_43815_n2259;
  wire _abc_43815_n2260;
  wire _abc_43815_n2261;
  wire _abc_43815_n2262_1;
  wire _abc_43815_n2263;
  wire _abc_43815_n2264;
  wire _abc_43815_n2265;
  wire _abc_43815_n2266;
  wire _abc_43815_n2267;
  wire _abc_43815_n2268;
  wire _abc_43815_n2269;
  wire _abc_43815_n2270;
  wire _abc_43815_n2271;
  wire _abc_43815_n2272_1;
  wire _abc_43815_n2273;
  wire _abc_43815_n2274;
  wire _abc_43815_n2276;
  wire _abc_43815_n2277;
  wire _abc_43815_n2278;
  wire _abc_43815_n2279;
  wire _abc_43815_n2280;
  wire _abc_43815_n2281;
  wire _abc_43815_n2282_1;
  wire _abc_43815_n2283;
  wire _abc_43815_n2284;
  wire _abc_43815_n2285;
  wire _abc_43815_n2286;
  wire _abc_43815_n2287;
  wire _abc_43815_n2288;
  wire _abc_43815_n2289;
  wire _abc_43815_n2290;
  wire _abc_43815_n2291;
  wire _abc_43815_n2292_1;
  wire _abc_43815_n2293;
  wire _abc_43815_n2294;
  wire _abc_43815_n2295;
  wire _abc_43815_n2296;
  wire _abc_43815_n2297;
  wire _abc_43815_n2298;
  wire _abc_43815_n2299;
  wire _abc_43815_n2300;
  wire _abc_43815_n2301;
  wire _abc_43815_n2302_1;
  wire _abc_43815_n2303;
  wire _abc_43815_n2304;
  wire _abc_43815_n2305;
  wire _abc_43815_n2306;
  wire _abc_43815_n2307;
  wire _abc_43815_n2308;
  wire _abc_43815_n2309;
  wire _abc_43815_n2310;
  wire _abc_43815_n2312_1;
  wire _abc_43815_n2313;
  wire _abc_43815_n2314;
  wire _abc_43815_n2315;
  wire _abc_43815_n2316;
  wire _abc_43815_n2317;
  wire _abc_43815_n2318;
  wire _abc_43815_n2319;
  wire _abc_43815_n2320;
  wire _abc_43815_n2321;
  wire _abc_43815_n2322_1;
  wire _abc_43815_n2323;
  wire _abc_43815_n2324;
  wire _abc_43815_n2325;
  wire _abc_43815_n2326;
  wire _abc_43815_n2327;
  wire _abc_43815_n2328;
  wire _abc_43815_n2329;
  wire _abc_43815_n2330;
  wire _abc_43815_n2331;
  wire _abc_43815_n2332_1;
  wire _abc_43815_n2333;
  wire _abc_43815_n2334;
  wire _abc_43815_n2335;
  wire _abc_43815_n2336;
  wire _abc_43815_n2337;
  wire _abc_43815_n2338;
  wire _abc_43815_n2339;
  wire _abc_43815_n2340;
  wire _abc_43815_n2341;
  wire _abc_43815_n2342_1;
  wire _abc_43815_n2343;
  wire _abc_43815_n2344;
  wire _abc_43815_n2345;
  wire _abc_43815_n2346;
  wire _abc_43815_n2347;
  wire _abc_43815_n2348;
  wire _abc_43815_n2349;
  wire _abc_43815_n2350;
  wire _abc_43815_n2351;
  wire _abc_43815_n2352_1;
  wire _abc_43815_n2353;
  wire _abc_43815_n2355;
  wire _abc_43815_n2356;
  wire _abc_43815_n2357;
  wire _abc_43815_n2358;
  wire _abc_43815_n2359;
  wire _abc_43815_n2360;
  wire _abc_43815_n2361;
  wire _abc_43815_n2362_1;
  wire _abc_43815_n2363;
  wire _abc_43815_n2364;
  wire _abc_43815_n2365;
  wire _abc_43815_n2366;
  wire _abc_43815_n2367;
  wire _abc_43815_n2368;
  wire _abc_43815_n2369;
  wire _abc_43815_n2370;
  wire _abc_43815_n2371;
  wire _abc_43815_n2372_1;
  wire _abc_43815_n2373;
  wire _abc_43815_n2374;
  wire _abc_43815_n2375;
  wire _abc_43815_n2376;
  wire _abc_43815_n2377;
  wire _abc_43815_n2378;
  wire _abc_43815_n2379;
  wire _abc_43815_n2380;
  wire _abc_43815_n2381;
  wire _abc_43815_n2382;
  wire _abc_43815_n2383;
  wire _abc_43815_n2384;
  wire _abc_43815_n2385;
  wire _abc_43815_n2386;
  wire _abc_43815_n2387;
  wire _abc_43815_n2388;
  wire _abc_43815_n2389;
  wire _abc_43815_n2390;
  wire _abc_43815_n2391;
  wire _abc_43815_n2392;
  wire _abc_43815_n2394;
  wire _abc_43815_n2395;
  wire _abc_43815_n2396_1;
  wire _abc_43815_n2397;
  wire _abc_43815_n2398;
  wire _abc_43815_n2399;
  wire _abc_43815_n2400;
  wire _abc_43815_n2401;
  wire _abc_43815_n2402;
  wire _abc_43815_n2403;
  wire _abc_43815_n2404;
  wire _abc_43815_n2405;
  wire _abc_43815_n2406;
  wire _abc_43815_n2407;
  wire _abc_43815_n2408;
  wire _abc_43815_n2409;
  wire _abc_43815_n2410;
  wire _abc_43815_n2411;
  wire _abc_43815_n2412;
  wire _abc_43815_n2413;
  wire _abc_43815_n2414;
  wire _abc_43815_n2415;
  wire _abc_43815_n2416;
  wire _abc_43815_n2417;
  wire _abc_43815_n2418;
  wire _abc_43815_n2419;
  wire _abc_43815_n2420_1;
  wire _abc_43815_n2421;
  wire _abc_43815_n2422;
  wire _abc_43815_n2423;
  wire _abc_43815_n2424;
  wire _abc_43815_n2425;
  wire _abc_43815_n2426;
  wire _abc_43815_n2427;
  wire _abc_43815_n2428;
  wire _abc_43815_n2429;
  wire _abc_43815_n2431;
  wire _abc_43815_n2432;
  wire _abc_43815_n2433;
  wire _abc_43815_n2434;
  wire _abc_43815_n2435;
  wire _abc_43815_n2436;
  wire _abc_43815_n2437;
  wire _abc_43815_n2438;
  wire _abc_43815_n2439;
  wire _abc_43815_n2440;
  wire _abc_43815_n2441;
  wire _abc_43815_n2442;
  wire _abc_43815_n2443;
  wire _abc_43815_n2444;
  wire _abc_43815_n2445_1;
  wire _abc_43815_n2446;
  wire _abc_43815_n2447;
  wire _abc_43815_n2448;
  wire _abc_43815_n2449;
  wire _abc_43815_n2450;
  wire _abc_43815_n2451;
  wire _abc_43815_n2452;
  wire _abc_43815_n2453;
  wire _abc_43815_n2454;
  wire _abc_43815_n2455;
  wire _abc_43815_n2456;
  wire _abc_43815_n2457;
  wire _abc_43815_n2458;
  wire _abc_43815_n2459;
  wire _abc_43815_n2460;
  wire _abc_43815_n2461;
  wire _abc_43815_n2462;
  wire _abc_43815_n2463;
  wire _abc_43815_n2464;
  wire _abc_43815_n2465;
  wire _abc_43815_n2466;
  wire _abc_43815_n2467;
  wire _abc_43815_n2468;
  wire _abc_43815_n2470;
  wire _abc_43815_n2471;
  wire _abc_43815_n2472;
  wire _abc_43815_n2473;
  wire _abc_43815_n2474;
  wire _abc_43815_n2475;
  wire _abc_43815_n2476;
  wire _abc_43815_n2477;
  wire _abc_43815_n2478;
  wire _abc_43815_n2479;
  wire _abc_43815_n2480;
  wire _abc_43815_n2481;
  wire _abc_43815_n2482;
  wire _abc_43815_n2483;
  wire _abc_43815_n2484;
  wire _abc_43815_n2485;
  wire _abc_43815_n2486;
  wire _abc_43815_n2487;
  wire _abc_43815_n2488;
  wire _abc_43815_n2489;
  wire _abc_43815_n2490;
  wire _abc_43815_n2491;
  wire _abc_43815_n2492;
  wire _abc_43815_n2493_1;
  wire _abc_43815_n2494;
  wire _abc_43815_n2495;
  wire _abc_43815_n2496;
  wire _abc_43815_n2497;
  wire _abc_43815_n2498;
  wire _abc_43815_n2499;
  wire _abc_43815_n2500;
  wire _abc_43815_n2501;
  wire _abc_43815_n2502;
  wire _abc_43815_n2503;
  wire _abc_43815_n2504;
  wire _abc_43815_n2505;
  wire _abc_43815_n2506;
  wire _abc_43815_n2507;
  wire _abc_43815_n2508;
  wire _abc_43815_n2509;
  wire _abc_43815_n2511;
  wire _abc_43815_n2512;
  wire _abc_43815_n2513;
  wire _abc_43815_n2514;
  wire _abc_43815_n2515;
  wire _abc_43815_n2516;
  wire _abc_43815_n2517_1;
  wire _abc_43815_n2518;
  wire _abc_43815_n2519;
  wire _abc_43815_n2520;
  wire _abc_43815_n2521;
  wire _abc_43815_n2522;
  wire _abc_43815_n2523;
  wire _abc_43815_n2524;
  wire _abc_43815_n2525;
  wire _abc_43815_n2526;
  wire _abc_43815_n2527;
  wire _abc_43815_n2528;
  wire _abc_43815_n2529;
  wire _abc_43815_n2530;
  wire _abc_43815_n2531;
  wire _abc_43815_n2532;
  wire _abc_43815_n2533;
  wire _abc_43815_n2534;
  wire _abc_43815_n2535;
  wire _abc_43815_n2536;
  wire _abc_43815_n2537;
  wire _abc_43815_n2538;
  wire _abc_43815_n2539;
  wire _abc_43815_n2540;
  wire _abc_43815_n2541_1;
  wire _abc_43815_n2542;
  wire _abc_43815_n2543;
  wire _abc_43815_n2544;
  wire _abc_43815_n2545;
  wire _abc_43815_n2547;
  wire _abc_43815_n2548;
  wire _abc_43815_n2549;
  wire _abc_43815_n2550;
  wire _abc_43815_n2551;
  wire _abc_43815_n2552;
  wire _abc_43815_n2553;
  wire _abc_43815_n2554;
  wire _abc_43815_n2555;
  wire _abc_43815_n2556;
  wire _abc_43815_n2557;
  wire _abc_43815_n2558;
  wire _abc_43815_n2559;
  wire _abc_43815_n2560;
  wire _abc_43815_n2561;
  wire _abc_43815_n2562;
  wire _abc_43815_n2563;
  wire _abc_43815_n2564;
  wire _abc_43815_n2565_1;
  wire _abc_43815_n2566;
  wire _abc_43815_n2567;
  wire _abc_43815_n2568;
  wire _abc_43815_n2569;
  wire _abc_43815_n2570;
  wire _abc_43815_n2571;
  wire _abc_43815_n2572;
  wire _abc_43815_n2573;
  wire _abc_43815_n2574;
  wire _abc_43815_n2575;
  wire _abc_43815_n2576;
  wire _abc_43815_n2577;
  wire _abc_43815_n2578;
  wire _abc_43815_n2579;
  wire _abc_43815_n2580;
  wire _abc_43815_n2581;
  wire _abc_43815_n2582;
  wire _abc_43815_n2583;
  wire _abc_43815_n2584;
  wire _abc_43815_n2586;
  wire _abc_43815_n2587;
  wire _abc_43815_n2588;
  wire _abc_43815_n2589_1;
  wire _abc_43815_n2590;
  wire _abc_43815_n2591;
  wire _abc_43815_n2592;
  wire _abc_43815_n2593;
  wire _abc_43815_n2594;
  wire _abc_43815_n2595;
  wire _abc_43815_n2596;
  wire _abc_43815_n2597;
  wire _abc_43815_n2598;
  wire _abc_43815_n2599;
  wire _abc_43815_n2600;
  wire _abc_43815_n2601;
  wire _abc_43815_n2602;
  wire _abc_43815_n2603;
  wire _abc_43815_n2604;
  wire _abc_43815_n2605;
  wire _abc_43815_n2606;
  wire _abc_43815_n2607;
  wire _abc_43815_n2608;
  wire _abc_43815_n2609;
  wire _abc_43815_n2610;
  wire _abc_43815_n2611;
  wire _abc_43815_n2612;
  wire _abc_43815_n2613;
  wire _abc_43815_n2614_1;
  wire _abc_43815_n2615;
  wire _abc_43815_n2616;
  wire _abc_43815_n2617;
  wire _abc_43815_n2618;
  wire _abc_43815_n2619;
  wire _abc_43815_n2620;
  wire _abc_43815_n2622;
  wire _abc_43815_n2623;
  wire _abc_43815_n2624;
  wire _abc_43815_n2626;
  wire _abc_43815_n2627;
  wire _abc_43815_n2628;
  wire _abc_43815_n2630;
  wire _abc_43815_n2631;
  wire _abc_43815_n2632;
  wire _abc_43815_n2634;
  wire _abc_43815_n2635;
  wire _abc_43815_n2636;
  wire _abc_43815_n2638_1;
  wire _abc_43815_n2639;
  wire _abc_43815_n2640;
  wire _abc_43815_n2642;
  wire _abc_43815_n2643;
  wire _abc_43815_n2644;
  wire _abc_43815_n2646;
  wire _abc_43815_n2647;
  wire _abc_43815_n2648;
  wire _abc_43815_n2650;
  wire _abc_43815_n2651;
  wire _abc_43815_n2652;
  wire _abc_43815_n2654;
  wire _abc_43815_n2655;
  wire _abc_43815_n2656;
  wire _abc_43815_n2657;
  wire _abc_43815_n2658;
  wire _abc_43815_n2660;
  wire _abc_43815_n2661;
  wire _abc_43815_n2662_1;
  wire _abc_43815_n2663;
  wire _abc_43815_n2664;
  wire _abc_43815_n2665;
  wire _abc_43815_n2666;
  wire _abc_43815_n2668;
  wire _abc_43815_n2669;
  wire _abc_43815_n2670;
  wire _abc_43815_n2671;
  wire _abc_43815_n2672;
  wire _abc_43815_n2674;
  wire _abc_43815_n2675;
  wire _abc_43815_n2676;
  wire _abc_43815_n2677;
  wire _abc_43815_n2678;
  wire _abc_43815_n2679;
  wire _abc_43815_n2680;
  wire _abc_43815_n2682;
  wire _abc_43815_n2683;
  wire _abc_43815_n2684;
  wire _abc_43815_n2686_1;
  wire _abc_43815_n2687;
  wire _abc_43815_n2688;
  wire _abc_43815_n2690;
  wire _abc_43815_n2691;
  wire _abc_43815_n2692;
  wire _abc_43815_n2694;
  wire _abc_43815_n2695;
  wire _abc_43815_n2696;
  wire _abc_43815_n2698;
  wire _abc_43815_n2699;
  wire _abc_43815_n2700;
  wire _abc_43815_n2702;
  wire _abc_43815_n2703;
  wire _abc_43815_n2704;
  wire _abc_43815_n2706;
  wire _abc_43815_n2707;
  wire _abc_43815_n2708;
  wire _abc_43815_n2710_1;
  wire _abc_43815_n2711;
  wire _abc_43815_n2712;
  wire _abc_43815_n2714;
  wire _abc_43815_n2715;
  wire _abc_43815_n2716;
  wire _abc_43815_n2718;
  wire _abc_43815_n2719;
  wire _abc_43815_n2720;
  wire _abc_43815_n2722;
  wire _abc_43815_n2723;
  wire _abc_43815_n2724;
  wire _abc_43815_n2726;
  wire _abc_43815_n2727;
  wire _abc_43815_n2728;
  wire _abc_43815_n2730;
  wire _abc_43815_n2731;
  wire _abc_43815_n2732;
  wire _abc_43815_n2734_1;
  wire _abc_43815_n2735;
  wire _abc_43815_n2736;
  wire _abc_43815_n2738;
  wire _abc_43815_n2739;
  wire _abc_43815_n2740;
  wire _abc_43815_n2742;
  wire _abc_43815_n2743;
  wire _abc_43815_n2744;
  wire _abc_43815_n2746;
  wire _abc_43815_n2747;
  wire _abc_43815_n2748;
  wire _abc_43815_n2750;
  wire _abc_43815_n2751;
  wire _abc_43815_n2752;
  wire _abc_43815_n2754;
  wire _abc_43815_n2755;
  wire _abc_43815_n2756;
  wire _abc_43815_n2758_1;
  wire _abc_43815_n2759_1;
  wire _abc_43815_n2760;
  wire _abc_43815_n2762;
  wire _abc_43815_n2763;
  wire _abc_43815_n2764;
  wire _abc_43815_n2765;
  wire _abc_43815_n2766;
  wire _abc_43815_n2767;
  wire _abc_43815_n2768;
  wire _abc_43815_n2769;
  wire _abc_43815_n2770;
  wire _abc_43815_n2771;
  wire _abc_43815_n2772;
  wire _abc_43815_n2773;
  wire _abc_43815_n2774;
  wire _abc_43815_n2775;
  wire _abc_43815_n2776;
  wire _abc_43815_n2777;
  wire _abc_43815_n2778;
  wire _abc_43815_n2779;
  wire _abc_43815_n2780;
  wire _abc_43815_n2781;
  wire _abc_43815_n2782;
  wire _abc_43815_n2783;
  wire _abc_43815_n2784_1;
  wire _abc_43815_n2785_1;
  wire _abc_43815_n2786;
  wire _abc_43815_n2787;
  wire _abc_43815_n2788;
  wire _abc_43815_n2789;
  wire _abc_43815_n2790;
  wire _abc_43815_n2791;
  wire _abc_43815_n2792;
  wire _abc_43815_n2793;
  wire _abc_43815_n2794;
  wire _abc_43815_n2795;
  wire _abc_43815_n2796;
  wire _abc_43815_n2797;
  wire _abc_43815_n2798;
  wire _abc_43815_n2799;
  wire _abc_43815_n2801;
  wire _abc_43815_n2803;
  wire _abc_43815_n2805;
  wire _abc_43815_n2807;
  wire _abc_43815_n2809;
  wire _abc_43815_n2810_1;
  wire _abc_43815_n2811_1;
  wire _abc_43815_n2812;
  wire _abc_43815_n2813;
  wire _abc_43815_n2814;
  wire _abc_43815_n2815;
  wire _abc_43815_n2816;
  wire _abc_43815_n2817;
  wire _abc_43815_n2818;
  wire _abc_43815_n2819;
  wire _abc_43815_n2821;
  wire _abc_43815_n2822;
  wire _abc_43815_n2824;
  wire _abc_43815_n2825;
  wire _abc_43815_n2827;
  wire _abc_43815_n2828;
  wire _abc_43815_n2830;
  wire _abc_43815_n2831;
  wire _abc_43815_n2833;
  wire _abc_43815_n2834;
  wire _abc_43815_n2836_1;
  wire _abc_43815_n2837_1;
  wire _abc_43815_n2838;
  wire _abc_43815_n2839;
  wire _abc_43815_n2840;
  wire _abc_43815_n2840_bF_buf0;
  wire _abc_43815_n2840_bF_buf1;
  wire _abc_43815_n2840_bF_buf2;
  wire _abc_43815_n2840_bF_buf3;
  wire _abc_43815_n2840_bF_buf4;
  wire _abc_43815_n2841;
  wire _abc_43815_n2843;
  wire _abc_43815_n2844;
  wire _abc_43815_n2845;
  wire _abc_43815_n2846;
  wire _abc_43815_n2848;
  wire _abc_43815_n2849;
  wire _abc_43815_n2850;
  wire _abc_43815_n2851;
  wire _abc_43815_n2853;
  wire _abc_43815_n2854;
  wire _abc_43815_n2855;
  wire _abc_43815_n2856;
  wire _abc_43815_n2858;
  wire _abc_43815_n2859;
  wire _abc_43815_n2860;
  wire _abc_43815_n2861;
  wire _abc_43815_n2863_1;
  wire _abc_43815_n2864;
  wire _abc_43815_n2865;
  wire _abc_43815_n2866;
  wire _abc_43815_n2868;
  wire _abc_43815_n2869;
  wire _abc_43815_n2870;
  wire _abc_43815_n2871;
  wire _abc_43815_n2873;
  wire _abc_43815_n2874;
  wire _abc_43815_n2875;
  wire _abc_43815_n2876;
  wire _abc_43815_n2878;
  wire _abc_43815_n2879;
  wire _abc_43815_n2880;
  wire _abc_43815_n2881;
  wire _abc_43815_n2883;
  wire _abc_43815_n2884;
  wire _abc_43815_n2885;
  wire _abc_43815_n2886;
  wire _abc_43815_n2888_1;
  wire _abc_43815_n2889_1;
  wire _abc_43815_n2890;
  wire _abc_43815_n2891;
  wire _abc_43815_n2892;
  wire _abc_43815_n2893;
  wire _abc_43815_n2894;
  wire _abc_43815_n2895;
  wire _abc_43815_n2896;
  wire _abc_43815_n2897;
  wire _abc_43815_n2899;
  wire _abc_43815_n2900;
  wire _abc_43815_n2901;
  wire _abc_43815_n2902;
  wire _abc_43815_n2903;
  wire _abc_43815_n2905;
  wire _abc_43815_n2906;
  wire _abc_43815_n2907;
  wire _abc_43815_n2908;
  wire _abc_43815_n2909;
  wire _abc_43815_n2911;
  wire _abc_43815_n2912;
  wire _abc_43815_n2913;
  wire _abc_43815_n2914_1;
  wire _abc_43815_n2915_1;
  wire _abc_43815_n2917;
  wire _abc_43815_n2918;
  wire _abc_43815_n2919;
  wire _abc_43815_n2920;
  wire _abc_43815_n2921;
  wire _abc_43815_n2923;
  wire _abc_43815_n2924;
  wire _abc_43815_n2925;
  wire _abc_43815_n2926;
  wire _abc_43815_n2927;
  wire _abc_43815_n2929;
  wire _abc_43815_n2930;
  wire _abc_43815_n2931;
  wire _abc_43815_n2932;
  wire _abc_43815_n2933;
  wire _abc_43815_n2935;
  wire _abc_43815_n2936;
  wire _abc_43815_n2937;
  wire _abc_43815_n2938;
  wire _abc_43815_n2939;
  wire _abc_43815_n2941_1;
  wire _abc_43815_n2942;
  wire _abc_43815_n2943;
  wire _abc_43815_n2944;
  wire _abc_43815_n2945;
  wire _abc_43815_n2947;
  wire _abc_43815_n2948;
  wire _abc_43815_n2949;
  wire _abc_43815_n2950;
  wire _abc_43815_n2951;
  wire _abc_43815_n2953;
  wire _abc_43815_n2954;
  wire _abc_43815_n2955;
  wire _abc_43815_n2956;
  wire _abc_43815_n2957;
  wire _abc_43815_n2959;
  wire _abc_43815_n2960;
  wire _abc_43815_n2961;
  wire _abc_43815_n2962;
  wire _abc_43815_n2963;
  wire _abc_43815_n2965;
  wire _abc_43815_n2966_1;
  wire _abc_43815_n2967_1;
  wire _abc_43815_n2968;
  wire _abc_43815_n2969;
  wire _abc_43815_n2971;
  wire _abc_43815_n2972;
  wire _abc_43815_n2973;
  wire _abc_43815_n2974;
  wire _abc_43815_n2975;
  wire _abc_43815_n2977;
  wire _abc_43815_n2978;
  wire _abc_43815_n2979;
  wire _abc_43815_n2980;
  wire _abc_43815_n2981;
  wire _abc_43815_n2983;
  wire _abc_43815_n2984;
  wire _abc_43815_n2985;
  wire _abc_43815_n2986;
  wire _abc_43815_n2987;
  wire _abc_43815_n2989;
  wire _abc_43815_n2990;
  wire _abc_43815_n2991;
  wire _abc_43815_n2991_bF_buf0;
  wire _abc_43815_n2991_bF_buf1;
  wire _abc_43815_n2991_bF_buf2;
  wire _abc_43815_n2991_bF_buf3;
  wire _abc_43815_n2991_bF_buf4;
  wire _abc_43815_n2992_1;
  wire _abc_43815_n2993_1;
  wire _abc_43815_n2993_1_bF_buf0;
  wire _abc_43815_n2993_1_bF_buf1;
  wire _abc_43815_n2993_1_bF_buf2;
  wire _abc_43815_n2993_1_bF_buf3;
  wire _abc_43815_n2993_1_bF_buf4;
  wire _abc_43815_n2994;
  wire _abc_43815_n2995;
  wire _abc_43815_n2996;
  wire _abc_43815_n2997;
  wire _abc_43815_n2998;
  wire _abc_43815_n2999;
  wire _abc_43815_n3001;
  wire _abc_43815_n3002;
  wire _abc_43815_n3002_bF_buf0;
  wire _abc_43815_n3002_bF_buf1;
  wire _abc_43815_n3002_bF_buf2;
  wire _abc_43815_n3002_bF_buf3;
  wire _abc_43815_n3002_bF_buf4;
  wire _abc_43815_n3003;
  wire _abc_43815_n3005;
  wire _abc_43815_n3006;
  wire _abc_43815_n3007;
  wire _abc_43815_n3008;
  wire _abc_43815_n3009;
  wire _abc_43815_n3010;
  wire _abc_43815_n3011;
  wire _abc_43815_n3012;
  wire _abc_43815_n3014;
  wire _abc_43815_n3015;
  wire _abc_43815_n3016;
  wire _abc_43815_n3017;
  wire _abc_43815_n3018_1;
  wire _abc_43815_n3019_1;
  wire _abc_43815_n3020;
  wire _abc_43815_n3021;
  wire _abc_43815_n3022;
  wire _abc_43815_n3023;
  wire _abc_43815_n3024;
  wire _abc_43815_n3025;
  wire _abc_43815_n3027;
  wire _abc_43815_n3028;
  wire _abc_43815_n3029;
  wire _abc_43815_n3030;
  wire _abc_43815_n3031;
  wire _abc_43815_n3032;
  wire _abc_43815_n3033;
  wire _abc_43815_n3034;
  wire _abc_43815_n3036;
  wire _abc_43815_n3037;
  wire _abc_43815_n3038;
  wire _abc_43815_n3039;
  wire _abc_43815_n3040;
  wire _abc_43815_n3041;
  wire _abc_43815_n3042;
  wire _abc_43815_n3043;
  wire _abc_43815_n3045_1;
  wire _abc_43815_n3046;
  wire _abc_43815_n3047;
  wire _abc_43815_n3048;
  wire _abc_43815_n3049;
  wire _abc_43815_n3050;
  wire _abc_43815_n3051;
  wire _abc_43815_n3052;
  wire _abc_43815_n3054;
  wire _abc_43815_n3055;
  wire _abc_43815_n3056;
  wire _abc_43815_n3057;
  wire _abc_43815_n3058;
  wire _abc_43815_n3059;
  wire _abc_43815_n3060;
  wire _abc_43815_n3061;
  wire _abc_43815_n3063;
  wire _abc_43815_n3064;
  wire _abc_43815_n3065;
  wire _abc_43815_n3066;
  wire _abc_43815_n3067;
  wire _abc_43815_n3068;
  wire _abc_43815_n3069;
  wire _abc_43815_n3070_1;
  wire _abc_43815_n3072;
  wire _abc_43815_n3073;
  wire _abc_43815_n3074;
  wire _abc_43815_n3075;
  wire _abc_43815_n3076;
  wire _abc_43815_n3077;
  wire _abc_43815_n3079;
  wire _abc_43815_n3080;
  wire _abc_43815_n3081;
  wire _abc_43815_n3082;
  wire _abc_43815_n3083;
  wire _abc_43815_n3084;
  wire _abc_43815_n3085;
  wire _abc_43815_n3086;
  wire _abc_43815_n3087;
  wire _abc_43815_n3088;
  wire _abc_43815_n3089;
  wire _abc_43815_n3090;
  wire _abc_43815_n3092;
  wire _abc_43815_n3093;
  wire _abc_43815_n3094;
  wire _abc_43815_n3095;
  wire _abc_43815_n3096_1;
  wire _abc_43815_n3097_1;
  wire _abc_43815_n3098;
  wire _abc_43815_n3099;
  wire _abc_43815_n3100;
  wire _abc_43815_n3101;
  wire _abc_43815_n3102;
  wire _abc_43815_n3103;
  wire _abc_43815_n3105;
  wire _abc_43815_n3106;
  wire _abc_43815_n3107;
  wire _abc_43815_n3108;
  wire _abc_43815_n3109;
  wire _abc_43815_n3110;
  wire _abc_43815_n3112;
  wire _abc_43815_n3113;
  wire _abc_43815_n3114;
  wire _abc_43815_n3115;
  wire _abc_43815_n3116;
  wire _abc_43815_n3117;
  wire _abc_43815_n3119;
  wire _abc_43815_n3120;
  wire _abc_43815_n3121;
  wire _abc_43815_n3122_1;
  wire _abc_43815_n3123_1;
  wire _abc_43815_n3124;
  wire _abc_43815_n3126;
  wire _abc_43815_n3127;
  wire _abc_43815_n3128;
  wire _abc_43815_n3129;
  wire _abc_43815_n3130;
  wire _abc_43815_n3131;
  wire _abc_43815_n3133;
  wire _abc_43815_n3134;
  wire _abc_43815_n3135;
  wire _abc_43815_n3136;
  wire _abc_43815_n3137;
  wire _abc_43815_n3138;
  wire _abc_43815_n3139;
  wire _abc_43815_n3141;
  wire _abc_43815_n3142;
  wire _abc_43815_n3143;
  wire _abc_43815_n3144;
  wire _abc_43815_n3145;
  wire _abc_43815_n3146;
  wire _abc_43815_n3147;
  wire _abc_43815_n3148_1;
  wire _abc_43815_n3149_1;
  wire _abc_43815_n3151;
  wire _abc_43815_n3152;
  wire _abc_43815_n3153;
  wire _abc_43815_n3154;
  wire _abc_43815_n3155;
  wire _abc_43815_n3156;
  wire _abc_43815_n3157;
  wire _abc_43815_n3158;
  wire _abc_43815_n3159;
  wire _abc_43815_n3161;
  wire _abc_43815_n3162;
  wire _abc_43815_n3163;
  wire _abc_43815_n3164;
  wire _abc_43815_n3165;
  wire _abc_43815_n3166;
  wire _abc_43815_n3167;
  wire _abc_43815_n3168;
  wire _abc_43815_n3170;
  wire _abc_43815_n3171;
  wire _abc_43815_n3172;
  wire _abc_43815_n3173;
  wire _abc_43815_n3174_1;
  wire _abc_43815_n3175;
  wire _abc_43815_n3176;
  wire _abc_43815_n3177;
  wire _abc_43815_n3179;
  wire _abc_43815_n3180;
  wire _abc_43815_n3181;
  wire _abc_43815_n3182;
  wire _abc_43815_n3183;
  wire _abc_43815_n3184;
  wire _abc_43815_n3185;
  wire _abc_43815_n3186;
  wire _abc_43815_n3187;
  wire _abc_43815_n3189;
  wire _abc_43815_n3190;
  wire _abc_43815_n3191;
  wire _abc_43815_n3192;
  wire _abc_43815_n3193_1;
  wire _abc_43815_n3194;
  wire _abc_43815_n3195;
  wire _abc_43815_n3196;
  wire _abc_43815_n3197;
  wire _abc_43815_n3199;
  wire _abc_43815_n3200;
  wire _abc_43815_n3201;
  wire _abc_43815_n3202;
  wire _abc_43815_n3203;
  wire _abc_43815_n3204;
  wire _abc_43815_n3205;
  wire _abc_43815_n3206;
  wire _abc_43815_n3207;
  wire _abc_43815_n3209_1;
  wire _abc_43815_n3210;
  wire _abc_43815_n3211;
  wire _abc_43815_n3212;
  wire _abc_43815_n3213;
  wire _abc_43815_n3214;
  wire _abc_43815_n3215;
  wire _abc_43815_n3216;
  wire _abc_43815_n3217_1;
  wire _abc_43815_n3219;
  wire _abc_43815_n3220;
  wire _abc_43815_n3221;
  wire _abc_43815_n3222;
  wire _abc_43815_n3223;
  wire _abc_43815_n3224;
  wire _abc_43815_n3225;
  wire _abc_43815_n3226;
  wire _abc_43815_n3227;
  wire _abc_43815_n3229;
  wire _abc_43815_n3230;
  wire _abc_43815_n3231;
  wire _abc_43815_n3232;
  wire _abc_43815_n3233;
  wire _abc_43815_n3234;
  wire _abc_43815_n3235_1;
  wire _abc_43815_n3236;
  wire _abc_43815_n3237;
  wire _abc_43815_n3239;
  wire _abc_43815_n3240;
  wire _abc_43815_n3241;
  wire _abc_43815_n3242;
  wire _abc_43815_n3243;
  wire _abc_43815_n3244_1;
  wire _abc_43815_n3245;
  wire _abc_43815_n3246_1;
  wire _abc_43815_n3247;
  wire _abc_43815_n3249;
  wire _abc_43815_n3250_1;
  wire _abc_43815_n3251;
  wire _abc_43815_n3252_1;
  wire _abc_43815_n3253;
  wire _abc_43815_n3254_1;
  wire _abc_43815_n3255;
  wire _abc_43815_n3256_1;
  wire _abc_43815_n3257;
  wire _abc_43815_n3259;
  wire _abc_43815_n3260_1;
  wire _abc_43815_n3261;
  wire _abc_43815_n3262_1;
  wire _abc_43815_n3263;
  wire _abc_43815_n3264_1;
  wire _abc_43815_n3265;
  wire _abc_43815_n3266_1;
  wire _abc_43815_n3267;
  wire _abc_43815_n3269;
  wire _abc_43815_n3270_1;
  wire _abc_43815_n3271;
  wire _abc_43815_n3272_1;
  wire _abc_43815_n3273;
  wire _abc_43815_n3274_1;
  wire _abc_43815_n3275;
  wire _abc_43815_n3276_1;
  wire _abc_43815_n3277;
  wire _abc_43815_n3279;
  wire _abc_43815_n3280_1;
  wire _abc_43815_n3281;
  wire _abc_43815_n3282_1;
  wire _abc_43815_n3283;
  wire _abc_43815_n3284_1;
  wire _abc_43815_n3285;
  wire _abc_43815_n3286_1;
  wire _abc_43815_n3287;
  wire _abc_43815_n3289;
  wire _abc_43815_n3290_1;
  wire _abc_43815_n3291;
  wire _abc_43815_n3292_1;
  wire _abc_43815_n3293;
  wire _abc_43815_n3294_1;
  wire _abc_43815_n3295;
  wire _abc_43815_n3296_1;
  wire _abc_43815_n3297;
  wire _abc_43815_n3299;
  wire _abc_43815_n3300_1;
  wire _abc_43815_n3301;
  wire _abc_43815_n3302_1;
  wire _abc_43815_n3303;
  wire _abc_43815_n3304_1;
  wire _abc_43815_n3306_1;
  wire _abc_43815_n3307;
  wire _abc_43815_n3308_1;
  wire _abc_43815_n3309;
  wire _abc_43815_n3311;
  wire _abc_43815_n3313;
  wire _abc_43815_n3314;
  wire _abc_43815_n3315;
  wire _abc_43815_n3316_1;
  wire _abc_43815_n3317;
  wire _abc_43815_n3317_bF_buf0;
  wire _abc_43815_n3317_bF_buf1;
  wire _abc_43815_n3317_bF_buf2;
  wire _abc_43815_n3317_bF_buf3;
  wire _abc_43815_n3318;
  wire _abc_43815_n3320;
  wire _abc_43815_n3321;
  wire _abc_43815_n3322;
  wire _abc_43815_n3323_1;
  wire _abc_43815_n3324_1;
  wire _abc_43815_n3325;
  wire _abc_43815_n3326;
  wire _abc_43815_n3327;
  wire _abc_43815_n3328;
  wire _abc_43815_n3329;
  wire _abc_43815_n3332_1;
  wire _abc_43815_n3333;
  wire _abc_43815_n3334;
  wire _abc_43815_n3335;
  wire _abc_43815_n3337;
  wire _abc_43815_n3338;
  wire _abc_43815_n3339_1;
  wire _abc_43815_n3340_1;
  wire _abc_43815_n3342;
  wire _abc_43815_n3343;
  wire _abc_43815_n3344;
  wire _abc_43815_n3345;
  wire _abc_43815_n3347_1;
  wire _abc_43815_n3348_1;
  wire _abc_43815_n3349;
  wire _abc_43815_n3350;
  wire _abc_43815_n3352;
  wire _abc_43815_n3353;
  wire _abc_43815_n3354;
  wire _abc_43815_n3355;
  wire _abc_43815_n3357;
  wire _abc_43815_n3358;
  wire _abc_43815_n3359_1;
  wire _abc_43815_n3360_1;
  wire _abc_43815_n3362;
  wire _abc_43815_n3363;
  wire _abc_43815_n3364;
  wire _abc_43815_n3365;
  wire _abc_43815_n3367;
  wire _abc_43815_n3368;
  wire _abc_43815_n3369_1;
  wire _abc_43815_n3370_1;
  wire _abc_43815_n3372;
  wire _abc_43815_n3373;
  wire _abc_43815_n3374;
  wire _abc_43815_n3375;
  wire _abc_43815_n3377;
  wire _abc_43815_n3378;
  wire _abc_43815_n3379_1;
  wire _abc_43815_n3380_1;
  wire _abc_43815_n3382;
  wire _abc_43815_n3383;
  wire _abc_43815_n3384;
  wire _abc_43815_n3385;
  wire _abc_43815_n3387;
  wire _abc_43815_n3388;
  wire _abc_43815_n3389_1;
  wire _abc_43815_n3390_1;
  wire _abc_43815_n3392;
  wire _abc_43815_n3393;
  wire _abc_43815_n3394;
  wire _abc_43815_n3395;
  wire _abc_43815_n3397;
  wire _abc_43815_n3398;
  wire _abc_43815_n3399_1;
  wire _abc_43815_n3400_1;
  wire _abc_43815_n3402;
  wire _abc_43815_n3403;
  wire _abc_43815_n3404;
  wire _abc_43815_n3405;
  wire _abc_43815_n3407;
  wire _abc_43815_n3408;
  wire _abc_43815_n3409_1;
  wire _abc_43815_n3410_1;
  wire _abc_43815_n3412;
  wire _abc_43815_n3413;
  wire _abc_43815_n3414;
  wire _abc_43815_n3415;
  wire _abc_43815_n3417;
  wire _abc_43815_n3418;
  wire _abc_43815_n3419_1;
  wire _abc_43815_n3420_1;
  wire _abc_43815_n3422;
  wire _abc_43815_n3423;
  wire _abc_43815_n3424;
  wire _abc_43815_n3425;
  wire _abc_43815_n3427;
  wire _abc_43815_n3428;
  wire _abc_43815_n3429_1;
  wire _abc_43815_n3430_1;
  wire _abc_43815_n3432;
  wire _abc_43815_n3433;
  wire _abc_43815_n3434;
  wire _abc_43815_n3435;
  wire _abc_43815_n3437;
  wire _abc_43815_n3438_1;
  wire _abc_43815_n3439_1;
  wire _abc_43815_n3440;
  wire _abc_43815_n3442;
  wire _abc_43815_n3443;
  wire _abc_43815_n3444;
  wire _abc_43815_n3445;
  wire _abc_43815_n3447_1;
  wire _abc_43815_n3448_1;
  wire _abc_43815_n3449;
  wire _abc_43815_n3450;
  wire _abc_43815_n3452;
  wire _abc_43815_n3453;
  wire _abc_43815_n3454;
  wire _abc_43815_n3455;
  wire _abc_43815_n3457_1;
  wire _abc_43815_n3458;
  wire _abc_43815_n3459;
  wire _abc_43815_n3460;
  wire _abc_43815_n3462;
  wire _abc_43815_n3463;
  wire _abc_43815_n3464;
  wire _abc_43815_n3465_1;
  wire _abc_43815_n3467;
  wire _abc_43815_n3468;
  wire _abc_43815_n3469;
  wire _abc_43815_n3470;
  wire _abc_43815_n3472;
  wire _abc_43815_n3473;
  wire _abc_43815_n3474_1;
  wire _abc_43815_n3475_1;
  wire _abc_43815_n3477;
  wire _abc_43815_n3478;
  wire _abc_43815_n3479;
  wire _abc_43815_n3480;
  wire _abc_43815_n3482;
  wire _abc_43815_n3483_1;
  wire _abc_43815_n3484_1;
  wire _abc_43815_n3485;
  wire _abc_43815_n3487;
  wire _abc_43815_n3488;
  wire _abc_43815_n3489;
  wire _abc_43815_n3490;
  wire _abc_43815_n3492_1;
  wire _abc_43815_n3493_1;
  wire _abc_43815_n3494;
  wire _abc_43815_n3495;
  wire _abc_43815_n3496;
  wire _abc_43815_n3496_bF_buf0;
  wire _abc_43815_n3496_bF_buf1;
  wire _abc_43815_n3496_bF_buf2;
  wire _abc_43815_n3496_bF_buf3;
  wire _abc_43815_n3497;
  wire _abc_43815_n3498;
  wire _abc_43815_n3499;
  wire _abc_43815_n3500;
  wire _abc_43815_n3501_1;
  wire _abc_43815_n3502_1;
  wire _abc_43815_n3503;
  wire _abc_43815_n3504;
  wire _abc_43815_n3505;
  wire _abc_43815_n3506;
  wire _abc_43815_n3508;
  wire _abc_43815_n3509;
  wire _abc_43815_n3510;
  wire _abc_43815_n3511_1;
  wire _abc_43815_n3512_1;
  wire _abc_43815_n3513;
  wire _abc_43815_n3514;
  wire _abc_43815_n3515;
  wire _abc_43815_n3516;
  wire _abc_43815_n3518;
  wire _abc_43815_n3519;
  wire _abc_43815_n3520;
  wire _abc_43815_n3521_1;
  wire _abc_43815_n3521_1_bF_buf0;
  wire _abc_43815_n3521_1_bF_buf1;
  wire _abc_43815_n3521_1_bF_buf2;
  wire _abc_43815_n3521_1_bF_buf3;
  wire _abc_43815_n3522_1;
  wire _abc_43815_n3523;
  wire _abc_43815_n3524;
  wire _abc_43815_n3525;
  wire _abc_43815_n3526;
  wire _abc_43815_n3527;
  wire _abc_43815_n3528;
  wire _abc_43815_n3530;
  wire _abc_43815_n3531_1;
  wire _abc_43815_n3532_1;
  wire _abc_43815_n3533;
  wire _abc_43815_n3534;
  wire _abc_43815_n3535;
  wire _abc_43815_n3536;
  wire _abc_43815_n3538;
  wire _abc_43815_n3539;
  wire _abc_43815_n3540;
  wire _abc_43815_n3541_1;
  wire _abc_43815_n3542_1;
  wire _abc_43815_n3543;
  wire _abc_43815_n3544;
  wire _abc_43815_n3545;
  wire _abc_43815_n3546;
  wire _abc_43815_n3547;
  wire _abc_43815_n3548;
  wire _abc_43815_n3549;
  wire _abc_43815_n3549_bF_buf0;
  wire _abc_43815_n3549_bF_buf1;
  wire _abc_43815_n3549_bF_buf2;
  wire _abc_43815_n3549_bF_buf3;
  wire _abc_43815_n3549_bF_buf4;
  wire _abc_43815_n3550;
  wire _abc_43815_n3552_1;
  wire _abc_43815_n3553;
  wire _abc_43815_n3554;
  wire _abc_43815_n3555;
  wire _abc_43815_n3556;
  wire _abc_43815_n3557;
  wire _abc_43815_n3558;
  wire _abc_43815_n3559;
  wire _abc_43815_n3560;
  wire _abc_43815_n3562_1;
  wire _abc_43815_n3563;
  wire _abc_43815_n3564;
  wire _abc_43815_n3565;
  wire _abc_43815_n3566;
  wire _abc_43815_n3567;
  wire _abc_43815_n3568;
  wire _abc_43815_n3569;
  wire _abc_43815_n3570;
  wire _abc_43815_n3572_1;
  wire _abc_43815_n3573;
  wire _abc_43815_n3574;
  wire _abc_43815_n3575;
  wire _abc_43815_n3576;
  wire _abc_43815_n3577;
  wire _abc_43815_n3578;
  wire _abc_43815_n3579;
  wire _abc_43815_n3580;
  wire _abc_43815_n3582_1;
  wire _abc_43815_n3583;
  wire _abc_43815_n3584;
  wire _abc_43815_n3585;
  wire _abc_43815_n3586;
  wire _abc_43815_n3587;
  wire _abc_43815_n3588;
  wire _abc_43815_n3589;
  wire _abc_43815_n3590_1;
  wire _abc_43815_n3592;
  wire _abc_43815_n3593;
  wire _abc_43815_n3594;
  wire _abc_43815_n3595;
  wire _abc_43815_n3596;
  wire _abc_43815_n3597;
  wire _abc_43815_n3598;
  wire _abc_43815_n3599_1;
  wire _abc_43815_n3600_1;
  wire _abc_43815_n3602;
  wire _abc_43815_n3603;
  wire _abc_43815_n3604;
  wire _abc_43815_n3605;
  wire _abc_43815_n3606;
  wire _abc_43815_n3607;
  wire _abc_43815_n3608_1;
  wire _abc_43815_n3609_1;
  wire _abc_43815_n3610;
  wire _abc_43815_n3612;
  wire _abc_43815_n3613;
  wire _abc_43815_n3614;
  wire _abc_43815_n3615;
  wire _abc_43815_n3616;
  wire _abc_43815_n3617_1;
  wire _abc_43815_n3618_1;
  wire _abc_43815_n3619;
  wire _abc_43815_n3620;
  wire _abc_43815_n3622;
  wire _abc_43815_n3623;
  wire _abc_43815_n3624;
  wire _abc_43815_n3625;
  wire _abc_43815_n3626_1;
  wire _abc_43815_n3627_1;
  wire _abc_43815_n3628;
  wire _abc_43815_n3629;
  wire _abc_43815_n3630;
  wire _abc_43815_n3631;
  wire _abc_43815_n3632;
  wire _abc_43815_n3633;
  wire _abc_43815_n3634;
  wire _abc_43815_n3635_1;
  wire _abc_43815_n3637;
  wire _abc_43815_n3638;
  wire _abc_43815_n3639;
  wire _abc_43815_n3640;
  wire _abc_43815_n3641;
  wire _abc_43815_n3642;
  wire _abc_43815_n3643;
  wire _abc_43815_n3644_1;
  wire _abc_43815_n3645_1;
  wire _abc_43815_n3646;
  wire _abc_43815_n3647;
  wire _abc_43815_n3648;
  wire _abc_43815_n3649;
  wire _abc_43815_n3650;
  wire _abc_43815_n3652;
  wire _abc_43815_n3653_1;
  wire _abc_43815_n3654;
  wire _abc_43815_n3655_1;
  wire _abc_43815_n3656;
  wire _abc_43815_n3657;
  wire _abc_43815_n3658;
  wire _abc_43815_n3659;
  wire _abc_43815_n3660;
  wire _abc_43815_n3661;
  wire _abc_43815_n3662;
  wire _abc_43815_n3663;
  wire _abc_43815_n3664;
  wire _abc_43815_n3665;
  wire _abc_43815_n3667_1;
  wire _abc_43815_n3668_1;
  wire _abc_43815_n3669_1;
  wire _abc_43815_n3670;
  wire _abc_43815_n3671;
  wire _abc_43815_n3672;
  wire _abc_43815_n3673;
  wire _abc_43815_n3674;
  wire _abc_43815_n3675;
  wire _abc_43815_n3676;
  wire _abc_43815_n3677;
  wire _abc_43815_n3678;
  wire _abc_43815_n3679;
  wire _abc_43815_n3680_1;
  wire _abc_43815_n3682;
  wire _abc_43815_n3683_1;
  wire _abc_43815_n3684;
  wire _abc_43815_n3685;
  wire _abc_43815_n3686;
  wire _abc_43815_n3687;
  wire _abc_43815_n3688;
  wire _abc_43815_n3689;
  wire _abc_43815_n3690;
  wire _abc_43815_n3691;
  wire _abc_43815_n3692;
  wire _abc_43815_n3693;
  wire _abc_43815_n3694_1;
  wire _abc_43815_n3695_1;
  wire _abc_43815_n3697;
  wire _abc_43815_n3698;
  wire _abc_43815_n3699;
  wire _abc_43815_n3700;
  wire _abc_43815_n3701_1;
  wire _abc_43815_n3702_1;
  wire _abc_43815_n3703;
  wire _abc_43815_n3704;
  wire _abc_43815_n3705;
  wire _abc_43815_n3706;
  wire _abc_43815_n3707_1;
  wire _abc_43815_n3708;
  wire _abc_43815_n3709;
  wire _abc_43815_n3710;
  wire _abc_43815_n3712;
  wire _abc_43815_n3713_1;
  wire _abc_43815_n3714;
  wire _abc_43815_n3715;
  wire _abc_43815_n3716;
  wire _abc_43815_n3717;
  wire _abc_43815_n3718;
  wire _abc_43815_n3719;
  wire _abc_43815_n3720_1;
  wire _abc_43815_n3721;
  wire _abc_43815_n3722;
  wire _abc_43815_n3723;
  wire _abc_43815_n3724;
  wire _abc_43815_n3725;
  wire _abc_43815_n3727;
  wire _abc_43815_n3728;
  wire _abc_43815_n3729;
  wire _abc_43815_n3730;
  wire _abc_43815_n3731;
  wire _abc_43815_n3732;
  wire _abc_43815_n3733_1;
  wire _abc_43815_n3734;
  wire _abc_43815_n3735;
  wire _abc_43815_n3736;
  wire _abc_43815_n3737;
  wire _abc_43815_n3738;
  wire _abc_43815_n3739;
  wire _abc_43815_n3740;
  wire _abc_43815_n3742;
  wire _abc_43815_n3743_1;
  wire _abc_43815_n3744;
  wire _abc_43815_n3745;
  wire _abc_43815_n3746;
  wire _abc_43815_n3747;
  wire _abc_43815_n3748;
  wire _abc_43815_n3749;
  wire _abc_43815_n3750_1;
  wire _abc_43815_n3751;
  wire _abc_43815_n3752;
  wire _abc_43815_n3753;
  wire _abc_43815_n3755;
  wire _abc_43815_n3756_1;
  wire _abc_43815_n3757;
  wire _abc_43815_n3758;
  wire _abc_43815_n3759;
  wire _abc_43815_n3760;
  wire _abc_43815_n3761;
  wire _abc_43815_n3762;
  wire _abc_43815_n3763_1;
  wire _abc_43815_n3764;
  wire _abc_43815_n3765;
  wire _abc_43815_n3766;
  wire _abc_43815_n3768;
  wire _abc_43815_n3769;
  wire _abc_43815_n3770;
  wire _abc_43815_n3771;
  wire _abc_43815_n3772;
  wire _abc_43815_n3773_1;
  wire _abc_43815_n3774;
  wire _abc_43815_n3775;
  wire _abc_43815_n3776;
  wire _abc_43815_n3777;
  wire _abc_43815_n3778;
  wire _abc_43815_n3779;
  wire _abc_43815_n3781;
  wire _abc_43815_n3782;
  wire _abc_43815_n3783;
  wire _abc_43815_n3784;
  wire _abc_43815_n3785;
  wire _abc_43815_n3786_1;
  wire _abc_43815_n3787;
  wire _abc_43815_n3788;
  wire _abc_43815_n3789;
  wire _abc_43815_n3790;
  wire _abc_43815_n3791;
  wire _abc_43815_n3793_1;
  wire _abc_43815_n3794;
  wire _abc_43815_n3795;
  wire _abc_43815_n3796;
  wire _abc_43815_n3797;
  wire _abc_43815_n3798;
  wire _abc_43815_n3799;
  wire _abc_43815_n3800;
  wire _abc_43815_n3801;
  wire _abc_43815_n3802;
  wire _abc_43815_n3803;
  wire _abc_43815_n3804;
  wire _abc_43815_n3806;
  wire _abc_43815_n3807;
  wire _abc_43815_n3808;
  wire _abc_43815_n3809;
  wire _abc_43815_n3810;
  wire _abc_43815_n3811;
  wire _abc_43815_n3812_1;
  wire _abc_43815_n3813;
  wire _abc_43815_n3814;
  wire _abc_43815_n3815;
  wire _abc_43815_n3816;
  wire _abc_43815_n3817;
  wire _abc_43815_n3819;
  wire _abc_43815_n3820;
  wire _abc_43815_n3821;
  wire _abc_43815_n3822;
  wire _abc_43815_n3823;
  wire _abc_43815_n3824;
  wire _abc_43815_n3825_1;
  wire _abc_43815_n3826;
  wire _abc_43815_n3827;
  wire _abc_43815_n3828;
  wire _abc_43815_n3829;
  wire _abc_43815_n3830;
  wire _abc_43815_n3832;
  wire _abc_43815_n3833;
  wire _abc_43815_n3834;
  wire _abc_43815_n3835_1;
  wire _abc_43815_n3836;
  wire _abc_43815_n3837;
  wire _abc_43815_n3838;
  wire _abc_43815_n3839;
  wire _abc_43815_n3840;
  wire _abc_43815_n3841;
  wire _abc_43815_n3842_1;
  wire _abc_43815_n3844;
  wire _abc_43815_n3845;
  wire _abc_43815_n3846;
  wire _abc_43815_n3847;
  wire _abc_43815_n3848;
  wire _abc_43815_n3849_1;
  wire _abc_43815_n3850;
  wire _abc_43815_n3851;
  wire _abc_43815_n3852;
  wire _abc_43815_n3853;
  wire _abc_43815_n3854;
  wire _abc_43815_n3855;
  wire _abc_43815_n3856_1;
  wire _abc_43815_n3857;
  wire _abc_43815_n3859;
  wire _abc_43815_n3860;
  wire _abc_43815_n3861;
  wire _abc_43815_n3862;
  wire _abc_43815_n3863;
  wire _abc_43815_n3864;
  wire _abc_43815_n3865;
  wire _abc_43815_n3866;
  wire _abc_43815_n3867;
  wire _abc_43815_n3868;
  wire _abc_43815_n3869;
  wire _abc_43815_n3870_1;
  wire _abc_43815_n3871;
  wire _abc_43815_n3872;
  wire _abc_43815_n3874;
  wire _abc_43815_n3875;
  wire _abc_43815_n3876;
  wire _abc_43815_n3877_1;
  wire _abc_43815_n3878;
  wire _abc_43815_n3879;
  wire _abc_43815_n3880;
  wire _abc_43815_n3881;
  wire _abc_43815_n3882;
  wire _abc_43815_n3883;
  wire _abc_43815_n3884_1;
  wire _abc_43815_n3885;
  wire _abc_43815_n3886;
  wire _abc_43815_n3887;
  wire _abc_43815_n3889;
  wire _abc_43815_n3890;
  wire _abc_43815_n3891_1;
  wire _abc_43815_n3892;
  wire _abc_43815_n3893;
  wire _abc_43815_n3894;
  wire _abc_43815_n3895;
  wire _abc_43815_n3896;
  wire _abc_43815_n3897;
  wire _abc_43815_n3898;
  wire _abc_43815_n3899;
  wire _abc_43815_n3900;
  wire _abc_43815_n3901_1;
  wire _abc_43815_n3902;
  wire _abc_43815_n3904;
  wire _abc_43815_n3905;
  wire _abc_43815_n3906;
  wire _abc_43815_n3907;
  wire _abc_43815_n3908_1;
  wire _abc_43815_n3909;
  wire _abc_43815_n3910;
  wire _abc_43815_n3911;
  wire _abc_43815_n3912;
  wire _abc_43815_n3913;
  wire _abc_43815_n3914;
  wire _abc_43815_n3915;
  wire _abc_43815_n3916_1;
  wire _abc_43815_n3917;
  wire _abc_43815_n3919;
  wire _abc_43815_n3920;
  wire _abc_43815_n3921;
  wire _abc_43815_n3922;
  wire _abc_43815_n3923_1;
  wire _abc_43815_n3924;
  wire _abc_43815_n3925;
  wire _abc_43815_n3926;
  wire _abc_43815_n3927;
  wire _abc_43815_n3928;
  wire _abc_43815_n3929;
  wire _abc_43815_n3930;
  wire _abc_43815_n3931;
  wire _abc_43815_n3932;
  wire _abc_43815_n3934;
  wire _abc_43815_n3935;
  wire _abc_43815_n3936;
  wire _abc_43815_n3937;
  wire _abc_43815_n3938_1;
  wire _abc_43815_n3939;
  wire _abc_43815_n3940;
  wire _abc_43815_n3941;
  wire _abc_43815_n3942;
  wire _abc_43815_n3943;
  wire _abc_43815_n3944;
  wire _abc_43815_n3945_1;
  wire _abc_43815_n3946;
  wire _abc_43815_n3947;
  wire _abc_43815_n3949;
  wire _abc_43815_n3950;
  wire _abc_43815_n3951_1;
  wire _abc_43815_n3952;
  wire _abc_43815_n3953;
  wire _abc_43815_n3954;
  wire _abc_43815_n3955;
  wire _abc_43815_n3956;
  wire _abc_43815_n3957;
  wire _abc_43815_n3958_1;
  wire _abc_43815_n3959;
  wire _abc_43815_n3960;
  wire _abc_43815_n3961;
  wire _abc_43815_n3962;
  wire _abc_43815_n3964;
  wire _abc_43815_n3965;
  wire _abc_43815_n3966_1;
  wire _abc_43815_n3967;
  wire _abc_43815_n3968;
  wire _abc_43815_n3969;
  wire _abc_43815_n3970;
  wire _abc_43815_n3972;
  wire _abc_43815_n3973_1;
  wire _abc_43815_n3974;
  wire _abc_43815_n3975;
  wire _abc_43815_n3977;
  wire _abc_43815_n3978_1;
  wire _abc_43815_n3979;
  wire _abc_43815_n3980;
  wire _abc_43815_n3981;
  wire _abc_43815_n3982;
  wire _abc_43815_n3984;
  wire _abc_43815_n3985_1;
  wire _abc_43815_n3985_1_bF_buf0;
  wire _abc_43815_n3985_1_bF_buf1;
  wire _abc_43815_n3985_1_bF_buf2;
  wire _abc_43815_n3985_1_bF_buf3;
  wire _abc_43815_n3985_1_bF_buf4;
  wire _abc_43815_n3986;
  wire _abc_43815_n3988;
  wire _abc_43815_n3989;
  wire _abc_43815_n3991;
  wire _abc_43815_n3992;
  wire _abc_43815_n3993;
  wire _abc_43815_n3994;
  wire _abc_43815_n3995_1;
  wire _abc_43815_n3996;
  wire _abc_43815_n3997;
  wire _abc_43815_n3998;
  wire _abc_43815_n3999;
  wire _abc_43815_n4000;
  wire _abc_43815_n4001;
  wire _abc_43815_n4002_1;
  wire _abc_43815_n4003;
  wire _abc_43815_n4004;
  wire _abc_43815_n4005;
  wire _abc_43815_n4007;
  wire _abc_43815_n4008_1;
  wire _abc_43815_n4009;
  wire _abc_43815_n4010;
  wire _abc_43815_n4011;
  wire _abc_43815_n4012;
  wire _abc_43815_n4013;
  wire _abc_43815_n4014;
  wire _abc_43815_n4015_1;
  wire _abc_43815_n4016;
  wire _abc_43815_n4017;
  wire _abc_43815_n4018;
  wire _abc_43815_n4019;
  wire _abc_43815_n4021;
  wire _abc_43815_n4022_1;
  wire _abc_43815_n4023;
  wire _abc_43815_n4024;
  wire _abc_43815_n4025;
  wire _abc_43815_n4026;
  wire _abc_43815_n4027;
  wire _abc_43815_n4028;
  wire _abc_43815_n4029_1;
  wire _abc_43815_n4030;
  wire _abc_43815_n4031;
  wire _abc_43815_n4032;
  wire _abc_43815_n4033;
  wire _abc_43815_n4034_1;
  wire _abc_43815_n4035;
  wire _abc_43815_n4036;
  wire _abc_43815_n4038;
  wire _abc_43815_n4039;
  wire _abc_43815_n4040;
  wire _abc_43815_n4041_1;
  wire _abc_43815_n4042;
  wire _abc_43815_n4043;
  wire _abc_43815_n4044;
  wire _abc_43815_n4045;
  wire _abc_43815_n4046;
  wire _abc_43815_n4047;
  wire _abc_43815_n4048;
  wire _abc_43815_n4049;
  wire _abc_43815_n4050;
  wire _abc_43815_n4052;
  wire _abc_43815_n4053;
  wire _abc_43815_n4054;
  wire _abc_43815_n4055_1;
  wire _abc_43815_n4056;
  wire _abc_43815_n4057;
  wire _abc_43815_n4058;
  wire _abc_43815_n4059;
  wire _abc_43815_n4060;
  wire _abc_43815_n4061;
  wire _abc_43815_n4062_1;
  wire _abc_43815_n4063;
  wire _abc_43815_n4064;
  wire _abc_43815_n4066;
  wire _abc_43815_n4067;
  wire _abc_43815_n4068_1;
  wire _abc_43815_n4069;
  wire _abc_43815_n4070;
  wire _abc_43815_n4071;
  wire _abc_43815_n4072;
  wire _abc_43815_n4073;
  wire _abc_43815_n4074;
  wire _abc_43815_n4075_1;
  wire _abc_43815_n4076;
  wire _abc_43815_n4077;
  wire _abc_43815_n4078;
  wire _abc_43815_n4080;
  wire _abc_43815_n4081;
  wire _abc_43815_n4082_1;
  wire _abc_43815_n4083;
  wire _abc_43815_n4084;
  wire _abc_43815_n4085;
  wire _abc_43815_n4086;
  wire _abc_43815_n4087;
  wire _abc_43815_n4088;
  wire _abc_43815_n4089_1;
  wire _abc_43815_n4090;
  wire _abc_43815_n4091;
  wire _abc_43815_n4092;
  wire _abc_43815_n4093;
  wire _abc_43815_n4094_1;
  wire _abc_43815_n4095;
  wire _abc_43815_n4097;
  wire _abc_43815_n4098;
  wire _abc_43815_n4099;
  wire _abc_43815_n4100;
  wire _abc_43815_n4101_1;
  wire _abc_43815_n4102;
  wire _abc_43815_n4103;
  wire _abc_43815_n4104;
  wire _abc_43815_n4105;
  wire _abc_43815_n4106;
  wire _abc_43815_n4107;
  wire _abc_43815_n4108;
  wire _abc_43815_n4109;
  wire _abc_43815_n4110;
  wire _abc_43815_n4112_1;
  wire _abc_43815_n4113;
  wire _abc_43815_n4114;
  wire _abc_43815_n4115;
  wire _abc_43815_n4116;
  wire _abc_43815_n4117;
  wire _abc_43815_n4118;
  wire _abc_43815_n4119_1;
  wire _abc_43815_n4120;
  wire _abc_43815_n4121;
  wire _abc_43815_n4122;
  wire _abc_43815_n4123;
  wire _abc_43815_n4124_1;
  wire _abc_43815_n4125;
  wire _abc_43815_n4126;
  wire _abc_43815_n4127;
  wire _abc_43815_n4128;
  wire _abc_43815_n4129;
  wire _abc_43815_n4131_1;
  wire _abc_43815_n4132;
  wire _abc_43815_n4133;
  wire _abc_43815_n4134;
  wire _abc_43815_n4135;
  wire _abc_43815_n4136;
  wire _abc_43815_n4137;
  wire _abc_43815_n4138_1;
  wire _abc_43815_n4139;
  wire _abc_43815_n4140;
  wire _abc_43815_n4141;
  wire _abc_43815_n4142;
  wire _abc_43815_n4143;
  wire _abc_43815_n4144;
  wire _abc_43815_n4145_1;
  wire _abc_43815_n4146;
  wire _abc_43815_n4147;
  wire _abc_43815_n4148;
  wire _abc_43815_n4150_1;
  wire _abc_43815_n4151;
  wire _abc_43815_n4152;
  wire _abc_43815_n4153;
  wire _abc_43815_n4154;
  wire _abc_43815_n4155;
  wire _abc_43815_n4156;
  wire _abc_43815_n4157_1;
  wire _abc_43815_n4158_1;
  wire _abc_43815_n4159;
  wire _abc_43815_n4160;
  wire _abc_43815_n4161_1;
  wire _abc_43815_n4162_1;
  wire _abc_43815_n4163;
  wire _abc_43815_n4164_1;
  wire _abc_43815_n4165_1;
  wire _abc_43815_n4166_1;
  wire _abc_43815_n4167;
  wire _abc_43815_n4167_1;
  wire _abc_43815_n4167_bF_buf0;
  wire _abc_43815_n4167_bF_buf1;
  wire _abc_43815_n4167_bF_buf10;
  wire _abc_43815_n4167_bF_buf11;
  wire _abc_43815_n4167_bF_buf12;
  wire _abc_43815_n4167_bF_buf13;
  wire _abc_43815_n4167_bF_buf14;
  wire _abc_43815_n4167_bF_buf15;
  wire _abc_43815_n4167_bF_buf15_bF_buf0;
  wire _abc_43815_n4167_bF_buf15_bF_buf1;
  wire _abc_43815_n4167_bF_buf15_bF_buf2;
  wire _abc_43815_n4167_bF_buf15_bF_buf3;
  wire _abc_43815_n4167_bF_buf2;
  wire _abc_43815_n4167_bF_buf3;
  wire _abc_43815_n4167_bF_buf4;
  wire _abc_43815_n4167_bF_buf5;
  wire _abc_43815_n4167_bF_buf6;
  wire _abc_43815_n4167_bF_buf7;
  wire _abc_43815_n4167_bF_buf8;
  wire _abc_43815_n4167_bF_buf9;
  wire _abc_43815_n4168;
  wire _abc_43815_n4169;
  wire _abc_43815_n4170;
  wire _abc_43815_n4171;
  wire _abc_43815_n4172;
  wire _abc_43815_n4174;
  wire _abc_43815_n4175;
  wire _abc_43815_n4176;
  wire _abc_43815_n4177;
  wire _abc_43815_n4178;
  wire _abc_43815_n4179;
  wire _abc_43815_n4180;
  wire _abc_43815_n4181;
  wire _abc_43815_n4182;
  wire _abc_43815_n4183;
  wire _abc_43815_n4184;
  wire _abc_43815_n4185;
  wire _abc_43815_n4186;
  wire _abc_43815_n4187;
  wire _abc_43815_n4188;
  wire _abc_43815_n4189;
  wire _abc_43815_n4190;
  wire _abc_43815_n4191;
  wire _abc_43815_n4192;
  wire _abc_43815_n4193;
  wire _abc_43815_n4195;
  wire _abc_43815_n4196;
  wire _abc_43815_n4197;
  wire _abc_43815_n4198;
  wire _abc_43815_n4199;
  wire _abc_43815_n4200;
  wire _abc_43815_n4201;
  wire _abc_43815_n4202;
  wire _abc_43815_n4203;
  wire _abc_43815_n4204;
  wire _abc_43815_n4205;
  wire _abc_43815_n4206;
  wire _abc_43815_n4207;
  wire _abc_43815_n4208;
  wire _abc_43815_n4209;
  wire _abc_43815_n4210;
  wire _abc_43815_n4211;
  wire _abc_43815_n4212;
  wire _abc_43815_n4214;
  wire _abc_43815_n4215;
  wire _abc_43815_n4216;
  wire _abc_43815_n4217;
  wire _abc_43815_n4217_bF_buf0;
  wire _abc_43815_n4217_bF_buf1;
  wire _abc_43815_n4217_bF_buf2;
  wire _abc_43815_n4217_bF_buf3;
  wire _abc_43815_n4217_bF_buf4;
  wire _abc_43815_n4218;
  wire _abc_43815_n4219;
  wire _abc_43815_n4220;
  wire _abc_43815_n4221;
  wire _abc_43815_n4222;
  wire _abc_43815_n4223;
  wire _abc_43815_n4224;
  wire _abc_43815_n4225;
  wire _abc_43815_n4226;
  wire _abc_43815_n4227;
  wire _abc_43815_n4228;
  wire _abc_43815_n4229;
  wire _abc_43815_n4230;
  wire _abc_43815_n4231;
  wire _abc_43815_n4232;
  wire _abc_43815_n4234;
  wire _abc_43815_n4235;
  wire _abc_43815_n4236;
  wire _abc_43815_n4237;
  wire _abc_43815_n4238;
  wire _abc_43815_n4239;
  wire _abc_43815_n4240;
  wire _abc_43815_n4241;
  wire _abc_43815_n4242;
  wire _abc_43815_n4243;
  wire _abc_43815_n4244;
  wire _abc_43815_n4245;
  wire _abc_43815_n4246;
  wire _abc_43815_n4247;
  wire _abc_43815_n4248;
  wire _abc_43815_n4249;
  wire _abc_43815_n4250;
  wire _abc_43815_n4251;
  wire _abc_43815_n4252;
  wire _abc_43815_n4253;
  wire _abc_43815_n4254;
  wire _abc_43815_n4255;
  wire _abc_43815_n4256;
  wire _abc_43815_n4258;
  wire _abc_43815_n4259;
  wire _abc_43815_n4260;
  wire _abc_43815_n4261;
  wire _abc_43815_n4262;
  wire _abc_43815_n4263;
  wire _abc_43815_n4264;
  wire _abc_43815_n4265;
  wire _abc_43815_n4266;
  wire _abc_43815_n4267;
  wire _abc_43815_n4268;
  wire _abc_43815_n4269;
  wire _abc_43815_n4270;
  wire _abc_43815_n4271;
  wire _abc_43815_n4273;
  wire _abc_43815_n4274;
  wire _abc_43815_n4275;
  wire _abc_43815_n4276;
  wire _abc_43815_n4277;
  wire _abc_43815_n4278;
  wire _abc_43815_n4279;
  wire _abc_43815_n4280;
  wire _abc_43815_n4281;
  wire _abc_43815_n4282;
  wire _abc_43815_n4283;
  wire _abc_43815_n4284;
  wire _abc_43815_n4285;
  wire _abc_43815_n4286;
  wire _abc_43815_n4287;
  wire _abc_43815_n4288;
  wire _abc_43815_n4289;
  wire _abc_43815_n4291;
  wire _abc_43815_n4292;
  wire _abc_43815_n4293;
  wire _abc_43815_n4294;
  wire _abc_43815_n4295;
  wire _abc_43815_n4296;
  wire _abc_43815_n4297;
  wire _abc_43815_n4298;
  wire _abc_43815_n4299;
  wire _abc_43815_n4300;
  wire _abc_43815_n4301;
  wire _abc_43815_n4302;
  wire _abc_43815_n4303;
  wire _abc_43815_n4304;
  wire _abc_43815_n4306;
  wire _abc_43815_n4307;
  wire _abc_43815_n4308;
  wire _abc_43815_n4309;
  wire _abc_43815_n4310;
  wire _abc_43815_n4311;
  wire _abc_43815_n4312;
  wire _abc_43815_n4313;
  wire _abc_43815_n4314;
  wire _abc_43815_n4315;
  wire _abc_43815_n4316;
  wire _abc_43815_n4317;
  wire _abc_43815_n4318;
  wire _abc_43815_n4319;
  wire _abc_43815_n4320;
  wire _abc_43815_n4321;
  wire _abc_43815_n4322;
  wire _abc_43815_n4323;
  wire _abc_43815_n4324;
  wire _abc_43815_n4325;
  wire _abc_43815_n4326;
  wire _abc_43815_n4328;
  wire _abc_43815_n4329;
  wire _abc_43815_n4330;
  wire _abc_43815_n4331;
  wire _abc_43815_n4332;
  wire _abc_43815_n4333;
  wire _abc_43815_n4334;
  wire _abc_43815_n4335;
  wire _abc_43815_n4336;
  wire _abc_43815_n4337;
  wire _abc_43815_n4338;
  wire _abc_43815_n4339;
  wire _abc_43815_n4340;
  wire _abc_43815_n4341;
  wire _abc_43815_n4343;
  wire _abc_43815_n4344;
  wire _abc_43815_n4345;
  wire _abc_43815_n4346;
  wire _abc_43815_n4347;
  wire _abc_43815_n4348;
  wire _abc_43815_n4349;
  wire _abc_43815_n4350;
  wire _abc_43815_n4351;
  wire _abc_43815_n4352;
  wire _abc_43815_n4353;
  wire _abc_43815_n4354;
  wire _abc_43815_n4355;
  wire _abc_43815_n4356;
  wire _abc_43815_n4357;
  wire _abc_43815_n4358;
  wire _abc_43815_n4360;
  wire _abc_43815_n4361;
  wire _abc_43815_n4362;
  wire _abc_43815_n4363;
  wire _abc_43815_n4364;
  wire _abc_43815_n4365;
  wire _abc_43815_n4366;
  wire _abc_43815_n4367;
  wire _abc_43815_n4368;
  wire _abc_43815_n4369;
  wire _abc_43815_n4370;
  wire _abc_43815_n4371;
  wire _abc_43815_n4372;
  wire _abc_43815_n4373;
  wire _abc_43815_n4375;
  wire _abc_43815_n4376;
  wire _abc_43815_n4377;
  wire _abc_43815_n4378;
  wire _abc_43815_n4379;
  wire _abc_43815_n4380;
  wire _abc_43815_n4381;
  wire _abc_43815_n4382;
  wire _abc_43815_n4383;
  wire _abc_43815_n4384;
  wire _abc_43815_n4385;
  wire _abc_43815_n4386;
  wire _abc_43815_n4387;
  wire _abc_43815_n4388;
  wire _abc_43815_n4389;
  wire _abc_43815_n4390;
  wire _abc_43815_n4391;
  wire _abc_43815_n4392;
  wire _abc_43815_n4393;
  wire _abc_43815_n4394;
  wire _abc_43815_n4395;
  wire _abc_43815_n4397;
  wire _abc_43815_n4398;
  wire _abc_43815_n4399;
  wire _abc_43815_n4400;
  wire _abc_43815_n4401;
  wire _abc_43815_n4402;
  wire _abc_43815_n4403;
  wire _abc_43815_n4404;
  wire _abc_43815_n4405;
  wire _abc_43815_n4406;
  wire _abc_43815_n4407;
  wire _abc_43815_n4408;
  wire _abc_43815_n4409;
  wire _abc_43815_n4410;
  wire _abc_43815_n4412;
  wire _abc_43815_n4413;
  wire _abc_43815_n4414;
  wire _abc_43815_n4415;
  wire _abc_43815_n4416;
  wire _abc_43815_n4417;
  wire _abc_43815_n4418;
  wire _abc_43815_n4419;
  wire _abc_43815_n4420;
  wire _abc_43815_n4421;
  wire _abc_43815_n4422;
  wire _abc_43815_n4423;
  wire _abc_43815_n4424;
  wire _abc_43815_n4425;
  wire _abc_43815_n4426;
  wire _abc_43815_n4427;
  wire _abc_43815_n4428;
  wire _abc_43815_n4430;
  wire _abc_43815_n4431;
  wire _abc_43815_n4432;
  wire _abc_43815_n4433;
  wire _abc_43815_n4434;
  wire _abc_43815_n4435;
  wire _abc_43815_n4436;
  wire _abc_43815_n4437;
  wire _abc_43815_n4438;
  wire _abc_43815_n4439;
  wire _abc_43815_n4440;
  wire _abc_43815_n4441;
  wire _abc_43815_n4442;
  wire _abc_43815_n4443;
  wire _abc_43815_n4445;
  wire _abc_43815_n4446;
  wire _abc_43815_n4447;
  wire _abc_43815_n4448;
  wire _abc_43815_n4449;
  wire _abc_43815_n4450;
  wire _abc_43815_n4451;
  wire _abc_43815_n4452;
  wire _abc_43815_n4453;
  wire _abc_43815_n4454;
  wire _abc_43815_n4455;
  wire _abc_43815_n4456;
  wire _abc_43815_n4457;
  wire _abc_43815_n4458;
  wire _abc_43815_n4459;
  wire _abc_43815_n4460;
  wire _abc_43815_n4461;
  wire _abc_43815_n4462;
  wire _abc_43815_n4463;
  wire _abc_43815_n4464;
  wire _abc_43815_n4465;
  wire _abc_43815_n4466;
  wire _abc_43815_n4467;
  wire _abc_43815_n4468;
  wire _abc_43815_n4469;
  wire _abc_43815_n4471;
  wire _abc_43815_n4472;
  wire _abc_43815_n4473;
  wire _abc_43815_n4474;
  wire _abc_43815_n4475;
  wire _abc_43815_n4476;
  wire _abc_43815_n4477;
  wire _abc_43815_n4478;
  wire _abc_43815_n4479;
  wire _abc_43815_n4480;
  wire _abc_43815_n4481;
  wire _abc_43815_n4482;
  wire _abc_43815_n4483;
  wire _abc_43815_n4484;
  wire _abc_43815_n4486;
  wire _abc_43815_n4487;
  wire _abc_43815_n4488;
  wire _abc_43815_n4489;
  wire _abc_43815_n4490;
  wire _abc_43815_n4491;
  wire _abc_43815_n4492;
  wire _abc_43815_n4493;
  wire _abc_43815_n4494;
  wire _abc_43815_n4495;
  wire _abc_43815_n4496;
  wire _abc_43815_n4497;
  wire _abc_43815_n4498;
  wire _abc_43815_n4499;
  wire _abc_43815_n4500;
  wire _abc_43815_n4501;
  wire _abc_43815_n4502;
  wire _abc_43815_n4503;
  wire _abc_43815_n4504;
  wire _abc_43815_n4506;
  wire _abc_43815_n4507;
  wire _abc_43815_n4508;
  wire _abc_43815_n4509;
  wire _abc_43815_n4510;
  wire _abc_43815_n4511;
  wire _abc_43815_n4512;
  wire _abc_43815_n4513;
  wire _abc_43815_n4514;
  wire _abc_43815_n4515;
  wire _abc_43815_n4516;
  wire _abc_43815_n4517;
  wire _abc_43815_n4518;
  wire _abc_43815_n4519;
  wire _abc_43815_n4522;
  wire _abc_43815_n4524;
  wire _abc_43815_n617;
  wire _abc_43815_n618;
  wire _abc_43815_n619;
  wire _abc_43815_n621;
  wire _abc_43815_n622;
  wire _abc_43815_n623;
  wire _abc_43815_n624_1;
  wire _abc_43815_n625;
  wire _abc_43815_n626;
  wire _abc_43815_n627_1;
  wire _abc_43815_n628;
  wire _abc_43815_n629;
  wire _abc_43815_n630;
  wire _abc_43815_n631;
  wire _abc_43815_n632;
  wire _abc_43815_n634;
  wire _abc_43815_n635;
  wire _abc_43815_n636;
  wire _abc_43815_n637;
  wire _abc_43815_n638;
  wire _abc_43815_n639;
  wire _abc_43815_n640;
  wire _abc_43815_n641;
  wire _abc_43815_n641_bF_buf0;
  wire _abc_43815_n641_bF_buf1;
  wire _abc_43815_n641_bF_buf2;
  wire _abc_43815_n641_bF_buf3;
  wire _abc_43815_n642_1;
  wire _abc_43815_n642_1_bF_buf0;
  wire _abc_43815_n642_1_bF_buf1;
  wire _abc_43815_n642_1_bF_buf2;
  wire _abc_43815_n642_1_bF_buf3;
  wire _abc_43815_n642_1_bF_buf4;
  wire _abc_43815_n642_1_bF_buf5;
  wire _abc_43815_n643_1;
  wire _abc_43815_n644;
  wire _abc_43815_n645_1;
  wire _abc_43815_n645_1_bF_buf0;
  wire _abc_43815_n645_1_bF_buf1;
  wire _abc_43815_n645_1_bF_buf2;
  wire _abc_43815_n645_1_bF_buf3;
  wire _abc_43815_n645_1_bF_buf4;
  wire _abc_43815_n646_1;
  wire _abc_43815_n646_1_bF_buf0;
  wire _abc_43815_n646_1_bF_buf1;
  wire _abc_43815_n646_1_bF_buf2;
  wire _abc_43815_n646_1_bF_buf3;
  wire _abc_43815_n647_1;
  wire _abc_43815_n648;
  wire _abc_43815_n649;
  wire _abc_43815_n649_bF_buf0;
  wire _abc_43815_n649_bF_buf1;
  wire _abc_43815_n649_bF_buf2;
  wire _abc_43815_n649_bF_buf3;
  wire _abc_43815_n649_bF_buf4;
  wire _abc_43815_n650;
  wire _abc_43815_n650_bF_buf0;
  wire _abc_43815_n650_bF_buf1;
  wire _abc_43815_n650_bF_buf2;
  wire _abc_43815_n650_bF_buf3;
  wire _abc_43815_n650_bF_buf4;
  wire _abc_43815_n651_1;
  wire _abc_43815_n652;
  wire _abc_43815_n653;
  wire _abc_43815_n654;
  wire _abc_43815_n655;
  wire _abc_43815_n656;
  wire _abc_43815_n657;
  wire _abc_43815_n658;
  wire _abc_43815_n659;
  wire _abc_43815_n660;
  wire _abc_43815_n661;
  wire _abc_43815_n662;
  wire _abc_43815_n663;
  wire _abc_43815_n664_1;
  wire _abc_43815_n665;
  wire _abc_43815_n666;
  wire _abc_43815_n667;
  wire _abc_43815_n668;
  wire _abc_43815_n669;
  wire _abc_43815_n670_1;
  wire _abc_43815_n671;
  wire _abc_43815_n671_bF_buf0;
  wire _abc_43815_n671_bF_buf1;
  wire _abc_43815_n671_bF_buf2;
  wire _abc_43815_n671_bF_buf3;
  wire _abc_43815_n671_bF_buf4;
  wire _abc_43815_n672;
  wire _abc_43815_n674_1;
  wire _abc_43815_n675;
  wire _abc_43815_n677;
  wire _abc_43815_n678;
  wire _abc_43815_n679_1;
  wire _abc_43815_n680_1;
  wire _abc_43815_n680_1_bF_buf0;
  wire _abc_43815_n680_1_bF_buf1;
  wire _abc_43815_n680_1_bF_buf2;
  wire _abc_43815_n680_1_bF_buf3;
  wire _abc_43815_n680_1_bF_buf4;
  wire _abc_43815_n682;
  wire _abc_43815_n683;
  wire _abc_43815_n684;
  wire _abc_43815_n685;
  wire _abc_43815_n686_1;
  wire _abc_43815_n686_1_bF_buf0;
  wire _abc_43815_n686_1_bF_buf1;
  wire _abc_43815_n686_1_bF_buf2;
  wire _abc_43815_n686_1_bF_buf3;
  wire _abc_43815_n686_1_bF_buf4;
  wire _abc_43815_n687;
  wire _abc_43815_n688;
  wire _abc_43815_n689;
  wire _abc_43815_n690;
  wire _abc_43815_n691;
  wire _abc_43815_n692;
  wire _abc_43815_n692_bF_buf0;
  wire _abc_43815_n692_bF_buf1;
  wire _abc_43815_n692_bF_buf2;
  wire _abc_43815_n692_bF_buf3;
  wire _abc_43815_n693;
  wire _abc_43815_n694;
  wire _abc_43815_n695;
  wire _abc_43815_n696;
  wire _abc_43815_n697;
  wire _abc_43815_n698;
  wire _abc_43815_n699;
  wire _abc_43815_n700;
  wire _abc_43815_n701;
  wire _abc_43815_n702;
  wire _abc_43815_n703;
  wire _abc_43815_n704;
  wire _abc_43815_n705;
  wire _abc_43815_n706_1;
  wire _abc_43815_n707_1;
  wire _abc_43815_n708;
  wire _abc_43815_n709;
  wire _abc_43815_n710;
  wire _abc_43815_n711;
  wire _abc_43815_n712;
  wire _abc_43815_n714;
  wire _abc_43815_n715;
  wire _abc_43815_n716;
  wire _abc_43815_n717;
  wire _abc_43815_n718;
  wire _abc_43815_n719;
  wire _abc_43815_n720;
  wire _abc_43815_n721;
  wire _abc_43815_n722;
  wire _abc_43815_n723;
  wire _abc_43815_n724;
  wire _abc_43815_n725;
  wire _abc_43815_n726;
  wire _abc_43815_n727;
  wire _abc_43815_n728;
  wire _abc_43815_n730_1;
  wire _abc_43815_n731;
  wire _abc_43815_n732;
  wire _abc_43815_n733_1;
  wire _abc_43815_n734;
  wire _abc_43815_n735;
  wire _abc_43815_n736;
  wire _abc_43815_n737;
  wire _abc_43815_n738;
  wire _abc_43815_n739;
  wire _abc_43815_n740;
  wire _abc_43815_n741;
  wire _abc_43815_n742;
  wire _abc_43815_n743;
  wire _abc_43815_n744;
  wire _abc_43815_n746;
  wire _abc_43815_n747;
  wire _abc_43815_n748;
  wire _abc_43815_n749;
  wire _abc_43815_n750;
  wire _abc_43815_n751;
  wire _abc_43815_n752;
  wire _abc_43815_n753_1;
  wire _abc_43815_n754_1;
  wire _abc_43815_n755;
  wire _abc_43815_n756;
  wire _abc_43815_n757;
  wire _abc_43815_n758;
  wire _abc_43815_n759;
  wire _abc_43815_n760_1;
  wire _abc_43815_n762;
  wire _abc_43815_n763;
  wire _abc_43815_n764;
  wire _abc_43815_n765_1;
  wire _abc_43815_n766;
  wire _abc_43815_n767;
  wire _abc_43815_n768;
  wire _abc_43815_n769;
  wire _abc_43815_n770;
  wire _abc_43815_n771;
  wire _abc_43815_n772;
  wire _abc_43815_n773;
  wire _abc_43815_n774;
  wire _abc_43815_n775;
  wire _abc_43815_n776;
  wire _abc_43815_n778;
  wire _abc_43815_n779;
  wire _abc_43815_n780;
  wire _abc_43815_n781_1;
  wire _abc_43815_n782_1;
  wire _abc_43815_n783;
  wire _abc_43815_n784;
  wire _abc_43815_n785;
  wire _abc_43815_n786;
  wire _abc_43815_n787;
  wire _abc_43815_n788;
  wire _abc_43815_n789;
  wire _abc_43815_n790;
  wire _abc_43815_n791;
  wire _abc_43815_n792;
  wire _abc_43815_n794;
  wire _abc_43815_n795_1;
  wire _abc_43815_n796;
  wire _abc_43815_n797;
  wire _abc_43815_n798;
  wire _abc_43815_n799;
  wire _abc_43815_n800_1;
  wire _abc_43815_n801;
  wire _abc_43815_n802;
  wire _abc_43815_n803;
  wire _abc_43815_n804;
  wire _abc_43815_n805;
  wire _abc_43815_n806;
  wire _abc_43815_n807;
  wire _abc_43815_n808;
  wire _abc_43815_n810;
  wire _abc_43815_n811;
  wire _abc_43815_n812;
  wire _abc_43815_n813;
  wire _abc_43815_n814;
  wire _abc_43815_n815;
  wire _abc_43815_n816_1;
  wire _abc_43815_n817_1;
  wire _abc_43815_n818;
  wire _abc_43815_n819;
  wire _abc_43815_n820;
  wire _abc_43815_n821;
  wire _abc_43815_n822;
  wire _abc_43815_n823;
  wire _abc_43815_n824;
  wire _abc_43815_n826;
  wire _abc_43815_n827;
  wire _abc_43815_n828;
  wire _abc_43815_n829_1;
  wire _abc_43815_n830;
  wire _abc_43815_n831;
  wire _abc_43815_n832_1;
  wire _abc_43815_n832_1_bF_buf0;
  wire _abc_43815_n832_1_bF_buf1;
  wire _abc_43815_n832_1_bF_buf2;
  wire _abc_43815_n832_1_bF_buf3;
  wire _abc_43815_n833;
  wire _abc_43815_n835;
  wire _abc_43815_n836;
  wire _abc_43815_n837;
  wire _abc_43815_n838;
  wire _abc_43815_n839;
  wire _abc_43815_n840;
  wire _abc_43815_n842;
  wire _abc_43815_n843;
  wire _abc_43815_n844;
  wire _abc_43815_n845;
  wire _abc_43815_n846;
  wire _abc_43815_n847;
  wire _abc_43815_n849_1;
  wire _abc_43815_n850;
  wire _abc_43815_n851;
  wire _abc_43815_n852;
  wire _abc_43815_n853;
  wire _abc_43815_n854;
  wire _abc_43815_n856;
  wire _abc_43815_n857;
  wire _abc_43815_n858;
  wire _abc_43815_n859;
  wire _abc_43815_n860;
  wire _abc_43815_n861;
  wire _abc_43815_n863;
  wire _abc_43815_n864;
  wire _abc_43815_n865_1;
  wire _abc_43815_n866;
  wire _abc_43815_n867;
  wire _abc_43815_n868_1;
  wire _abc_43815_n870;
  wire _abc_43815_n871;
  wire _abc_43815_n872;
  wire _abc_43815_n873;
  wire _abc_43815_n874;
  wire _abc_43815_n875;
  wire _abc_43815_n877;
  wire _abc_43815_n878;
  wire _abc_43815_n879;
  wire _abc_43815_n880;
  wire _abc_43815_n881;
  wire _abc_43815_n882;
  wire _abc_43815_n884_1;
  wire _abc_43815_n885_1;
  wire _abc_43815_n886;
  wire _abc_43815_n887;
  wire _abc_43815_n888;
  wire _abc_43815_n889;
  wire _abc_43815_n890;
  wire _abc_43815_n892;
  wire _abc_43815_n893;
  wire _abc_43815_n894;
  wire _abc_43815_n895;
  wire _abc_43815_n896;
  wire _abc_43815_n898;
  wire _abc_43815_n899;
  wire _abc_43815_n900_1;
  wire _abc_43815_n901;
  wire _abc_43815_n902;
  wire _abc_43815_n904;
  wire _abc_43815_n905;
  wire _abc_43815_n906;
  wire _abc_43815_n907;
  wire _abc_43815_n908;
  wire _abc_43815_n910;
  wire _abc_43815_n911;
  wire _abc_43815_n912;
  wire _abc_43815_n913;
  wire _abc_43815_n914;
  wire _abc_43815_n916_1;
  wire _abc_43815_n917_1;
  wire _abc_43815_n918;
  wire _abc_43815_n919;
  wire _abc_43815_n920;
  wire _abc_43815_n922;
  wire _abc_43815_n923;
  wire _abc_43815_n924;
  wire _abc_43815_n925;
  wire _abc_43815_n926;
  wire _abc_43815_n928;
  wire _abc_43815_n929;
  wire _abc_43815_n930;
  wire _abc_43815_n931;
  wire _abc_43815_n932;
  wire _abc_43815_n934_1;
  wire _abc_43815_n935;
  wire _abc_43815_n936;
  wire _abc_43815_n937_1;
  wire _abc_43815_n938;
  wire _abc_43815_n940;
  wire _abc_43815_n941;
  wire _abc_43815_n942;
  wire _abc_43815_n943;
  wire _abc_43815_n944;
  wire _abc_43815_n946;
  wire _abc_43815_n947;
  wire _abc_43815_n948;
  wire _abc_43815_n949;
  wire _abc_43815_n950;
  wire _abc_43815_n952;
  wire _abc_43815_n953;
  wire _abc_43815_n954;
  wire _abc_43815_n955_1;
  wire _abc_43815_n956_1;
  wire _abc_43815_n958;
  wire _abc_43815_n959;
  wire _abc_43815_n960;
  wire _abc_43815_n961;
  wire _abc_43815_n962;
  wire _abc_43815_n964_1;
  wire _abc_43815_n965;
  wire _abc_43815_n966;
  wire _abc_43815_n967;
  wire _abc_43815_n968;
  wire _abc_43815_n970;
  wire _abc_43815_n971;
  wire _abc_43815_n972;
  wire _abc_43815_n973;
  wire _abc_43815_n974;
  wire _abc_43815_n976;
  wire _abc_43815_n977;
  wire _abc_43815_n978;
  wire _abc_43815_n979;
  wire _abc_43815_n980;
  wire _abc_43815_n983;
  wire _abc_43815_n984;
  wire _abc_43815_n985;
  wire _abc_43815_n986;
  wire _abc_43815_n986_bF_buf0;
  wire _abc_43815_n986_bF_buf1;
  wire _abc_43815_n986_bF_buf2;
  wire _abc_43815_n986_bF_buf3;
  wire _abc_43815_n986_bF_buf4;
  wire _abc_43815_n987;
  wire _abc_43815_n988;
  wire _abc_43815_n989;
  wire _abc_43815_n990;
  wire _abc_43815_n991;
  wire _abc_43815_n992;
  wire _abc_43815_n993_1;
  wire _abc_43815_n994_1;
  wire _abc_43815_n995;
  wire _abc_43815_n996;
  wire _abc_43815_n997;
  wire _abc_43815_n998;
  wire _abc_43815_n999;
  wire _auto_iopadmap_cc_313_execute_47726;
  wire _auto_iopadmap_cc_313_execute_47728;
  wire _auto_iopadmap_cc_313_execute_47730_0_;
  wire _auto_iopadmap_cc_313_execute_47730_10_;
  wire _auto_iopadmap_cc_313_execute_47730_11_;
  wire _auto_iopadmap_cc_313_execute_47730_12_;
  wire _auto_iopadmap_cc_313_execute_47730_13_;
  wire _auto_iopadmap_cc_313_execute_47730_14_;
  wire _auto_iopadmap_cc_313_execute_47730_15_;
  wire _auto_iopadmap_cc_313_execute_47730_16_;
  wire _auto_iopadmap_cc_313_execute_47730_17_;
  wire _auto_iopadmap_cc_313_execute_47730_18_;
  wire _auto_iopadmap_cc_313_execute_47730_19_;
  wire _auto_iopadmap_cc_313_execute_47730_1_;
  wire _auto_iopadmap_cc_313_execute_47730_20_;
  wire _auto_iopadmap_cc_313_execute_47730_21_;
  wire _auto_iopadmap_cc_313_execute_47730_22_;
  wire _auto_iopadmap_cc_313_execute_47730_23_;
  wire _auto_iopadmap_cc_313_execute_47730_24_;
  wire _auto_iopadmap_cc_313_execute_47730_25_;
  wire _auto_iopadmap_cc_313_execute_47730_26_;
  wire _auto_iopadmap_cc_313_execute_47730_27_;
  wire _auto_iopadmap_cc_313_execute_47730_28_;
  wire _auto_iopadmap_cc_313_execute_47730_29_;
  wire _auto_iopadmap_cc_313_execute_47730_2_;
  wire _auto_iopadmap_cc_313_execute_47730_30_;
  wire _auto_iopadmap_cc_313_execute_47730_31_;
  wire _auto_iopadmap_cc_313_execute_47730_3_;
  wire _auto_iopadmap_cc_313_execute_47730_4_;
  wire _auto_iopadmap_cc_313_execute_47730_5_;
  wire _auto_iopadmap_cc_313_execute_47730_6_;
  wire _auto_iopadmap_cc_313_execute_47730_7_;
  wire _auto_iopadmap_cc_313_execute_47730_8_;
  wire _auto_iopadmap_cc_313_execute_47730_9_;
  wire _auto_iopadmap_cc_313_execute_47767;
  wire _auto_iopadmap_cc_313_execute_47769_0_;
  wire _auto_iopadmap_cc_313_execute_47769_10_;
  wire _auto_iopadmap_cc_313_execute_47769_11_;
  wire _auto_iopadmap_cc_313_execute_47769_12_;
  wire _auto_iopadmap_cc_313_execute_47769_13_;
  wire _auto_iopadmap_cc_313_execute_47769_14_;
  wire _auto_iopadmap_cc_313_execute_47769_15_;
  wire _auto_iopadmap_cc_313_execute_47769_16_;
  wire _auto_iopadmap_cc_313_execute_47769_17_;
  wire _auto_iopadmap_cc_313_execute_47769_18_;
  wire _auto_iopadmap_cc_313_execute_47769_19_;
  wire _auto_iopadmap_cc_313_execute_47769_1_;
  wire _auto_iopadmap_cc_313_execute_47769_20_;
  wire _auto_iopadmap_cc_313_execute_47769_21_;
  wire _auto_iopadmap_cc_313_execute_47769_22_;
  wire _auto_iopadmap_cc_313_execute_47769_23_;
  wire _auto_iopadmap_cc_313_execute_47769_24_;
  wire _auto_iopadmap_cc_313_execute_47769_25_;
  wire _auto_iopadmap_cc_313_execute_47769_26_;
  wire _auto_iopadmap_cc_313_execute_47769_27_;
  wire _auto_iopadmap_cc_313_execute_47769_28_;
  wire _auto_iopadmap_cc_313_execute_47769_29_;
  wire _auto_iopadmap_cc_313_execute_47769_2_;
  wire _auto_iopadmap_cc_313_execute_47769_30_;
  wire _auto_iopadmap_cc_313_execute_47769_31_;
  wire _auto_iopadmap_cc_313_execute_47769_3_;
  wire _auto_iopadmap_cc_313_execute_47769_4_;
  wire _auto_iopadmap_cc_313_execute_47769_5_;
  wire _auto_iopadmap_cc_313_execute_47769_6_;
  wire _auto_iopadmap_cc_313_execute_47769_7_;
  wire _auto_iopadmap_cc_313_execute_47769_8_;
  wire _auto_iopadmap_cc_313_execute_47769_9_;
  wire _auto_iopadmap_cc_313_execute_47802_0_;
  wire _auto_iopadmap_cc_313_execute_47802_1_;
  wire _auto_iopadmap_cc_313_execute_47802_2_;
  wire _auto_iopadmap_cc_313_execute_47802_3_;
  wire _auto_iopadmap_cc_313_execute_47807;
  wire _auto_iopadmap_cc_313_execute_47809;
  wire alu__abc_41358_n1000;
  wire alu__abc_41358_n1001_1;
  wire alu__abc_41358_n1002;
  wire alu__abc_41358_n1003;
  wire alu__abc_41358_n1004;
  wire alu__abc_41358_n1005;
  wire alu__abc_41358_n1006;
  wire alu__abc_41358_n1007;
  wire alu__abc_41358_n1008;
  wire alu__abc_41358_n1009;
  wire alu__abc_41358_n1010;
  wire alu__abc_41358_n1011;
  wire alu__abc_41358_n1012;
  wire alu__abc_41358_n1013;
  wire alu__abc_41358_n1014;
  wire alu__abc_41358_n1015;
  wire alu__abc_41358_n1016;
  wire alu__abc_41358_n1017;
  wire alu__abc_41358_n1018;
  wire alu__abc_41358_n1019;
  wire alu__abc_41358_n1020;
  wire alu__abc_41358_n1021;
  wire alu__abc_41358_n1022;
  wire alu__abc_41358_n1023;
  wire alu__abc_41358_n1024_1;
  wire alu__abc_41358_n1025;
  wire alu__abc_41358_n1026;
  wire alu__abc_41358_n1027;
  wire alu__abc_41358_n1028;
  wire alu__abc_41358_n1029;
  wire alu__abc_41358_n1030;
  wire alu__abc_41358_n1031;
  wire alu__abc_41358_n1032;
  wire alu__abc_41358_n1033;
  wire alu__abc_41358_n1034;
  wire alu__abc_41358_n1035;
  wire alu__abc_41358_n1036;
  wire alu__abc_41358_n1037;
  wire alu__abc_41358_n1038;
  wire alu__abc_41358_n1039;
  wire alu__abc_41358_n1040;
  wire alu__abc_41358_n1041;
  wire alu__abc_41358_n1042;
  wire alu__abc_41358_n1043;
  wire alu__abc_41358_n1044;
  wire alu__abc_41358_n1045;
  wire alu__abc_41358_n1046;
  wire alu__abc_41358_n1047;
  wire alu__abc_41358_n1048;
  wire alu__abc_41358_n1049;
  wire alu__abc_41358_n1050_1;
  wire alu__abc_41358_n1051;
  wire alu__abc_41358_n1052;
  wire alu__abc_41358_n1053;
  wire alu__abc_41358_n1054;
  wire alu__abc_41358_n1055;
  wire alu__abc_41358_n1056;
  wire alu__abc_41358_n1057;
  wire alu__abc_41358_n1057_bF_buf0;
  wire alu__abc_41358_n1057_bF_buf1;
  wire alu__abc_41358_n1057_bF_buf2;
  wire alu__abc_41358_n1057_bF_buf3;
  wire alu__abc_41358_n1057_bF_buf4;
  wire alu__abc_41358_n1058;
  wire alu__abc_41358_n1059;
  wire alu__abc_41358_n1060;
  wire alu__abc_41358_n1061;
  wire alu__abc_41358_n1061_bF_buf0;
  wire alu__abc_41358_n1061_bF_buf1;
  wire alu__abc_41358_n1061_bF_buf2;
  wire alu__abc_41358_n1061_bF_buf3;
  wire alu__abc_41358_n1061_bF_buf4;
  wire alu__abc_41358_n1062;
  wire alu__abc_41358_n1063;
  wire alu__abc_41358_n1064;
  wire alu__abc_41358_n1065;
  wire alu__abc_41358_n1066;
  wire alu__abc_41358_n1067;
  wire alu__abc_41358_n1068;
  wire alu__abc_41358_n1069;
  wire alu__abc_41358_n1070;
  wire alu__abc_41358_n1071;
  wire alu__abc_41358_n1072;
  wire alu__abc_41358_n1073;
  wire alu__abc_41358_n1074_1;
  wire alu__abc_41358_n1075;
  wire alu__abc_41358_n1076;
  wire alu__abc_41358_n1077;
  wire alu__abc_41358_n1078;
  wire alu__abc_41358_n1079;
  wire alu__abc_41358_n1080;
  wire alu__abc_41358_n1081;
  wire alu__abc_41358_n1082;
  wire alu__abc_41358_n1083;
  wire alu__abc_41358_n1084;
  wire alu__abc_41358_n1086;
  wire alu__abc_41358_n1087;
  wire alu__abc_41358_n1088;
  wire alu__abc_41358_n1089;
  wire alu__abc_41358_n1090;
  wire alu__abc_41358_n1091;
  wire alu__abc_41358_n1092;
  wire alu__abc_41358_n1093;
  wire alu__abc_41358_n1094;
  wire alu__abc_41358_n1095;
  wire alu__abc_41358_n1096;
  wire alu__abc_41358_n1097_1;
  wire alu__abc_41358_n1098;
  wire alu__abc_41358_n1099;
  wire alu__abc_41358_n110;
  wire alu__abc_41358_n1100;
  wire alu__abc_41358_n1101;
  wire alu__abc_41358_n1102;
  wire alu__abc_41358_n1103;
  wire alu__abc_41358_n1104;
  wire alu__abc_41358_n1105;
  wire alu__abc_41358_n1106;
  wire alu__abc_41358_n1107;
  wire alu__abc_41358_n1108;
  wire alu__abc_41358_n1109;
  wire alu__abc_41358_n111;
  wire alu__abc_41358_n1110;
  wire alu__abc_41358_n1111;
  wire alu__abc_41358_n1112;
  wire alu__abc_41358_n1113;
  wire alu__abc_41358_n1114;
  wire alu__abc_41358_n1115;
  wire alu__abc_41358_n1116;
  wire alu__abc_41358_n1117_1;
  wire alu__abc_41358_n1118;
  wire alu__abc_41358_n1119;
  wire alu__abc_41358_n1120;
  wire alu__abc_41358_n1121;
  wire alu__abc_41358_n1122;
  wire alu__abc_41358_n1123;
  wire alu__abc_41358_n1124;
  wire alu__abc_41358_n1125;
  wire alu__abc_41358_n1126;
  wire alu__abc_41358_n1127;
  wire alu__abc_41358_n1128;
  wire alu__abc_41358_n1129;
  wire alu__abc_41358_n112_1;
  wire alu__abc_41358_n1130;
  wire alu__abc_41358_n1131;
  wire alu__abc_41358_n1132;
  wire alu__abc_41358_n1133;
  wire alu__abc_41358_n1134;
  wire alu__abc_41358_n1135;
  wire alu__abc_41358_n1136;
  wire alu__abc_41358_n1137_1;
  wire alu__abc_41358_n1138;
  wire alu__abc_41358_n1139;
  wire alu__abc_41358_n113_1;
  wire alu__abc_41358_n114;
  wire alu__abc_41358_n1140;
  wire alu__abc_41358_n1141;
  wire alu__abc_41358_n1142;
  wire alu__abc_41358_n1143;
  wire alu__abc_41358_n1144;
  wire alu__abc_41358_n1145;
  wire alu__abc_41358_n1146;
  wire alu__abc_41358_n1147;
  wire alu__abc_41358_n1148;
  wire alu__abc_41358_n1149;
  wire alu__abc_41358_n115;
  wire alu__abc_41358_n1150;
  wire alu__abc_41358_n1151;
  wire alu__abc_41358_n1152;
  wire alu__abc_41358_n1153;
  wire alu__abc_41358_n1154;
  wire alu__abc_41358_n1155;
  wire alu__abc_41358_n1156;
  wire alu__abc_41358_n1157;
  wire alu__abc_41358_n1158_1;
  wire alu__abc_41358_n1159;
  wire alu__abc_41358_n116;
  wire alu__abc_41358_n1160;
  wire alu__abc_41358_n1161;
  wire alu__abc_41358_n1163;
  wire alu__abc_41358_n1164;
  wire alu__abc_41358_n1165;
  wire alu__abc_41358_n1166;
  wire alu__abc_41358_n1167;
  wire alu__abc_41358_n1168;
  wire alu__abc_41358_n1169;
  wire alu__abc_41358_n117;
  wire alu__abc_41358_n1170;
  wire alu__abc_41358_n1171;
  wire alu__abc_41358_n1172;
  wire alu__abc_41358_n1173;
  wire alu__abc_41358_n1174;
  wire alu__abc_41358_n1175;
  wire alu__abc_41358_n1176;
  wire alu__abc_41358_n1177;
  wire alu__abc_41358_n1178;
  wire alu__abc_41358_n1179;
  wire alu__abc_41358_n118;
  wire alu__abc_41358_n1180;
  wire alu__abc_41358_n1181_1;
  wire alu__abc_41358_n1182;
  wire alu__abc_41358_n1183;
  wire alu__abc_41358_n1184;
  wire alu__abc_41358_n1185;
  wire alu__abc_41358_n1186;
  wire alu__abc_41358_n1187;
  wire alu__abc_41358_n1188;
  wire alu__abc_41358_n1189;
  wire alu__abc_41358_n1190;
  wire alu__abc_41358_n1191;
  wire alu__abc_41358_n1192;
  wire alu__abc_41358_n1193;
  wire alu__abc_41358_n1194;
  wire alu__abc_41358_n1195;
  wire alu__abc_41358_n1196;
  wire alu__abc_41358_n1197;
  wire alu__abc_41358_n1198;
  wire alu__abc_41358_n1199;
  wire alu__abc_41358_n119_1;
  wire alu__abc_41358_n1200;
  wire alu__abc_41358_n1201;
  wire alu__abc_41358_n1202_1;
  wire alu__abc_41358_n1203;
  wire alu__abc_41358_n1204;
  wire alu__abc_41358_n1205;
  wire alu__abc_41358_n1206;
  wire alu__abc_41358_n1207;
  wire alu__abc_41358_n1208;
  wire alu__abc_41358_n1209;
  wire alu__abc_41358_n120_1;
  wire alu__abc_41358_n121;
  wire alu__abc_41358_n1210;
  wire alu__abc_41358_n1211;
  wire alu__abc_41358_n1212;
  wire alu__abc_41358_n1213;
  wire alu__abc_41358_n1214;
  wire alu__abc_41358_n1215;
  wire alu__abc_41358_n1216;
  wire alu__abc_41358_n1217;
  wire alu__abc_41358_n1218;
  wire alu__abc_41358_n1219;
  wire alu__abc_41358_n122;
  wire alu__abc_41358_n1220;
  wire alu__abc_41358_n1221;
  wire alu__abc_41358_n1222;
  wire alu__abc_41358_n1223_1;
  wire alu__abc_41358_n1224;
  wire alu__abc_41358_n1225;
  wire alu__abc_41358_n1226;
  wire alu__abc_41358_n1227;
  wire alu__abc_41358_n1228;
  wire alu__abc_41358_n1229;
  wire alu__abc_41358_n123;
  wire alu__abc_41358_n1230;
  wire alu__abc_41358_n1231;
  wire alu__abc_41358_n1232;
  wire alu__abc_41358_n1233;
  wire alu__abc_41358_n1234;
  wire alu__abc_41358_n1235;
  wire alu__abc_41358_n1236;
  wire alu__abc_41358_n1237;
  wire alu__abc_41358_n1239;
  wire alu__abc_41358_n1240;
  wire alu__abc_41358_n1241;
  wire alu__abc_41358_n1242;
  wire alu__abc_41358_n1243_1;
  wire alu__abc_41358_n1244;
  wire alu__abc_41358_n1245;
  wire alu__abc_41358_n1246;
  wire alu__abc_41358_n1247;
  wire alu__abc_41358_n1248;
  wire alu__abc_41358_n1249;
  wire alu__abc_41358_n124_1;
  wire alu__abc_41358_n1250;
  wire alu__abc_41358_n1251;
  wire alu__abc_41358_n1252;
  wire alu__abc_41358_n1253;
  wire alu__abc_41358_n1254;
  wire alu__abc_41358_n1255;
  wire alu__abc_41358_n1256;
  wire alu__abc_41358_n1257;
  wire alu__abc_41358_n1258;
  wire alu__abc_41358_n1259;
  wire alu__abc_41358_n125_1;
  wire alu__abc_41358_n126;
  wire alu__abc_41358_n1260;
  wire alu__abc_41358_n1261;
  wire alu__abc_41358_n1262;
  wire alu__abc_41358_n1263;
  wire alu__abc_41358_n1264_1;
  wire alu__abc_41358_n1265;
  wire alu__abc_41358_n1266;
  wire alu__abc_41358_n1267;
  wire alu__abc_41358_n1268;
  wire alu__abc_41358_n1269;
  wire alu__abc_41358_n127;
  wire alu__abc_41358_n1270;
  wire alu__abc_41358_n1271;
  wire alu__abc_41358_n1272;
  wire alu__abc_41358_n1273;
  wire alu__abc_41358_n1274;
  wire alu__abc_41358_n1275;
  wire alu__abc_41358_n1276;
  wire alu__abc_41358_n1277;
  wire alu__abc_41358_n1278;
  wire alu__abc_41358_n1279;
  wire alu__abc_41358_n128;
  wire alu__abc_41358_n1280;
  wire alu__abc_41358_n1281;
  wire alu__abc_41358_n1282;
  wire alu__abc_41358_n1283;
  wire alu__abc_41358_n1284_1;
  wire alu__abc_41358_n1285;
  wire alu__abc_41358_n1286;
  wire alu__abc_41358_n1287;
  wire alu__abc_41358_n1288;
  wire alu__abc_41358_n1289;
  wire alu__abc_41358_n129;
  wire alu__abc_41358_n1290;
  wire alu__abc_41358_n1292;
  wire alu__abc_41358_n1293;
  wire alu__abc_41358_n1294;
  wire alu__abc_41358_n1295;
  wire alu__abc_41358_n1296;
  wire alu__abc_41358_n1297;
  wire alu__abc_41358_n1298;
  wire alu__abc_41358_n1299;
  wire alu__abc_41358_n1300;
  wire alu__abc_41358_n1301;
  wire alu__abc_41358_n1302;
  wire alu__abc_41358_n1303;
  wire alu__abc_41358_n1304_1;
  wire alu__abc_41358_n1305;
  wire alu__abc_41358_n1306;
  wire alu__abc_41358_n1307;
  wire alu__abc_41358_n1308;
  wire alu__abc_41358_n1309;
  wire alu__abc_41358_n130_1;
  wire alu__abc_41358_n1310;
  wire alu__abc_41358_n1311;
  wire alu__abc_41358_n1312;
  wire alu__abc_41358_n1313;
  wire alu__abc_41358_n1314;
  wire alu__abc_41358_n1315;
  wire alu__abc_41358_n1316;
  wire alu__abc_41358_n1317;
  wire alu__abc_41358_n1318;
  wire alu__abc_41358_n1319;
  wire alu__abc_41358_n131_1;
  wire alu__abc_41358_n132;
  wire alu__abc_41358_n1320;
  wire alu__abc_41358_n1321;
  wire alu__abc_41358_n1322;
  wire alu__abc_41358_n1323_1;
  wire alu__abc_41358_n1324;
  wire alu__abc_41358_n1325;
  wire alu__abc_41358_n1326;
  wire alu__abc_41358_n1327;
  wire alu__abc_41358_n1328;
  wire alu__abc_41358_n1329;
  wire alu__abc_41358_n133;
  wire alu__abc_41358_n1330;
  wire alu__abc_41358_n1331;
  wire alu__abc_41358_n1332;
  wire alu__abc_41358_n1333;
  wire alu__abc_41358_n1334;
  wire alu__abc_41358_n1335;
  wire alu__abc_41358_n1336;
  wire alu__abc_41358_n1337;
  wire alu__abc_41358_n1338;
  wire alu__abc_41358_n1339;
  wire alu__abc_41358_n134;
  wire alu__abc_41358_n1340;
  wire alu__abc_41358_n1341;
  wire alu__abc_41358_n1342;
  wire alu__abc_41358_n1343;
  wire alu__abc_41358_n1344_1;
  wire alu__abc_41358_n1346;
  wire alu__abc_41358_n1347;
  wire alu__abc_41358_n1348;
  wire alu__abc_41358_n1349;
  wire alu__abc_41358_n1350;
  wire alu__abc_41358_n1351;
  wire alu__abc_41358_n1352;
  wire alu__abc_41358_n1353;
  wire alu__abc_41358_n1354;
  wire alu__abc_41358_n1355;
  wire alu__abc_41358_n1356;
  wire alu__abc_41358_n1357;
  wire alu__abc_41358_n1358;
  wire alu__abc_41358_n1359;
  wire alu__abc_41358_n135_1;
  wire alu__abc_41358_n1360;
  wire alu__abc_41358_n1361;
  wire alu__abc_41358_n1362_1;
  wire alu__abc_41358_n1363;
  wire alu__abc_41358_n1364;
  wire alu__abc_41358_n1365;
  wire alu__abc_41358_n1366;
  wire alu__abc_41358_n1367;
  wire alu__abc_41358_n1368;
  wire alu__abc_41358_n1369;
  wire alu__abc_41358_n136_1;
  wire alu__abc_41358_n137;
  wire alu__abc_41358_n1370;
  wire alu__abc_41358_n1371;
  wire alu__abc_41358_n1372;
  wire alu__abc_41358_n1373;
  wire alu__abc_41358_n1374;
  wire alu__abc_41358_n1375;
  wire alu__abc_41358_n1376;
  wire alu__abc_41358_n1377;
  wire alu__abc_41358_n1378;
  wire alu__abc_41358_n1379;
  wire alu__abc_41358_n138;
  wire alu__abc_41358_n1380;
  wire alu__abc_41358_n1381;
  wire alu__abc_41358_n1382_1;
  wire alu__abc_41358_n1383;
  wire alu__abc_41358_n1384;
  wire alu__abc_41358_n1385;
  wire alu__abc_41358_n1386;
  wire alu__abc_41358_n1387;
  wire alu__abc_41358_n1388;
  wire alu__abc_41358_n1389;
  wire alu__abc_41358_n139;
  wire alu__abc_41358_n1390;
  wire alu__abc_41358_n1391;
  wire alu__abc_41358_n1392;
  wire alu__abc_41358_n1393;
  wire alu__abc_41358_n1394;
  wire alu__abc_41358_n1395;
  wire alu__abc_41358_n1396;
  wire alu__abc_41358_n1398;
  wire alu__abc_41358_n1399;
  wire alu__abc_41358_n140;
  wire alu__abc_41358_n1400;
  wire alu__abc_41358_n1401_1;
  wire alu__abc_41358_n1402;
  wire alu__abc_41358_n1403;
  wire alu__abc_41358_n1404;
  wire alu__abc_41358_n1405;
  wire alu__abc_41358_n1406;
  wire alu__abc_41358_n1407;
  wire alu__abc_41358_n1408;
  wire alu__abc_41358_n1409;
  wire alu__abc_41358_n141;
  wire alu__abc_41358_n1410;
  wire alu__abc_41358_n1411;
  wire alu__abc_41358_n1412;
  wire alu__abc_41358_n1413;
  wire alu__abc_41358_n1414;
  wire alu__abc_41358_n1415;
  wire alu__abc_41358_n1416;
  wire alu__abc_41358_n1417;
  wire alu__abc_41358_n1418;
  wire alu__abc_41358_n1419_1;
  wire alu__abc_41358_n142;
  wire alu__abc_41358_n1420;
  wire alu__abc_41358_n1421;
  wire alu__abc_41358_n1422;
  wire alu__abc_41358_n1423;
  wire alu__abc_41358_n1424;
  wire alu__abc_41358_n1425;
  wire alu__abc_41358_n1426;
  wire alu__abc_41358_n1427;
  wire alu__abc_41358_n1428;
  wire alu__abc_41358_n1429;
  wire alu__abc_41358_n1430;
  wire alu__abc_41358_n1431;
  wire alu__abc_41358_n1432;
  wire alu__abc_41358_n1433;
  wire alu__abc_41358_n1434;
  wire alu__abc_41358_n1435_1;
  wire alu__abc_41358_n1436;
  wire alu__abc_41358_n1437;
  wire alu__abc_41358_n1438;
  wire alu__abc_41358_n1439;
  wire alu__abc_41358_n143_1;
  wire alu__abc_41358_n1440;
  wire alu__abc_41358_n1441;
  wire alu__abc_41358_n1442;
  wire alu__abc_41358_n1443;
  wire alu__abc_41358_n1444;
  wire alu__abc_41358_n1445;
  wire alu__abc_41358_n1446;
  wire alu__abc_41358_n1447;
  wire alu__abc_41358_n1448;
  wire alu__abc_41358_n1449;
  wire alu__abc_41358_n144_1;
  wire alu__abc_41358_n145;
  wire alu__abc_41358_n1450;
  wire alu__abc_41358_n1452;
  wire alu__abc_41358_n1453;
  wire alu__abc_41358_n1454;
  wire alu__abc_41358_n1455;
  wire alu__abc_41358_n1456;
  wire alu__abc_41358_n1457;
  wire alu__abc_41358_n1458;
  wire alu__abc_41358_n1459;
  wire alu__abc_41358_n146;
  wire alu__abc_41358_n1460;
  wire alu__abc_41358_n1461;
  wire alu__abc_41358_n1462;
  wire alu__abc_41358_n1463;
  wire alu__abc_41358_n1464;
  wire alu__abc_41358_n1465;
  wire alu__abc_41358_n1466;
  wire alu__abc_41358_n1467;
  wire alu__abc_41358_n1468;
  wire alu__abc_41358_n1469;
  wire alu__abc_41358_n147;
  wire alu__abc_41358_n1470;
  wire alu__abc_41358_n1471;
  wire alu__abc_41358_n1472;
  wire alu__abc_41358_n1473;
  wire alu__abc_41358_n1474;
  wire alu__abc_41358_n1475;
  wire alu__abc_41358_n1476;
  wire alu__abc_41358_n1477;
  wire alu__abc_41358_n1478;
  wire alu__abc_41358_n1479;
  wire alu__abc_41358_n1480;
  wire alu__abc_41358_n1481;
  wire alu__abc_41358_n1482;
  wire alu__abc_41358_n1483;
  wire alu__abc_41358_n1484;
  wire alu__abc_41358_n1485;
  wire alu__abc_41358_n1486;
  wire alu__abc_41358_n1487;
  wire alu__abc_41358_n1488;
  wire alu__abc_41358_n1489_1;
  wire alu__abc_41358_n148_1;
  wire alu__abc_41358_n1490_1;
  wire alu__abc_41358_n1491_1;
  wire alu__abc_41358_n1492;
  wire alu__abc_41358_n1493;
  wire alu__abc_41358_n1494;
  wire alu__abc_41358_n1496;
  wire alu__abc_41358_n1497;
  wire alu__abc_41358_n1498;
  wire alu__abc_41358_n1499;
  wire alu__abc_41358_n149_1;
  wire alu__abc_41358_n150;
  wire alu__abc_41358_n1500;
  wire alu__abc_41358_n1501;
  wire alu__abc_41358_n1502;
  wire alu__abc_41358_n1503;
  wire alu__abc_41358_n1504;
  wire alu__abc_41358_n1505;
  wire alu__abc_41358_n1506;
  wire alu__abc_41358_n1507;
  wire alu__abc_41358_n1508;
  wire alu__abc_41358_n1509;
  wire alu__abc_41358_n151;
  wire alu__abc_41358_n1510;
  wire alu__abc_41358_n1511;
  wire alu__abc_41358_n1512;
  wire alu__abc_41358_n1513;
  wire alu__abc_41358_n1514;
  wire alu__abc_41358_n1515;
  wire alu__abc_41358_n1516;
  wire alu__abc_41358_n1517;
  wire alu__abc_41358_n1518;
  wire alu__abc_41358_n1519;
  wire alu__abc_41358_n152;
  wire alu__abc_41358_n1520;
  wire alu__abc_41358_n1521;
  wire alu__abc_41358_n1522;
  wire alu__abc_41358_n1523;
  wire alu__abc_41358_n1524;
  wire alu__abc_41358_n1525;
  wire alu__abc_41358_n1526;
  wire alu__abc_41358_n1527;
  wire alu__abc_41358_n1528;
  wire alu__abc_41358_n1529;
  wire alu__abc_41358_n153;
  wire alu__abc_41358_n1530;
  wire alu__abc_41358_n1531;
  wire alu__abc_41358_n1532;
  wire alu__abc_41358_n1533;
  wire alu__abc_41358_n1534;
  wire alu__abc_41358_n1535;
  wire alu__abc_41358_n1536;
  wire alu__abc_41358_n1537;
  wire alu__abc_41358_n1538;
  wire alu__abc_41358_n1539;
  wire alu__abc_41358_n1540;
  wire alu__abc_41358_n1542;
  wire alu__abc_41358_n1543;
  wire alu__abc_41358_n1544;
  wire alu__abc_41358_n1545;
  wire alu__abc_41358_n1546;
  wire alu__abc_41358_n1547;
  wire alu__abc_41358_n1548;
  wire alu__abc_41358_n1549;
  wire alu__abc_41358_n154_1;
  wire alu__abc_41358_n1550;
  wire alu__abc_41358_n1551;
  wire alu__abc_41358_n1552;
  wire alu__abc_41358_n1553;
  wire alu__abc_41358_n1554;
  wire alu__abc_41358_n1555;
  wire alu__abc_41358_n1556;
  wire alu__abc_41358_n1557;
  wire alu__abc_41358_n1558;
  wire alu__abc_41358_n1559;
  wire alu__abc_41358_n155_1;
  wire alu__abc_41358_n156;
  wire alu__abc_41358_n1560;
  wire alu__abc_41358_n1561;
  wire alu__abc_41358_n1562;
  wire alu__abc_41358_n1563;
  wire alu__abc_41358_n1564;
  wire alu__abc_41358_n1565;
  wire alu__abc_41358_n1566;
  wire alu__abc_41358_n1567;
  wire alu__abc_41358_n1568;
  wire alu__abc_41358_n1569;
  wire alu__abc_41358_n157;
  wire alu__abc_41358_n1570;
  wire alu__abc_41358_n1571;
  wire alu__abc_41358_n1572;
  wire alu__abc_41358_n1573;
  wire alu__abc_41358_n1574;
  wire alu__abc_41358_n1575;
  wire alu__abc_41358_n1576;
  wire alu__abc_41358_n1577;
  wire alu__abc_41358_n1578;
  wire alu__abc_41358_n1579;
  wire alu__abc_41358_n158;
  wire alu__abc_41358_n1580;
  wire alu__abc_41358_n1581;
  wire alu__abc_41358_n1582;
  wire alu__abc_41358_n1583;
  wire alu__abc_41358_n1584;
  wire alu__abc_41358_n1585;
  wire alu__abc_41358_n1586;
  wire alu__abc_41358_n1588;
  wire alu__abc_41358_n1589;
  wire alu__abc_41358_n1590;
  wire alu__abc_41358_n1591;
  wire alu__abc_41358_n1592;
  wire alu__abc_41358_n1593;
  wire alu__abc_41358_n1594;
  wire alu__abc_41358_n1595;
  wire alu__abc_41358_n1596;
  wire alu__abc_41358_n1597;
  wire alu__abc_41358_n1598;
  wire alu__abc_41358_n1599;
  wire alu__abc_41358_n159_1;
  wire alu__abc_41358_n1600;
  wire alu__abc_41358_n1601;
  wire alu__abc_41358_n1602;
  wire alu__abc_41358_n1603;
  wire alu__abc_41358_n1604;
  wire alu__abc_41358_n1605;
  wire alu__abc_41358_n1606;
  wire alu__abc_41358_n1607;
  wire alu__abc_41358_n1608;
  wire alu__abc_41358_n1609;
  wire alu__abc_41358_n160_1;
  wire alu__abc_41358_n161;
  wire alu__abc_41358_n1610;
  wire alu__abc_41358_n1611;
  wire alu__abc_41358_n1612;
  wire alu__abc_41358_n1613;
  wire alu__abc_41358_n1614;
  wire alu__abc_41358_n1615;
  wire alu__abc_41358_n1616;
  wire alu__abc_41358_n1617;
  wire alu__abc_41358_n1618;
  wire alu__abc_41358_n1619;
  wire alu__abc_41358_n162;
  wire alu__abc_41358_n1620;
  wire alu__abc_41358_n1621;
  wire alu__abc_41358_n1622;
  wire alu__abc_41358_n1623;
  wire alu__abc_41358_n1624;
  wire alu__abc_41358_n1625;
  wire alu__abc_41358_n1626;
  wire alu__abc_41358_n1627;
  wire alu__abc_41358_n1628;
  wire alu__abc_41358_n1629;
  wire alu__abc_41358_n163;
  wire alu__abc_41358_n1630;
  wire alu__abc_41358_n1631;
  wire alu__abc_41358_n1633;
  wire alu__abc_41358_n1634;
  wire alu__abc_41358_n1635;
  wire alu__abc_41358_n1636;
  wire alu__abc_41358_n1637;
  wire alu__abc_41358_n1638;
  wire alu__abc_41358_n1639;
  wire alu__abc_41358_n164;
  wire alu__abc_41358_n1640;
  wire alu__abc_41358_n1641;
  wire alu__abc_41358_n1642;
  wire alu__abc_41358_n1643;
  wire alu__abc_41358_n1644;
  wire alu__abc_41358_n1645;
  wire alu__abc_41358_n1646;
  wire alu__abc_41358_n1647;
  wire alu__abc_41358_n1648;
  wire alu__abc_41358_n1649;
  wire alu__abc_41358_n165;
  wire alu__abc_41358_n1650;
  wire alu__abc_41358_n1651;
  wire alu__abc_41358_n1652;
  wire alu__abc_41358_n1653;
  wire alu__abc_41358_n1654;
  wire alu__abc_41358_n1655;
  wire alu__abc_41358_n1656;
  wire alu__abc_41358_n1657;
  wire alu__abc_41358_n1658;
  wire alu__abc_41358_n1659;
  wire alu__abc_41358_n1660;
  wire alu__abc_41358_n1661;
  wire alu__abc_41358_n1662;
  wire alu__abc_41358_n1663;
  wire alu__abc_41358_n1664;
  wire alu__abc_41358_n1665;
  wire alu__abc_41358_n1666;
  wire alu__abc_41358_n1667;
  wire alu__abc_41358_n1668;
  wire alu__abc_41358_n1669;
  wire alu__abc_41358_n166_1;
  wire alu__abc_41358_n1670;
  wire alu__abc_41358_n1671;
  wire alu__abc_41358_n1672;
  wire alu__abc_41358_n1673;
  wire alu__abc_41358_n1674;
  wire alu__abc_41358_n1675;
  wire alu__abc_41358_n1676;
  wire alu__abc_41358_n1677;
  wire alu__abc_41358_n1679;
  wire alu__abc_41358_n167_1;
  wire alu__abc_41358_n168;
  wire alu__abc_41358_n1680;
  wire alu__abc_41358_n1681;
  wire alu__abc_41358_n1682;
  wire alu__abc_41358_n1683;
  wire alu__abc_41358_n1684;
  wire alu__abc_41358_n1685;
  wire alu__abc_41358_n1686;
  wire alu__abc_41358_n1687;
  wire alu__abc_41358_n1688;
  wire alu__abc_41358_n1689;
  wire alu__abc_41358_n169;
  wire alu__abc_41358_n1690;
  wire alu__abc_41358_n1691;
  wire alu__abc_41358_n1692;
  wire alu__abc_41358_n1693;
  wire alu__abc_41358_n1694;
  wire alu__abc_41358_n1695;
  wire alu__abc_41358_n1696;
  wire alu__abc_41358_n1697;
  wire alu__abc_41358_n1698;
  wire alu__abc_41358_n1699;
  wire alu__abc_41358_n170;
  wire alu__abc_41358_n1700;
  wire alu__abc_41358_n1701;
  wire alu__abc_41358_n1702;
  wire alu__abc_41358_n1703;
  wire alu__abc_41358_n1704;
  wire alu__abc_41358_n1705;
  wire alu__abc_41358_n1706;
  wire alu__abc_41358_n1707;
  wire alu__abc_41358_n1708;
  wire alu__abc_41358_n1709;
  wire alu__abc_41358_n1710;
  wire alu__abc_41358_n1711;
  wire alu__abc_41358_n1712;
  wire alu__abc_41358_n1713;
  wire alu__abc_41358_n1714;
  wire alu__abc_41358_n1715;
  wire alu__abc_41358_n1716;
  wire alu__abc_41358_n1717;
  wire alu__abc_41358_n1718;
  wire alu__abc_41358_n1719;
  wire alu__abc_41358_n171_1;
  wire alu__abc_41358_n1720;
  wire alu__abc_41358_n1721;
  wire alu__abc_41358_n1722;
  wire alu__abc_41358_n1724;
  wire alu__abc_41358_n1725;
  wire alu__abc_41358_n1726;
  wire alu__abc_41358_n1727;
  wire alu__abc_41358_n1728;
  wire alu__abc_41358_n1729;
  wire alu__abc_41358_n172_1;
  wire alu__abc_41358_n173;
  wire alu__abc_41358_n1730;
  wire alu__abc_41358_n1731;
  wire alu__abc_41358_n1732;
  wire alu__abc_41358_n1733;
  wire alu__abc_41358_n1734;
  wire alu__abc_41358_n1735;
  wire alu__abc_41358_n1736;
  wire alu__abc_41358_n1737;
  wire alu__abc_41358_n1738;
  wire alu__abc_41358_n1739;
  wire alu__abc_41358_n174;
  wire alu__abc_41358_n1740;
  wire alu__abc_41358_n1741;
  wire alu__abc_41358_n1742;
  wire alu__abc_41358_n1743;
  wire alu__abc_41358_n1744;
  wire alu__abc_41358_n1745;
  wire alu__abc_41358_n1746;
  wire alu__abc_41358_n1747;
  wire alu__abc_41358_n1748;
  wire alu__abc_41358_n1749;
  wire alu__abc_41358_n175;
  wire alu__abc_41358_n1750;
  wire alu__abc_41358_n1751;
  wire alu__abc_41358_n1752;
  wire alu__abc_41358_n1753;
  wire alu__abc_41358_n1754;
  wire alu__abc_41358_n1755;
  wire alu__abc_41358_n1756;
  wire alu__abc_41358_n1757;
  wire alu__abc_41358_n1758;
  wire alu__abc_41358_n1759;
  wire alu__abc_41358_n176;
  wire alu__abc_41358_n1760;
  wire alu__abc_41358_n1761;
  wire alu__abc_41358_n1762;
  wire alu__abc_41358_n1763;
  wire alu__abc_41358_n1764;
  wire alu__abc_41358_n1765;
  wire alu__abc_41358_n1766;
  wire alu__abc_41358_n1767;
  wire alu__abc_41358_n1768;
  wire alu__abc_41358_n1769;
  wire alu__abc_41358_n1770;
  wire alu__abc_41358_n1772;
  wire alu__abc_41358_n1773;
  wire alu__abc_41358_n1774;
  wire alu__abc_41358_n1775;
  wire alu__abc_41358_n1776;
  wire alu__abc_41358_n1777;
  wire alu__abc_41358_n1778;
  wire alu__abc_41358_n1779;
  wire alu__abc_41358_n177_1;
  wire alu__abc_41358_n1780;
  wire alu__abc_41358_n1781;
  wire alu__abc_41358_n1782;
  wire alu__abc_41358_n1783;
  wire alu__abc_41358_n1784;
  wire alu__abc_41358_n1785;
  wire alu__abc_41358_n1786;
  wire alu__abc_41358_n1787;
  wire alu__abc_41358_n1788;
  wire alu__abc_41358_n1789;
  wire alu__abc_41358_n178_1;
  wire alu__abc_41358_n179;
  wire alu__abc_41358_n1790;
  wire alu__abc_41358_n1791;
  wire alu__abc_41358_n1792;
  wire alu__abc_41358_n1793;
  wire alu__abc_41358_n1794;
  wire alu__abc_41358_n1795;
  wire alu__abc_41358_n1796;
  wire alu__abc_41358_n1797;
  wire alu__abc_41358_n1798;
  wire alu__abc_41358_n1799;
  wire alu__abc_41358_n180;
  wire alu__abc_41358_n1800;
  wire alu__abc_41358_n1801;
  wire alu__abc_41358_n1802;
  wire alu__abc_41358_n1803;
  wire alu__abc_41358_n1804;
  wire alu__abc_41358_n1805;
  wire alu__abc_41358_n1806;
  wire alu__abc_41358_n1807;
  wire alu__abc_41358_n1808;
  wire alu__abc_41358_n1809;
  wire alu__abc_41358_n181;
  wire alu__abc_41358_n1810;
  wire alu__abc_41358_n1811;
  wire alu__abc_41358_n1812;
  wire alu__abc_41358_n1813;
  wire alu__abc_41358_n1814;
  wire alu__abc_41358_n1815;
  wire alu__abc_41358_n1817;
  wire alu__abc_41358_n1818;
  wire alu__abc_41358_n1819;
  wire alu__abc_41358_n1820;
  wire alu__abc_41358_n1821;
  wire alu__abc_41358_n1822;
  wire alu__abc_41358_n1823;
  wire alu__abc_41358_n1824;
  wire alu__abc_41358_n1825;
  wire alu__abc_41358_n1826;
  wire alu__abc_41358_n1827;
  wire alu__abc_41358_n1828;
  wire alu__abc_41358_n1829;
  wire alu__abc_41358_n182_1;
  wire alu__abc_41358_n1830;
  wire alu__abc_41358_n1831;
  wire alu__abc_41358_n1832;
  wire alu__abc_41358_n1833;
  wire alu__abc_41358_n1834;
  wire alu__abc_41358_n1835;
  wire alu__abc_41358_n1836;
  wire alu__abc_41358_n1837;
  wire alu__abc_41358_n1838;
  wire alu__abc_41358_n1839;
  wire alu__abc_41358_n183_1;
  wire alu__abc_41358_n184;
  wire alu__abc_41358_n1840;
  wire alu__abc_41358_n1841;
  wire alu__abc_41358_n1842;
  wire alu__abc_41358_n1843;
  wire alu__abc_41358_n1844;
  wire alu__abc_41358_n1845;
  wire alu__abc_41358_n1846;
  wire alu__abc_41358_n1847;
  wire alu__abc_41358_n1848;
  wire alu__abc_41358_n1849;
  wire alu__abc_41358_n185;
  wire alu__abc_41358_n1850;
  wire alu__abc_41358_n1851;
  wire alu__abc_41358_n1852;
  wire alu__abc_41358_n1853;
  wire alu__abc_41358_n1854;
  wire alu__abc_41358_n1855;
  wire alu__abc_41358_n1856;
  wire alu__abc_41358_n1857;
  wire alu__abc_41358_n1859;
  wire alu__abc_41358_n186;
  wire alu__abc_41358_n1860;
  wire alu__abc_41358_n1861;
  wire alu__abc_41358_n1862;
  wire alu__abc_41358_n1863;
  wire alu__abc_41358_n1864;
  wire alu__abc_41358_n1865;
  wire alu__abc_41358_n1866;
  wire alu__abc_41358_n1867;
  wire alu__abc_41358_n1868;
  wire alu__abc_41358_n1869;
  wire alu__abc_41358_n187;
  wire alu__abc_41358_n1870;
  wire alu__abc_41358_n1871;
  wire alu__abc_41358_n1872;
  wire alu__abc_41358_n1873;
  wire alu__abc_41358_n1874;
  wire alu__abc_41358_n1875;
  wire alu__abc_41358_n1876;
  wire alu__abc_41358_n1877;
  wire alu__abc_41358_n1878;
  wire alu__abc_41358_n1879;
  wire alu__abc_41358_n188;
  wire alu__abc_41358_n1880;
  wire alu__abc_41358_n1881;
  wire alu__abc_41358_n1882;
  wire alu__abc_41358_n1883;
  wire alu__abc_41358_n1884;
  wire alu__abc_41358_n1885;
  wire alu__abc_41358_n1886;
  wire alu__abc_41358_n1887;
  wire alu__abc_41358_n1888;
  wire alu__abc_41358_n1889;
  wire alu__abc_41358_n189;
  wire alu__abc_41358_n1890;
  wire alu__abc_41358_n1891;
  wire alu__abc_41358_n1892;
  wire alu__abc_41358_n1893;
  wire alu__abc_41358_n1894;
  wire alu__abc_41358_n1895;
  wire alu__abc_41358_n1896;
  wire alu__abc_41358_n1897;
  wire alu__abc_41358_n1898;
  wire alu__abc_41358_n1899;
  wire alu__abc_41358_n190;
  wire alu__abc_41358_n1901;
  wire alu__abc_41358_n1902;
  wire alu__abc_41358_n1903;
  wire alu__abc_41358_n1904;
  wire alu__abc_41358_n1905;
  wire alu__abc_41358_n1906;
  wire alu__abc_41358_n1907;
  wire alu__abc_41358_n1908;
  wire alu__abc_41358_n1909;
  wire alu__abc_41358_n1910;
  wire alu__abc_41358_n1911;
  wire alu__abc_41358_n1912;
  wire alu__abc_41358_n1913;
  wire alu__abc_41358_n1914;
  wire alu__abc_41358_n1915;
  wire alu__abc_41358_n1916;
  wire alu__abc_41358_n1917;
  wire alu__abc_41358_n1918;
  wire alu__abc_41358_n1919;
  wire alu__abc_41358_n191_1;
  wire alu__abc_41358_n1920;
  wire alu__abc_41358_n1921;
  wire alu__abc_41358_n1922;
  wire alu__abc_41358_n1923;
  wire alu__abc_41358_n1924;
  wire alu__abc_41358_n1925;
  wire alu__abc_41358_n1926;
  wire alu__abc_41358_n1927;
  wire alu__abc_41358_n1928;
  wire alu__abc_41358_n1929;
  wire alu__abc_41358_n192_1;
  wire alu__abc_41358_n193;
  wire alu__abc_41358_n1930;
  wire alu__abc_41358_n1931;
  wire alu__abc_41358_n1932;
  wire alu__abc_41358_n1933;
  wire alu__abc_41358_n1934;
  wire alu__abc_41358_n1935;
  wire alu__abc_41358_n1936;
  wire alu__abc_41358_n1937;
  wire alu__abc_41358_n1938;
  wire alu__abc_41358_n1939;
  wire alu__abc_41358_n1940;
  wire alu__abc_41358_n1941;
  wire alu__abc_41358_n1942;
  wire alu__abc_41358_n1943;
  wire alu__abc_41358_n1945;
  wire alu__abc_41358_n1946;
  wire alu__abc_41358_n1947;
  wire alu__abc_41358_n1948;
  wire alu__abc_41358_n1949;
  wire alu__abc_41358_n194_1;
  wire alu__abc_41358_n195;
  wire alu__abc_41358_n1950;
  wire alu__abc_41358_n1951;
  wire alu__abc_41358_n1952;
  wire alu__abc_41358_n1953;
  wire alu__abc_41358_n1954;
  wire alu__abc_41358_n1955;
  wire alu__abc_41358_n1956;
  wire alu__abc_41358_n1957;
  wire alu__abc_41358_n1958;
  wire alu__abc_41358_n1959;
  wire alu__abc_41358_n1960;
  wire alu__abc_41358_n1961;
  wire alu__abc_41358_n1962;
  wire alu__abc_41358_n1963;
  wire alu__abc_41358_n1964;
  wire alu__abc_41358_n1965;
  wire alu__abc_41358_n1966;
  wire alu__abc_41358_n1967;
  wire alu__abc_41358_n1968;
  wire alu__abc_41358_n1969;
  wire alu__abc_41358_n196_1;
  wire alu__abc_41358_n197;
  wire alu__abc_41358_n1970;
  wire alu__abc_41358_n1971;
  wire alu__abc_41358_n1972;
  wire alu__abc_41358_n1973;
  wire alu__abc_41358_n1974;
  wire alu__abc_41358_n1975;
  wire alu__abc_41358_n1976;
  wire alu__abc_41358_n1977;
  wire alu__abc_41358_n1978;
  wire alu__abc_41358_n1979;
  wire alu__abc_41358_n1980;
  wire alu__abc_41358_n1981;
  wire alu__abc_41358_n1982;
  wire alu__abc_41358_n1983;
  wire alu__abc_41358_n1984;
  wire alu__abc_41358_n1985;
  wire alu__abc_41358_n1987;
  wire alu__abc_41358_n1988;
  wire alu__abc_41358_n1989;
  wire alu__abc_41358_n198_1;
  wire alu__abc_41358_n199;
  wire alu__abc_41358_n1990;
  wire alu__abc_41358_n1991;
  wire alu__abc_41358_n1992;
  wire alu__abc_41358_n1993;
  wire alu__abc_41358_n1994;
  wire alu__abc_41358_n1995;
  wire alu__abc_41358_n1996;
  wire alu__abc_41358_n1997;
  wire alu__abc_41358_n1998;
  wire alu__abc_41358_n1999;
  wire alu__abc_41358_n200;
  wire alu__abc_41358_n2000;
  wire alu__abc_41358_n2001;
  wire alu__abc_41358_n2002;
  wire alu__abc_41358_n2003;
  wire alu__abc_41358_n2004;
  wire alu__abc_41358_n2005;
  wire alu__abc_41358_n2006;
  wire alu__abc_41358_n2007;
  wire alu__abc_41358_n2008;
  wire alu__abc_41358_n2009;
  wire alu__abc_41358_n201;
  wire alu__abc_41358_n2010;
  wire alu__abc_41358_n2011;
  wire alu__abc_41358_n2012;
  wire alu__abc_41358_n2013;
  wire alu__abc_41358_n2014;
  wire alu__abc_41358_n2015;
  wire alu__abc_41358_n2016;
  wire alu__abc_41358_n2017;
  wire alu__abc_41358_n2018;
  wire alu__abc_41358_n2019;
  wire alu__abc_41358_n202;
  wire alu__abc_41358_n2020;
  wire alu__abc_41358_n2021;
  wire alu__abc_41358_n2022;
  wire alu__abc_41358_n2023;
  wire alu__abc_41358_n2024;
  wire alu__abc_41358_n2025;
  wire alu__abc_41358_n2026;
  wire alu__abc_41358_n2028;
  wire alu__abc_41358_n2029;
  wire alu__abc_41358_n2030;
  wire alu__abc_41358_n2031;
  wire alu__abc_41358_n2032;
  wire alu__abc_41358_n2033;
  wire alu__abc_41358_n2034;
  wire alu__abc_41358_n2035;
  wire alu__abc_41358_n2036;
  wire alu__abc_41358_n2037;
  wire alu__abc_41358_n2038;
  wire alu__abc_41358_n2039;
  wire alu__abc_41358_n203_1;
  wire alu__abc_41358_n204;
  wire alu__abc_41358_n2040;
  wire alu__abc_41358_n2041;
  wire alu__abc_41358_n2042;
  wire alu__abc_41358_n2043;
  wire alu__abc_41358_n2044;
  wire alu__abc_41358_n2045;
  wire alu__abc_41358_n2046;
  wire alu__abc_41358_n2047;
  wire alu__abc_41358_n2048;
  wire alu__abc_41358_n2049;
  wire alu__abc_41358_n205;
  wire alu__abc_41358_n2050;
  wire alu__abc_41358_n2051;
  wire alu__abc_41358_n2052;
  wire alu__abc_41358_n2053;
  wire alu__abc_41358_n2054;
  wire alu__abc_41358_n2055;
  wire alu__abc_41358_n2056;
  wire alu__abc_41358_n2057;
  wire alu__abc_41358_n2058;
  wire alu__abc_41358_n2059;
  wire alu__abc_41358_n2060;
  wire alu__abc_41358_n2061;
  wire alu__abc_41358_n2062;
  wire alu__abc_41358_n2063;
  wire alu__abc_41358_n2064;
  wire alu__abc_41358_n2065;
  wire alu__abc_41358_n2066;
  wire alu__abc_41358_n2067;
  wire alu__abc_41358_n2068;
  wire alu__abc_41358_n206_1;
  wire alu__abc_41358_n207;
  wire alu__abc_41358_n2070;
  wire alu__abc_41358_n2071;
  wire alu__abc_41358_n2072;
  wire alu__abc_41358_n2073;
  wire alu__abc_41358_n2074;
  wire alu__abc_41358_n2075;
  wire alu__abc_41358_n2076;
  wire alu__abc_41358_n2077;
  wire alu__abc_41358_n2078;
  wire alu__abc_41358_n2079;
  wire alu__abc_41358_n208;
  wire alu__abc_41358_n2080;
  wire alu__abc_41358_n2081;
  wire alu__abc_41358_n2082;
  wire alu__abc_41358_n2083;
  wire alu__abc_41358_n2084;
  wire alu__abc_41358_n2085;
  wire alu__abc_41358_n2086;
  wire alu__abc_41358_n2087;
  wire alu__abc_41358_n2088;
  wire alu__abc_41358_n2089;
  wire alu__abc_41358_n209;
  wire alu__abc_41358_n2090;
  wire alu__abc_41358_n2091;
  wire alu__abc_41358_n2092;
  wire alu__abc_41358_n2093;
  wire alu__abc_41358_n2094;
  wire alu__abc_41358_n2095;
  wire alu__abc_41358_n2096;
  wire alu__abc_41358_n2097;
  wire alu__abc_41358_n2098;
  wire alu__abc_41358_n2099;
  wire alu__abc_41358_n210;
  wire alu__abc_41358_n2100;
  wire alu__abc_41358_n2101;
  wire alu__abc_41358_n2102;
  wire alu__abc_41358_n2103;
  wire alu__abc_41358_n2104;
  wire alu__abc_41358_n2105;
  wire alu__abc_41358_n2106;
  wire alu__abc_41358_n2107;
  wire alu__abc_41358_n2108;
  wire alu__abc_41358_n2109;
  wire alu__abc_41358_n211;
  wire alu__abc_41358_n2110;
  wire alu__abc_41358_n2111;
  wire alu__abc_41358_n2113;
  wire alu__abc_41358_n2114;
  wire alu__abc_41358_n2115;
  wire alu__abc_41358_n2116;
  wire alu__abc_41358_n2117;
  wire alu__abc_41358_n2118;
  wire alu__abc_41358_n2119;
  wire alu__abc_41358_n212;
  wire alu__abc_41358_n2120;
  wire alu__abc_41358_n2121;
  wire alu__abc_41358_n2122;
  wire alu__abc_41358_n2123;
  wire alu__abc_41358_n2124;
  wire alu__abc_41358_n2125;
  wire alu__abc_41358_n2126;
  wire alu__abc_41358_n2127;
  wire alu__abc_41358_n2128;
  wire alu__abc_41358_n2129;
  wire alu__abc_41358_n213;
  wire alu__abc_41358_n2130;
  wire alu__abc_41358_n2131;
  wire alu__abc_41358_n2132;
  wire alu__abc_41358_n2133;
  wire alu__abc_41358_n2134;
  wire alu__abc_41358_n2135;
  wire alu__abc_41358_n2136;
  wire alu__abc_41358_n2137;
  wire alu__abc_41358_n2138;
  wire alu__abc_41358_n2139;
  wire alu__abc_41358_n214;
  wire alu__abc_41358_n2140;
  wire alu__abc_41358_n2141;
  wire alu__abc_41358_n2142;
  wire alu__abc_41358_n2143;
  wire alu__abc_41358_n2144;
  wire alu__abc_41358_n2145;
  wire alu__abc_41358_n2146;
  wire alu__abc_41358_n2147;
  wire alu__abc_41358_n2148;
  wire alu__abc_41358_n2149;
  wire alu__abc_41358_n215;
  wire alu__abc_41358_n2150;
  wire alu__abc_41358_n2151;
  wire alu__abc_41358_n2152;
  wire alu__abc_41358_n2153;
  wire alu__abc_41358_n2155;
  wire alu__abc_41358_n2156;
  wire alu__abc_41358_n2157;
  wire alu__abc_41358_n2158;
  wire alu__abc_41358_n2159;
  wire alu__abc_41358_n216;
  wire alu__abc_41358_n2160;
  wire alu__abc_41358_n2161;
  wire alu__abc_41358_n2162;
  wire alu__abc_41358_n2163;
  wire alu__abc_41358_n2164;
  wire alu__abc_41358_n2165;
  wire alu__abc_41358_n2166;
  wire alu__abc_41358_n2167;
  wire alu__abc_41358_n2168;
  wire alu__abc_41358_n2169;
  wire alu__abc_41358_n217;
  wire alu__abc_41358_n2170;
  wire alu__abc_41358_n2171;
  wire alu__abc_41358_n2172;
  wire alu__abc_41358_n2173;
  wire alu__abc_41358_n2174;
  wire alu__abc_41358_n2175;
  wire alu__abc_41358_n2176;
  wire alu__abc_41358_n2177;
  wire alu__abc_41358_n2178;
  wire alu__abc_41358_n2179;
  wire alu__abc_41358_n218;
  wire alu__abc_41358_n2180;
  wire alu__abc_41358_n2181;
  wire alu__abc_41358_n2182;
  wire alu__abc_41358_n2183;
  wire alu__abc_41358_n2184;
  wire alu__abc_41358_n2185;
  wire alu__abc_41358_n2186;
  wire alu__abc_41358_n2187;
  wire alu__abc_41358_n2188;
  wire alu__abc_41358_n2189;
  wire alu__abc_41358_n219;
  wire alu__abc_41358_n2190;
  wire alu__abc_41358_n2191;
  wire alu__abc_41358_n2192;
  wire alu__abc_41358_n2194;
  wire alu__abc_41358_n2195;
  wire alu__abc_41358_n2196;
  wire alu__abc_41358_n2197;
  wire alu__abc_41358_n2198;
  wire alu__abc_41358_n2199;
  wire alu__abc_41358_n220;
  wire alu__abc_41358_n2200;
  wire alu__abc_41358_n2201;
  wire alu__abc_41358_n2202;
  wire alu__abc_41358_n2203;
  wire alu__abc_41358_n2204;
  wire alu__abc_41358_n2205;
  wire alu__abc_41358_n2206;
  wire alu__abc_41358_n2207;
  wire alu__abc_41358_n2208;
  wire alu__abc_41358_n2209;
  wire alu__abc_41358_n221;
  wire alu__abc_41358_n2210;
  wire alu__abc_41358_n2211;
  wire alu__abc_41358_n2212;
  wire alu__abc_41358_n2213;
  wire alu__abc_41358_n2214;
  wire alu__abc_41358_n2215;
  wire alu__abc_41358_n2216;
  wire alu__abc_41358_n2217;
  wire alu__abc_41358_n2218;
  wire alu__abc_41358_n2219;
  wire alu__abc_41358_n222;
  wire alu__abc_41358_n2220;
  wire alu__abc_41358_n2221;
  wire alu__abc_41358_n2222;
  wire alu__abc_41358_n2223;
  wire alu__abc_41358_n2224;
  wire alu__abc_41358_n2225;
  wire alu__abc_41358_n2226;
  wire alu__abc_41358_n2227;
  wire alu__abc_41358_n2228;
  wire alu__abc_41358_n2229;
  wire alu__abc_41358_n223;
  wire alu__abc_41358_n2230;
  wire alu__abc_41358_n2231;
  wire alu__abc_41358_n2232;
  wire alu__abc_41358_n2233;
  wire alu__abc_41358_n2235;
  wire alu__abc_41358_n2236;
  wire alu__abc_41358_n2237;
  wire alu__abc_41358_n2238;
  wire alu__abc_41358_n2239;
  wire alu__abc_41358_n224;
  wire alu__abc_41358_n2240;
  wire alu__abc_41358_n2241;
  wire alu__abc_41358_n2242;
  wire alu__abc_41358_n2243;
  wire alu__abc_41358_n2244;
  wire alu__abc_41358_n2245;
  wire alu__abc_41358_n2246;
  wire alu__abc_41358_n2247;
  wire alu__abc_41358_n2248;
  wire alu__abc_41358_n2249;
  wire alu__abc_41358_n225;
  wire alu__abc_41358_n2250;
  wire alu__abc_41358_n2251;
  wire alu__abc_41358_n2252;
  wire alu__abc_41358_n2253;
  wire alu__abc_41358_n2254;
  wire alu__abc_41358_n2255;
  wire alu__abc_41358_n2256;
  wire alu__abc_41358_n2257;
  wire alu__abc_41358_n2258;
  wire alu__abc_41358_n2259;
  wire alu__abc_41358_n226;
  wire alu__abc_41358_n2260;
  wire alu__abc_41358_n2261;
  wire alu__abc_41358_n2262;
  wire alu__abc_41358_n2263;
  wire alu__abc_41358_n2264;
  wire alu__abc_41358_n2265;
  wire alu__abc_41358_n2266;
  wire alu__abc_41358_n2267;
  wire alu__abc_41358_n2268;
  wire alu__abc_41358_n2269;
  wire alu__abc_41358_n227;
  wire alu__abc_41358_n2270;
  wire alu__abc_41358_n2271;
  wire alu__abc_41358_n2272;
  wire alu__abc_41358_n2273;
  wire alu__abc_41358_n2274;
  wire alu__abc_41358_n2275;
  wire alu__abc_41358_n2276;
  wire alu__abc_41358_n2278;
  wire alu__abc_41358_n2279;
  wire alu__abc_41358_n228;
  wire alu__abc_41358_n2280;
  wire alu__abc_41358_n2281;
  wire alu__abc_41358_n2282;
  wire alu__abc_41358_n2283;
  wire alu__abc_41358_n2284;
  wire alu__abc_41358_n2285;
  wire alu__abc_41358_n2286;
  wire alu__abc_41358_n2287;
  wire alu__abc_41358_n2288;
  wire alu__abc_41358_n2289;
  wire alu__abc_41358_n229;
  wire alu__abc_41358_n2290;
  wire alu__abc_41358_n2291;
  wire alu__abc_41358_n2292;
  wire alu__abc_41358_n2293;
  wire alu__abc_41358_n2294;
  wire alu__abc_41358_n2295;
  wire alu__abc_41358_n2296;
  wire alu__abc_41358_n2297;
  wire alu__abc_41358_n2298;
  wire alu__abc_41358_n2299;
  wire alu__abc_41358_n230;
  wire alu__abc_41358_n2300;
  wire alu__abc_41358_n2301;
  wire alu__abc_41358_n2302;
  wire alu__abc_41358_n2303;
  wire alu__abc_41358_n2304;
  wire alu__abc_41358_n2305;
  wire alu__abc_41358_n2306;
  wire alu__abc_41358_n2307;
  wire alu__abc_41358_n2308;
  wire alu__abc_41358_n2309;
  wire alu__abc_41358_n231;
  wire alu__abc_41358_n2310;
  wire alu__abc_41358_n2311;
  wire alu__abc_41358_n2312;
  wire alu__abc_41358_n2313;
  wire alu__abc_41358_n2314;
  wire alu__abc_41358_n2315;
  wire alu__abc_41358_n2316;
  wire alu__abc_41358_n2317;
  wire alu__abc_41358_n2319;
  wire alu__abc_41358_n232;
  wire alu__abc_41358_n2320;
  wire alu__abc_41358_n2321;
  wire alu__abc_41358_n2322;
  wire alu__abc_41358_n2323;
  wire alu__abc_41358_n2324;
  wire alu__abc_41358_n2325;
  wire alu__abc_41358_n2326;
  wire alu__abc_41358_n2327;
  wire alu__abc_41358_n2328;
  wire alu__abc_41358_n2329;
  wire alu__abc_41358_n233;
  wire alu__abc_41358_n2330;
  wire alu__abc_41358_n2331;
  wire alu__abc_41358_n2332;
  wire alu__abc_41358_n2333;
  wire alu__abc_41358_n2334;
  wire alu__abc_41358_n2335;
  wire alu__abc_41358_n2336;
  wire alu__abc_41358_n2337;
  wire alu__abc_41358_n2338;
  wire alu__abc_41358_n2339;
  wire alu__abc_41358_n234;
  wire alu__abc_41358_n2340;
  wire alu__abc_41358_n2341;
  wire alu__abc_41358_n2342;
  wire alu__abc_41358_n2343;
  wire alu__abc_41358_n2344;
  wire alu__abc_41358_n2345;
  wire alu__abc_41358_n2346;
  wire alu__abc_41358_n2347;
  wire alu__abc_41358_n2348;
  wire alu__abc_41358_n2349;
  wire alu__abc_41358_n235;
  wire alu__abc_41358_n2350;
  wire alu__abc_41358_n2351;
  wire alu__abc_41358_n2352;
  wire alu__abc_41358_n2353;
  wire alu__abc_41358_n2354;
  wire alu__abc_41358_n2355;
  wire alu__abc_41358_n2356;
  wire alu__abc_41358_n2358;
  wire alu__abc_41358_n2359;
  wire alu__abc_41358_n236;
  wire alu__abc_41358_n2360;
  wire alu__abc_41358_n2361;
  wire alu__abc_41358_n2362;
  wire alu__abc_41358_n2363;
  wire alu__abc_41358_n2364;
  wire alu__abc_41358_n2365;
  wire alu__abc_41358_n2366;
  wire alu__abc_41358_n2367;
  wire alu__abc_41358_n2368;
  wire alu__abc_41358_n2369;
  wire alu__abc_41358_n237;
  wire alu__abc_41358_n2370;
  wire alu__abc_41358_n2371;
  wire alu__abc_41358_n2372;
  wire alu__abc_41358_n2373;
  wire alu__abc_41358_n2374;
  wire alu__abc_41358_n2375;
  wire alu__abc_41358_n2376;
  wire alu__abc_41358_n2377;
  wire alu__abc_41358_n2378;
  wire alu__abc_41358_n2379;
  wire alu__abc_41358_n238;
  wire alu__abc_41358_n2380;
  wire alu__abc_41358_n2381;
  wire alu__abc_41358_n2382;
  wire alu__abc_41358_n2383;
  wire alu__abc_41358_n2384;
  wire alu__abc_41358_n2385;
  wire alu__abc_41358_n2386;
  wire alu__abc_41358_n2387;
  wire alu__abc_41358_n2388;
  wire alu__abc_41358_n2389;
  wire alu__abc_41358_n239;
  wire alu__abc_41358_n2390;
  wire alu__abc_41358_n2391;
  wire alu__abc_41358_n2392;
  wire alu__abc_41358_n2393;
  wire alu__abc_41358_n2394;
  wire alu__abc_41358_n2395;
  wire alu__abc_41358_n2396;
  wire alu__abc_41358_n2397;
  wire alu__abc_41358_n2398;
  wire alu__abc_41358_n2399;
  wire alu__abc_41358_n240;
  wire alu__abc_41358_n2401;
  wire alu__abc_41358_n2402;
  wire alu__abc_41358_n2403;
  wire alu__abc_41358_n2404;
  wire alu__abc_41358_n2405;
  wire alu__abc_41358_n2406;
  wire alu__abc_41358_n2407;
  wire alu__abc_41358_n2408;
  wire alu__abc_41358_n2409;
  wire alu__abc_41358_n241;
  wire alu__abc_41358_n2410;
  wire alu__abc_41358_n2411;
  wire alu__abc_41358_n2412;
  wire alu__abc_41358_n2413;
  wire alu__abc_41358_n2414;
  wire alu__abc_41358_n2415;
  wire alu__abc_41358_n2416;
  wire alu__abc_41358_n2417;
  wire alu__abc_41358_n2418;
  wire alu__abc_41358_n2419;
  wire alu__abc_41358_n242;
  wire alu__abc_41358_n2420;
  wire alu__abc_41358_n2421;
  wire alu__abc_41358_n2422;
  wire alu__abc_41358_n2423;
  wire alu__abc_41358_n2424;
  wire alu__abc_41358_n2425;
  wire alu__abc_41358_n2426;
  wire alu__abc_41358_n2427;
  wire alu__abc_41358_n2428;
  wire alu__abc_41358_n2429;
  wire alu__abc_41358_n243;
  wire alu__abc_41358_n2430;
  wire alu__abc_41358_n2431;
  wire alu__abc_41358_n2432;
  wire alu__abc_41358_n2433;
  wire alu__abc_41358_n2434;
  wire alu__abc_41358_n2435;
  wire alu__abc_41358_n2436;
  wire alu__abc_41358_n2437;
  wire alu__abc_41358_n2439;
  wire alu__abc_41358_n244;
  wire alu__abc_41358_n2440;
  wire alu__abc_41358_n2441;
  wire alu__abc_41358_n2442;
  wire alu__abc_41358_n2443;
  wire alu__abc_41358_n2444;
  wire alu__abc_41358_n2445;
  wire alu__abc_41358_n2446;
  wire alu__abc_41358_n2447;
  wire alu__abc_41358_n2448;
  wire alu__abc_41358_n2449;
  wire alu__abc_41358_n245;
  wire alu__abc_41358_n2450;
  wire alu__abc_41358_n2451;
  wire alu__abc_41358_n2452;
  wire alu__abc_41358_n2453;
  wire alu__abc_41358_n2454;
  wire alu__abc_41358_n2455;
  wire alu__abc_41358_n2456;
  wire alu__abc_41358_n2457;
  wire alu__abc_41358_n2458;
  wire alu__abc_41358_n2459;
  wire alu__abc_41358_n246;
  wire alu__abc_41358_n2460;
  wire alu__abc_41358_n2461;
  wire alu__abc_41358_n2462;
  wire alu__abc_41358_n2463;
  wire alu__abc_41358_n2464;
  wire alu__abc_41358_n2465;
  wire alu__abc_41358_n2466;
  wire alu__abc_41358_n2467;
  wire alu__abc_41358_n2468;
  wire alu__abc_41358_n2469;
  wire alu__abc_41358_n247;
  wire alu__abc_41358_n2470;
  wire alu__abc_41358_n2471;
  wire alu__abc_41358_n2472;
  wire alu__abc_41358_n2473;
  wire alu__abc_41358_n2474;
  wire alu__abc_41358_n2475;
  wire alu__abc_41358_n2477;
  wire alu__abc_41358_n2478;
  wire alu__abc_41358_n2479;
  wire alu__abc_41358_n248;
  wire alu__abc_41358_n2480;
  wire alu__abc_41358_n2481;
  wire alu__abc_41358_n2482;
  wire alu__abc_41358_n2483;
  wire alu__abc_41358_n2484;
  wire alu__abc_41358_n2485;
  wire alu__abc_41358_n2486;
  wire alu__abc_41358_n2487;
  wire alu__abc_41358_n2488;
  wire alu__abc_41358_n2489;
  wire alu__abc_41358_n249;
  wire alu__abc_41358_n2490;
  wire alu__abc_41358_n2491;
  wire alu__abc_41358_n2492;
  wire alu__abc_41358_n2493;
  wire alu__abc_41358_n2494;
  wire alu__abc_41358_n2495;
  wire alu__abc_41358_n2496;
  wire alu__abc_41358_n2497;
  wire alu__abc_41358_n2498;
  wire alu__abc_41358_n2499;
  wire alu__abc_41358_n250;
  wire alu__abc_41358_n2500;
  wire alu__abc_41358_n2501;
  wire alu__abc_41358_n2502;
  wire alu__abc_41358_n2503;
  wire alu__abc_41358_n2504;
  wire alu__abc_41358_n2505;
  wire alu__abc_41358_n2506;
  wire alu__abc_41358_n2507;
  wire alu__abc_41358_n2508;
  wire alu__abc_41358_n2509;
  wire alu__abc_41358_n251;
  wire alu__abc_41358_n2510;
  wire alu__abc_41358_n2511;
  wire alu__abc_41358_n2512;
  wire alu__abc_41358_n2513;
  wire alu__abc_41358_n2514;
  wire alu__abc_41358_n2515;
  wire alu__abc_41358_n2516;
  wire alu__abc_41358_n2517;
  wire alu__abc_41358_n2518;
  wire alu__abc_41358_n2519;
  wire alu__abc_41358_n252;
  wire alu__abc_41358_n2520;
  wire alu__abc_41358_n2521;
  wire alu__abc_41358_n2522;
  wire alu__abc_41358_n2523;
  wire alu__abc_41358_n2524;
  wire alu__abc_41358_n2525;
  wire alu__abc_41358_n2526;
  wire alu__abc_41358_n2527;
  wire alu__abc_41358_n2528;
  wire alu__abc_41358_n2529;
  wire alu__abc_41358_n252_bF_buf0;
  wire alu__abc_41358_n252_bF_buf1;
  wire alu__abc_41358_n252_bF_buf2;
  wire alu__abc_41358_n252_bF_buf3;
  wire alu__abc_41358_n252_bF_buf4;
  wire alu__abc_41358_n252_bF_buf5;
  wire alu__abc_41358_n252_bF_buf6;
  wire alu__abc_41358_n253;
  wire alu__abc_41358_n2530;
  wire alu__abc_41358_n2531;
  wire alu__abc_41358_n2532;
  wire alu__abc_41358_n2533;
  wire alu__abc_41358_n2534;
  wire alu__abc_41358_n2535;
  wire alu__abc_41358_n2536;
  wire alu__abc_41358_n2537;
  wire alu__abc_41358_n2538;
  wire alu__abc_41358_n2539;
  wire alu__abc_41358_n254;
  wire alu__abc_41358_n2540;
  wire alu__abc_41358_n2541;
  wire alu__abc_41358_n2542;
  wire alu__abc_41358_n2543;
  wire alu__abc_41358_n2544;
  wire alu__abc_41358_n2545;
  wire alu__abc_41358_n2546;
  wire alu__abc_41358_n2547;
  wire alu__abc_41358_n2548;
  wire alu__abc_41358_n2549;
  wire alu__abc_41358_n255;
  wire alu__abc_41358_n2550;
  wire alu__abc_41358_n2551;
  wire alu__abc_41358_n2552;
  wire alu__abc_41358_n2553;
  wire alu__abc_41358_n2554;
  wire alu__abc_41358_n2555;
  wire alu__abc_41358_n2556;
  wire alu__abc_41358_n2557;
  wire alu__abc_41358_n2558;
  wire alu__abc_41358_n2559;
  wire alu__abc_41358_n256;
  wire alu__abc_41358_n2560;
  wire alu__abc_41358_n2562;
  wire alu__abc_41358_n2563;
  wire alu__abc_41358_n257;
  wire alu__abc_41358_n258;
  wire alu__abc_41358_n259;
  wire alu__abc_41358_n259_bF_buf0;
  wire alu__abc_41358_n259_bF_buf1;
  wire alu__abc_41358_n259_bF_buf2;
  wire alu__abc_41358_n259_bF_buf3;
  wire alu__abc_41358_n259_bF_buf4;
  wire alu__abc_41358_n260;
  wire alu__abc_41358_n261;
  wire alu__abc_41358_n262;
  wire alu__abc_41358_n263;
  wire alu__abc_41358_n264;
  wire alu__abc_41358_n265;
  wire alu__abc_41358_n266;
  wire alu__abc_41358_n267;
  wire alu__abc_41358_n268;
  wire alu__abc_41358_n269;
  wire alu__abc_41358_n270;
  wire alu__abc_41358_n271;
  wire alu__abc_41358_n272;
  wire alu__abc_41358_n273;
  wire alu__abc_41358_n274;
  wire alu__abc_41358_n275;
  wire alu__abc_41358_n276;
  wire alu__abc_41358_n277;
  wire alu__abc_41358_n278;
  wire alu__abc_41358_n279;
  wire alu__abc_41358_n279_bF_buf0;
  wire alu__abc_41358_n279_bF_buf1;
  wire alu__abc_41358_n279_bF_buf2;
  wire alu__abc_41358_n279_bF_buf3;
  wire alu__abc_41358_n279_bF_buf4;
  wire alu__abc_41358_n279_bF_buf5;
  wire alu__abc_41358_n280;
  wire alu__abc_41358_n281;
  wire alu__abc_41358_n282;
  wire alu__abc_41358_n283;
  wire alu__abc_41358_n284;
  wire alu__abc_41358_n285;
  wire alu__abc_41358_n286;
  wire alu__abc_41358_n287;
  wire alu__abc_41358_n288;
  wire alu__abc_41358_n289;
  wire alu__abc_41358_n290;
  wire alu__abc_41358_n291;
  wire alu__abc_41358_n292;
  wire alu__abc_41358_n293;
  wire alu__abc_41358_n294;
  wire alu__abc_41358_n294_bF_buf0;
  wire alu__abc_41358_n294_bF_buf1;
  wire alu__abc_41358_n294_bF_buf2;
  wire alu__abc_41358_n294_bF_buf3;
  wire alu__abc_41358_n294_bF_buf4;
  wire alu__abc_41358_n294_bF_buf5;
  wire alu__abc_41358_n294_bF_buf6;
  wire alu__abc_41358_n294_bF_buf7;
  wire alu__abc_41358_n295;
  wire alu__abc_41358_n296;
  wire alu__abc_41358_n297;
  wire alu__abc_41358_n298;
  wire alu__abc_41358_n299;
  wire alu__abc_41358_n299_bF_buf0;
  wire alu__abc_41358_n299_bF_buf1;
  wire alu__abc_41358_n299_bF_buf2;
  wire alu__abc_41358_n299_bF_buf3;
  wire alu__abc_41358_n299_bF_buf4;
  wire alu__abc_41358_n299_bF_buf5;
  wire alu__abc_41358_n299_bF_buf6;
  wire alu__abc_41358_n299_bF_buf7;
  wire alu__abc_41358_n300;
  wire alu__abc_41358_n301;
  wire alu__abc_41358_n302;
  wire alu__abc_41358_n303;
  wire alu__abc_41358_n304;
  wire alu__abc_41358_n305;
  wire alu__abc_41358_n306;
  wire alu__abc_41358_n307;
  wire alu__abc_41358_n308;
  wire alu__abc_41358_n309;
  wire alu__abc_41358_n310;
  wire alu__abc_41358_n311;
  wire alu__abc_41358_n312;
  wire alu__abc_41358_n313;
  wire alu__abc_41358_n314;
  wire alu__abc_41358_n315;
  wire alu__abc_41358_n316;
  wire alu__abc_41358_n317;
  wire alu__abc_41358_n318;
  wire alu__abc_41358_n319;
  wire alu__abc_41358_n320;
  wire alu__abc_41358_n321;
  wire alu__abc_41358_n322;
  wire alu__abc_41358_n323;
  wire alu__abc_41358_n324;
  wire alu__abc_41358_n325;
  wire alu__abc_41358_n326;
  wire alu__abc_41358_n327;
  wire alu__abc_41358_n328;
  wire alu__abc_41358_n329_1;
  wire alu__abc_41358_n330;
  wire alu__abc_41358_n331;
  wire alu__abc_41358_n332;
  wire alu__abc_41358_n333;
  wire alu__abc_41358_n334;
  wire alu__abc_41358_n335;
  wire alu__abc_41358_n336;
  wire alu__abc_41358_n337;
  wire alu__abc_41358_n338;
  wire alu__abc_41358_n339;
  wire alu__abc_41358_n340;
  wire alu__abc_41358_n341;
  wire alu__abc_41358_n342;
  wire alu__abc_41358_n343;
  wire alu__abc_41358_n344;
  wire alu__abc_41358_n345;
  wire alu__abc_41358_n346;
  wire alu__abc_41358_n347;
  wire alu__abc_41358_n348;
  wire alu__abc_41358_n349;
  wire alu__abc_41358_n350;
  wire alu__abc_41358_n351;
  wire alu__abc_41358_n352;
  wire alu__abc_41358_n353;
  wire alu__abc_41358_n354;
  wire alu__abc_41358_n355;
  wire alu__abc_41358_n356;
  wire alu__abc_41358_n357;
  wire alu__abc_41358_n358;
  wire alu__abc_41358_n359;
  wire alu__abc_41358_n360;
  wire alu__abc_41358_n361;
  wire alu__abc_41358_n362;
  wire alu__abc_41358_n363;
  wire alu__abc_41358_n364;
  wire alu__abc_41358_n365;
  wire alu__abc_41358_n366;
  wire alu__abc_41358_n367;
  wire alu__abc_41358_n368;
  wire alu__abc_41358_n369;
  wire alu__abc_41358_n370;
  wire alu__abc_41358_n371;
  wire alu__abc_41358_n372;
  wire alu__abc_41358_n373;
  wire alu__abc_41358_n374;
  wire alu__abc_41358_n375;
  wire alu__abc_41358_n376;
  wire alu__abc_41358_n378;
  wire alu__abc_41358_n379;
  wire alu__abc_41358_n380;
  wire alu__abc_41358_n382;
  wire alu__abc_41358_n383;
  wire alu__abc_41358_n384;
  wire alu__abc_41358_n385;
  wire alu__abc_41358_n387;
  wire alu__abc_41358_n388;
  wire alu__abc_41358_n389;
  wire alu__abc_41358_n390;
  wire alu__abc_41358_n391;
  wire alu__abc_41358_n392;
  wire alu__abc_41358_n393;
  wire alu__abc_41358_n394;
  wire alu__abc_41358_n395;
  wire alu__abc_41358_n396;
  wire alu__abc_41358_n397;
  wire alu__abc_41358_n398;
  wire alu__abc_41358_n399;
  wire alu__abc_41358_n400;
  wire alu__abc_41358_n401;
  wire alu__abc_41358_n402;
  wire alu__abc_41358_n403;
  wire alu__abc_41358_n404;
  wire alu__abc_41358_n405;
  wire alu__abc_41358_n406;
  wire alu__abc_41358_n407;
  wire alu__abc_41358_n408;
  wire alu__abc_41358_n409;
  wire alu__abc_41358_n410;
  wire alu__abc_41358_n411;
  wire alu__abc_41358_n412;
  wire alu__abc_41358_n413;
  wire alu__abc_41358_n414;
  wire alu__abc_41358_n415;
  wire alu__abc_41358_n416;
  wire alu__abc_41358_n417;
  wire alu__abc_41358_n418;
  wire alu__abc_41358_n419;
  wire alu__abc_41358_n420;
  wire alu__abc_41358_n421;
  wire alu__abc_41358_n422;
  wire alu__abc_41358_n423;
  wire alu__abc_41358_n424;
  wire alu__abc_41358_n425;
  wire alu__abc_41358_n426;
  wire alu__abc_41358_n427;
  wire alu__abc_41358_n428;
  wire alu__abc_41358_n429;
  wire alu__abc_41358_n430;
  wire alu__abc_41358_n431;
  wire alu__abc_41358_n432;
  wire alu__abc_41358_n433;
  wire alu__abc_41358_n434;
  wire alu__abc_41358_n435;
  wire alu__abc_41358_n436;
  wire alu__abc_41358_n437;
  wire alu__abc_41358_n438;
  wire alu__abc_41358_n439;
  wire alu__abc_41358_n440;
  wire alu__abc_41358_n441;
  wire alu__abc_41358_n442;
  wire alu__abc_41358_n443;
  wire alu__abc_41358_n444;
  wire alu__abc_41358_n445;
  wire alu__abc_41358_n446;
  wire alu__abc_41358_n447;
  wire alu__abc_41358_n448;
  wire alu__abc_41358_n449;
  wire alu__abc_41358_n450;
  wire alu__abc_41358_n451;
  wire alu__abc_41358_n452;
  wire alu__abc_41358_n453;
  wire alu__abc_41358_n454;
  wire alu__abc_41358_n455;
  wire alu__abc_41358_n456;
  wire alu__abc_41358_n457;
  wire alu__abc_41358_n458;
  wire alu__abc_41358_n459;
  wire alu__abc_41358_n460;
  wire alu__abc_41358_n461;
  wire alu__abc_41358_n462;
  wire alu__abc_41358_n463;
  wire alu__abc_41358_n464;
  wire alu__abc_41358_n465;
  wire alu__abc_41358_n466;
  wire alu__abc_41358_n467;
  wire alu__abc_41358_n468;
  wire alu__abc_41358_n469;
  wire alu__abc_41358_n470;
  wire alu__abc_41358_n471;
  wire alu__abc_41358_n472;
  wire alu__abc_41358_n473;
  wire alu__abc_41358_n474;
  wire alu__abc_41358_n475;
  wire alu__abc_41358_n476;
  wire alu__abc_41358_n477;
  wire alu__abc_41358_n478;
  wire alu__abc_41358_n479;
  wire alu__abc_41358_n480;
  wire alu__abc_41358_n481;
  wire alu__abc_41358_n482;
  wire alu__abc_41358_n483;
  wire alu__abc_41358_n484;
  wire alu__abc_41358_n485;
  wire alu__abc_41358_n486;
  wire alu__abc_41358_n487;
  wire alu__abc_41358_n488;
  wire alu__abc_41358_n489;
  wire alu__abc_41358_n490;
  wire alu__abc_41358_n491;
  wire alu__abc_41358_n492;
  wire alu__abc_41358_n493;
  wire alu__abc_41358_n494;
  wire alu__abc_41358_n495;
  wire alu__abc_41358_n496;
  wire alu__abc_41358_n497;
  wire alu__abc_41358_n498;
  wire alu__abc_41358_n499;
  wire alu__abc_41358_n500;
  wire alu__abc_41358_n501;
  wire alu__abc_41358_n502;
  wire alu__abc_41358_n503;
  wire alu__abc_41358_n504;
  wire alu__abc_41358_n505;
  wire alu__abc_41358_n506;
  wire alu__abc_41358_n507;
  wire alu__abc_41358_n508;
  wire alu__abc_41358_n509;
  wire alu__abc_41358_n510;
  wire alu__abc_41358_n511;
  wire alu__abc_41358_n513;
  wire alu__abc_41358_n514;
  wire alu__abc_41358_n515;
  wire alu__abc_41358_n516;
  wire alu__abc_41358_n517;
  wire alu__abc_41358_n518;
  wire alu__abc_41358_n519;
  wire alu__abc_41358_n520;
  wire alu__abc_41358_n521;
  wire alu__abc_41358_n522;
  wire alu__abc_41358_n523;
  wire alu__abc_41358_n524;
  wire alu__abc_41358_n525;
  wire alu__abc_41358_n526;
  wire alu__abc_41358_n527;
  wire alu__abc_41358_n528;
  wire alu__abc_41358_n529;
  wire alu__abc_41358_n530;
  wire alu__abc_41358_n531;
  wire alu__abc_41358_n532;
  wire alu__abc_41358_n533;
  wire alu__abc_41358_n534;
  wire alu__abc_41358_n535;
  wire alu__abc_41358_n536;
  wire alu__abc_41358_n537;
  wire alu__abc_41358_n538;
  wire alu__abc_41358_n539;
  wire alu__abc_41358_n540;
  wire alu__abc_41358_n541;
  wire alu__abc_41358_n542;
  wire alu__abc_41358_n543;
  wire alu__abc_41358_n544;
  wire alu__abc_41358_n545;
  wire alu__abc_41358_n546;
  wire alu__abc_41358_n547;
  wire alu__abc_41358_n548;
  wire alu__abc_41358_n549;
  wire alu__abc_41358_n550;
  wire alu__abc_41358_n551;
  wire alu__abc_41358_n552;
  wire alu__abc_41358_n553;
  wire alu__abc_41358_n554;
  wire alu__abc_41358_n555;
  wire alu__abc_41358_n556;
  wire alu__abc_41358_n557;
  wire alu__abc_41358_n558;
  wire alu__abc_41358_n559;
  wire alu__abc_41358_n560;
  wire alu__abc_41358_n561;
  wire alu__abc_41358_n562;
  wire alu__abc_41358_n563;
  wire alu__abc_41358_n564;
  wire alu__abc_41358_n565_1;
  wire alu__abc_41358_n566;
  wire alu__abc_41358_n567;
  wire alu__abc_41358_n568;
  wire alu__abc_41358_n569;
  wire alu__abc_41358_n570;
  wire alu__abc_41358_n571;
  wire alu__abc_41358_n572;
  wire alu__abc_41358_n573;
  wire alu__abc_41358_n574;
  wire alu__abc_41358_n575;
  wire alu__abc_41358_n576;
  wire alu__abc_41358_n577;
  wire alu__abc_41358_n578;
  wire alu__abc_41358_n579;
  wire alu__abc_41358_n580;
  wire alu__abc_41358_n581;
  wire alu__abc_41358_n582;
  wire alu__abc_41358_n583;
  wire alu__abc_41358_n584;
  wire alu__abc_41358_n585;
  wire alu__abc_41358_n586;
  wire alu__abc_41358_n587;
  wire alu__abc_41358_n588;
  wire alu__abc_41358_n589;
  wire alu__abc_41358_n590;
  wire alu__abc_41358_n591;
  wire alu__abc_41358_n592;
  wire alu__abc_41358_n593;
  wire alu__abc_41358_n594;
  wire alu__abc_41358_n595;
  wire alu__abc_41358_n596;
  wire alu__abc_41358_n597;
  wire alu__abc_41358_n598;
  wire alu__abc_41358_n599;
  wire alu__abc_41358_n600;
  wire alu__abc_41358_n601;
  wire alu__abc_41358_n602;
  wire alu__abc_41358_n603;
  wire alu__abc_41358_n604;
  wire alu__abc_41358_n605;
  wire alu__abc_41358_n606;
  wire alu__abc_41358_n607;
  wire alu__abc_41358_n608;
  wire alu__abc_41358_n609;
  wire alu__abc_41358_n610;
  wire alu__abc_41358_n611;
  wire alu__abc_41358_n612;
  wire alu__abc_41358_n613;
  wire alu__abc_41358_n614;
  wire alu__abc_41358_n615;
  wire alu__abc_41358_n616;
  wire alu__abc_41358_n617;
  wire alu__abc_41358_n618;
  wire alu__abc_41358_n619;
  wire alu__abc_41358_n620_1;
  wire alu__abc_41358_n621;
  wire alu__abc_41358_n622;
  wire alu__abc_41358_n623;
  wire alu__abc_41358_n624;
  wire alu__abc_41358_n625;
  wire alu__abc_41358_n626;
  wire alu__abc_41358_n627;
  wire alu__abc_41358_n628;
  wire alu__abc_41358_n629;
  wire alu__abc_41358_n630;
  wire alu__abc_41358_n631;
  wire alu__abc_41358_n632;
  wire alu__abc_41358_n633;
  wire alu__abc_41358_n634;
  wire alu__abc_41358_n635;
  wire alu__abc_41358_n636;
  wire alu__abc_41358_n637;
  wire alu__abc_41358_n638;
  wire alu__abc_41358_n639;
  wire alu__abc_41358_n640;
  wire alu__abc_41358_n641;
  wire alu__abc_41358_n642;
  wire alu__abc_41358_n643;
  wire alu__abc_41358_n644;
  wire alu__abc_41358_n645;
  wire alu__abc_41358_n646;
  wire alu__abc_41358_n647;
  wire alu__abc_41358_n648;
  wire alu__abc_41358_n649;
  wire alu__abc_41358_n650;
  wire alu__abc_41358_n651;
  wire alu__abc_41358_n652;
  wire alu__abc_41358_n653;
  wire alu__abc_41358_n654;
  wire alu__abc_41358_n655;
  wire alu__abc_41358_n656;
  wire alu__abc_41358_n657;
  wire alu__abc_41358_n658;
  wire alu__abc_41358_n659;
  wire alu__abc_41358_n660;
  wire alu__abc_41358_n661;
  wire alu__abc_41358_n662;
  wire alu__abc_41358_n663;
  wire alu__abc_41358_n664;
  wire alu__abc_41358_n665;
  wire alu__abc_41358_n666;
  wire alu__abc_41358_n667;
  wire alu__abc_41358_n668;
  wire alu__abc_41358_n669;
  wire alu__abc_41358_n670;
  wire alu__abc_41358_n671;
  wire alu__abc_41358_n672;
  wire alu__abc_41358_n673;
  wire alu__abc_41358_n674;
  wire alu__abc_41358_n675;
  wire alu__abc_41358_n676;
  wire alu__abc_41358_n677;
  wire alu__abc_41358_n678;
  wire alu__abc_41358_n679;
  wire alu__abc_41358_n680;
  wire alu__abc_41358_n681;
  wire alu__abc_41358_n682;
  wire alu__abc_41358_n683;
  wire alu__abc_41358_n684;
  wire alu__abc_41358_n685;
  wire alu__abc_41358_n686;
  wire alu__abc_41358_n687;
  wire alu__abc_41358_n688;
  wire alu__abc_41358_n689;
  wire alu__abc_41358_n690;
  wire alu__abc_41358_n691;
  wire alu__abc_41358_n692;
  wire alu__abc_41358_n693;
  wire alu__abc_41358_n694;
  wire alu__abc_41358_n695;
  wire alu__abc_41358_n696;
  wire alu__abc_41358_n697;
  wire alu__abc_41358_n698;
  wire alu__abc_41358_n699;
  wire alu__abc_41358_n700;
  wire alu__abc_41358_n701;
  wire alu__abc_41358_n702;
  wire alu__abc_41358_n703;
  wire alu__abc_41358_n704_1;
  wire alu__abc_41358_n705;
  wire alu__abc_41358_n706;
  wire alu__abc_41358_n707;
  wire alu__abc_41358_n708;
  wire alu__abc_41358_n709;
  wire alu__abc_41358_n710;
  wire alu__abc_41358_n711;
  wire alu__abc_41358_n712;
  wire alu__abc_41358_n713;
  wire alu__abc_41358_n714;
  wire alu__abc_41358_n715;
  wire alu__abc_41358_n716;
  wire alu__abc_41358_n717;
  wire alu__abc_41358_n718;
  wire alu__abc_41358_n719;
  wire alu__abc_41358_n720;
  wire alu__abc_41358_n721;
  wire alu__abc_41358_n722;
  wire alu__abc_41358_n723;
  wire alu__abc_41358_n724;
  wire alu__abc_41358_n725;
  wire alu__abc_41358_n726;
  wire alu__abc_41358_n727;
  wire alu__abc_41358_n728;
  wire alu__abc_41358_n729;
  wire alu__abc_41358_n730;
  wire alu__abc_41358_n731;
  wire alu__abc_41358_n732;
  wire alu__abc_41358_n733;
  wire alu__abc_41358_n734;
  wire alu__abc_41358_n735;
  wire alu__abc_41358_n736;
  wire alu__abc_41358_n737;
  wire alu__abc_41358_n738;
  wire alu__abc_41358_n739;
  wire alu__abc_41358_n740;
  wire alu__abc_41358_n741;
  wire alu__abc_41358_n742;
  wire alu__abc_41358_n743;
  wire alu__abc_41358_n744;
  wire alu__abc_41358_n745;
  wire alu__abc_41358_n746;
  wire alu__abc_41358_n747;
  wire alu__abc_41358_n748;
  wire alu__abc_41358_n749;
  wire alu__abc_41358_n750;
  wire alu__abc_41358_n751;
  wire alu__abc_41358_n752;
  wire alu__abc_41358_n753;
  wire alu__abc_41358_n754;
  wire alu__abc_41358_n755_1;
  wire alu__abc_41358_n756;
  wire alu__abc_41358_n757;
  wire alu__abc_41358_n758;
  wire alu__abc_41358_n759;
  wire alu__abc_41358_n760;
  wire alu__abc_41358_n761;
  wire alu__abc_41358_n762;
  wire alu__abc_41358_n763;
  wire alu__abc_41358_n764;
  wire alu__abc_41358_n765;
  wire alu__abc_41358_n766;
  wire alu__abc_41358_n767;
  wire alu__abc_41358_n768;
  wire alu__abc_41358_n769;
  wire alu__abc_41358_n770;
  wire alu__abc_41358_n771;
  wire alu__abc_41358_n772;
  wire alu__abc_41358_n773;
  wire alu__abc_41358_n774;
  wire alu__abc_41358_n775;
  wire alu__abc_41358_n776;
  wire alu__abc_41358_n777;
  wire alu__abc_41358_n778;
  wire alu__abc_41358_n779;
  wire alu__abc_41358_n780;
  wire alu__abc_41358_n781;
  wire alu__abc_41358_n782;
  wire alu__abc_41358_n783;
  wire alu__abc_41358_n784;
  wire alu__abc_41358_n785;
  wire alu__abc_41358_n786;
  wire alu__abc_41358_n787_1;
  wire alu__abc_41358_n788;
  wire alu__abc_41358_n789;
  wire alu__abc_41358_n790;
  wire alu__abc_41358_n791;
  wire alu__abc_41358_n792;
  wire alu__abc_41358_n793;
  wire alu__abc_41358_n794;
  wire alu__abc_41358_n795;
  wire alu__abc_41358_n796;
  wire alu__abc_41358_n797;
  wire alu__abc_41358_n798;
  wire alu__abc_41358_n799;
  wire alu__abc_41358_n800;
  wire alu__abc_41358_n801;
  wire alu__abc_41358_n802;
  wire alu__abc_41358_n803;
  wire alu__abc_41358_n804;
  wire alu__abc_41358_n805;
  wire alu__abc_41358_n806;
  wire alu__abc_41358_n807;
  wire alu__abc_41358_n808;
  wire alu__abc_41358_n809;
  wire alu__abc_41358_n810;
  wire alu__abc_41358_n811;
  wire alu__abc_41358_n812;
  wire alu__abc_41358_n813;
  wire alu__abc_41358_n814;
  wire alu__abc_41358_n815;
  wire alu__abc_41358_n816;
  wire alu__abc_41358_n817;
  wire alu__abc_41358_n818_1;
  wire alu__abc_41358_n819;
  wire alu__abc_41358_n820;
  wire alu__abc_41358_n821;
  wire alu__abc_41358_n822;
  wire alu__abc_41358_n823;
  wire alu__abc_41358_n824;
  wire alu__abc_41358_n825;
  wire alu__abc_41358_n826;
  wire alu__abc_41358_n827;
  wire alu__abc_41358_n828;
  wire alu__abc_41358_n829;
  wire alu__abc_41358_n830;
  wire alu__abc_41358_n832;
  wire alu__abc_41358_n833;
  wire alu__abc_41358_n833_bF_buf0;
  wire alu__abc_41358_n833_bF_buf1;
  wire alu__abc_41358_n833_bF_buf2;
  wire alu__abc_41358_n833_bF_buf3;
  wire alu__abc_41358_n833_bF_buf4;
  wire alu__abc_41358_n834;
  wire alu__abc_41358_n835;
  wire alu__abc_41358_n836;
  wire alu__abc_41358_n837;
  wire alu__abc_41358_n838;
  wire alu__abc_41358_n839;
  wire alu__abc_41358_n840;
  wire alu__abc_41358_n841;
  wire alu__abc_41358_n842;
  wire alu__abc_41358_n843;
  wire alu__abc_41358_n844;
  wire alu__abc_41358_n845;
  wire alu__abc_41358_n846;
  wire alu__abc_41358_n847_1;
  wire alu__abc_41358_n848;
  wire alu__abc_41358_n849;
  wire alu__abc_41358_n850;
  wire alu__abc_41358_n851;
  wire alu__abc_41358_n852;
  wire alu__abc_41358_n853;
  wire alu__abc_41358_n854;
  wire alu__abc_41358_n855;
  wire alu__abc_41358_n856;
  wire alu__abc_41358_n857;
  wire alu__abc_41358_n858;
  wire alu__abc_41358_n859;
  wire alu__abc_41358_n860;
  wire alu__abc_41358_n861;
  wire alu__abc_41358_n862;
  wire alu__abc_41358_n863;
  wire alu__abc_41358_n864;
  wire alu__abc_41358_n865;
  wire alu__abc_41358_n866;
  wire alu__abc_41358_n867;
  wire alu__abc_41358_n868;
  wire alu__abc_41358_n869;
  wire alu__abc_41358_n870;
  wire alu__abc_41358_n871;
  wire alu__abc_41358_n872_1;
  wire alu__abc_41358_n873;
  wire alu__abc_41358_n874;
  wire alu__abc_41358_n875;
  wire alu__abc_41358_n876;
  wire alu__abc_41358_n877;
  wire alu__abc_41358_n878;
  wire alu__abc_41358_n879;
  wire alu__abc_41358_n880;
  wire alu__abc_41358_n881;
  wire alu__abc_41358_n882;
  wire alu__abc_41358_n883;
  wire alu__abc_41358_n884;
  wire alu__abc_41358_n885;
  wire alu__abc_41358_n886;
  wire alu__abc_41358_n887;
  wire alu__abc_41358_n888;
  wire alu__abc_41358_n889;
  wire alu__abc_41358_n890;
  wire alu__abc_41358_n891;
  wire alu__abc_41358_n892;
  wire alu__abc_41358_n893;
  wire alu__abc_41358_n894;
  wire alu__abc_41358_n895;
  wire alu__abc_41358_n896;
  wire alu__abc_41358_n897;
  wire alu__abc_41358_n898;
  wire alu__abc_41358_n899;
  wire alu__abc_41358_n900;
  wire alu__abc_41358_n901;
  wire alu__abc_41358_n902;
  wire alu__abc_41358_n903_1;
  wire alu__abc_41358_n904;
  wire alu__abc_41358_n905;
  wire alu__abc_41358_n906;
  wire alu__abc_41358_n907;
  wire alu__abc_41358_n908;
  wire alu__abc_41358_n909;
  wire alu__abc_41358_n910;
  wire alu__abc_41358_n911;
  wire alu__abc_41358_n912;
  wire alu__abc_41358_n913;
  wire alu__abc_41358_n914;
  wire alu__abc_41358_n915;
  wire alu__abc_41358_n916;
  wire alu__abc_41358_n917;
  wire alu__abc_41358_n918;
  wire alu__abc_41358_n919;
  wire alu__abc_41358_n920;
  wire alu__abc_41358_n921;
  wire alu__abc_41358_n922;
  wire alu__abc_41358_n923;
  wire alu__abc_41358_n924;
  wire alu__abc_41358_n925;
  wire alu__abc_41358_n926;
  wire alu__abc_41358_n927;
  wire alu__abc_41358_n927_bF_buf0;
  wire alu__abc_41358_n927_bF_buf1;
  wire alu__abc_41358_n927_bF_buf2;
  wire alu__abc_41358_n927_bF_buf3;
  wire alu__abc_41358_n927_bF_buf4;
  wire alu__abc_41358_n928;
  wire alu__abc_41358_n929;
  wire alu__abc_41358_n930;
  wire alu__abc_41358_n931;
  wire alu__abc_41358_n932;
  wire alu__abc_41358_n932_bF_buf0;
  wire alu__abc_41358_n932_bF_buf1;
  wire alu__abc_41358_n932_bF_buf2;
  wire alu__abc_41358_n932_bF_buf3;
  wire alu__abc_41358_n932_bF_buf4;
  wire alu__abc_41358_n933_1;
  wire alu__abc_41358_n934;
  wire alu__abc_41358_n935;
  wire alu__abc_41358_n935_bF_buf0;
  wire alu__abc_41358_n935_bF_buf1;
  wire alu__abc_41358_n935_bF_buf2;
  wire alu__abc_41358_n935_bF_buf3;
  wire alu__abc_41358_n935_bF_buf4;
  wire alu__abc_41358_n936;
  wire alu__abc_41358_n937;
  wire alu__abc_41358_n938;
  wire alu__abc_41358_n939;
  wire alu__abc_41358_n940;
  wire alu__abc_41358_n941;
  wire alu__abc_41358_n942;
  wire alu__abc_41358_n942_bF_buf0;
  wire alu__abc_41358_n942_bF_buf1;
  wire alu__abc_41358_n942_bF_buf2;
  wire alu__abc_41358_n942_bF_buf3;
  wire alu__abc_41358_n942_bF_buf4;
  wire alu__abc_41358_n943;
  wire alu__abc_41358_n944;
  wire alu__abc_41358_n945;
  wire alu__abc_41358_n946;
  wire alu__abc_41358_n947;
  wire alu__abc_41358_n948;
  wire alu__abc_41358_n948_bF_buf0;
  wire alu__abc_41358_n948_bF_buf1;
  wire alu__abc_41358_n948_bF_buf2;
  wire alu__abc_41358_n948_bF_buf3;
  wire alu__abc_41358_n948_bF_buf4;
  wire alu__abc_41358_n949;
  wire alu__abc_41358_n950;
  wire alu__abc_41358_n951;
  wire alu__abc_41358_n952;
  wire alu__abc_41358_n953_1;
  wire alu__abc_41358_n954;
  wire alu__abc_41358_n955;
  wire alu__abc_41358_n956;
  wire alu__abc_41358_n957;
  wire alu__abc_41358_n958;
  wire alu__abc_41358_n959;
  wire alu__abc_41358_n961;
  wire alu__abc_41358_n962;
  wire alu__abc_41358_n963;
  wire alu__abc_41358_n964;
  wire alu__abc_41358_n965;
  wire alu__abc_41358_n966;
  wire alu__abc_41358_n967;
  wire alu__abc_41358_n968;
  wire alu__abc_41358_n969;
  wire alu__abc_41358_n970;
  wire alu__abc_41358_n971;
  wire alu__abc_41358_n972;
  wire alu__abc_41358_n973;
  wire alu__abc_41358_n974;
  wire alu__abc_41358_n975_1;
  wire alu__abc_41358_n976;
  wire alu__abc_41358_n977;
  wire alu__abc_41358_n978;
  wire alu__abc_41358_n979;
  wire alu__abc_41358_n980;
  wire alu__abc_41358_n981;
  wire alu__abc_41358_n982;
  wire alu__abc_41358_n983;
  wire alu__abc_41358_n984;
  wire alu__abc_41358_n985;
  wire alu__abc_41358_n986;
  wire alu__abc_41358_n987;
  wire alu__abc_41358_n988;
  wire alu__abc_41358_n989;
  wire alu__abc_41358_n990;
  wire alu__abc_41358_n991;
  wire alu__abc_41358_n992;
  wire alu__abc_41358_n993;
  wire alu__abc_41358_n994;
  wire alu__abc_41358_n995;
  wire alu__abc_41358_n996;
  wire alu__abc_41358_n997;
  wire alu__abc_41358_n998;
  wire alu__abc_41358_n999;
  wire alu_a_i_0_;
  wire alu_a_i_10_;
  wire alu_a_i_11_;
  wire alu_a_i_12_;
  wire alu_a_i_13_;
  wire alu_a_i_14_;
  wire alu_a_i_15_;
  wire alu_a_i_16_;
  wire alu_a_i_17_;
  wire alu_a_i_18_;
  wire alu_a_i_19_;
  wire alu_a_i_1_;
  wire alu_a_i_20_;
  wire alu_a_i_21_;
  wire alu_a_i_22_;
  wire alu_a_i_23_;
  wire alu_a_i_24_;
  wire alu_a_i_25_;
  wire alu_a_i_26_;
  wire alu_a_i_27_;
  wire alu_a_i_28_;
  wire alu_a_i_29_;
  wire alu_a_i_2_;
  wire alu_a_i_30_;
  wire alu_a_i_31_;
  wire alu_a_i_3_;
  wire alu_a_i_4_;
  wire alu_a_i_5_;
  wire alu_a_i_6_;
  wire alu_a_i_7_;
  wire alu_a_i_8_;
  wire alu_a_i_9_;
  wire alu_b_i_0_;
  wire alu_b_i_0_bF_buf0;
  wire alu_b_i_0_bF_buf1;
  wire alu_b_i_0_bF_buf2;
  wire alu_b_i_0_bF_buf3;
  wire alu_b_i_0_bF_buf4;
  wire alu_b_i_10_;
  wire alu_b_i_11_;
  wire alu_b_i_12_;
  wire alu_b_i_13_;
  wire alu_b_i_14_;
  wire alu_b_i_15_;
  wire alu_b_i_16_;
  wire alu_b_i_17_;
  wire alu_b_i_18_;
  wire alu_b_i_19_;
  wire alu_b_i_1_;
  wire alu_b_i_1_bF_buf0;
  wire alu_b_i_1_bF_buf1;
  wire alu_b_i_1_bF_buf2;
  wire alu_b_i_1_bF_buf3;
  wire alu_b_i_1_bF_buf4;
  wire alu_b_i_1_bF_buf5;
  wire alu_b_i_1_bF_buf6;
  wire alu_b_i_1_bF_buf7;
  wire alu_b_i_20_;
  wire alu_b_i_21_;
  wire alu_b_i_22_;
  wire alu_b_i_23_;
  wire alu_b_i_24_;
  wire alu_b_i_25_;
  wire alu_b_i_26_;
  wire alu_b_i_27_;
  wire alu_b_i_28_;
  wire alu_b_i_29_;
  wire alu_b_i_2_;
  wire alu_b_i_2_bF_buf0;
  wire alu_b_i_2_bF_buf1;
  wire alu_b_i_2_bF_buf2;
  wire alu_b_i_2_bF_buf3;
  wire alu_b_i_2_bF_buf4;
  wire alu_b_i_2_bF_buf5;
  wire alu_b_i_2_bF_buf6;
  wire alu_b_i_30_;
  wire alu_b_i_31_;
  wire alu_b_i_3_;
  wire alu_b_i_3_bF_buf0;
  wire alu_b_i_3_bF_buf1;
  wire alu_b_i_3_bF_buf2;
  wire alu_b_i_3_bF_buf3;
  wire alu_b_i_3_bF_buf4;
  wire alu_b_i_3_bF_buf5;
  wire alu_b_i_3_bF_buf6;
  wire alu_b_i_4_;
  wire alu_b_i_4_bF_buf0;
  wire alu_b_i_4_bF_buf1;
  wire alu_b_i_4_bF_buf2;
  wire alu_b_i_4_bF_buf3;
  wire alu_b_i_4_bF_buf4;
  wire alu_b_i_5_;
  wire alu_b_i_6_;
  wire alu_b_i_7_;
  wire alu_b_i_8_;
  wire alu_b_i_9_;
  wire alu_c_i;
  wire alu_c_o;
  wire alu_c_update_o;
  wire alu_equal_o;
  wire alu_flag_update_o;
  wire alu_func_r_0_;
  wire alu_func_r_1_;
  wire alu_func_r_2_;
  wire alu_func_r_3_;
  wire alu_greater_than_o;
  wire alu_greater_than_signed_o;
  wire alu_input_a_r_0_;
  wire alu_input_a_r_10_;
  wire alu_input_a_r_11_;
  wire alu_input_a_r_12_;
  wire alu_input_a_r_13_;
  wire alu_input_a_r_14_;
  wire alu_input_a_r_15_;
  wire alu_input_a_r_16_;
  wire alu_input_a_r_17_;
  wire alu_input_a_r_18_;
  wire alu_input_a_r_19_;
  wire alu_input_a_r_1_;
  wire alu_input_a_r_20_;
  wire alu_input_a_r_21_;
  wire alu_input_a_r_22_;
  wire alu_input_a_r_23_;
  wire alu_input_a_r_24_;
  wire alu_input_a_r_25_;
  wire alu_input_a_r_26_;
  wire alu_input_a_r_27_;
  wire alu_input_a_r_28_;
  wire alu_input_a_r_29_;
  wire alu_input_a_r_2_;
  wire alu_input_a_r_30_;
  wire alu_input_a_r_31_;
  wire alu_input_a_r_3_;
  wire alu_input_a_r_4_;
  wire alu_input_a_r_5_;
  wire alu_input_a_r_6_;
  wire alu_input_a_r_7_;
  wire alu_input_a_r_8_;
  wire alu_input_a_r_9_;
  wire alu_input_b_r_0_;
  wire alu_input_b_r_10_;
  wire alu_input_b_r_11_;
  wire alu_input_b_r_12_;
  wire alu_input_b_r_13_;
  wire alu_input_b_r_14_;
  wire alu_input_b_r_15_;
  wire alu_input_b_r_16_;
  wire alu_input_b_r_17_;
  wire alu_input_b_r_18_;
  wire alu_input_b_r_19_;
  wire alu_input_b_r_1_;
  wire alu_input_b_r_20_;
  wire alu_input_b_r_21_;
  wire alu_input_b_r_22_;
  wire alu_input_b_r_23_;
  wire alu_input_b_r_24_;
  wire alu_input_b_r_25_;
  wire alu_input_b_r_26_;
  wire alu_input_b_r_27_;
  wire alu_input_b_r_28_;
  wire alu_input_b_r_29_;
  wire alu_input_b_r_2_;
  wire alu_input_b_r_30_;
  wire alu_input_b_r_31_;
  wire alu_input_b_r_3_;
  wire alu_input_b_r_4_;
  wire alu_input_b_r_5_;
  wire alu_input_b_r_6_;
  wire alu_input_b_r_7_;
  wire alu_input_b_r_8_;
  wire alu_input_b_r_9_;
  wire alu_less_than_o;
  wire alu_less_than_signed_o;
  wire alu_op_i_0_;
  wire alu_op_i_0_bF_buf0;
  wire alu_op_i_0_bF_buf1;
  wire alu_op_i_0_bF_buf2;
  wire alu_op_i_0_bF_buf3;
  wire alu_op_i_0_bF_buf4;
  wire alu_op_i_0_bF_buf5;
  wire alu_op_i_1_;
  wire alu_op_i_2_;
  wire alu_op_i_3_;
  wire alu_op_r_0_;
  wire alu_op_r_1_;
  wire alu_op_r_2_;
  wire alu_op_r_3_;
  wire alu_op_r_4_;
  wire alu_op_r_5_;
  wire alu_op_r_6_;
  wire alu_op_r_7_;
  wire alu_p_o_0_;
  wire alu_p_o_10_;
  wire alu_p_o_11_;
  wire alu_p_o_12_;
  wire alu_p_o_13_;
  wire alu_p_o_14_;
  wire alu_p_o_15_;
  wire alu_p_o_16_;
  wire alu_p_o_17_;
  wire alu_p_o_18_;
  wire alu_p_o_19_;
  wire alu_p_o_1_;
  wire alu_p_o_20_;
  wire alu_p_o_21_;
  wire alu_p_o_22_;
  wire alu_p_o_23_;
  wire alu_p_o_24_;
  wire alu_p_o_25_;
  wire alu_p_o_26_;
  wire alu_p_o_27_;
  wire alu_p_o_28_;
  wire alu_p_o_29_;
  wire alu_p_o_2_;
  wire alu_p_o_30_;
  wire alu_p_o_31_;
  wire alu_p_o_3_;
  wire alu_p_o_4_;
  wire alu_p_o_5_;
  wire alu_p_o_6_;
  wire alu_p_o_7_;
  wire alu_p_o_8_;
  wire alu_p_o_9_;
  output break_o;
  input clk_i;
  wire clk_i_bF_buf0;
  wire clk_i_bF_buf1;
  wire clk_i_bF_buf10;
  wire clk_i_bF_buf100;
  wire clk_i_bF_buf101;
  wire clk_i_bF_buf102;
  wire clk_i_bF_buf103;
  wire clk_i_bF_buf104;
  wire clk_i_bF_buf105;
  wire clk_i_bF_buf106;
  wire clk_i_bF_buf107;
  wire clk_i_bF_buf108;
  wire clk_i_bF_buf109;
  wire clk_i_bF_buf11;
  wire clk_i_bF_buf110;
  wire clk_i_bF_buf111;
  wire clk_i_bF_buf112;
  wire clk_i_bF_buf113;
  wire clk_i_bF_buf114;
  wire clk_i_bF_buf12;
  wire clk_i_bF_buf13;
  wire clk_i_bF_buf14;
  wire clk_i_bF_buf15;
  wire clk_i_bF_buf16;
  wire clk_i_bF_buf17;
  wire clk_i_bF_buf18;
  wire clk_i_bF_buf19;
  wire clk_i_bF_buf2;
  wire clk_i_bF_buf20;
  wire clk_i_bF_buf21;
  wire clk_i_bF_buf22;
  wire clk_i_bF_buf23;
  wire clk_i_bF_buf24;
  wire clk_i_bF_buf25;
  wire clk_i_bF_buf26;
  wire clk_i_bF_buf27;
  wire clk_i_bF_buf28;
  wire clk_i_bF_buf29;
  wire clk_i_bF_buf3;
  wire clk_i_bF_buf30;
  wire clk_i_bF_buf31;
  wire clk_i_bF_buf32;
  wire clk_i_bF_buf33;
  wire clk_i_bF_buf34;
  wire clk_i_bF_buf35;
  wire clk_i_bF_buf36;
  wire clk_i_bF_buf37;
  wire clk_i_bF_buf38;
  wire clk_i_bF_buf39;
  wire clk_i_bF_buf4;
  wire clk_i_bF_buf40;
  wire clk_i_bF_buf41;
  wire clk_i_bF_buf42;
  wire clk_i_bF_buf43;
  wire clk_i_bF_buf44;
  wire clk_i_bF_buf45;
  wire clk_i_bF_buf46;
  wire clk_i_bF_buf47;
  wire clk_i_bF_buf48;
  wire clk_i_bF_buf49;
  wire clk_i_bF_buf5;
  wire clk_i_bF_buf50;
  wire clk_i_bF_buf51;
  wire clk_i_bF_buf52;
  wire clk_i_bF_buf53;
  wire clk_i_bF_buf54;
  wire clk_i_bF_buf55;
  wire clk_i_bF_buf56;
  wire clk_i_bF_buf57;
  wire clk_i_bF_buf58;
  wire clk_i_bF_buf59;
  wire clk_i_bF_buf6;
  wire clk_i_bF_buf60;
  wire clk_i_bF_buf61;
  wire clk_i_bF_buf62;
  wire clk_i_bF_buf63;
  wire clk_i_bF_buf64;
  wire clk_i_bF_buf65;
  wire clk_i_bF_buf66;
  wire clk_i_bF_buf67;
  wire clk_i_bF_buf68;
  wire clk_i_bF_buf69;
  wire clk_i_bF_buf7;
  wire clk_i_bF_buf70;
  wire clk_i_bF_buf71;
  wire clk_i_bF_buf72;
  wire clk_i_bF_buf73;
  wire clk_i_bF_buf74;
  wire clk_i_bF_buf75;
  wire clk_i_bF_buf76;
  wire clk_i_bF_buf77;
  wire clk_i_bF_buf78;
  wire clk_i_bF_buf79;
  wire clk_i_bF_buf8;
  wire clk_i_bF_buf80;
  wire clk_i_bF_buf81;
  wire clk_i_bF_buf82;
  wire clk_i_bF_buf83;
  wire clk_i_bF_buf84;
  wire clk_i_bF_buf85;
  wire clk_i_bF_buf86;
  wire clk_i_bF_buf87;
  wire clk_i_bF_buf88;
  wire clk_i_bF_buf89;
  wire clk_i_bF_buf9;
  wire clk_i_bF_buf90;
  wire clk_i_bF_buf91;
  wire clk_i_bF_buf92;
  wire clk_i_bF_buf93;
  wire clk_i_bF_buf94;
  wire clk_i_bF_buf95;
  wire clk_i_bF_buf96;
  wire clk_i_bF_buf97;
  wire clk_i_bF_buf98;
  wire clk_i_bF_buf99;
  wire clk_i_hier0_bF_buf0;
  wire clk_i_hier0_bF_buf1;
  wire clk_i_hier0_bF_buf2;
  wire clk_i_hier0_bF_buf3;
  wire clk_i_hier0_bF_buf4;
  wire clk_i_hier0_bF_buf5;
  wire clk_i_hier0_bF_buf6;
  wire clk_i_hier0_bF_buf7;
  wire clk_i_hier0_bF_buf8;
  wire clk_i_hier0_bF_buf9;
  input enable_i;
  wire enable_i_bF_buf0;
  wire enable_i_bF_buf1;
  wire enable_i_bF_buf2;
  wire enable_i_bF_buf3;
  wire enable_i_bF_buf4;
  wire enable_i_bF_buf5;
  wire enable_i_bF_buf6;
  wire enable_i_bF_buf7;
  wire epc_q_0_;
  wire epc_q_0__FF_INPUT;
  wire epc_q_10_;
  wire epc_q_10__FF_INPUT;
  wire epc_q_11_;
  wire epc_q_11__FF_INPUT;
  wire epc_q_12_;
  wire epc_q_12__FF_INPUT;
  wire epc_q_13_;
  wire epc_q_13__FF_INPUT;
  wire epc_q_14_;
  wire epc_q_14__FF_INPUT;
  wire epc_q_15_;
  wire epc_q_15__FF_INPUT;
  wire epc_q_16_;
  wire epc_q_16__FF_INPUT;
  wire epc_q_17_;
  wire epc_q_17__FF_INPUT;
  wire epc_q_18_;
  wire epc_q_18__FF_INPUT;
  wire epc_q_19_;
  wire epc_q_19__FF_INPUT;
  wire epc_q_1_;
  wire epc_q_1__FF_INPUT;
  wire epc_q_20_;
  wire epc_q_20__FF_INPUT;
  wire epc_q_21_;
  wire epc_q_21__FF_INPUT;
  wire epc_q_22_;
  wire epc_q_22__FF_INPUT;
  wire epc_q_23_;
  wire epc_q_23__FF_INPUT;
  wire epc_q_24_;
  wire epc_q_24__FF_INPUT;
  wire epc_q_25_;
  wire epc_q_25__FF_INPUT;
  wire epc_q_26_;
  wire epc_q_26__FF_INPUT;
  wire epc_q_27_;
  wire epc_q_27__FF_INPUT;
  wire epc_q_28_;
  wire epc_q_28__FF_INPUT;
  wire epc_q_29_;
  wire epc_q_29__FF_INPUT;
  wire epc_q_2_;
  wire epc_q_2__FF_INPUT;
  wire epc_q_30_;
  wire epc_q_30__FF_INPUT;
  wire epc_q_31_;
  wire epc_q_31__FF_INPUT;
  wire epc_q_3_;
  wire epc_q_3__FF_INPUT;
  wire epc_q_4_;
  wire epc_q_4__FF_INPUT;
  wire epc_q_5_;
  wire epc_q_5__FF_INPUT;
  wire epc_q_6_;
  wire epc_q_6__FF_INPUT;
  wire epc_q_7_;
  wire epc_q_7__FF_INPUT;
  wire epc_q_8_;
  wire epc_q_8__FF_INPUT;
  wire epc_q_9_;
  wire epc_q_9__FF_INPUT;
  wire esr_q_10_;
  wire esr_q_10__FF_INPUT;
  wire esr_q_2_;
  wire esr_q_2__FF_INPUT;
  wire esr_q_9_;
  wire esr_q_9__FF_INPUT;
  wire ex_rd_q_0__FF_INPUT;
  wire ex_rd_q_1__FF_INPUT;
  wire ex_rd_q_2__FF_INPUT;
  wire ex_rd_q_3__FF_INPUT;
  wire ex_rd_q_4__FF_INPUT;
  output fault_o;
  wire fault_o_FF_INPUT;
  wire inst_r_0_;
  wire inst_r_1_;
  wire inst_r_2_;
  wire inst_r_3_;
  wire inst_r_4_;
  wire inst_r_5_;
  wire inst_trap_w;
  wire int32_r_10_;
  wire int32_r_4_;
  wire int32_r_5_;
  input intr_i;
  input mem_ack_i;
  output \mem_addr_o[0] ;
  output \mem_addr_o[10] ;
  output \mem_addr_o[11] ;
  output \mem_addr_o[12] ;
  output \mem_addr_o[13] ;
  output \mem_addr_o[14] ;
  output \mem_addr_o[15] ;
  output \mem_addr_o[16] ;
  output \mem_addr_o[17] ;
  output \mem_addr_o[18] ;
  output \mem_addr_o[19] ;
  output \mem_addr_o[1] ;
  output \mem_addr_o[20] ;
  output \mem_addr_o[21] ;
  output \mem_addr_o[22] ;
  output \mem_addr_o[23] ;
  output \mem_addr_o[24] ;
  output \mem_addr_o[25] ;
  output \mem_addr_o[26] ;
  output \mem_addr_o[27] ;
  output \mem_addr_o[28] ;
  output \mem_addr_o[29] ;
  output \mem_addr_o[2] ;
  output \mem_addr_o[30] ;
  output \mem_addr_o[31] ;
  output \mem_addr_o[3] ;
  output \mem_addr_o[4] ;
  output \mem_addr_o[5] ;
  output \mem_addr_o[6] ;
  output \mem_addr_o[7] ;
  output \mem_addr_o[8] ;
  output \mem_addr_o[9] ;
  wire mem_addr_o_0__FF_INPUT;
  wire mem_addr_o_10__FF_INPUT;
  wire mem_addr_o_11__FF_INPUT;
  wire mem_addr_o_12__FF_INPUT;
  wire mem_addr_o_13__FF_INPUT;
  wire mem_addr_o_14__FF_INPUT;
  wire mem_addr_o_15__FF_INPUT;
  wire mem_addr_o_16__FF_INPUT;
  wire mem_addr_o_17__FF_INPUT;
  wire mem_addr_o_18__FF_INPUT;
  wire mem_addr_o_19__FF_INPUT;
  wire mem_addr_o_1__FF_INPUT;
  wire mem_addr_o_20__FF_INPUT;
  wire mem_addr_o_21__FF_INPUT;
  wire mem_addr_o_22__FF_INPUT;
  wire mem_addr_o_23__FF_INPUT;
  wire mem_addr_o_24__FF_INPUT;
  wire mem_addr_o_25__FF_INPUT;
  wire mem_addr_o_26__FF_INPUT;
  wire mem_addr_o_27__FF_INPUT;
  wire mem_addr_o_28__FF_INPUT;
  wire mem_addr_o_29__FF_INPUT;
  wire mem_addr_o_2__FF_INPUT;
  wire mem_addr_o_30__FF_INPUT;
  wire mem_addr_o_31__FF_INPUT;
  wire mem_addr_o_3__FF_INPUT;
  wire mem_addr_o_4__FF_INPUT;
  wire mem_addr_o_5__FF_INPUT;
  wire mem_addr_o_6__FF_INPUT;
  wire mem_addr_o_7__FF_INPUT;
  wire mem_addr_o_8__FF_INPUT;
  wire mem_addr_o_9__FF_INPUT;
  output \mem_cti_o[0] ;
  output \mem_cti_o[1] ;
  output \mem_cti_o[2] ;
  output mem_cyc_o;
  wire mem_cyc_o_FF_INPUT;
  input \mem_dat_i[0] ;
  input \mem_dat_i[10] ;
  input \mem_dat_i[11] ;
  input \mem_dat_i[12] ;
  input \mem_dat_i[13] ;
  input \mem_dat_i[14] ;
  input \mem_dat_i[15] ;
  input \mem_dat_i[16] ;
  input \mem_dat_i[17] ;
  input \mem_dat_i[18] ;
  input \mem_dat_i[19] ;
  input \mem_dat_i[1] ;
  input \mem_dat_i[20] ;
  input \mem_dat_i[21] ;
  input \mem_dat_i[22] ;
  input \mem_dat_i[23] ;
  input \mem_dat_i[24] ;
  input \mem_dat_i[25] ;
  input \mem_dat_i[26] ;
  input \mem_dat_i[27] ;
  input \mem_dat_i[28] ;
  input \mem_dat_i[29] ;
  input \mem_dat_i[2] ;
  input \mem_dat_i[30] ;
  input \mem_dat_i[31] ;
  input \mem_dat_i[3] ;
  input \mem_dat_i[4] ;
  input \mem_dat_i[5] ;
  input \mem_dat_i[6] ;
  input \mem_dat_i[7] ;
  input \mem_dat_i[8] ;
  input \mem_dat_i[9] ;
  output \mem_dat_o[0] ;
  output \mem_dat_o[10] ;
  output \mem_dat_o[11] ;
  output \mem_dat_o[12] ;
  output \mem_dat_o[13] ;
  output \mem_dat_o[14] ;
  output \mem_dat_o[15] ;
  output \mem_dat_o[16] ;
  output \mem_dat_o[17] ;
  output \mem_dat_o[18] ;
  output \mem_dat_o[19] ;
  output \mem_dat_o[1] ;
  output \mem_dat_o[20] ;
  output \mem_dat_o[21] ;
  output \mem_dat_o[22] ;
  output \mem_dat_o[23] ;
  output \mem_dat_o[24] ;
  output \mem_dat_o[25] ;
  output \mem_dat_o[26] ;
  output \mem_dat_o[27] ;
  output \mem_dat_o[28] ;
  output \mem_dat_o[29] ;
  output \mem_dat_o[2] ;
  output \mem_dat_o[30] ;
  output \mem_dat_o[31] ;
  output \mem_dat_o[3] ;
  output \mem_dat_o[4] ;
  output \mem_dat_o[5] ;
  output \mem_dat_o[6] ;
  output \mem_dat_o[7] ;
  output \mem_dat_o[8] ;
  output \mem_dat_o[9] ;
  wire mem_dat_o_0__FF_INPUT;
  wire mem_dat_o_10__FF_INPUT;
  wire mem_dat_o_11__FF_INPUT;
  wire mem_dat_o_12__FF_INPUT;
  wire mem_dat_o_13__FF_INPUT;
  wire mem_dat_o_14__FF_INPUT;
  wire mem_dat_o_15__FF_INPUT;
  wire mem_dat_o_16__FF_INPUT;
  wire mem_dat_o_17__FF_INPUT;
  wire mem_dat_o_18__FF_INPUT;
  wire mem_dat_o_19__FF_INPUT;
  wire mem_dat_o_1__FF_INPUT;
  wire mem_dat_o_20__FF_INPUT;
  wire mem_dat_o_21__FF_INPUT;
  wire mem_dat_o_22__FF_INPUT;
  wire mem_dat_o_23__FF_INPUT;
  wire mem_dat_o_24__FF_INPUT;
  wire mem_dat_o_25__FF_INPUT;
  wire mem_dat_o_26__FF_INPUT;
  wire mem_dat_o_27__FF_INPUT;
  wire mem_dat_o_28__FF_INPUT;
  wire mem_dat_o_29__FF_INPUT;
  wire mem_dat_o_2__FF_INPUT;
  wire mem_dat_o_30__FF_INPUT;
  wire mem_dat_o_31__FF_INPUT;
  wire mem_dat_o_3__FF_INPUT;
  wire mem_dat_o_4__FF_INPUT;
  wire mem_dat_o_5__FF_INPUT;
  wire mem_dat_o_6__FF_INPUT;
  wire mem_dat_o_7__FF_INPUT;
  wire mem_dat_o_8__FF_INPUT;
  wire mem_dat_o_9__FF_INPUT;
  wire mem_offset_q_0_;
  wire mem_offset_q_0__FF_INPUT;
  wire mem_offset_q_1_;
  wire mem_offset_q_1__FF_INPUT;
  output \mem_sel_o[0] ;
  output \mem_sel_o[1] ;
  output \mem_sel_o[2] ;
  output \mem_sel_o[3] ;
  wire mem_sel_o_0__FF_INPUT;
  wire mem_sel_o_1__FF_INPUT;
  wire mem_sel_o_2__FF_INPUT;
  wire mem_sel_o_3__FF_INPUT;
  input mem_stall_i;
  output mem_stb_o;
  wire mem_stb_o_FF_INPUT;
  output mem_we_o;
  wire mem_we_o_FF_INPUT;
  wire next_pc_r_0_;
  wire next_pc_r_1_;
  input nmi_i;
  wire nmi_q;
  wire nmi_q_FF_INPUT;
  wire opcode_q_0__FF_INPUT;
  wire opcode_q_10__FF_INPUT;
  wire opcode_q_11__FF_INPUT;
  wire opcode_q_12__FF_INPUT;
  wire opcode_q_13__FF_INPUT;
  wire opcode_q_14__FF_INPUT;
  wire opcode_q_15__FF_INPUT;
  wire opcode_q_16__FF_INPUT;
  wire opcode_q_17__FF_INPUT;
  wire opcode_q_18__FF_INPUT;
  wire opcode_q_19__FF_INPUT;
  wire opcode_q_1__FF_INPUT;
  wire opcode_q_20__FF_INPUT;
  wire opcode_q_21_;
  wire opcode_q_21__FF_INPUT;
  wire opcode_q_22_;
  wire opcode_q_22__FF_INPUT;
  wire opcode_q_23_;
  wire opcode_q_23__FF_INPUT;
  wire opcode_q_24_;
  wire opcode_q_24__FF_INPUT;
  wire opcode_q_25_;
  wire opcode_q_25__FF_INPUT;
  wire opcode_q_26__FF_INPUT;
  wire opcode_q_27__FF_INPUT;
  wire opcode_q_28__FF_INPUT;
  wire opcode_q_29__FF_INPUT;
  wire opcode_q_2__FF_INPUT;
  wire opcode_q_30__FF_INPUT;
  wire opcode_q_31__FF_INPUT;
  wire opcode_q_3__FF_INPUT;
  wire opcode_q_4__FF_INPUT;
  wire opcode_q_5__FF_INPUT;
  wire opcode_q_6__FF_INPUT;
  wire opcode_q_7__FF_INPUT;
  wire opcode_q_8__FF_INPUT;
  wire opcode_q_9__FF_INPUT;
  wire pc_q_0__FF_INPUT;
  wire pc_q_10_;
  wire pc_q_10__FF_INPUT;
  wire pc_q_11_;
  wire pc_q_11__FF_INPUT;
  wire pc_q_12_;
  wire pc_q_12__FF_INPUT;
  wire pc_q_13_;
  wire pc_q_13__FF_INPUT;
  wire pc_q_14_;
  wire pc_q_14__FF_INPUT;
  wire pc_q_15_;
  wire pc_q_15__FF_INPUT;
  wire pc_q_16_;
  wire pc_q_16__FF_INPUT;
  wire pc_q_17_;
  wire pc_q_17__FF_INPUT;
  wire pc_q_18_;
  wire pc_q_18__FF_INPUT;
  wire pc_q_19_;
  wire pc_q_19__FF_INPUT;
  wire pc_q_1__FF_INPUT;
  wire pc_q_20_;
  wire pc_q_20__FF_INPUT;
  wire pc_q_21_;
  wire pc_q_21__FF_INPUT;
  wire pc_q_22_;
  wire pc_q_22__FF_INPUT;
  wire pc_q_23_;
  wire pc_q_23__FF_INPUT;
  wire pc_q_24_;
  wire pc_q_24__FF_INPUT;
  wire pc_q_25_;
  wire pc_q_25__FF_INPUT;
  wire pc_q_26_;
  wire pc_q_26__FF_INPUT;
  wire pc_q_27_;
  wire pc_q_27__FF_INPUT;
  wire pc_q_28_;
  wire pc_q_28__FF_INPUT;
  wire pc_q_29_;
  wire pc_q_29__FF_INPUT;
  wire pc_q_2_;
  wire pc_q_2__FF_INPUT;
  wire pc_q_30_;
  wire pc_q_30__FF_INPUT;
  wire pc_q_31_;
  wire pc_q_31__FF_INPUT;
  wire pc_q_3_;
  wire pc_q_3__FF_INPUT;
  wire pc_q_4_;
  wire pc_q_4__FF_INPUT;
  wire pc_q_5_;
  wire pc_q_5__FF_INPUT;
  wire pc_q_6_;
  wire pc_q_6__FF_INPUT;
  wire pc_q_7_;
  wire pc_q_7__FF_INPUT;
  wire pc_q_8_;
  wire pc_q_8__FF_INPUT;
  wire pc_q_9_;
  wire pc_q_9__FF_INPUT;
  input rst_i;
  wire sr_q_10__FF_INPUT;
  wire sr_q_2_;
  wire sr_q_2__FF_INPUT;
  wire sr_q_9_;
  wire sr_q_9__FF_INPUT;
  wire state_q_0_;
  wire state_q_1_;
  wire state_q_1_bF_buf0;
  wire state_q_1_bF_buf1;
  wire state_q_1_bF_buf2;
  wire state_q_1_bF_buf3;
  wire state_q_1_bF_buf4;
  wire state_q_2_;
  wire state_q_3_;
  wire state_q_3_bF_buf0;
  wire state_q_3_bF_buf1;
  wire state_q_3_bF_buf2;
  wire state_q_3_bF_buf3;
  wire state_q_3_bF_buf4;
  wire state_q_3_bF_buf5;
  wire state_q_4_;
  wire state_q_5_;
  AND2X2 AND2X2_1 ( .A(mem_ack_i), .B(state_q_1_bF_buf4), .Y(_abc_43815_n617) );
  AND2X2 AND2X2_10 ( .A(_abc_43815_n634), .B(state_q_4_), .Y(_abc_43815_n635) );
  AND2X2 AND2X2_100 ( .A(_abc_43815_n781_1), .B(_abc_43815_n686_1_bF_buf4), .Y(_abc_43815_n782_1) );
  AND2X2 AND2X2_1000 ( .A(_abc_43815_n2543), .B(_abc_43815_n2545), .Y(epc_q_29__FF_INPUT) );
  AND2X2 AND2X2_1001 ( .A(_abc_43815_n2512), .B(pc_q_30_), .Y(_abc_43815_n2548) );
  AND2X2 AND2X2_1002 ( .A(_abc_43815_n2549), .B(_abc_43815_n2547), .Y(_abc_43815_n2550) );
  AND2X2 AND2X2_1003 ( .A(_abc_43815_n2550), .B(_abc_43815_n1461_bF_buf0), .Y(_abc_43815_n2551) );
  AND2X2 AND2X2_1004 ( .A(_abc_43815_n2486), .B(_abc_43815_n2522), .Y(_abc_43815_n2553) );
  AND2X2 AND2X2_1005 ( .A(_abc_43815_n2482), .B(_abc_43815_n2553), .Y(_abc_43815_n2554) );
  AND2X2 AND2X2_1006 ( .A(_abc_43815_n2485), .B(_abc_43815_n2521), .Y(_abc_43815_n2555) );
  AND2X2 AND2X2_1007 ( .A(opcode_q_25_), .B(pc_q_30_), .Y(_abc_43815_n2559) );
  AND2X2 AND2X2_1008 ( .A(_abc_43815_n2560), .B(_abc_43815_n2558), .Y(_abc_43815_n2561) );
  AND2X2 AND2X2_1009 ( .A(_abc_43815_n2557), .B(_abc_43815_n2561), .Y(_abc_43815_n2562) );
  AND2X2 AND2X2_101 ( .A(_abc_43815_n689), .B(\mem_dat_i[29] ), .Y(_abc_43815_n783) );
  AND2X2 AND2X2_1010 ( .A(_abc_43815_n2564), .B(_abc_43815_n1425_1_bF_buf0), .Y(_abc_43815_n2565_1) );
  AND2X2 AND2X2_1011 ( .A(_abc_43815_n2565_1), .B(_abc_43815_n2563), .Y(_abc_43815_n2566) );
  AND2X2 AND2X2_1012 ( .A(_abc_43815_n1065_1_bF_buf1), .B(epc_q_30_), .Y(_abc_43815_n2567) );
  AND2X2 AND2X2_1013 ( .A(_abc_43815_n2569), .B(_abc_43815_n2570), .Y(_abc_43815_n2571) );
  AND2X2 AND2X2_1014 ( .A(_abc_43815_n2573), .B(_abc_43815_n2572), .Y(_abc_43815_n2574) );
  AND2X2 AND2X2_1015 ( .A(_abc_43815_n1418_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_43815_n2576) );
  AND2X2 AND2X2_1016 ( .A(_abc_43815_n1489_bF_buf0), .B(epc_q_30_), .Y(_abc_43815_n2577) );
  AND2X2 AND2X2_1017 ( .A(_abc_43815_n2579), .B(_abc_43815_n1351_bF_buf1), .Y(_abc_43815_n2580) );
  AND2X2 AND2X2_1018 ( .A(_abc_43815_n2575), .B(_abc_43815_n2580), .Y(_abc_43815_n2581) );
  AND2X2 AND2X2_1019 ( .A(_abc_43815_n2583), .B(enable_i_bF_buf1), .Y(_abc_43815_n2584) );
  AND2X2 AND2X2_102 ( .A(_abc_43815_n696), .B(\mem_dat_i[13] ), .Y(_abc_43815_n784) );
  AND2X2 AND2X2_1020 ( .A(_abc_43815_n2582), .B(_abc_43815_n2584), .Y(epc_q_30__FF_INPUT) );
  AND2X2 AND2X2_1021 ( .A(_abc_43815_n2548), .B(pc_q_31_), .Y(_abc_43815_n2587) );
  AND2X2 AND2X2_1022 ( .A(_abc_43815_n2588), .B(_abc_43815_n2586), .Y(_abc_43815_n2589_1) );
  AND2X2 AND2X2_1023 ( .A(_abc_43815_n2589_1), .B(_abc_43815_n1461_bF_buf3), .Y(_abc_43815_n2590) );
  AND2X2 AND2X2_1024 ( .A(_abc_43815_n2594), .B(_abc_43815_n2596), .Y(_abc_43815_n2597) );
  AND2X2 AND2X2_1025 ( .A(_abc_43815_n2600), .B(_abc_43815_n1425_1_bF_buf4), .Y(_abc_43815_n2601) );
  AND2X2 AND2X2_1026 ( .A(_abc_43815_n2601), .B(_abc_43815_n2598), .Y(_abc_43815_n2602) );
  AND2X2 AND2X2_1027 ( .A(_abc_43815_n1065_1_bF_buf0), .B(epc_q_31_), .Y(_abc_43815_n2603) );
  AND2X2 AND2X2_1028 ( .A(_abc_43815_n2605), .B(_abc_43815_n2606), .Y(_abc_43815_n2607) );
  AND2X2 AND2X2_1029 ( .A(_abc_43815_n2609), .B(_abc_43815_n2608), .Y(_abc_43815_n2610) );
  AND2X2 AND2X2_103 ( .A(_abc_43815_n704), .B(\mem_dat_i[21] ), .Y(_abc_43815_n786) );
  AND2X2 AND2X2_1030 ( .A(_abc_43815_n1418_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_43815_n2612) );
  AND2X2 AND2X2_1031 ( .A(_abc_43815_n1489_bF_buf4), .B(epc_q_31_), .Y(_abc_43815_n2613) );
  AND2X2 AND2X2_1032 ( .A(_abc_43815_n2615), .B(_abc_43815_n1351_bF_buf0), .Y(_abc_43815_n2616) );
  AND2X2 AND2X2_1033 ( .A(_abc_43815_n2611), .B(_abc_43815_n2616), .Y(_abc_43815_n2617) );
  AND2X2 AND2X2_1034 ( .A(_abc_43815_n2619), .B(enable_i_bF_buf0), .Y(_abc_43815_n2620) );
  AND2X2 AND2X2_1035 ( .A(_abc_43815_n2618), .B(_abc_43815_n2620), .Y(epc_q_31__FF_INPUT) );
  AND2X2 AND2X2_1036 ( .A(_abc_43815_n1278_bF_buf1), .B(next_pc_r_0_), .Y(_abc_43815_n2622) );
  AND2X2 AND2X2_1037 ( .A(_abc_43815_n1399_bF_buf1), .B(_abc_43815_n1433), .Y(_abc_43815_n2623) );
  AND2X2 AND2X2_1038 ( .A(_abc_43815_n2624), .B(enable_i_bF_buf7), .Y(pc_q_0__FF_INPUT) );
  AND2X2 AND2X2_1039 ( .A(_abc_43815_n1278_bF_buf0), .B(next_pc_r_1_), .Y(_abc_43815_n2626) );
  AND2X2 AND2X2_104 ( .A(_abc_43815_n706_1), .B(\mem_dat_i[5] ), .Y(_abc_43815_n787) );
  AND2X2 AND2X2_1040 ( .A(_abc_43815_n1399_bF_buf0), .B(_abc_43815_n1452), .Y(_abc_43815_n2627) );
  AND2X2 AND2X2_1041 ( .A(_abc_43815_n2628), .B(enable_i_bF_buf6), .Y(pc_q_1__FF_INPUT) );
  AND2X2 AND2X2_1042 ( .A(_abc_43815_n1399_bF_buf4), .B(_abc_43815_n1487), .Y(_abc_43815_n2630) );
  AND2X2 AND2X2_1043 ( .A(_abc_43815_n1278_bF_buf7), .B(pc_q_2_), .Y(_abc_43815_n2631) );
  AND2X2 AND2X2_1044 ( .A(_abc_43815_n2632), .B(enable_i_bF_buf5), .Y(pc_q_2__FF_INPUT) );
  AND2X2 AND2X2_1045 ( .A(_abc_43815_n1399_bF_buf3), .B(_abc_43815_n1528), .Y(_abc_43815_n2634) );
  AND2X2 AND2X2_1046 ( .A(_abc_43815_n1278_bF_buf6), .B(pc_q_3_), .Y(_abc_43815_n2635) );
  AND2X2 AND2X2_1047 ( .A(_abc_43815_n2636), .B(enable_i_bF_buf4), .Y(pc_q_3__FF_INPUT) );
  AND2X2 AND2X2_1048 ( .A(_abc_43815_n1399_bF_buf2), .B(_abc_43815_n1565), .Y(_abc_43815_n2638_1) );
  AND2X2 AND2X2_1049 ( .A(_abc_43815_n1278_bF_buf5), .B(pc_q_4_), .Y(_abc_43815_n2639) );
  AND2X2 AND2X2_105 ( .A(_abc_43815_n789), .B(_abc_43815_n685), .Y(_abc_43815_n790) );
  AND2X2 AND2X2_1050 ( .A(_abc_43815_n2640), .B(enable_i_bF_buf3), .Y(pc_q_4__FF_INPUT) );
  AND2X2 AND2X2_1051 ( .A(_abc_43815_n1399_bF_buf1), .B(_abc_43815_n1605), .Y(_abc_43815_n2642) );
  AND2X2 AND2X2_1052 ( .A(_abc_43815_n1278_bF_buf4), .B(pc_q_5_), .Y(_abc_43815_n2643) );
  AND2X2 AND2X2_1053 ( .A(_abc_43815_n2644), .B(enable_i_bF_buf2), .Y(pc_q_5__FF_INPUT) );
  AND2X2 AND2X2_1054 ( .A(_abc_43815_n1399_bF_buf0), .B(_abc_43815_n1637), .Y(_abc_43815_n2646) );
  AND2X2 AND2X2_1055 ( .A(_abc_43815_n1278_bF_buf3), .B(pc_q_6_), .Y(_abc_43815_n2647) );
  AND2X2 AND2X2_1056 ( .A(_abc_43815_n2648), .B(enable_i_bF_buf1), .Y(pc_q_6__FF_INPUT) );
  AND2X2 AND2X2_1057 ( .A(_abc_43815_n1278_bF_buf2), .B(pc_q_7_), .Y(_abc_43815_n2650) );
  AND2X2 AND2X2_1058 ( .A(_abc_43815_n1399_bF_buf4), .B(_abc_43815_n1682), .Y(_abc_43815_n2651) );
  AND2X2 AND2X2_1059 ( .A(_abc_43815_n2652), .B(enable_i_bF_buf0), .Y(pc_q_7__FF_INPUT) );
  AND2X2 AND2X2_106 ( .A(_abc_43815_n791), .B(state_q_1_bF_buf1), .Y(_abc_43815_n792) );
  AND2X2 AND2X2_1060 ( .A(_abc_43815_n2655), .B(_abc_43815_n1398), .Y(_abc_43815_n2656) );
  AND2X2 AND2X2_1061 ( .A(_abc_43815_n1278_bF_buf1), .B(pc_q_8_), .Y(_abc_43815_n2657) );
  AND2X2 AND2X2_1062 ( .A(_abc_43815_n2660), .B(_abc_43815_n1740), .Y(_abc_43815_n2661) );
  AND2X2 AND2X2_1063 ( .A(_abc_43815_n2661), .B(_abc_43815_n1193), .Y(_abc_43815_n2662_1) );
  AND2X2 AND2X2_1064 ( .A(_abc_43815_n2665), .B(enable_i_bF_buf7), .Y(_abc_43815_n2666) );
  AND2X2 AND2X2_1065 ( .A(_abc_43815_n2664), .B(_abc_43815_n2666), .Y(pc_q_9__FF_INPUT) );
  AND2X2 AND2X2_1066 ( .A(_abc_43815_n1802_1), .B(_abc_43815_n1349), .Y(_abc_43815_n2668) );
  AND2X2 AND2X2_1067 ( .A(_abc_43815_n2669), .B(_abc_43815_n1194), .Y(_abc_43815_n2670) );
  AND2X2 AND2X2_1068 ( .A(_abc_43815_n1278_bF_buf7), .B(pc_q_10_), .Y(_abc_43815_n2671) );
  AND2X2 AND2X2_1069 ( .A(_abc_43815_n2672), .B(enable_i_bF_buf6), .Y(pc_q_10__FF_INPUT) );
  AND2X2 AND2X2_107 ( .A(_abc_43815_n682), .B(alu_p_o_6_), .Y(_abc_43815_n794) );
  AND2X2 AND2X2_1070 ( .A(_abc_43815_n1834), .B(_abc_43815_n1352_1), .Y(_abc_43815_n2674) );
  AND2X2 AND2X2_1071 ( .A(_abc_43815_n1192), .B(_abc_43815_n2675), .Y(_abc_43815_n2676) );
  AND2X2 AND2X2_1072 ( .A(_abc_43815_n2679), .B(enable_i_bF_buf5), .Y(_abc_43815_n2680) );
  AND2X2 AND2X2_1073 ( .A(_abc_43815_n2678), .B(_abc_43815_n2680), .Y(pc_q_11__FF_INPUT) );
  AND2X2 AND2X2_1074 ( .A(_abc_43815_n1882), .B(_abc_43815_n1399_bF_buf3), .Y(_abc_43815_n2682) );
  AND2X2 AND2X2_1075 ( .A(_abc_43815_n1278_bF_buf5), .B(pc_q_12_), .Y(_abc_43815_n2683) );
  AND2X2 AND2X2_1076 ( .A(_abc_43815_n2684), .B(enable_i_bF_buf4), .Y(pc_q_12__FF_INPUT) );
  AND2X2 AND2X2_1077 ( .A(_abc_43815_n1921), .B(_abc_43815_n1399_bF_buf2), .Y(_abc_43815_n2686_1) );
  AND2X2 AND2X2_1078 ( .A(_abc_43815_n1278_bF_buf4), .B(pc_q_13_), .Y(_abc_43815_n2687) );
  AND2X2 AND2X2_1079 ( .A(_abc_43815_n2688), .B(enable_i_bF_buf3), .Y(pc_q_13__FF_INPUT) );
  AND2X2 AND2X2_108 ( .A(_abc_43815_n694), .B(\mem_dat_i[22] ), .Y(_abc_43815_n795_1) );
  AND2X2 AND2X2_1080 ( .A(_abc_43815_n1958), .B(_abc_43815_n1399_bF_buf1), .Y(_abc_43815_n2690) );
  AND2X2 AND2X2_1081 ( .A(_abc_43815_n1278_bF_buf3), .B(pc_q_14_), .Y(_abc_43815_n2691) );
  AND2X2 AND2X2_1082 ( .A(_abc_43815_n2692), .B(enable_i_bF_buf2), .Y(pc_q_14__FF_INPUT) );
  AND2X2 AND2X2_1083 ( .A(_abc_43815_n1990), .B(_abc_43815_n1399_bF_buf0), .Y(_abc_43815_n2694) );
  AND2X2 AND2X2_1084 ( .A(_abc_43815_n1278_bF_buf2), .B(pc_q_15_), .Y(_abc_43815_n2695) );
  AND2X2 AND2X2_1085 ( .A(_abc_43815_n2696), .B(enable_i_bF_buf1), .Y(pc_q_15__FF_INPUT) );
  AND2X2 AND2X2_1086 ( .A(_abc_43815_n2039), .B(_abc_43815_n1399_bF_buf4), .Y(_abc_43815_n2698) );
  AND2X2 AND2X2_1087 ( .A(_abc_43815_n1278_bF_buf1), .B(pc_q_16_), .Y(_abc_43815_n2699) );
  AND2X2 AND2X2_1088 ( .A(_abc_43815_n2700), .B(enable_i_bF_buf0), .Y(pc_q_16__FF_INPUT) );
  AND2X2 AND2X2_1089 ( .A(_abc_43815_n2078), .B(_abc_43815_n1399_bF_buf3), .Y(_abc_43815_n2702) );
  AND2X2 AND2X2_109 ( .A(_abc_43815_n697), .B(\mem_dat_i[6] ), .Y(_abc_43815_n796) );
  AND2X2 AND2X2_1090 ( .A(_abc_43815_n1278_bF_buf0), .B(pc_q_17_), .Y(_abc_43815_n2703) );
  AND2X2 AND2X2_1091 ( .A(_abc_43815_n2704), .B(enable_i_bF_buf7), .Y(pc_q_17__FF_INPUT) );
  AND2X2 AND2X2_1092 ( .A(_abc_43815_n2111), .B(_abc_43815_n1399_bF_buf2), .Y(_abc_43815_n2706) );
  AND2X2 AND2X2_1093 ( .A(_abc_43815_n1278_bF_buf7), .B(pc_q_18_), .Y(_abc_43815_n2707) );
  AND2X2 AND2X2_1094 ( .A(_abc_43815_n2708), .B(enable_i_bF_buf6), .Y(pc_q_18__FF_INPUT) );
  AND2X2 AND2X2_1095 ( .A(_abc_43815_n2147), .B(_abc_43815_n1399_bF_buf1), .Y(_abc_43815_n2710_1) );
  AND2X2 AND2X2_1096 ( .A(_abc_43815_n1278_bF_buf6), .B(pc_q_19_), .Y(_abc_43815_n2711) );
  AND2X2 AND2X2_1097 ( .A(_abc_43815_n2712), .B(enable_i_bF_buf5), .Y(pc_q_19__FF_INPUT) );
  AND2X2 AND2X2_1098 ( .A(_abc_43815_n2190), .B(_abc_43815_n1399_bF_buf0), .Y(_abc_43815_n2714) );
  AND2X2 AND2X2_1099 ( .A(_abc_43815_n1278_bF_buf5), .B(pc_q_20_), .Y(_abc_43815_n2715) );
  AND2X2 AND2X2_11 ( .A(inst_r_4_), .B(inst_r_5_), .Y(_abc_43815_n636) );
  AND2X2 AND2X2_110 ( .A(_abc_43815_n706_1), .B(\mem_dat_i[6] ), .Y(_abc_43815_n799) );
  AND2X2 AND2X2_1100 ( .A(_abc_43815_n2716), .B(enable_i_bF_buf4), .Y(pc_q_20__FF_INPUT) );
  AND2X2 AND2X2_1101 ( .A(_abc_43815_n2228), .B(_abc_43815_n1399_bF_buf4), .Y(_abc_43815_n2718) );
  AND2X2 AND2X2_1102 ( .A(_abc_43815_n1278_bF_buf4), .B(pc_q_21_), .Y(_abc_43815_n2719) );
  AND2X2 AND2X2_1103 ( .A(_abc_43815_n2720), .B(enable_i_bF_buf3), .Y(pc_q_21__FF_INPUT) );
  AND2X2 AND2X2_1104 ( .A(_abc_43815_n2264), .B(_abc_43815_n1399_bF_buf3), .Y(_abc_43815_n2722) );
  AND2X2 AND2X2_1105 ( .A(_abc_43815_n1278_bF_buf3), .B(pc_q_22_), .Y(_abc_43815_n2723) );
  AND2X2 AND2X2_1106 ( .A(_abc_43815_n2724), .B(enable_i_bF_buf2), .Y(pc_q_22__FF_INPUT) );
  AND2X2 AND2X2_1107 ( .A(_abc_43815_n2300), .B(_abc_43815_n1399_bF_buf2), .Y(_abc_43815_n2726) );
  AND2X2 AND2X2_1108 ( .A(_abc_43815_n1278_bF_buf2), .B(pc_q_23_), .Y(_abc_43815_n2727) );
  AND2X2 AND2X2_1109 ( .A(_abc_43815_n2728), .B(enable_i_bF_buf1), .Y(pc_q_23__FF_INPUT) );
  AND2X2 AND2X2_111 ( .A(_abc_43815_n696), .B(\mem_dat_i[14] ), .Y(_abc_43815_n800_1) );
  AND2X2 AND2X2_1110 ( .A(_abc_43815_n2343), .B(_abc_43815_n1399_bF_buf1), .Y(_abc_43815_n2730) );
  AND2X2 AND2X2_1111 ( .A(_abc_43815_n1278_bF_buf1), .B(pc_q_24_), .Y(_abc_43815_n2731) );
  AND2X2 AND2X2_1112 ( .A(_abc_43815_n2732), .B(enable_i_bF_buf0), .Y(pc_q_24__FF_INPUT) );
  AND2X2 AND2X2_1113 ( .A(_abc_43815_n2382), .B(_abc_43815_n1399_bF_buf0), .Y(_abc_43815_n2734_1) );
  AND2X2 AND2X2_1114 ( .A(_abc_43815_n1278_bF_buf0), .B(pc_q_25_), .Y(_abc_43815_n2735) );
  AND2X2 AND2X2_1115 ( .A(_abc_43815_n2736), .B(enable_i_bF_buf7), .Y(pc_q_25__FF_INPUT) );
  AND2X2 AND2X2_1116 ( .A(_abc_43815_n2419), .B(_abc_43815_n1399_bF_buf4), .Y(_abc_43815_n2738) );
  AND2X2 AND2X2_1117 ( .A(_abc_43815_n1278_bF_buf7), .B(pc_q_26_), .Y(_abc_43815_n2739) );
  AND2X2 AND2X2_1118 ( .A(_abc_43815_n2740), .B(enable_i_bF_buf6), .Y(pc_q_26__FF_INPUT) );
  AND2X2 AND2X2_1119 ( .A(_abc_43815_n2458), .B(_abc_43815_n1399_bF_buf3), .Y(_abc_43815_n2742) );
  AND2X2 AND2X2_112 ( .A(_abc_43815_n689), .B(\mem_dat_i[30] ), .Y(_abc_43815_n802) );
  AND2X2 AND2X2_1120 ( .A(_abc_43815_n1278_bF_buf6), .B(pc_q_27_), .Y(_abc_43815_n2743) );
  AND2X2 AND2X2_1121 ( .A(_abc_43815_n2744), .B(enable_i_bF_buf5), .Y(pc_q_27__FF_INPUT) );
  AND2X2 AND2X2_1122 ( .A(_abc_43815_n2499), .B(_abc_43815_n1399_bF_buf2), .Y(_abc_43815_n2746) );
  AND2X2 AND2X2_1123 ( .A(_abc_43815_n1278_bF_buf5), .B(pc_q_28_), .Y(_abc_43815_n2747) );
  AND2X2 AND2X2_1124 ( .A(_abc_43815_n2748), .B(enable_i_bF_buf4), .Y(pc_q_28__FF_INPUT) );
  AND2X2 AND2X2_1125 ( .A(_abc_43815_n2535), .B(_abc_43815_n1399_bF_buf1), .Y(_abc_43815_n2750) );
  AND2X2 AND2X2_1126 ( .A(_abc_43815_n1278_bF_buf4), .B(pc_q_29_), .Y(_abc_43815_n2751) );
  AND2X2 AND2X2_1127 ( .A(_abc_43815_n2752), .B(enable_i_bF_buf3), .Y(pc_q_29__FF_INPUT) );
  AND2X2 AND2X2_1128 ( .A(_abc_43815_n1278_bF_buf3), .B(pc_q_30_), .Y(_abc_43815_n2754) );
  AND2X2 AND2X2_1129 ( .A(_abc_43815_n2574), .B(_abc_43815_n1399_bF_buf0), .Y(_abc_43815_n2755) );
  AND2X2 AND2X2_113 ( .A(_abc_43815_n704), .B(\mem_dat_i[22] ), .Y(_abc_43815_n803) );
  AND2X2 AND2X2_1130 ( .A(_abc_43815_n2756), .B(enable_i_bF_buf2), .Y(pc_q_30__FF_INPUT) );
  AND2X2 AND2X2_1131 ( .A(_abc_43815_n2610), .B(_abc_43815_n1399_bF_buf4), .Y(_abc_43815_n2758_1) );
  AND2X2 AND2X2_1132 ( .A(_abc_43815_n1278_bF_buf2), .B(pc_q_31_), .Y(_abc_43815_n2759_1) );
  AND2X2 AND2X2_1133 ( .A(_abc_43815_n2760), .B(enable_i_bF_buf1), .Y(pc_q_31__FF_INPUT) );
  AND2X2 AND2X2_1134 ( .A(_abc_43815_n1156_1), .B(_abc_43815_n1131), .Y(_abc_43815_n2766) );
  AND2X2 AND2X2_1135 ( .A(_abc_43815_n1115), .B(_abc_43815_n1161), .Y(_abc_43815_n2767) );
  AND2X2 AND2X2_1136 ( .A(alu_op_r_7_), .B(alu_op_r_6_), .Y(_abc_43815_n2769) );
  AND2X2 AND2X2_1137 ( .A(_abc_43815_n1112), .B(_abc_43815_n2769), .Y(_abc_43815_n2770) );
  AND2X2 AND2X2_1138 ( .A(_abc_43815_n1106), .B(_abc_43815_n2770), .Y(_abc_43815_n2771) );
  AND2X2 AND2X2_1139 ( .A(_abc_43815_n2771), .B(_abc_43815_n2768), .Y(_abc_43815_n2772) );
  AND2X2 AND2X2_114 ( .A(_abc_43815_n806), .B(state_q_1_bF_buf0), .Y(_abc_43815_n807) );
  AND2X2 AND2X2_1140 ( .A(_abc_43815_n1179), .B(_abc_43815_n1110), .Y(_abc_43815_n2775) );
  AND2X2 AND2X2_1141 ( .A(_abc_43815_n1113), .B(_abc_43815_n1130), .Y(_abc_43815_n2781) );
  AND2X2 AND2X2_1142 ( .A(_abc_43815_n1106), .B(_abc_43815_n1161), .Y(_abc_43815_n2782) );
  AND2X2 AND2X2_1143 ( .A(_abc_43815_n2782), .B(_abc_43815_n2781), .Y(_abc_43815_n2783) );
  AND2X2 AND2X2_1144 ( .A(_abc_43815_n2781), .B(_abc_43815_n1106), .Y(_abc_43815_n2784_1) );
  AND2X2 AND2X2_1145 ( .A(_abc_43815_n2784_1), .B(_abc_43815_n1116_1), .Y(_abc_43815_n2785_1) );
  AND2X2 AND2X2_1146 ( .A(_abc_43815_n1106), .B(_abc_43815_n1119_1), .Y(_abc_43815_n2787) );
  AND2X2 AND2X2_1147 ( .A(_abc_43815_n2787), .B(_abc_43815_n1113), .Y(_abc_43815_n2788) );
  AND2X2 AND2X2_1148 ( .A(_abc_43815_n2787), .B(_abc_43815_n2789), .Y(_abc_43815_n2790) );
  AND2X2 AND2X2_1149 ( .A(_abc_43815_n2795), .B(_abc_43815_n1058), .Y(_abc_43815_n2796) );
  AND2X2 AND2X2_115 ( .A(_abc_43815_n798), .B(_abc_43815_n807), .Y(_abc_43815_n808) );
  AND2X2 AND2X2_1150 ( .A(_abc_43815_n2798), .B(opcode_q_21_), .Y(_abc_43815_n2799) );
  AND2X2 AND2X2_1151 ( .A(_abc_43815_n1172_1_bF_buf2), .B(opcode_q_22_), .Y(_abc_43815_n2801) );
  AND2X2 AND2X2_1152 ( .A(_abc_43815_n2798), .B(_abc_43815_n2801), .Y(ex_rd_q_1__FF_INPUT) );
  AND2X2 AND2X2_1153 ( .A(_abc_43815_n1172_1_bF_buf1), .B(opcode_q_23_), .Y(_abc_43815_n2803) );
  AND2X2 AND2X2_1154 ( .A(_abc_43815_n2798), .B(_abc_43815_n2803), .Y(ex_rd_q_2__FF_INPUT) );
  AND2X2 AND2X2_1155 ( .A(_abc_43815_n2798), .B(opcode_q_24_), .Y(_abc_43815_n2805) );
  AND2X2 AND2X2_1156 ( .A(_abc_43815_n1172_1_bF_buf0), .B(opcode_q_25_), .Y(_abc_43815_n2807) );
  AND2X2 AND2X2_1157 ( .A(_abc_43815_n2798), .B(_abc_43815_n2807), .Y(ex_rd_q_4__FF_INPUT) );
  AND2X2 AND2X2_1158 ( .A(_abc_43815_n2813), .B(alu_op_r_0_), .Y(_abc_43815_n2814) );
  AND2X2 AND2X2_1159 ( .A(_abc_43815_n2784_1), .B(_abc_43815_n1131), .Y(_abc_43815_n2815) );
  AND2X2 AND2X2_116 ( .A(_abc_43815_n689), .B(\mem_dat_i[31] ), .Y(_abc_43815_n810) );
  AND2X2 AND2X2_1160 ( .A(_abc_43815_n2818), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_43815_n2819) );
  AND2X2 AND2X2_1161 ( .A(_abc_43815_n2813), .B(alu_op_r_1_), .Y(_abc_43815_n2821) );
  AND2X2 AND2X2_1162 ( .A(_abc_43815_n2818), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_43815_n2822) );
  AND2X2 AND2X2_1163 ( .A(_abc_43815_n2813), .B(alu_op_r_2_), .Y(_abc_43815_n2824) );
  AND2X2 AND2X2_1164 ( .A(_abc_43815_n2818), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n2825) );
  AND2X2 AND2X2_1165 ( .A(_abc_43815_n2813), .B(alu_op_r_3_), .Y(_abc_43815_n2827) );
  AND2X2 AND2X2_1166 ( .A(_abc_43815_n2818), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_43815_n2828) );
  AND2X2 AND2X2_1167 ( .A(_abc_43815_n2813), .B(int32_r_4_), .Y(_abc_43815_n2830) );
  AND2X2 AND2X2_1168 ( .A(_abc_43815_n2818), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_43815_n2831) );
  AND2X2 AND2X2_1169 ( .A(_abc_43815_n2813), .B(int32_r_5_), .Y(_abc_43815_n2833) );
  AND2X2 AND2X2_117 ( .A(_abc_43815_n696), .B(\mem_dat_i[15] ), .Y(_abc_43815_n811) );
  AND2X2 AND2X2_1170 ( .A(_abc_43815_n2818), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_43815_n2834) );
  AND2X2 AND2X2_1171 ( .A(_abc_43815_n986_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_43815_n2836_1) );
  AND2X2 AND2X2_1172 ( .A(_abc_43815_n2812), .B(alu_op_r_4_), .Y(_abc_43815_n2837_1) );
  AND2X2 AND2X2_1173 ( .A(_abc_43815_n2840_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_43815_n2841) );
  AND2X2 AND2X2_1174 ( .A(_abc_43815_n986_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_43815_n2843) );
  AND2X2 AND2X2_1175 ( .A(_abc_43815_n2812), .B(alu_op_r_5_), .Y(_abc_43815_n2844) );
  AND2X2 AND2X2_1176 ( .A(_abc_43815_n2840_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_43815_n2846) );
  AND2X2 AND2X2_1177 ( .A(_abc_43815_n986_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_43815_n2848) );
  AND2X2 AND2X2_1178 ( .A(_abc_43815_n2812), .B(alu_op_r_6_), .Y(_abc_43815_n2849) );
  AND2X2 AND2X2_1179 ( .A(_abc_43815_n2840_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_43815_n2851) );
  AND2X2 AND2X2_118 ( .A(_abc_43815_n704), .B(\mem_dat_i[23] ), .Y(_abc_43815_n813) );
  AND2X2 AND2X2_1180 ( .A(_abc_43815_n986_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n2853) );
  AND2X2 AND2X2_1181 ( .A(_abc_43815_n2812), .B(alu_op_r_7_), .Y(_abc_43815_n2854) );
  AND2X2 AND2X2_1182 ( .A(_abc_43815_n2840_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n2856) );
  AND2X2 AND2X2_1183 ( .A(_abc_43815_n986_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_43815_n2858) );
  AND2X2 AND2X2_1184 ( .A(_abc_43815_n2812), .B(int32_r_10_), .Y(_abc_43815_n2859) );
  AND2X2 AND2X2_1185 ( .A(_abc_43815_n2840_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_43815_n2861) );
  AND2X2 AND2X2_1186 ( .A(_abc_43815_n986_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_43815_n2863_1) );
  AND2X2 AND2X2_1187 ( .A(_abc_43815_n2812), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_43815_n2864) );
  AND2X2 AND2X2_1188 ( .A(_abc_43815_n2840_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_43815_n2866) );
  AND2X2 AND2X2_1189 ( .A(_abc_43815_n986_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_43815_n2868) );
  AND2X2 AND2X2_119 ( .A(_abc_43815_n706_1), .B(\mem_dat_i[7] ), .Y(_abc_43815_n814) );
  AND2X2 AND2X2_1190 ( .A(_abc_43815_n2812), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_43815_n2869) );
  AND2X2 AND2X2_1191 ( .A(_abc_43815_n2840_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_43815_n2871) );
  AND2X2 AND2X2_1192 ( .A(_abc_43815_n986_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_43815_n2873) );
  AND2X2 AND2X2_1193 ( .A(_abc_43815_n2812), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_43815_n2874) );
  AND2X2 AND2X2_1194 ( .A(_abc_43815_n2840_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_43815_n2876) );
  AND2X2 AND2X2_1195 ( .A(_abc_43815_n986_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_43815_n2878) );
  AND2X2 AND2X2_1196 ( .A(_abc_43815_n2812), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_43815_n2879) );
  AND2X2 AND2X2_1197 ( .A(_abc_43815_n2840_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_43815_n2881) );
  AND2X2 AND2X2_1198 ( .A(_abc_43815_n986_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_43815_n2883) );
  AND2X2 AND2X2_1199 ( .A(_abc_43815_n2812), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1), .Y(_abc_43815_n2884) );
  AND2X2 AND2X2_12 ( .A(_abc_43815_n637), .B(inst_r_2_), .Y(_abc_43815_n638) );
  AND2X2 AND2X2_120 ( .A(_abc_43815_n697), .B(\mem_dat_i[7] ), .Y(_abc_43815_n818) );
  AND2X2 AND2X2_1200 ( .A(_abc_43815_n2840_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_43815_n2886) );
  AND2X2 AND2X2_1201 ( .A(_abc_43815_n1054), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0), .Y(_abc_43815_n2888_1) );
  AND2X2 AND2X2_1202 ( .A(_abc_43815_n986_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_43815_n2889_1) );
  AND2X2 AND2X2_1203 ( .A(_abc_43815_n1050), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3), .Y(_abc_43815_n2890) );
  AND2X2 AND2X2_1204 ( .A(_abc_43815_n2892), .B(_abc_43815_n2894), .Y(_abc_43815_n2895) );
  AND2X2 AND2X2_1205 ( .A(_abc_43815_n2840_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_43815_n2897) );
  AND2X2 AND2X2_1206 ( .A(_abc_43815_n986_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_43815_n2899) );
  AND2X2 AND2X2_1207 ( .A(_abc_43815_n2900), .B(_abc_43815_n2894), .Y(_abc_43815_n2901) );
  AND2X2 AND2X2_1208 ( .A(_abc_43815_n2840_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_43815_n2903) );
  AND2X2 AND2X2_1209 ( .A(_abc_43815_n986_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_43815_n2905) );
  AND2X2 AND2X2_121 ( .A(_abc_43815_n694), .B(\mem_dat_i[23] ), .Y(_abc_43815_n819) );
  AND2X2 AND2X2_1210 ( .A(_abc_43815_n2906), .B(_abc_43815_n2894), .Y(_abc_43815_n2907) );
  AND2X2 AND2X2_1211 ( .A(_abc_43815_n2840_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_43815_n2909) );
  AND2X2 AND2X2_1212 ( .A(_abc_43815_n986_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_43815_n2911) );
  AND2X2 AND2X2_1213 ( .A(_abc_43815_n2912), .B(_abc_43815_n2894), .Y(_abc_43815_n2913) );
  AND2X2 AND2X2_1214 ( .A(_abc_43815_n2840_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_43815_n2915_1) );
  AND2X2 AND2X2_1215 ( .A(_abc_43815_n986_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_43815_n2917) );
  AND2X2 AND2X2_1216 ( .A(_abc_43815_n2918), .B(_abc_43815_n2894), .Y(_abc_43815_n2919) );
  AND2X2 AND2X2_1217 ( .A(_abc_43815_n2840_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_43815_n2921) );
  AND2X2 AND2X2_1218 ( .A(_abc_43815_n986_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_43815_n2923) );
  AND2X2 AND2X2_1219 ( .A(_abc_43815_n2924), .B(_abc_43815_n2894), .Y(_abc_43815_n2925) );
  AND2X2 AND2X2_122 ( .A(_abc_43815_n821), .B(_abc_43815_n817_1), .Y(_abc_43815_n822) );
  AND2X2 AND2X2_1220 ( .A(_abc_43815_n2840_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_43815_n2927) );
  AND2X2 AND2X2_1221 ( .A(_abc_43815_n986_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_43815_n2929) );
  AND2X2 AND2X2_1222 ( .A(_abc_43815_n2930), .B(_abc_43815_n2894), .Y(_abc_43815_n2931) );
  AND2X2 AND2X2_1223 ( .A(_abc_43815_n2840_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_43815_n2933) );
  AND2X2 AND2X2_1224 ( .A(_abc_43815_n986_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_43815_n2935) );
  AND2X2 AND2X2_1225 ( .A(_abc_43815_n2936), .B(_abc_43815_n2894), .Y(_abc_43815_n2937) );
  AND2X2 AND2X2_1226 ( .A(_abc_43815_n2840_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_43815_n2939) );
  AND2X2 AND2X2_1227 ( .A(_abc_43815_n986_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_43815_n2941_1) );
  AND2X2 AND2X2_1228 ( .A(_abc_43815_n2942), .B(_abc_43815_n2894), .Y(_abc_43815_n2943) );
  AND2X2 AND2X2_1229 ( .A(_abc_43815_n2840_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_43815_n2945) );
  AND2X2 AND2X2_123 ( .A(_abc_43815_n823), .B(_abc_43815_n824), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_) );
  AND2X2 AND2X2_1230 ( .A(_abc_43815_n986_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_43815_n2947) );
  AND2X2 AND2X2_1231 ( .A(_abc_43815_n2948), .B(_abc_43815_n2894), .Y(_abc_43815_n2949) );
  AND2X2 AND2X2_1232 ( .A(_abc_43815_n2840_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_43815_n2951) );
  AND2X2 AND2X2_1233 ( .A(_abc_43815_n986_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_43815_n2953) );
  AND2X2 AND2X2_1234 ( .A(_abc_43815_n2954), .B(_abc_43815_n2894), .Y(_abc_43815_n2955) );
  AND2X2 AND2X2_1235 ( .A(_abc_43815_n2840_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_43815_n2957) );
  AND2X2 AND2X2_1236 ( .A(_abc_43815_n986_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_43815_n2959) );
  AND2X2 AND2X2_1237 ( .A(_abc_43815_n2960), .B(_abc_43815_n2894), .Y(_abc_43815_n2961) );
  AND2X2 AND2X2_1238 ( .A(_abc_43815_n2840_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_43815_n2963) );
  AND2X2 AND2X2_1239 ( .A(_abc_43815_n986_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_43815_n2965) );
  AND2X2 AND2X2_124 ( .A(_abc_43815_n828), .B(_abc_43815_n686_1_bF_buf1), .Y(_abc_43815_n829_1) );
  AND2X2 AND2X2_1240 ( .A(_abc_43815_n2966_1), .B(_abc_43815_n2894), .Y(_abc_43815_n2967_1) );
  AND2X2 AND2X2_1241 ( .A(_abc_43815_n2840_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_43815_n2969) );
  AND2X2 AND2X2_1242 ( .A(_abc_43815_n986_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_43815_n2971) );
  AND2X2 AND2X2_1243 ( .A(_abc_43815_n2972), .B(_abc_43815_n2894), .Y(_abc_43815_n2973) );
  AND2X2 AND2X2_1244 ( .A(_abc_43815_n2840_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_43815_n2975) );
  AND2X2 AND2X2_1245 ( .A(_abc_43815_n986_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_43815_n2977) );
  AND2X2 AND2X2_1246 ( .A(_abc_43815_n2978), .B(_abc_43815_n2894), .Y(_abc_43815_n2979) );
  AND2X2 AND2X2_1247 ( .A(_abc_43815_n2840_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_43815_n2981) );
  AND2X2 AND2X2_1248 ( .A(_abc_43815_n986_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_43815_n2983) );
  AND2X2 AND2X2_1249 ( .A(_abc_43815_n2984), .B(_abc_43815_n2894), .Y(_abc_43815_n2985) );
  AND2X2 AND2X2_125 ( .A(_abc_43815_n829_1), .B(_abc_43815_n827), .Y(_abc_43815_n830) );
  AND2X2 AND2X2_1250 ( .A(_abc_43815_n2840_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_43815_n2987) );
  AND2X2 AND2X2_1251 ( .A(_abc_43815_n2991_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_0_), .Y(_abc_43815_n2992_1) );
  AND2X2 AND2X2_1252 ( .A(_abc_43815_n1417), .B(_abc_43815_n1058), .Y(_abc_43815_n2993_1) );
  AND2X2 AND2X2_1253 ( .A(_abc_43815_n2993_1_bF_buf4), .B(epc_q_0_), .Y(_abc_43815_n2994) );
  AND2X2 AND2X2_1254 ( .A(_abc_43815_n2997), .B(_abc_43815_n1057), .Y(_abc_43815_n2998) );
  AND2X2 AND2X2_1255 ( .A(_abc_43815_n2996), .B(_abc_43815_n2998), .Y(_abc_43815_n2999) );
  AND2X2 AND2X2_1256 ( .A(_abc_43815_n3002_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_0_), .Y(_abc_43815_n3003) );
  AND2X2 AND2X2_1257 ( .A(_abc_43815_n2993_1_bF_buf3), .B(epc_q_1_), .Y(_abc_43815_n3005) );
  AND2X2 AND2X2_1258 ( .A(_abc_43815_n2991_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_1_), .Y(_abc_43815_n3006) );
  AND2X2 AND2X2_1259 ( .A(_abc_43815_n3009), .B(_abc_43815_n1057), .Y(_abc_43815_n3010) );
  AND2X2 AND2X2_126 ( .A(_abc_43815_n816_1), .B(_abc_43815_n684), .Y(_abc_43815_n831) );
  AND2X2 AND2X2_1260 ( .A(_abc_43815_n3008), .B(_abc_43815_n3010), .Y(_abc_43815_n3011) );
  AND2X2 AND2X2_1261 ( .A(_abc_43815_n3002_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_1_), .Y(_abc_43815_n3012) );
  AND2X2 AND2X2_1262 ( .A(_abc_43815_n2991_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_2_), .Y(_abc_43815_n3014) );
  AND2X2 AND2X2_1263 ( .A(_abc_43815_n1272), .B(_abc_43815_n1264), .Y(_abc_43815_n3016) );
  AND2X2 AND2X2_1264 ( .A(_abc_43815_n1417), .B(epc_q_2_), .Y(_abc_43815_n3017) );
  AND2X2 AND2X2_1265 ( .A(_abc_43815_n1239), .B(esr_q_2_), .Y(_abc_43815_n3018_1) );
  AND2X2 AND2X2_1266 ( .A(_abc_43815_n3020), .B(_abc_43815_n2796), .Y(_abc_43815_n3021) );
  AND2X2 AND2X2_1267 ( .A(_abc_43815_n3022), .B(_abc_43815_n3023), .Y(_abc_43815_n3024) );
  AND2X2 AND2X2_1268 ( .A(_abc_43815_n3002_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_2_), .Y(_abc_43815_n3025) );
  AND2X2 AND2X2_1269 ( .A(_abc_43815_n2993_1_bF_buf2), .B(epc_q_3_), .Y(_abc_43815_n3027) );
  AND2X2 AND2X2_127 ( .A(_abc_43815_n833), .B(_abc_43815_n826), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_) );
  AND2X2 AND2X2_1270 ( .A(_abc_43815_n2991_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_3_), .Y(_abc_43815_n3028) );
  AND2X2 AND2X2_1271 ( .A(_abc_43815_n3031), .B(_abc_43815_n1057), .Y(_abc_43815_n3032) );
  AND2X2 AND2X2_1272 ( .A(_abc_43815_n3030), .B(_abc_43815_n3032), .Y(_abc_43815_n3033) );
  AND2X2 AND2X2_1273 ( .A(_abc_43815_n3002_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_3_), .Y(_abc_43815_n3034) );
  AND2X2 AND2X2_1274 ( .A(_abc_43815_n2993_1_bF_buf1), .B(epc_q_4_), .Y(_abc_43815_n3036) );
  AND2X2 AND2X2_1275 ( .A(_abc_43815_n2991_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_4_), .Y(_abc_43815_n3037) );
  AND2X2 AND2X2_1276 ( .A(_abc_43815_n3040), .B(_abc_43815_n1057), .Y(_abc_43815_n3041) );
  AND2X2 AND2X2_1277 ( .A(_abc_43815_n3039), .B(_abc_43815_n3041), .Y(_abc_43815_n3042) );
  AND2X2 AND2X2_1278 ( .A(_abc_43815_n3002_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_4_), .Y(_abc_43815_n3043) );
  AND2X2 AND2X2_1279 ( .A(_abc_43815_n2993_1_bF_buf0), .B(epc_q_5_), .Y(_abc_43815_n3045_1) );
  AND2X2 AND2X2_128 ( .A(_abc_43815_n697), .B(\mem_dat_i[9] ), .Y(_abc_43815_n835) );
  AND2X2 AND2X2_1280 ( .A(_abc_43815_n2991_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_5_), .Y(_abc_43815_n3046) );
  AND2X2 AND2X2_1281 ( .A(_abc_43815_n3049), .B(_abc_43815_n1057), .Y(_abc_43815_n3050) );
  AND2X2 AND2X2_1282 ( .A(_abc_43815_n3048), .B(_abc_43815_n3050), .Y(_abc_43815_n3051) );
  AND2X2 AND2X2_1283 ( .A(_abc_43815_n3002_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_5_), .Y(_abc_43815_n3052) );
  AND2X2 AND2X2_1284 ( .A(_abc_43815_n2993_1_bF_buf4), .B(epc_q_6_), .Y(_abc_43815_n3054) );
  AND2X2 AND2X2_1285 ( .A(_abc_43815_n2991_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_6_), .Y(_abc_43815_n3055) );
  AND2X2 AND2X2_1286 ( .A(_abc_43815_n3058), .B(_abc_43815_n1057), .Y(_abc_43815_n3059) );
  AND2X2 AND2X2_1287 ( .A(_abc_43815_n3057), .B(_abc_43815_n3059), .Y(_abc_43815_n3060) );
  AND2X2 AND2X2_1288 ( .A(_abc_43815_n3002_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_6_), .Y(_abc_43815_n3061) );
  AND2X2 AND2X2_1289 ( .A(_abc_43815_n2993_1_bF_buf3), .B(epc_q_7_), .Y(_abc_43815_n3063) );
  AND2X2 AND2X2_129 ( .A(_abc_43815_n693), .B(_abc_43815_n722), .Y(_abc_43815_n836) );
  AND2X2 AND2X2_1290 ( .A(_abc_43815_n2991_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_7_), .Y(_abc_43815_n3064) );
  AND2X2 AND2X2_1291 ( .A(_abc_43815_n3067), .B(_abc_43815_n1057), .Y(_abc_43815_n3068) );
  AND2X2 AND2X2_1292 ( .A(_abc_43815_n3066), .B(_abc_43815_n3068), .Y(_abc_43815_n3069) );
  AND2X2 AND2X2_1293 ( .A(_abc_43815_n3002_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_7_), .Y(_abc_43815_n3070_1) );
  AND2X2 AND2X2_1294 ( .A(_abc_43815_n2991_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_8_), .Y(_abc_43815_n3072) );
  AND2X2 AND2X2_1295 ( .A(_abc_43815_n2993_1_bF_buf2), .B(epc_q_8_), .Y(_abc_43815_n3073) );
  AND2X2 AND2X2_1296 ( .A(_abc_43815_n1696), .B(_abc_43815_n1171_bF_buf5), .Y(_abc_43815_n3075) );
  AND2X2 AND2X2_1297 ( .A(_abc_43815_n3002_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_8_), .Y(_abc_43815_n3077) );
  AND2X2 AND2X2_1298 ( .A(_abc_43815_n2991_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_9_), .Y(_abc_43815_n3079) );
  AND2X2 AND2X2_1299 ( .A(_abc_43815_n1347), .B(_abc_43815_n1264), .Y(_abc_43815_n3081) );
  AND2X2 AND2X2_13 ( .A(_abc_43815_n630), .B(inst_r_1_), .Y(_abc_43815_n639) );
  AND2X2 AND2X2_130 ( .A(_abc_43815_n837), .B(_abc_43815_n686_1_bF_buf0), .Y(_abc_43815_n838) );
  AND2X2 AND2X2_1300 ( .A(_abc_43815_n1417), .B(epc_q_9_), .Y(_abc_43815_n3082) );
  AND2X2 AND2X2_1301 ( .A(_abc_43815_n1239), .B(esr_q_9_), .Y(_abc_43815_n3083) );
  AND2X2 AND2X2_1302 ( .A(_abc_43815_n3085), .B(_abc_43815_n2796), .Y(_abc_43815_n3086) );
  AND2X2 AND2X2_1303 ( .A(_abc_43815_n3087), .B(_abc_43815_n3088), .Y(_abc_43815_n3089) );
  AND2X2 AND2X2_1304 ( .A(_abc_43815_n3002_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_9_), .Y(_abc_43815_n3090) );
  AND2X2 AND2X2_1305 ( .A(_abc_43815_n2991_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_10_), .Y(_abc_43815_n3092) );
  AND2X2 AND2X2_1306 ( .A(_abc_43815_n1386), .B(_abc_43815_n1379), .Y(_abc_43815_n3094) );
  AND2X2 AND2X2_1307 ( .A(_abc_43815_n1417), .B(epc_q_10_), .Y(_abc_43815_n3095) );
  AND2X2 AND2X2_1308 ( .A(_abc_43815_n1239), .B(esr_q_10_), .Y(_abc_43815_n3096_1) );
  AND2X2 AND2X2_1309 ( .A(_abc_43815_n3098), .B(_abc_43815_n2796), .Y(_abc_43815_n3099) );
  AND2X2 AND2X2_131 ( .A(_abc_43815_n839), .B(_abc_43815_n840), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_) );
  AND2X2 AND2X2_1310 ( .A(_abc_43815_n3100), .B(_abc_43815_n3101), .Y(_abc_43815_n3102) );
  AND2X2 AND2X2_1311 ( .A(_abc_43815_n3002_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_10_), .Y(_abc_43815_n3103) );
  AND2X2 AND2X2_1312 ( .A(_abc_43815_n2991_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_43815_n3105) );
  AND2X2 AND2X2_1313 ( .A(_abc_43815_n2993_1_bF_buf1), .B(epc_q_11_), .Y(_abc_43815_n3106) );
  AND2X2 AND2X2_1314 ( .A(_abc_43815_n1813), .B(_abc_43815_n1171_bF_buf2), .Y(_abc_43815_n3108) );
  AND2X2 AND2X2_1315 ( .A(_abc_43815_n3002_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_43815_n3110) );
  AND2X2 AND2X2_1316 ( .A(_abc_43815_n2991_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_43815_n3112) );
  AND2X2 AND2X2_1317 ( .A(_abc_43815_n2993_1_bF_buf0), .B(epc_q_12_), .Y(_abc_43815_n3113) );
  AND2X2 AND2X2_1318 ( .A(_abc_43815_n1849), .B(_abc_43815_n1171_bF_buf1), .Y(_abc_43815_n3115) );
  AND2X2 AND2X2_1319 ( .A(_abc_43815_n3002_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_43815_n3117) );
  AND2X2 AND2X2_132 ( .A(_abc_43815_n844), .B(_abc_43815_n686_1_bF_buf4), .Y(_abc_43815_n845) );
  AND2X2 AND2X2_1320 ( .A(_abc_43815_n2991_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_43815_n3119) );
  AND2X2 AND2X2_1321 ( .A(_abc_43815_n2993_1_bF_buf4), .B(epc_q_13_), .Y(_abc_43815_n3120) );
  AND2X2 AND2X2_1322 ( .A(_abc_43815_n1893), .B(_abc_43815_n1171_bF_buf0), .Y(_abc_43815_n3122_1) );
  AND2X2 AND2X2_1323 ( .A(_abc_43815_n3002_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_43815_n3124) );
  AND2X2 AND2X2_1324 ( .A(_abc_43815_n2991_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_43815_n3126) );
  AND2X2 AND2X2_1325 ( .A(_abc_43815_n2993_1_bF_buf3), .B(epc_q_14_), .Y(_abc_43815_n3127) );
  AND2X2 AND2X2_1326 ( .A(_abc_43815_n1932), .B(_abc_43815_n1171_bF_buf5), .Y(_abc_43815_n3129) );
  AND2X2 AND2X2_1327 ( .A(_abc_43815_n3002_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_43815_n3131) );
  AND2X2 AND2X2_1328 ( .A(_abc_43815_n2993_1_bF_buf2), .B(epc_q_15_), .Y(_abc_43815_n3134) );
  AND2X2 AND2X2_1329 ( .A(_abc_43815_n2991_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_43815_n3135) );
  AND2X2 AND2X2_133 ( .A(_abc_43815_n845), .B(_abc_43815_n843), .Y(_abc_43815_n846) );
  AND2X2 AND2X2_1330 ( .A(_abc_43815_n3133), .B(_abc_43815_n3137), .Y(_abc_43815_n3138) );
  AND2X2 AND2X2_1331 ( .A(_abc_43815_n3002_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_43815_n3139) );
  AND2X2 AND2X2_1332 ( .A(_abc_43815_n2993_1_bF_buf1), .B(epc_q_16_), .Y(_abc_43815_n3142) );
  AND2X2 AND2X2_1333 ( .A(_abc_43815_n2991_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_43815_n3143) );
  AND2X2 AND2X2_1334 ( .A(_abc_43815_n1060_bF_buf1), .B(alu_op_r_0_), .Y(_abc_43815_n3144) );
  AND2X2 AND2X2_1335 ( .A(_abc_43815_n3141), .B(_abc_43815_n3147), .Y(_abc_43815_n3148_1) );
  AND2X2 AND2X2_1336 ( .A(_abc_43815_n3002_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_43815_n3149_1) );
  AND2X2 AND2X2_1337 ( .A(_abc_43815_n2991_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_43815_n3152) );
  AND2X2 AND2X2_1338 ( .A(_abc_43815_n2993_1_bF_buf0), .B(epc_q_17_), .Y(_abc_43815_n3153) );
  AND2X2 AND2X2_1339 ( .A(_abc_43815_n1060_bF_buf0), .B(alu_op_r_1_), .Y(_abc_43815_n3154) );
  AND2X2 AND2X2_134 ( .A(_abc_43815_n847), .B(_abc_43815_n842), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_) );
  AND2X2 AND2X2_1340 ( .A(_abc_43815_n3151), .B(_abc_43815_n3157), .Y(_abc_43815_n3158) );
  AND2X2 AND2X2_1341 ( .A(_abc_43815_n3002_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_43815_n3159) );
  AND2X2 AND2X2_1342 ( .A(_abc_43815_n2991_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_43815_n3161) );
  AND2X2 AND2X2_1343 ( .A(_abc_43815_n1060_bF_buf3), .B(alu_op_r_2_), .Y(_abc_43815_n3162) );
  AND2X2 AND2X2_1344 ( .A(_abc_43815_n2993_1_bF_buf4), .B(epc_q_18_), .Y(_abc_43815_n3164) );
  AND2X2 AND2X2_1345 ( .A(_abc_43815_n2089), .B(_abc_43815_n1171_bF_buf1), .Y(_abc_43815_n3166) );
  AND2X2 AND2X2_1346 ( .A(_abc_43815_n3002_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_43815_n3168) );
  AND2X2 AND2X2_1347 ( .A(_abc_43815_n2991_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_43815_n3170) );
  AND2X2 AND2X2_1348 ( .A(_abc_43815_n1060_bF_buf2), .B(alu_op_r_3_), .Y(_abc_43815_n3171) );
  AND2X2 AND2X2_1349 ( .A(_abc_43815_n2993_1_bF_buf3), .B(epc_q_19_), .Y(_abc_43815_n3172) );
  AND2X2 AND2X2_135 ( .A(_abc_43815_n851), .B(_abc_43815_n686_1_bF_buf3), .Y(_abc_43815_n852) );
  AND2X2 AND2X2_1350 ( .A(_abc_43815_n2126), .B(_abc_43815_n1171_bF_buf0), .Y(_abc_43815_n3175) );
  AND2X2 AND2X2_1351 ( .A(_abc_43815_n3002_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_43815_n3177) );
  AND2X2 AND2X2_1352 ( .A(_abc_43815_n2991_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_43815_n3180) );
  AND2X2 AND2X2_1353 ( .A(_abc_43815_n2993_1_bF_buf2), .B(epc_q_20_), .Y(_abc_43815_n3181) );
  AND2X2 AND2X2_1354 ( .A(_abc_43815_n1060_bF_buf1), .B(int32_r_4_), .Y(_abc_43815_n3182) );
  AND2X2 AND2X2_1355 ( .A(_abc_43815_n3179), .B(_abc_43815_n3185), .Y(_abc_43815_n3186) );
  AND2X2 AND2X2_1356 ( .A(_abc_43815_n3002_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_43815_n3187) );
  AND2X2 AND2X2_1357 ( .A(_abc_43815_n2991_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_43815_n3190) );
  AND2X2 AND2X2_1358 ( .A(_abc_43815_n2993_1_bF_buf1), .B(epc_q_21_), .Y(_abc_43815_n3191) );
  AND2X2 AND2X2_1359 ( .A(_abc_43815_n1060_bF_buf0), .B(int32_r_5_), .Y(_abc_43815_n3192) );
  AND2X2 AND2X2_136 ( .A(_abc_43815_n852), .B(_abc_43815_n850), .Y(_abc_43815_n853) );
  AND2X2 AND2X2_1360 ( .A(_abc_43815_n3189), .B(_abc_43815_n3195), .Y(_abc_43815_n3196) );
  AND2X2 AND2X2_1361 ( .A(_abc_43815_n3002_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_43815_n3197) );
  AND2X2 AND2X2_1362 ( .A(_abc_43815_n2993_1_bF_buf0), .B(epc_q_22_), .Y(_abc_43815_n3200) );
  AND2X2 AND2X2_1363 ( .A(_abc_43815_n2991_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_43815_n3201) );
  AND2X2 AND2X2_1364 ( .A(_abc_43815_n1060_bF_buf3), .B(alu_op_r_4_), .Y(_abc_43815_n3202) );
  AND2X2 AND2X2_1365 ( .A(_abc_43815_n3199), .B(_abc_43815_n3205), .Y(_abc_43815_n3206) );
  AND2X2 AND2X2_1366 ( .A(_abc_43815_n3002_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_43815_n3207) );
  AND2X2 AND2X2_1367 ( .A(_abc_43815_n2993_1_bF_buf4), .B(epc_q_23_), .Y(_abc_43815_n3210) );
  AND2X2 AND2X2_1368 ( .A(_abc_43815_n2991_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_43815_n3211) );
  AND2X2 AND2X2_1369 ( .A(_abc_43815_n1060_bF_buf2), .B(alu_op_r_5_), .Y(_abc_43815_n3212) );
  AND2X2 AND2X2_137 ( .A(_abc_43815_n854), .B(_abc_43815_n849_1), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_) );
  AND2X2 AND2X2_1370 ( .A(_abc_43815_n3209_1), .B(_abc_43815_n3215), .Y(_abc_43815_n3216) );
  AND2X2 AND2X2_1371 ( .A(_abc_43815_n3002_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_43815_n3217_1) );
  AND2X2 AND2X2_1372 ( .A(_abc_43815_n2993_1_bF_buf3), .B(epc_q_24_), .Y(_abc_43815_n3220) );
  AND2X2 AND2X2_1373 ( .A(_abc_43815_n2991_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_43815_n3221) );
  AND2X2 AND2X2_1374 ( .A(_abc_43815_n1060_bF_buf1), .B(alu_op_r_6_), .Y(_abc_43815_n3222) );
  AND2X2 AND2X2_1375 ( .A(_abc_43815_n3219), .B(_abc_43815_n3225), .Y(_abc_43815_n3226) );
  AND2X2 AND2X2_1376 ( .A(_abc_43815_n3002_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_43815_n3227) );
  AND2X2 AND2X2_1377 ( .A(_abc_43815_n2991_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_43815_n3230) );
  AND2X2 AND2X2_1378 ( .A(_abc_43815_n2993_1_bF_buf2), .B(epc_q_25_), .Y(_abc_43815_n3231) );
  AND2X2 AND2X2_1379 ( .A(_abc_43815_n1060_bF_buf0), .B(alu_op_r_7_), .Y(_abc_43815_n3232) );
  AND2X2 AND2X2_138 ( .A(_abc_43815_n858), .B(_abc_43815_n686_1_bF_buf2), .Y(_abc_43815_n859) );
  AND2X2 AND2X2_1380 ( .A(_abc_43815_n3229), .B(_abc_43815_n3235_1), .Y(_abc_43815_n3236) );
  AND2X2 AND2X2_1381 ( .A(_abc_43815_n3002_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_43815_n3237) );
  AND2X2 AND2X2_1382 ( .A(_abc_43815_n2991_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_43815_n3240) );
  AND2X2 AND2X2_1383 ( .A(_abc_43815_n2993_1_bF_buf1), .B(epc_q_26_), .Y(_abc_43815_n3241) );
  AND2X2 AND2X2_1384 ( .A(_abc_43815_n1060_bF_buf3), .B(int32_r_10_), .Y(_abc_43815_n3242) );
  AND2X2 AND2X2_1385 ( .A(_abc_43815_n3239), .B(_abc_43815_n3245), .Y(_abc_43815_n3246_1) );
  AND2X2 AND2X2_1386 ( .A(_abc_43815_n3002_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_43815_n3247) );
  AND2X2 AND2X2_1387 ( .A(_abc_43815_n2991_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_43815_n3250_1) );
  AND2X2 AND2X2_1388 ( .A(_abc_43815_n2993_1_bF_buf0), .B(epc_q_27_), .Y(_abc_43815_n3251) );
  AND2X2 AND2X2_1389 ( .A(_abc_43815_n1060_bF_buf2), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_43815_n3252_1) );
  AND2X2 AND2X2_139 ( .A(_abc_43815_n859), .B(_abc_43815_n857), .Y(_abc_43815_n860) );
  AND2X2 AND2X2_1390 ( .A(_abc_43815_n3249), .B(_abc_43815_n3255), .Y(_abc_43815_n3256_1) );
  AND2X2 AND2X2_1391 ( .A(_abc_43815_n3002_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_43815_n3257) );
  AND2X2 AND2X2_1392 ( .A(_abc_43815_n2993_1_bF_buf4), .B(epc_q_28_), .Y(_abc_43815_n3260_1) );
  AND2X2 AND2X2_1393 ( .A(_abc_43815_n2991_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_43815_n3261) );
  AND2X2 AND2X2_1394 ( .A(_abc_43815_n1060_bF_buf1), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_43815_n3262_1) );
  AND2X2 AND2X2_1395 ( .A(_abc_43815_n3259), .B(_abc_43815_n3265), .Y(_abc_43815_n3266_1) );
  AND2X2 AND2X2_1396 ( .A(_abc_43815_n3002_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_43815_n3267) );
  AND2X2 AND2X2_1397 ( .A(_abc_43815_n2993_1_bF_buf3), .B(epc_q_29_), .Y(_abc_43815_n3270_1) );
  AND2X2 AND2X2_1398 ( .A(_abc_43815_n2991_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_43815_n3271) );
  AND2X2 AND2X2_1399 ( .A(_abc_43815_n1060_bF_buf0), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_43815_n3272_1) );
  AND2X2 AND2X2_14 ( .A(_abc_43815_n638), .B(_abc_43815_n639), .Y(_abc_43815_n640) );
  AND2X2 AND2X2_140 ( .A(_abc_43815_n861), .B(_abc_43815_n856), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_) );
  AND2X2 AND2X2_1400 ( .A(_abc_43815_n3269), .B(_abc_43815_n3275), .Y(_abc_43815_n3276_1) );
  AND2X2 AND2X2_1401 ( .A(_abc_43815_n3002_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_43815_n3277) );
  AND2X2 AND2X2_1402 ( .A(_abc_43815_n2991_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_43815_n3280_1) );
  AND2X2 AND2X2_1403 ( .A(_abc_43815_n2993_1_bF_buf2), .B(epc_q_30_), .Y(_abc_43815_n3281) );
  AND2X2 AND2X2_1404 ( .A(_abc_43815_n1060_bF_buf3), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_43815_n3282_1) );
  AND2X2 AND2X2_1405 ( .A(_abc_43815_n3279), .B(_abc_43815_n3285), .Y(_abc_43815_n3286_1) );
  AND2X2 AND2X2_1406 ( .A(_abc_43815_n3002_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_43815_n3287) );
  AND2X2 AND2X2_1407 ( .A(_abc_43815_n2991_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_43815_n3290_1) );
  AND2X2 AND2X2_1408 ( .A(_abc_43815_n2993_1_bF_buf1), .B(epc_q_31_), .Y(_abc_43815_n3291) );
  AND2X2 AND2X2_1409 ( .A(_abc_43815_n1060_bF_buf2), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1), .Y(_abc_43815_n3292_1) );
  AND2X2 AND2X2_141 ( .A(_abc_43815_n865_1), .B(_abc_43815_n686_1_bF_buf1), .Y(_abc_43815_n866) );
  AND2X2 AND2X2_1410 ( .A(_abc_43815_n3289), .B(_abc_43815_n3295), .Y(_abc_43815_n3296_1) );
  AND2X2 AND2X2_1411 ( .A(_abc_43815_n3002_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_43815_n3297) );
  AND2X2 AND2X2_1412 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_0_), .B(alu_op_r_0_), .Y(_abc_43815_n3315) );
  AND2X2 AND2X2_1413 ( .A(_abc_43815_n3316_1), .B(_abc_43815_n1222), .Y(_abc_43815_n3317) );
  AND2X2 AND2X2_1414 ( .A(_abc_43815_n3318), .B(_abc_43815_n3313), .Y(mem_offset_q_0__FF_INPUT) );
  AND2X2 AND2X2_1415 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_1_), .B(alu_op_r_1_), .Y(_abc_43815_n3321) );
  AND2X2 AND2X2_1416 ( .A(_abc_43815_n3322), .B(_abc_43815_n1224), .Y(_abc_43815_n3323_1) );
  AND2X2 AND2X2_1417 ( .A(_abc_43815_n3324_1), .B(_abc_43815_n3316_1), .Y(_abc_43815_n3325) );
  AND2X2 AND2X2_1418 ( .A(_abc_43815_n3323_1), .B(_abc_43815_n3315), .Y(_abc_43815_n3326) );
  AND2X2 AND2X2_1419 ( .A(_abc_43815_n3329), .B(_abc_43815_n3320), .Y(mem_offset_q_1__FF_INPUT) );
  AND2X2 AND2X2_142 ( .A(_abc_43815_n866), .B(_abc_43815_n864), .Y(_abc_43815_n867) );
  AND2X2 AND2X2_1420 ( .A(mem_ack_i), .B(state_q_2_), .Y(_abc_27555_n4367) );
  AND2X2 AND2X2_1421 ( .A(_abc_27555_n4367_bF_buf6), .B(_abc_43815_n3333), .Y(_abc_43815_n3334) );
  AND2X2 AND2X2_1422 ( .A(_abc_43815_n3335), .B(_abc_43815_n3332_1), .Y(opcode_q_0__FF_INPUT) );
  AND2X2 AND2X2_1423 ( .A(_abc_27555_n4367_bF_buf4), .B(_abc_43815_n3338), .Y(_abc_43815_n3339_1) );
  AND2X2 AND2X2_1424 ( .A(_abc_43815_n3340_1), .B(_abc_43815_n3337), .Y(opcode_q_1__FF_INPUT) );
  AND2X2 AND2X2_1425 ( .A(_abc_27555_n4367_bF_buf2), .B(_abc_43815_n3343), .Y(_abc_43815_n3344) );
  AND2X2 AND2X2_1426 ( .A(_abc_43815_n3345), .B(_abc_43815_n3342), .Y(opcode_q_2__FF_INPUT) );
  AND2X2 AND2X2_1427 ( .A(_abc_27555_n4367_bF_buf0), .B(_abc_43815_n3348_1), .Y(_abc_43815_n3349) );
  AND2X2 AND2X2_1428 ( .A(_abc_43815_n3350), .B(_abc_43815_n3347_1), .Y(opcode_q_3__FF_INPUT) );
  AND2X2 AND2X2_1429 ( .A(_abc_27555_n4367_bF_buf6), .B(_abc_43815_n3353), .Y(_abc_43815_n3354) );
  AND2X2 AND2X2_143 ( .A(_abc_43815_n868_1), .B(_abc_43815_n863), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_) );
  AND2X2 AND2X2_1430 ( .A(_abc_43815_n3355), .B(_abc_43815_n3352), .Y(opcode_q_4__FF_INPUT) );
  AND2X2 AND2X2_1431 ( .A(_abc_27555_n4367_bF_buf4), .B(_abc_43815_n3358), .Y(_abc_43815_n3359_1) );
  AND2X2 AND2X2_1432 ( .A(_abc_43815_n3360_1), .B(_abc_43815_n3357), .Y(opcode_q_5__FF_INPUT) );
  AND2X2 AND2X2_1433 ( .A(_abc_27555_n4367_bF_buf2), .B(_abc_43815_n3363), .Y(_abc_43815_n3364) );
  AND2X2 AND2X2_1434 ( .A(_abc_43815_n3365), .B(_abc_43815_n3362), .Y(opcode_q_6__FF_INPUT) );
  AND2X2 AND2X2_1435 ( .A(_abc_27555_n4367_bF_buf0), .B(_abc_43815_n3368), .Y(_abc_43815_n3369_1) );
  AND2X2 AND2X2_1436 ( .A(_abc_43815_n3370_1), .B(_abc_43815_n3367), .Y(opcode_q_7__FF_INPUT) );
  AND2X2 AND2X2_1437 ( .A(_abc_27555_n4367_bF_buf6), .B(_abc_43815_n3373), .Y(_abc_43815_n3374) );
  AND2X2 AND2X2_1438 ( .A(_abc_43815_n3375), .B(_abc_43815_n3372), .Y(opcode_q_8__FF_INPUT) );
  AND2X2 AND2X2_1439 ( .A(_abc_27555_n4367_bF_buf4), .B(_abc_43815_n3378), .Y(_abc_43815_n3379_1) );
  AND2X2 AND2X2_144 ( .A(_abc_43815_n697), .B(\mem_dat_i[14] ), .Y(_abc_43815_n870) );
  AND2X2 AND2X2_1440 ( .A(_abc_43815_n3380_1), .B(_abc_43815_n3377), .Y(opcode_q_9__FF_INPUT) );
  AND2X2 AND2X2_1441 ( .A(_abc_27555_n4367_bF_buf2), .B(_abc_43815_n3383), .Y(_abc_43815_n3384) );
  AND2X2 AND2X2_1442 ( .A(_abc_43815_n3385), .B(_abc_43815_n3382), .Y(opcode_q_10__FF_INPUT) );
  AND2X2 AND2X2_1443 ( .A(_abc_27555_n4367_bF_buf0), .B(_abc_43815_n3388), .Y(_abc_43815_n3389_1) );
  AND2X2 AND2X2_1444 ( .A(_abc_43815_n3390_1), .B(_abc_43815_n3387), .Y(opcode_q_11__FF_INPUT) );
  AND2X2 AND2X2_1445 ( .A(_abc_27555_n4367_bF_buf6), .B(_abc_43815_n3393), .Y(_abc_43815_n3394) );
  AND2X2 AND2X2_1446 ( .A(_abc_43815_n3395), .B(_abc_43815_n3392), .Y(opcode_q_12__FF_INPUT) );
  AND2X2 AND2X2_1447 ( .A(_abc_27555_n4367_bF_buf4), .B(_abc_43815_n3398), .Y(_abc_43815_n3399_1) );
  AND2X2 AND2X2_1448 ( .A(_abc_43815_n3400_1), .B(_abc_43815_n3397), .Y(opcode_q_13__FF_INPUT) );
  AND2X2 AND2X2_1449 ( .A(_abc_27555_n4367_bF_buf2), .B(_abc_43815_n3403), .Y(_abc_43815_n3404) );
  AND2X2 AND2X2_145 ( .A(_abc_43815_n693), .B(_abc_43815_n802), .Y(_abc_43815_n871) );
  AND2X2 AND2X2_1450 ( .A(_abc_43815_n3405), .B(_abc_43815_n3402), .Y(opcode_q_14__FF_INPUT) );
  AND2X2 AND2X2_1451 ( .A(_abc_27555_n4367_bF_buf0), .B(_abc_43815_n3408), .Y(_abc_43815_n3409_1) );
  AND2X2 AND2X2_1452 ( .A(_abc_43815_n3410_1), .B(_abc_43815_n3407), .Y(opcode_q_15__FF_INPUT) );
  AND2X2 AND2X2_1453 ( .A(_abc_27555_n4367_bF_buf6), .B(_abc_43815_n3413), .Y(_abc_43815_n3414) );
  AND2X2 AND2X2_1454 ( .A(_abc_43815_n3415), .B(_abc_43815_n3412), .Y(opcode_q_16__FF_INPUT) );
  AND2X2 AND2X2_1455 ( .A(_abc_27555_n4367_bF_buf4), .B(_abc_43815_n3418), .Y(_abc_43815_n3419_1) );
  AND2X2 AND2X2_1456 ( .A(_abc_43815_n3420_1), .B(_abc_43815_n3417), .Y(opcode_q_17__FF_INPUT) );
  AND2X2 AND2X2_1457 ( .A(_abc_27555_n4367_bF_buf2), .B(_abc_43815_n3423), .Y(_abc_43815_n3424) );
  AND2X2 AND2X2_1458 ( .A(_abc_43815_n3425), .B(_abc_43815_n3422), .Y(opcode_q_18__FF_INPUT) );
  AND2X2 AND2X2_1459 ( .A(_abc_27555_n4367_bF_buf0), .B(_abc_43815_n3428), .Y(_abc_43815_n3429_1) );
  AND2X2 AND2X2_146 ( .A(_abc_43815_n872), .B(_abc_43815_n686_1_bF_buf0), .Y(_abc_43815_n873) );
  AND2X2 AND2X2_1460 ( .A(_abc_43815_n3430_1), .B(_abc_43815_n3427), .Y(opcode_q_19__FF_INPUT) );
  AND2X2 AND2X2_1461 ( .A(_abc_27555_n4367_bF_buf6), .B(_abc_43815_n3433), .Y(_abc_43815_n3434) );
  AND2X2 AND2X2_1462 ( .A(_abc_43815_n3435), .B(_abc_43815_n3432), .Y(opcode_q_20__FF_INPUT) );
  AND2X2 AND2X2_1463 ( .A(_abc_27555_n4367_bF_buf4), .B(_abc_43815_n3438_1), .Y(_abc_43815_n3439_1) );
  AND2X2 AND2X2_1464 ( .A(_abc_43815_n3440), .B(_abc_43815_n3437), .Y(opcode_q_21__FF_INPUT) );
  AND2X2 AND2X2_1465 ( .A(_abc_27555_n4367_bF_buf2), .B(_abc_43815_n3443), .Y(_abc_43815_n3444) );
  AND2X2 AND2X2_1466 ( .A(_abc_43815_n3445), .B(_abc_43815_n3442), .Y(opcode_q_22__FF_INPUT) );
  AND2X2 AND2X2_1467 ( .A(_abc_27555_n4367_bF_buf0), .B(_abc_43815_n3448_1), .Y(_abc_43815_n3449) );
  AND2X2 AND2X2_1468 ( .A(_abc_43815_n3450), .B(_abc_43815_n3447_1), .Y(opcode_q_23__FF_INPUT) );
  AND2X2 AND2X2_1469 ( .A(_abc_27555_n4367_bF_buf6), .B(_abc_43815_n3453), .Y(_abc_43815_n3454) );
  AND2X2 AND2X2_147 ( .A(_abc_43815_n874), .B(_abc_43815_n875), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_) );
  AND2X2 AND2X2_1470 ( .A(_abc_43815_n3455), .B(_abc_43815_n3452), .Y(opcode_q_24__FF_INPUT) );
  AND2X2 AND2X2_1471 ( .A(_abc_27555_n4367_bF_buf4), .B(_abc_43815_n3458), .Y(_abc_43815_n3459) );
  AND2X2 AND2X2_1472 ( .A(_abc_43815_n3460), .B(_abc_43815_n3457_1), .Y(opcode_q_25__FF_INPUT) );
  AND2X2 AND2X2_1473 ( .A(_abc_27555_n4367_bF_buf2), .B(_abc_43815_n3463), .Y(_abc_43815_n3464) );
  AND2X2 AND2X2_1474 ( .A(_abc_43815_n3465_1), .B(_abc_43815_n3462), .Y(opcode_q_26__FF_INPUT) );
  AND2X2 AND2X2_1475 ( .A(_abc_27555_n4367_bF_buf0), .B(_abc_43815_n3468), .Y(_abc_43815_n3469) );
  AND2X2 AND2X2_1476 ( .A(_abc_43815_n3470), .B(_abc_43815_n3467), .Y(opcode_q_27__FF_INPUT) );
  AND2X2 AND2X2_1477 ( .A(_abc_27555_n4367_bF_buf6), .B(_abc_43815_n3473), .Y(_abc_43815_n3474_1) );
  AND2X2 AND2X2_1478 ( .A(_abc_43815_n3475_1), .B(_abc_43815_n3472), .Y(opcode_q_28__FF_INPUT) );
  AND2X2 AND2X2_1479 ( .A(_abc_27555_n4367_bF_buf4), .B(_abc_43815_n3478), .Y(_abc_43815_n3479) );
  AND2X2 AND2X2_148 ( .A(_abc_43815_n879), .B(_abc_43815_n686_1_bF_buf4), .Y(_abc_43815_n880) );
  AND2X2 AND2X2_1480 ( .A(_abc_43815_n3480), .B(_abc_43815_n3477), .Y(opcode_q_29__FF_INPUT) );
  AND2X2 AND2X2_1481 ( .A(_abc_27555_n4367_bF_buf2), .B(_abc_43815_n3483_1), .Y(_abc_43815_n3484_1) );
  AND2X2 AND2X2_1482 ( .A(_abc_43815_n3485), .B(_abc_43815_n3482), .Y(opcode_q_30__FF_INPUT) );
  AND2X2 AND2X2_1483 ( .A(_abc_27555_n4367_bF_buf0), .B(_abc_43815_n3488), .Y(_abc_43815_n3489) );
  AND2X2 AND2X2_1484 ( .A(_abc_43815_n3490), .B(_abc_43815_n3487), .Y(opcode_q_31__FF_INPUT) );
  AND2X2 AND2X2_1485 ( .A(_abc_43815_n3328), .B(_abc_43815_n3495), .Y(_abc_43815_n3496) );
  AND2X2 AND2X2_1486 ( .A(_abc_43815_n3317_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47802_0_), .Y(_abc_43815_n3497) );
  AND2X2 AND2X2_1487 ( .A(_abc_43815_n3499), .B(_abc_43815_n3494), .Y(_abc_43815_n3500) );
  AND2X2 AND2X2_1488 ( .A(_abc_43815_n3500), .B(_abc_43815_n642_1_bF_buf3), .Y(_abc_43815_n3501_1) );
  AND2X2 AND2X2_1489 ( .A(_abc_43815_n641_bF_buf2), .B(_abc_43815_n3317_bF_buf0), .Y(_abc_43815_n3503) );
  AND2X2 AND2X2_149 ( .A(_abc_43815_n880), .B(_abc_43815_n878), .Y(_abc_43815_n881) );
  AND2X2 AND2X2_1490 ( .A(_abc_43815_n3503), .B(_abc_43815_n3323_1), .Y(_abc_43815_n3504) );
  AND2X2 AND2X2_1491 ( .A(_abc_43815_n3506), .B(_abc_43815_n3492_1), .Y(mem_sel_o_0__FF_INPUT) );
  AND2X2 AND2X2_1492 ( .A(_abc_43815_n642_1_bF_buf2), .B(_abc_43815_n3317_bF_buf3), .Y(_abc_43815_n3511_1) );
  AND2X2 AND2X2_1493 ( .A(_abc_43815_n3511_1), .B(_auto_iopadmap_cc_313_execute_47802_1_), .Y(_abc_43815_n3512_1) );
  AND2X2 AND2X2_1494 ( .A(_abc_43815_n3514), .B(_abc_43815_n3510), .Y(_abc_43815_n3515) );
  AND2X2 AND2X2_1495 ( .A(_abc_43815_n3516), .B(_abc_43815_n3508), .Y(mem_sel_o_1__FF_INPUT) );
  AND2X2 AND2X2_1496 ( .A(_abc_43815_n3519), .B(_abc_43815_n642_1_bF_buf1), .Y(_abc_43815_n3520) );
  AND2X2 AND2X2_1497 ( .A(_abc_43815_n3327), .B(_abc_43815_n3495), .Y(_abc_43815_n3521_1) );
  AND2X2 AND2X2_1498 ( .A(_abc_43815_n3317_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47802_2_), .Y(_abc_43815_n3522_1) );
  AND2X2 AND2X2_1499 ( .A(_abc_43815_n3520), .B(_abc_43815_n3524), .Y(_abc_43815_n3525) );
  AND2X2 AND2X2_15 ( .A(_abc_43815_n640), .B(_abc_43815_n636), .Y(_abc_43815_n641) );
  AND2X2 AND2X2_150 ( .A(_abc_43815_n882), .B(_abc_43815_n877), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_) );
  AND2X2 AND2X2_1500 ( .A(_abc_43815_n3503), .B(_abc_43815_n3324_1), .Y(_abc_43815_n3526) );
  AND2X2 AND2X2_1501 ( .A(_abc_43815_n3528), .B(_abc_43815_n3518), .Y(mem_sel_o_2__FF_INPUT) );
  AND2X2 AND2X2_1502 ( .A(_abc_43815_n3511_1), .B(_auto_iopadmap_cc_313_execute_47802_3_), .Y(_abc_43815_n3532_1) );
  AND2X2 AND2X2_1503 ( .A(_abc_43815_n3534), .B(_abc_43815_n3531_1), .Y(_abc_43815_n3535) );
  AND2X2 AND2X2_1504 ( .A(_abc_43815_n3536), .B(_abc_43815_n3530), .Y(mem_sel_o_3__FF_INPUT) );
  AND2X2 AND2X2_1505 ( .A(_abc_43815_n3538), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_43815_n3539) );
  AND2X2 AND2X2_1506 ( .A(_abc_43815_n649_bF_buf3), .B(_abc_43815_n3317_bF_buf1), .Y(_abc_43815_n3540) );
  AND2X2 AND2X2_1507 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_0_), .Y(_abc_43815_n3542_1) );
  AND2X2 AND2X2_1508 ( .A(_abc_43815_n3496_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_43815_n3543) );
  AND2X2 AND2X2_1509 ( .A(_abc_43815_n3543), .B(_abc_43815_n649_bF_buf2), .Y(_abc_43815_n3544) );
  AND2X2 AND2X2_151 ( .A(_abc_43815_n640), .B(_abc_43815_n653), .Y(_abc_43815_n884_1) );
  AND2X2 AND2X2_1510 ( .A(_abc_43815_n3545), .B(_abc_43815_n642_1_bF_buf0), .Y(_abc_43815_n3546) );
  AND2X2 AND2X2_1511 ( .A(_abc_43815_n3547), .B(_abc_43815_n671_bF_buf2), .Y(_abc_43815_n3548) );
  AND2X2 AND2X2_1512 ( .A(_abc_43815_n3549_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47769_0_), .Y(_abc_43815_n3550) );
  AND2X2 AND2X2_1513 ( .A(_abc_43815_n3538), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_43815_n3552_1) );
  AND2X2 AND2X2_1514 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_1_), .Y(_abc_43815_n3553) );
  AND2X2 AND2X2_1515 ( .A(_abc_43815_n3496_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_43815_n3554) );
  AND2X2 AND2X2_1516 ( .A(_abc_43815_n3554), .B(_abc_43815_n649_bF_buf1), .Y(_abc_43815_n3555) );
  AND2X2 AND2X2_1517 ( .A(_abc_43815_n3556), .B(_abc_43815_n642_1_bF_buf5), .Y(_abc_43815_n3557) );
  AND2X2 AND2X2_1518 ( .A(_abc_43815_n3558), .B(_abc_43815_n671_bF_buf1), .Y(_abc_43815_n3559) );
  AND2X2 AND2X2_1519 ( .A(_abc_43815_n3549_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_1_), .Y(_abc_43815_n3560) );
  AND2X2 AND2X2_152 ( .A(_abc_43815_n812), .B(_abc_43815_n884_1), .Y(_abc_43815_n885_1) );
  AND2X2 AND2X2_1520 ( .A(_abc_43815_n3538), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n3562_1) );
  AND2X2 AND2X2_1521 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_2_), .Y(_abc_43815_n3563) );
  AND2X2 AND2X2_1522 ( .A(_abc_43815_n3496_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n3564) );
  AND2X2 AND2X2_1523 ( .A(_abc_43815_n3564), .B(_abc_43815_n649_bF_buf0), .Y(_abc_43815_n3565) );
  AND2X2 AND2X2_1524 ( .A(_abc_43815_n3566), .B(_abc_43815_n642_1_bF_buf4), .Y(_abc_43815_n3567) );
  AND2X2 AND2X2_1525 ( .A(_abc_43815_n3568), .B(_abc_43815_n671_bF_buf0), .Y(_abc_43815_n3569) );
  AND2X2 AND2X2_1526 ( .A(_abc_43815_n3549_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_2_), .Y(_abc_43815_n3570) );
  AND2X2 AND2X2_1527 ( .A(_abc_43815_n3538), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_43815_n3572_1) );
  AND2X2 AND2X2_1528 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_3_), .Y(_abc_43815_n3573) );
  AND2X2 AND2X2_1529 ( .A(_abc_43815_n3496_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_43815_n3574) );
  AND2X2 AND2X2_153 ( .A(_abc_43815_n692_bF_buf3), .B(\mem_dat_i[16] ), .Y(_abc_43815_n886) );
  AND2X2 AND2X2_1530 ( .A(_abc_43815_n3574), .B(_abc_43815_n649_bF_buf4), .Y(_abc_43815_n3575) );
  AND2X2 AND2X2_1531 ( .A(_abc_43815_n3576), .B(_abc_43815_n642_1_bF_buf3), .Y(_abc_43815_n3577) );
  AND2X2 AND2X2_1532 ( .A(_abc_43815_n3578), .B(_abc_43815_n671_bF_buf4), .Y(_abc_43815_n3579) );
  AND2X2 AND2X2_1533 ( .A(_abc_43815_n3549_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_3_), .Y(_abc_43815_n3580) );
  AND2X2 AND2X2_1534 ( .A(_abc_43815_n3538), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_43815_n3582_1) );
  AND2X2 AND2X2_1535 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_4_), .Y(_abc_43815_n3583) );
  AND2X2 AND2X2_1536 ( .A(_abc_43815_n3496_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_43815_n3584) );
  AND2X2 AND2X2_1537 ( .A(_abc_43815_n3584), .B(_abc_43815_n649_bF_buf3), .Y(_abc_43815_n3585) );
  AND2X2 AND2X2_1538 ( .A(_abc_43815_n3586), .B(_abc_43815_n642_1_bF_buf2), .Y(_abc_43815_n3587) );
  AND2X2 AND2X2_1539 ( .A(_abc_43815_n3588), .B(_abc_43815_n671_bF_buf3), .Y(_abc_43815_n3589) );
  AND2X2 AND2X2_154 ( .A(_abc_43815_n887), .B(_abc_43815_n686_1_bF_buf3), .Y(_abc_43815_n888) );
  AND2X2 AND2X2_1540 ( .A(_abc_43815_n3549_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_4_), .Y(_abc_43815_n3590_1) );
  AND2X2 AND2X2_1541 ( .A(_abc_43815_n3538), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_43815_n3592) );
  AND2X2 AND2X2_1542 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_5_), .Y(_abc_43815_n3593) );
  AND2X2 AND2X2_1543 ( .A(_abc_43815_n3496_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_43815_n3594) );
  AND2X2 AND2X2_1544 ( .A(_abc_43815_n3594), .B(_abc_43815_n649_bF_buf2), .Y(_abc_43815_n3595) );
  AND2X2 AND2X2_1545 ( .A(_abc_43815_n3596), .B(_abc_43815_n642_1_bF_buf1), .Y(_abc_43815_n3597) );
  AND2X2 AND2X2_1546 ( .A(_abc_43815_n3598), .B(_abc_43815_n671_bF_buf2), .Y(_abc_43815_n3599_1) );
  AND2X2 AND2X2_1547 ( .A(_abc_43815_n3549_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47769_5_), .Y(_abc_43815_n3600_1) );
  AND2X2 AND2X2_1548 ( .A(_abc_43815_n3538), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_43815_n3602) );
  AND2X2 AND2X2_1549 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_6_), .Y(_abc_43815_n3603) );
  AND2X2 AND2X2_155 ( .A(_abc_43815_n889), .B(_abc_43815_n890), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_) );
  AND2X2 AND2X2_1550 ( .A(_abc_43815_n3496_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_43815_n3604) );
  AND2X2 AND2X2_1551 ( .A(_abc_43815_n3604), .B(_abc_43815_n649_bF_buf1), .Y(_abc_43815_n3605) );
  AND2X2 AND2X2_1552 ( .A(_abc_43815_n3606), .B(_abc_43815_n642_1_bF_buf0), .Y(_abc_43815_n3607) );
  AND2X2 AND2X2_1553 ( .A(_abc_43815_n3608_1), .B(_abc_43815_n671_bF_buf1), .Y(_abc_43815_n3609_1) );
  AND2X2 AND2X2_1554 ( .A(_abc_43815_n3549_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_6_), .Y(_abc_43815_n3610) );
  AND2X2 AND2X2_1555 ( .A(_abc_43815_n3538), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_43815_n3612) );
  AND2X2 AND2X2_1556 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_7_), .Y(_abc_43815_n3613) );
  AND2X2 AND2X2_1557 ( .A(_abc_43815_n3496_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_43815_n3614) );
  AND2X2 AND2X2_1558 ( .A(_abc_43815_n3614), .B(_abc_43815_n649_bF_buf0), .Y(_abc_43815_n3615) );
  AND2X2 AND2X2_1559 ( .A(_abc_43815_n3616), .B(_abc_43815_n642_1_bF_buf5), .Y(_abc_43815_n3617_1) );
  AND2X2 AND2X2_156 ( .A(_abc_43815_n692_bF_buf2), .B(\mem_dat_i[17] ), .Y(_abc_43815_n892) );
  AND2X2 AND2X2_1560 ( .A(_abc_43815_n3618_1), .B(_abc_43815_n671_bF_buf0), .Y(_abc_43815_n3619) );
  AND2X2 AND2X2_1561 ( .A(_abc_43815_n3549_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_7_), .Y(_abc_43815_n3620) );
  AND2X2 AND2X2_1562 ( .A(_abc_43815_n3549_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_8_), .Y(_abc_43815_n3622) );
  AND2X2 AND2X2_1563 ( .A(_abc_43815_n3496_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_43815_n3623) );
  AND2X2 AND2X2_1564 ( .A(_abc_43815_n3317_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_8_), .Y(_abc_43815_n3624) );
  AND2X2 AND2X2_1565 ( .A(_abc_43815_n645_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_43815_n3627_1) );
  AND2X2 AND2X2_1566 ( .A(_abc_43815_n646_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_8_), .Y(_abc_43815_n3628) );
  AND2X2 AND2X2_1567 ( .A(_abc_43815_n3626_1), .B(_abc_43815_n3630), .Y(_abc_43815_n3631) );
  AND2X2 AND2X2_1568 ( .A(_abc_43815_n3633), .B(_abc_43815_n671_bF_buf4), .Y(_abc_43815_n3634) );
  AND2X2 AND2X2_1569 ( .A(_abc_43815_n3632), .B(_abc_43815_n3634), .Y(_abc_43815_n3635_1) );
  AND2X2 AND2X2_157 ( .A(_abc_43815_n893), .B(_abc_43815_n686_1_bF_buf2), .Y(_abc_43815_n894) );
  AND2X2 AND2X2_1570 ( .A(_abc_43815_n3549_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_9_), .Y(_abc_43815_n3637) );
  AND2X2 AND2X2_1571 ( .A(_abc_43815_n3496_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n3638) );
  AND2X2 AND2X2_1572 ( .A(_abc_43815_n3317_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_9_), .Y(_abc_43815_n3639) );
  AND2X2 AND2X2_1573 ( .A(_abc_43815_n645_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n3642) );
  AND2X2 AND2X2_1574 ( .A(_abc_43815_n646_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_9_), .Y(_abc_43815_n3643) );
  AND2X2 AND2X2_1575 ( .A(_abc_43815_n3641), .B(_abc_43815_n3645_1), .Y(_abc_43815_n3646) );
  AND2X2 AND2X2_1576 ( .A(_abc_43815_n3648), .B(_abc_43815_n671_bF_buf3), .Y(_abc_43815_n3649) );
  AND2X2 AND2X2_1577 ( .A(_abc_43815_n3647), .B(_abc_43815_n3649), .Y(_abc_43815_n3650) );
  AND2X2 AND2X2_1578 ( .A(_abc_43815_n3549_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47769_10_), .Y(_abc_43815_n3652) );
  AND2X2 AND2X2_1579 ( .A(_abc_43815_n3496_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_43815_n3653_1) );
  AND2X2 AND2X2_158 ( .A(_abc_43815_n895), .B(_abc_43815_n896), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_) );
  AND2X2 AND2X2_1580 ( .A(_abc_43815_n3317_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_10_), .Y(_abc_43815_n3654) );
  AND2X2 AND2X2_1581 ( .A(_abc_43815_n645_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_43815_n3657) );
  AND2X2 AND2X2_1582 ( .A(_abc_43815_n646_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_10_), .Y(_abc_43815_n3658) );
  AND2X2 AND2X2_1583 ( .A(_abc_43815_n3656), .B(_abc_43815_n3660), .Y(_abc_43815_n3661) );
  AND2X2 AND2X2_1584 ( .A(_abc_43815_n3663), .B(_abc_43815_n671_bF_buf2), .Y(_abc_43815_n3664) );
  AND2X2 AND2X2_1585 ( .A(_abc_43815_n3662), .B(_abc_43815_n3664), .Y(_abc_43815_n3665) );
  AND2X2 AND2X2_1586 ( .A(_abc_43815_n3549_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_11_), .Y(_abc_43815_n3667_1) );
  AND2X2 AND2X2_1587 ( .A(_abc_43815_n3496_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_43815_n3668_1) );
  AND2X2 AND2X2_1588 ( .A(_abc_43815_n3317_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_11_), .Y(_abc_43815_n3669_1) );
  AND2X2 AND2X2_1589 ( .A(_abc_43815_n645_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_43815_n3672) );
  AND2X2 AND2X2_159 ( .A(_abc_43815_n692_bF_buf1), .B(\mem_dat_i[18] ), .Y(_abc_43815_n898) );
  AND2X2 AND2X2_1590 ( .A(_abc_43815_n646_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_11_), .Y(_abc_43815_n3673) );
  AND2X2 AND2X2_1591 ( .A(_abc_43815_n3671), .B(_abc_43815_n3675), .Y(_abc_43815_n3676) );
  AND2X2 AND2X2_1592 ( .A(_abc_43815_n3678), .B(_abc_43815_n671_bF_buf1), .Y(_abc_43815_n3679) );
  AND2X2 AND2X2_1593 ( .A(_abc_43815_n3677), .B(_abc_43815_n3679), .Y(_abc_43815_n3680_1) );
  AND2X2 AND2X2_1594 ( .A(_abc_43815_n3549_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_12_), .Y(_abc_43815_n3682) );
  AND2X2 AND2X2_1595 ( .A(_abc_43815_n3496_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_43815_n3683_1) );
  AND2X2 AND2X2_1596 ( .A(_abc_43815_n3317_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_12_), .Y(_abc_43815_n3684) );
  AND2X2 AND2X2_1597 ( .A(_abc_43815_n645_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_43815_n3687) );
  AND2X2 AND2X2_1598 ( .A(_abc_43815_n646_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_12_), .Y(_abc_43815_n3688) );
  AND2X2 AND2X2_1599 ( .A(_abc_43815_n3686), .B(_abc_43815_n3690), .Y(_abc_43815_n3691) );
  AND2X2 AND2X2_16 ( .A(_abc_43815_n629), .B(inst_r_0_), .Y(_abc_43815_n643_1) );
  AND2X2 AND2X2_160 ( .A(_abc_43815_n899), .B(_abc_43815_n686_1_bF_buf1), .Y(_abc_43815_n900_1) );
  AND2X2 AND2X2_1600 ( .A(_abc_43815_n3693), .B(_abc_43815_n671_bF_buf0), .Y(_abc_43815_n3694_1) );
  AND2X2 AND2X2_1601 ( .A(_abc_43815_n3692), .B(_abc_43815_n3694_1), .Y(_abc_43815_n3695_1) );
  AND2X2 AND2X2_1602 ( .A(_abc_43815_n3549_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_13_), .Y(_abc_43815_n3697) );
  AND2X2 AND2X2_1603 ( .A(_abc_43815_n3496_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_43815_n3698) );
  AND2X2 AND2X2_1604 ( .A(_abc_43815_n3317_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_13_), .Y(_abc_43815_n3699) );
  AND2X2 AND2X2_1605 ( .A(_abc_43815_n645_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_43815_n3702_1) );
  AND2X2 AND2X2_1606 ( .A(_abc_43815_n646_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_13_), .Y(_abc_43815_n3703) );
  AND2X2 AND2X2_1607 ( .A(_abc_43815_n3701_1), .B(_abc_43815_n3705), .Y(_abc_43815_n3706) );
  AND2X2 AND2X2_1608 ( .A(_abc_43815_n3708), .B(_abc_43815_n671_bF_buf4), .Y(_abc_43815_n3709) );
  AND2X2 AND2X2_1609 ( .A(_abc_43815_n3707_1), .B(_abc_43815_n3709), .Y(_abc_43815_n3710) );
  AND2X2 AND2X2_161 ( .A(_abc_43815_n901), .B(_abc_43815_n902), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_) );
  AND2X2 AND2X2_1610 ( .A(_abc_43815_n3549_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_14_), .Y(_abc_43815_n3712) );
  AND2X2 AND2X2_1611 ( .A(_abc_43815_n3496_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_43815_n3713_1) );
  AND2X2 AND2X2_1612 ( .A(_abc_43815_n3317_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_14_), .Y(_abc_43815_n3714) );
  AND2X2 AND2X2_1613 ( .A(_abc_43815_n645_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_43815_n3717) );
  AND2X2 AND2X2_1614 ( .A(_abc_43815_n646_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_14_), .Y(_abc_43815_n3718) );
  AND2X2 AND2X2_1615 ( .A(_abc_43815_n3716), .B(_abc_43815_n3720_1), .Y(_abc_43815_n3721) );
  AND2X2 AND2X2_1616 ( .A(_abc_43815_n3723), .B(_abc_43815_n671_bF_buf3), .Y(_abc_43815_n3724) );
  AND2X2 AND2X2_1617 ( .A(_abc_43815_n3722), .B(_abc_43815_n3724), .Y(_abc_43815_n3725) );
  AND2X2 AND2X2_1618 ( .A(_abc_43815_n3549_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47769_15_), .Y(_abc_43815_n3727) );
  AND2X2 AND2X2_1619 ( .A(_abc_43815_n3496_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_43815_n3728) );
  AND2X2 AND2X2_162 ( .A(_abc_43815_n692_bF_buf0), .B(\mem_dat_i[19] ), .Y(_abc_43815_n904) );
  AND2X2 AND2X2_1620 ( .A(_abc_43815_n3317_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_15_), .Y(_abc_43815_n3729) );
  AND2X2 AND2X2_1621 ( .A(_abc_43815_n645_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_43815_n3732) );
  AND2X2 AND2X2_1622 ( .A(_abc_43815_n646_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_15_), .Y(_abc_43815_n3733_1) );
  AND2X2 AND2X2_1623 ( .A(_abc_43815_n3731), .B(_abc_43815_n3735), .Y(_abc_43815_n3736) );
  AND2X2 AND2X2_1624 ( .A(_abc_43815_n3738), .B(_abc_43815_n671_bF_buf2), .Y(_abc_43815_n3739) );
  AND2X2 AND2X2_1625 ( .A(_abc_43815_n3737), .B(_abc_43815_n3739), .Y(_abc_43815_n3740) );
  AND2X2 AND2X2_1626 ( .A(_abc_43815_n3549_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_16_), .Y(_abc_43815_n3742) );
  AND2X2 AND2X2_1627 ( .A(_abc_43815_n3526), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_43815_n3743_1) );
  AND2X2 AND2X2_1628 ( .A(_abc_43815_n3521_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_43815_n3744) );
  AND2X2 AND2X2_1629 ( .A(_abc_43815_n3744), .B(_abc_43815_n649_bF_buf1), .Y(_abc_43815_n3745) );
  AND2X2 AND2X2_163 ( .A(_abc_43815_n905), .B(_abc_43815_n686_1_bF_buf0), .Y(_abc_43815_n906) );
  AND2X2 AND2X2_1630 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_16_), .Y(_abc_43815_n3746) );
  AND2X2 AND2X2_1631 ( .A(_abc_43815_n650_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_43815_n3747) );
  AND2X2 AND2X2_1632 ( .A(_abc_43815_n3747), .B(_abc_43815_n645_1_bF_buf4), .Y(_abc_43815_n3748) );
  AND2X2 AND2X2_1633 ( .A(_abc_43815_n3750_1), .B(_abc_43815_n642_1_bF_buf2), .Y(_abc_43815_n3751) );
  AND2X2 AND2X2_1634 ( .A(_abc_43815_n3752), .B(_abc_43815_n671_bF_buf1), .Y(_abc_43815_n3753) );
  AND2X2 AND2X2_1635 ( .A(_abc_43815_n3549_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_17_), .Y(_abc_43815_n3755) );
  AND2X2 AND2X2_1636 ( .A(_abc_43815_n3526), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_43815_n3756_1) );
  AND2X2 AND2X2_1637 ( .A(_abc_43815_n3521_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_43815_n3757) );
  AND2X2 AND2X2_1638 ( .A(_abc_43815_n3757), .B(_abc_43815_n649_bF_buf0), .Y(_abc_43815_n3758) );
  AND2X2 AND2X2_1639 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_17_), .Y(_abc_43815_n3759) );
  AND2X2 AND2X2_164 ( .A(_abc_43815_n907), .B(_abc_43815_n908), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_) );
  AND2X2 AND2X2_1640 ( .A(_abc_43815_n650_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_43815_n3760) );
  AND2X2 AND2X2_1641 ( .A(_abc_43815_n3760), .B(_abc_43815_n645_1_bF_buf3), .Y(_abc_43815_n3761) );
  AND2X2 AND2X2_1642 ( .A(_abc_43815_n3763_1), .B(_abc_43815_n642_1_bF_buf1), .Y(_abc_43815_n3764) );
  AND2X2 AND2X2_1643 ( .A(_abc_43815_n3765), .B(_abc_43815_n671_bF_buf0), .Y(_abc_43815_n3766) );
  AND2X2 AND2X2_1644 ( .A(_abc_43815_n3549_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_18_), .Y(_abc_43815_n3768) );
  AND2X2 AND2X2_1645 ( .A(_abc_43815_n3526), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n3769) );
  AND2X2 AND2X2_1646 ( .A(_abc_43815_n3521_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n3770) );
  AND2X2 AND2X2_1647 ( .A(_abc_43815_n3770), .B(_abc_43815_n649_bF_buf4), .Y(_abc_43815_n3771) );
  AND2X2 AND2X2_1648 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_18_), .Y(_abc_43815_n3772) );
  AND2X2 AND2X2_1649 ( .A(_abc_43815_n650_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_43815_n3773_1) );
  AND2X2 AND2X2_165 ( .A(_abc_43815_n692_bF_buf3), .B(\mem_dat_i[20] ), .Y(_abc_43815_n910) );
  AND2X2 AND2X2_1650 ( .A(_abc_43815_n3773_1), .B(_abc_43815_n645_1_bF_buf2), .Y(_abc_43815_n3774) );
  AND2X2 AND2X2_1651 ( .A(_abc_43815_n3776), .B(_abc_43815_n642_1_bF_buf0), .Y(_abc_43815_n3777) );
  AND2X2 AND2X2_1652 ( .A(_abc_43815_n3778), .B(_abc_43815_n671_bF_buf4), .Y(_abc_43815_n3779) );
  AND2X2 AND2X2_1653 ( .A(_abc_43815_n3549_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_19_), .Y(_abc_43815_n3781) );
  AND2X2 AND2X2_1654 ( .A(_abc_43815_n3526), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_43815_n3782) );
  AND2X2 AND2X2_1655 ( .A(_abc_43815_n3521_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_43815_n3783) );
  AND2X2 AND2X2_1656 ( .A(_abc_43815_n3783), .B(_abc_43815_n649_bF_buf3), .Y(_abc_43815_n3784) );
  AND2X2 AND2X2_1657 ( .A(_abc_43815_n645_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_43815_n3785) );
  AND2X2 AND2X2_1658 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_19_), .Y(_abc_43815_n3786_1) );
  AND2X2 AND2X2_1659 ( .A(_abc_43815_n3788), .B(_abc_43815_n642_1_bF_buf5), .Y(_abc_43815_n3789) );
  AND2X2 AND2X2_166 ( .A(_abc_43815_n911), .B(_abc_43815_n686_1_bF_buf4), .Y(_abc_43815_n912) );
  AND2X2 AND2X2_1660 ( .A(_abc_43815_n3790), .B(_abc_43815_n671_bF_buf3), .Y(_abc_43815_n3791) );
  AND2X2 AND2X2_1661 ( .A(_abc_43815_n3549_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47769_20_), .Y(_abc_43815_n3793_1) );
  AND2X2 AND2X2_1662 ( .A(_abc_43815_n3526), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_43815_n3794) );
  AND2X2 AND2X2_1663 ( .A(_abc_43815_n3521_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_43815_n3795) );
  AND2X2 AND2X2_1664 ( .A(_abc_43815_n3795), .B(_abc_43815_n649_bF_buf2), .Y(_abc_43815_n3796) );
  AND2X2 AND2X2_1665 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_20_), .Y(_abc_43815_n3797) );
  AND2X2 AND2X2_1666 ( .A(_abc_43815_n650_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_43815_n3798) );
  AND2X2 AND2X2_1667 ( .A(_abc_43815_n3798), .B(_abc_43815_n645_1_bF_buf0), .Y(_abc_43815_n3799) );
  AND2X2 AND2X2_1668 ( .A(_abc_43815_n3801), .B(_abc_43815_n642_1_bF_buf4), .Y(_abc_43815_n3802) );
  AND2X2 AND2X2_1669 ( .A(_abc_43815_n3803), .B(_abc_43815_n671_bF_buf2), .Y(_abc_43815_n3804) );
  AND2X2 AND2X2_167 ( .A(_abc_43815_n913), .B(_abc_43815_n914), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_) );
  AND2X2 AND2X2_1670 ( .A(_abc_43815_n3549_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_21_), .Y(_abc_43815_n3806) );
  AND2X2 AND2X2_1671 ( .A(_abc_43815_n3526), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_43815_n3807) );
  AND2X2 AND2X2_1672 ( .A(_abc_43815_n3521_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_43815_n3808) );
  AND2X2 AND2X2_1673 ( .A(_abc_43815_n3808), .B(_abc_43815_n649_bF_buf1), .Y(_abc_43815_n3809) );
  AND2X2 AND2X2_1674 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_21_), .Y(_abc_43815_n3810) );
  AND2X2 AND2X2_1675 ( .A(_abc_43815_n650_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_43815_n3811) );
  AND2X2 AND2X2_1676 ( .A(_abc_43815_n3811), .B(_abc_43815_n645_1_bF_buf4), .Y(_abc_43815_n3812_1) );
  AND2X2 AND2X2_1677 ( .A(_abc_43815_n3814), .B(_abc_43815_n642_1_bF_buf3), .Y(_abc_43815_n3815) );
  AND2X2 AND2X2_1678 ( .A(_abc_43815_n3816), .B(_abc_43815_n671_bF_buf1), .Y(_abc_43815_n3817) );
  AND2X2 AND2X2_1679 ( .A(_abc_43815_n3549_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_22_), .Y(_abc_43815_n3819) );
  AND2X2 AND2X2_168 ( .A(_abc_43815_n692_bF_buf2), .B(\mem_dat_i[21] ), .Y(_abc_43815_n916_1) );
  AND2X2 AND2X2_1680 ( .A(_abc_43815_n3526), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_43815_n3820) );
  AND2X2 AND2X2_1681 ( .A(_abc_43815_n3521_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_43815_n3821) );
  AND2X2 AND2X2_1682 ( .A(_abc_43815_n3821), .B(_abc_43815_n649_bF_buf0), .Y(_abc_43815_n3822) );
  AND2X2 AND2X2_1683 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_22_), .Y(_abc_43815_n3823) );
  AND2X2 AND2X2_1684 ( .A(_abc_43815_n650_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_43815_n3824) );
  AND2X2 AND2X2_1685 ( .A(_abc_43815_n3824), .B(_abc_43815_n645_1_bF_buf3), .Y(_abc_43815_n3825_1) );
  AND2X2 AND2X2_1686 ( .A(_abc_43815_n3827), .B(_abc_43815_n642_1_bF_buf2), .Y(_abc_43815_n3828) );
  AND2X2 AND2X2_1687 ( .A(_abc_43815_n3829), .B(_abc_43815_n671_bF_buf0), .Y(_abc_43815_n3830) );
  AND2X2 AND2X2_1688 ( .A(_abc_43815_n3549_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_23_), .Y(_abc_43815_n3832) );
  AND2X2 AND2X2_1689 ( .A(_abc_43815_n3526), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_43815_n3833) );
  AND2X2 AND2X2_169 ( .A(_abc_43815_n917_1), .B(_abc_43815_n686_1_bF_buf3), .Y(_abc_43815_n918) );
  AND2X2 AND2X2_1690 ( .A(_abc_43815_n3521_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_43815_n3834) );
  AND2X2 AND2X2_1691 ( .A(_abc_43815_n3834), .B(_abc_43815_n649_bF_buf4), .Y(_abc_43815_n3835_1) );
  AND2X2 AND2X2_1692 ( .A(_abc_43815_n645_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_43815_n3836) );
  AND2X2 AND2X2_1693 ( .A(_abc_43815_n3541_1), .B(_auto_iopadmap_cc_313_execute_47769_23_), .Y(_abc_43815_n3837) );
  AND2X2 AND2X2_1694 ( .A(_abc_43815_n3839), .B(_abc_43815_n642_1_bF_buf1), .Y(_abc_43815_n3840) );
  AND2X2 AND2X2_1695 ( .A(_abc_43815_n3841), .B(_abc_43815_n671_bF_buf4), .Y(_abc_43815_n3842_1) );
  AND2X2 AND2X2_1696 ( .A(_abc_43815_n3549_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_24_), .Y(_abc_43815_n3844) );
  AND2X2 AND2X2_1697 ( .A(_abc_43815_n646_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_24_), .Y(_abc_43815_n3846) );
  AND2X2 AND2X2_1698 ( .A(_abc_43815_n645_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_43815_n3847) );
  AND2X2 AND2X2_1699 ( .A(_abc_43815_n3521_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_43815_n3850) );
  AND2X2 AND2X2_17 ( .A(_abc_43815_n638), .B(_abc_43815_n643_1), .Y(_abc_43815_n644) );
  AND2X2 AND2X2_170 ( .A(_abc_43815_n919), .B(_abc_43815_n920), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_) );
  AND2X2 AND2X2_1700 ( .A(_abc_43815_n3317_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_24_), .Y(_abc_43815_n3851) );
  AND2X2 AND2X2_1701 ( .A(_abc_43815_n3853), .B(_abc_43815_n3849_1), .Y(_abc_43815_n3854) );
  AND2X2 AND2X2_1702 ( .A(_abc_43815_n3855), .B(_abc_43815_n3845), .Y(_abc_43815_n3856_1) );
  AND2X2 AND2X2_1703 ( .A(_abc_43815_n3856_1), .B(_abc_43815_n671_bF_buf3), .Y(_abc_43815_n3857) );
  AND2X2 AND2X2_1704 ( .A(_abc_43815_n3549_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47769_25_), .Y(_abc_43815_n3859) );
  AND2X2 AND2X2_1705 ( .A(_abc_43815_n646_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_25_), .Y(_abc_43815_n3861) );
  AND2X2 AND2X2_1706 ( .A(_abc_43815_n645_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_43815_n3862) );
  AND2X2 AND2X2_1707 ( .A(_abc_43815_n3521_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n3865) );
  AND2X2 AND2X2_1708 ( .A(_abc_43815_n3317_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_25_), .Y(_abc_43815_n3866) );
  AND2X2 AND2X2_1709 ( .A(_abc_43815_n3868), .B(_abc_43815_n3864), .Y(_abc_43815_n3869) );
  AND2X2 AND2X2_171 ( .A(_abc_43815_n692_bF_buf1), .B(\mem_dat_i[22] ), .Y(_abc_43815_n922) );
  AND2X2 AND2X2_1710 ( .A(_abc_43815_n3870_1), .B(_abc_43815_n3860), .Y(_abc_43815_n3871) );
  AND2X2 AND2X2_1711 ( .A(_abc_43815_n3871), .B(_abc_43815_n671_bF_buf2), .Y(_abc_43815_n3872) );
  AND2X2 AND2X2_1712 ( .A(_abc_43815_n3549_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_26_), .Y(_abc_43815_n3874) );
  AND2X2 AND2X2_1713 ( .A(_abc_43815_n646_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_26_), .Y(_abc_43815_n3876) );
  AND2X2 AND2X2_1714 ( .A(_abc_43815_n645_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_43815_n3877_1) );
  AND2X2 AND2X2_1715 ( .A(_abc_43815_n3521_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_43815_n3880) );
  AND2X2 AND2X2_1716 ( .A(_abc_43815_n3317_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_26_), .Y(_abc_43815_n3881) );
  AND2X2 AND2X2_1717 ( .A(_abc_43815_n3883), .B(_abc_43815_n3879), .Y(_abc_43815_n3884_1) );
  AND2X2 AND2X2_1718 ( .A(_abc_43815_n3885), .B(_abc_43815_n3875), .Y(_abc_43815_n3886) );
  AND2X2 AND2X2_1719 ( .A(_abc_43815_n3886), .B(_abc_43815_n671_bF_buf1), .Y(_abc_43815_n3887) );
  AND2X2 AND2X2_172 ( .A(_abc_43815_n923), .B(_abc_43815_n686_1_bF_buf2), .Y(_abc_43815_n924) );
  AND2X2 AND2X2_1720 ( .A(_abc_43815_n3549_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_27_), .Y(_abc_43815_n3889) );
  AND2X2 AND2X2_1721 ( .A(_abc_43815_n646_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_27_), .Y(_abc_43815_n3891_1) );
  AND2X2 AND2X2_1722 ( .A(_abc_43815_n645_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_43815_n3892) );
  AND2X2 AND2X2_1723 ( .A(_abc_43815_n3521_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_43815_n3895) );
  AND2X2 AND2X2_1724 ( .A(_abc_43815_n3317_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_27_), .Y(_abc_43815_n3896) );
  AND2X2 AND2X2_1725 ( .A(_abc_43815_n3898), .B(_abc_43815_n3894), .Y(_abc_43815_n3899) );
  AND2X2 AND2X2_1726 ( .A(_abc_43815_n3900), .B(_abc_43815_n3890), .Y(_abc_43815_n3901_1) );
  AND2X2 AND2X2_1727 ( .A(_abc_43815_n3901_1), .B(_abc_43815_n671_bF_buf0), .Y(_abc_43815_n3902) );
  AND2X2 AND2X2_1728 ( .A(_abc_43815_n3549_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_28_), .Y(_abc_43815_n3904) );
  AND2X2 AND2X2_1729 ( .A(_abc_43815_n646_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_28_), .Y(_abc_43815_n3906) );
  AND2X2 AND2X2_173 ( .A(_abc_43815_n925), .B(_abc_43815_n926), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_) );
  AND2X2 AND2X2_1730 ( .A(_abc_43815_n645_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_43815_n3907) );
  AND2X2 AND2X2_1731 ( .A(_abc_43815_n3521_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_43815_n3910) );
  AND2X2 AND2X2_1732 ( .A(_abc_43815_n3317_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_28_), .Y(_abc_43815_n3911) );
  AND2X2 AND2X2_1733 ( .A(_abc_43815_n3913), .B(_abc_43815_n3909), .Y(_abc_43815_n3914) );
  AND2X2 AND2X2_1734 ( .A(_abc_43815_n3915), .B(_abc_43815_n3905), .Y(_abc_43815_n3916_1) );
  AND2X2 AND2X2_1735 ( .A(_abc_43815_n3916_1), .B(_abc_43815_n671_bF_buf4), .Y(_abc_43815_n3917) );
  AND2X2 AND2X2_1736 ( .A(_abc_43815_n3549_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_29_), .Y(_abc_43815_n3919) );
  AND2X2 AND2X2_1737 ( .A(_abc_43815_n646_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47769_29_), .Y(_abc_43815_n3921) );
  AND2X2 AND2X2_1738 ( .A(_abc_43815_n645_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_43815_n3922) );
  AND2X2 AND2X2_1739 ( .A(_abc_43815_n3521_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_43815_n3925) );
  AND2X2 AND2X2_174 ( .A(_abc_43815_n692_bF_buf0), .B(\mem_dat_i[23] ), .Y(_abc_43815_n928) );
  AND2X2 AND2X2_1740 ( .A(_abc_43815_n3317_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_29_), .Y(_abc_43815_n3926) );
  AND2X2 AND2X2_1741 ( .A(_abc_43815_n3928), .B(_abc_43815_n3924), .Y(_abc_43815_n3929) );
  AND2X2 AND2X2_1742 ( .A(_abc_43815_n3930), .B(_abc_43815_n3920), .Y(_abc_43815_n3931) );
  AND2X2 AND2X2_1743 ( .A(_abc_43815_n3931), .B(_abc_43815_n671_bF_buf3), .Y(_abc_43815_n3932) );
  AND2X2 AND2X2_1744 ( .A(_abc_43815_n3549_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47769_30_), .Y(_abc_43815_n3934) );
  AND2X2 AND2X2_1745 ( .A(_abc_43815_n646_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_30_), .Y(_abc_43815_n3936) );
  AND2X2 AND2X2_1746 ( .A(_abc_43815_n645_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_43815_n3937) );
  AND2X2 AND2X2_1747 ( .A(_abc_43815_n3521_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_43815_n3940) );
  AND2X2 AND2X2_1748 ( .A(_abc_43815_n3317_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_30_), .Y(_abc_43815_n3941) );
  AND2X2 AND2X2_1749 ( .A(_abc_43815_n3943), .B(_abc_43815_n3939), .Y(_abc_43815_n3944) );
  AND2X2 AND2X2_175 ( .A(_abc_43815_n929), .B(_abc_43815_n686_1_bF_buf1), .Y(_abc_43815_n930) );
  AND2X2 AND2X2_1750 ( .A(_abc_43815_n3945_1), .B(_abc_43815_n3935), .Y(_abc_43815_n3946) );
  AND2X2 AND2X2_1751 ( .A(_abc_43815_n3946), .B(_abc_43815_n671_bF_buf2), .Y(_abc_43815_n3947) );
  AND2X2 AND2X2_1752 ( .A(_abc_43815_n3549_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47769_31_), .Y(_abc_43815_n3949) );
  AND2X2 AND2X2_1753 ( .A(_abc_43815_n646_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47769_31_), .Y(_abc_43815_n3951_1) );
  AND2X2 AND2X2_1754 ( .A(_abc_43815_n645_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_43815_n3952) );
  AND2X2 AND2X2_1755 ( .A(_abc_43815_n3521_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_43815_n3955) );
  AND2X2 AND2X2_1756 ( .A(_abc_43815_n3317_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47769_31_), .Y(_abc_43815_n3956) );
  AND2X2 AND2X2_1757 ( .A(_abc_43815_n3958_1), .B(_abc_43815_n3954), .Y(_abc_43815_n3959) );
  AND2X2 AND2X2_1758 ( .A(_abc_43815_n3960), .B(_abc_43815_n3950), .Y(_abc_43815_n3961) );
  AND2X2 AND2X2_1759 ( .A(_abc_43815_n3961), .B(_abc_43815_n671_bF_buf1), .Y(_abc_43815_n3962) );
  AND2X2 AND2X2_176 ( .A(_abc_43815_n931), .B(_abc_43815_n932), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_) );
  AND2X2 AND2X2_1760 ( .A(_abc_43815_n3509), .B(_abc_43815_n3964), .Y(_abc_43815_n3965) );
  AND2X2 AND2X2_1761 ( .A(_abc_43815_n3549_bF_buf2), .B(_abc_43815_n3967), .Y(_abc_43815_n3968) );
  AND2X2 AND2X2_1762 ( .A(_abc_43815_n3968), .B(_auto_iopadmap_cc_313_execute_47809), .Y(_abc_43815_n3969) );
  AND2X2 AND2X2_1763 ( .A(_abc_43815_n3970), .B(_abc_43815_n3966_1), .Y(mem_we_o_FF_INPUT) );
  AND2X2 AND2X2_1764 ( .A(_abc_43815_n3972), .B(state_q_5_), .Y(_abc_43815_n3973_1) );
  AND2X2 AND2X2_1765 ( .A(_auto_iopadmap_cc_313_execute_47807), .B(mem_stall_i), .Y(_abc_43815_n3974) );
  AND2X2 AND2X2_1766 ( .A(_abc_43815_n682), .B(_abc_43815_n3977), .Y(_abc_43815_n3978_1) );
  AND2X2 AND2X2_1767 ( .A(_abc_43815_n3980), .B(_auto_iopadmap_cc_313_execute_47767), .Y(_abc_43815_n3981) );
  AND2X2 AND2X2_1768 ( .A(state_q_3_bF_buf1), .B(next_pc_r_0_), .Y(_abc_43815_n3984) );
  AND2X2 AND2X2_1769 ( .A(_abc_43815_n3985_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47730_0_), .Y(_abc_43815_n3986) );
  AND2X2 AND2X2_177 ( .A(_abc_43815_n692_bF_buf3), .B(\mem_dat_i[24] ), .Y(_abc_43815_n934_1) );
  AND2X2 AND2X2_1770 ( .A(state_q_3_bF_buf0), .B(next_pc_r_1_), .Y(_abc_43815_n3988) );
  AND2X2 AND2X2_1771 ( .A(_abc_43815_n3985_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47730_1_), .Y(_abc_43815_n3989) );
  AND2X2 AND2X2_1772 ( .A(alu_op_r_2_), .B(REGFILE_SIM_reg_bank_reg_ra_o_2_), .Y(_abc_43815_n3992) );
  AND2X2 AND2X2_1773 ( .A(_abc_43815_n3993), .B(_abc_43815_n1217), .Y(_abc_43815_n3994) );
  AND2X2 AND2X2_1774 ( .A(_abc_43815_n3991), .B(_abc_43815_n3994), .Y(_abc_43815_n3995_1) );
  AND2X2 AND2X2_1775 ( .A(_abc_43815_n3996), .B(_abc_43815_n3997), .Y(_abc_43815_n3998) );
  AND2X2 AND2X2_1776 ( .A(_abc_43815_n679_1), .B(_abc_43815_n3998), .Y(_abc_43815_n3999) );
  AND2X2 AND2X2_1777 ( .A(_abc_43815_n678), .B(_auto_iopadmap_cc_313_execute_47730_2_), .Y(_abc_43815_n4000) );
  AND2X2 AND2X2_1778 ( .A(_abc_43815_n4001), .B(state_q_5_), .Y(_abc_43815_n4002_1) );
  AND2X2 AND2X2_1779 ( .A(_abc_43815_n3968), .B(_auto_iopadmap_cc_313_execute_47730_2_), .Y(_abc_43815_n4003) );
  AND2X2 AND2X2_178 ( .A(_abc_43815_n935), .B(_abc_43815_n686_1_bF_buf0), .Y(_abc_43815_n936) );
  AND2X2 AND2X2_1780 ( .A(state_q_3_bF_buf5), .B(pc_q_2_), .Y(_abc_43815_n4004) );
  AND2X2 AND2X2_1781 ( .A(_abc_43815_n3985_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47730_3_), .Y(_abc_43815_n4007) );
  AND2X2 AND2X2_1782 ( .A(state_q_3_bF_buf4), .B(pc_q_3_), .Y(_abc_43815_n4008_1) );
  AND2X2 AND2X2_1783 ( .A(alu_op_r_3_), .B(REGFILE_SIM_reg_bank_reg_ra_o_3_), .Y(_abc_43815_n4010) );
  AND2X2 AND2X2_1784 ( .A(_abc_43815_n4011), .B(_abc_43815_n1219), .Y(_abc_43815_n4012) );
  AND2X2 AND2X2_1785 ( .A(_abc_43815_n4016), .B(_abc_43815_n4013), .Y(_abc_43815_n4017) );
  AND2X2 AND2X2_1786 ( .A(_abc_43815_n680_1_bF_buf0), .B(_abc_43815_n4017), .Y(_abc_43815_n4018) );
  AND2X2 AND2X2_1787 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_4_), .B(int32_r_4_), .Y(_abc_43815_n4021) );
  AND2X2 AND2X2_1788 ( .A(_abc_43815_n4022_1), .B(_abc_43815_n1228), .Y(_abc_43815_n4023) );
  AND2X2 AND2X2_1789 ( .A(_abc_43815_n4009), .B(_abc_43815_n1219), .Y(_abc_43815_n4024) );
  AND2X2 AND2X2_179 ( .A(_abc_43815_n937_1), .B(_abc_43815_n938), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_) );
  AND2X2 AND2X2_1790 ( .A(_abc_43815_n4025), .B(_abc_43815_n4023), .Y(_abc_43815_n4026) );
  AND2X2 AND2X2_1791 ( .A(_abc_43815_n4028), .B(_abc_43815_n679_1), .Y(_abc_43815_n4029_1) );
  AND2X2 AND2X2_1792 ( .A(_abc_43815_n4029_1), .B(_abc_43815_n4027), .Y(_abc_43815_n4030) );
  AND2X2 AND2X2_1793 ( .A(_abc_43815_n678), .B(_auto_iopadmap_cc_313_execute_47730_4_), .Y(_abc_43815_n4031) );
  AND2X2 AND2X2_1794 ( .A(_abc_43815_n4032), .B(state_q_5_), .Y(_abc_43815_n4033) );
  AND2X2 AND2X2_1795 ( .A(_abc_43815_n3968), .B(_auto_iopadmap_cc_313_execute_47730_4_), .Y(_abc_43815_n4034_1) );
  AND2X2 AND2X2_1796 ( .A(state_q_3_bF_buf3), .B(pc_q_4_), .Y(_abc_43815_n4035) );
  AND2X2 AND2X2_1797 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_5_), .B(int32_r_5_), .Y(_abc_43815_n4039) );
  AND2X2 AND2X2_1798 ( .A(_abc_43815_n4040), .B(_abc_43815_n1234), .Y(_abc_43815_n4041_1) );
  AND2X2 AND2X2_1799 ( .A(_abc_43815_n4038), .B(_abc_43815_n4042), .Y(_abc_43815_n4043) );
  AND2X2 AND2X2_18 ( .A(_abc_43815_n644), .B(_abc_43815_n636), .Y(_abc_43815_n645_1) );
  AND2X2 AND2X2_180 ( .A(_abc_43815_n692_bF_buf2), .B(\mem_dat_i[25] ), .Y(_abc_43815_n940) );
  AND2X2 AND2X2_1800 ( .A(_abc_43815_n4044), .B(_abc_43815_n4041_1), .Y(_abc_43815_n4045) );
  AND2X2 AND2X2_1801 ( .A(_abc_43815_n4046), .B(_abc_43815_n680_1_bF_buf4), .Y(_abc_43815_n4047) );
  AND2X2 AND2X2_1802 ( .A(state_q_3_bF_buf2), .B(pc_q_5_), .Y(_abc_43815_n4048) );
  AND2X2 AND2X2_1803 ( .A(_abc_43815_n3985_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47730_5_), .Y(_abc_43815_n4049) );
  AND2X2 AND2X2_1804 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_6_), .B(alu_op_r_4_), .Y(_abc_43815_n4052) );
  AND2X2 AND2X2_1805 ( .A(_abc_43815_n4053), .B(_abc_43815_n1233_1), .Y(_abc_43815_n4054) );
  AND2X2 AND2X2_1806 ( .A(_abc_43815_n4038), .B(_abc_43815_n1234), .Y(_abc_43815_n4055_1) );
  AND2X2 AND2X2_1807 ( .A(_abc_43815_n4056), .B(_abc_43815_n4054), .Y(_abc_43815_n4058) );
  AND2X2 AND2X2_1808 ( .A(_abc_43815_n4059), .B(_abc_43815_n4057), .Y(_abc_43815_n4060) );
  AND2X2 AND2X2_1809 ( .A(_abc_43815_n4060), .B(_abc_43815_n680_1_bF_buf3), .Y(_abc_43815_n4061) );
  AND2X2 AND2X2_181 ( .A(_abc_43815_n941), .B(_abc_43815_n686_1_bF_buf4), .Y(_abc_43815_n942) );
  AND2X2 AND2X2_1810 ( .A(state_q_3_bF_buf1), .B(pc_q_6_), .Y(_abc_43815_n4062_1) );
  AND2X2 AND2X2_1811 ( .A(_abc_43815_n3985_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47730_6_), .Y(_abc_43815_n4063) );
  AND2X2 AND2X2_1812 ( .A(_abc_43815_n4059), .B(_abc_43815_n4053), .Y(_abc_43815_n4066) );
  AND2X2 AND2X2_1813 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_7_), .B(alu_op_r_5_), .Y(_abc_43815_n4067) );
  AND2X2 AND2X2_1814 ( .A(_abc_43815_n4068_1), .B(_abc_43815_n1230_1), .Y(_abc_43815_n4069) );
  AND2X2 AND2X2_1815 ( .A(_abc_43815_n4073), .B(_abc_43815_n4071), .Y(_abc_43815_n4074) );
  AND2X2 AND2X2_1816 ( .A(_abc_43815_n4074), .B(_abc_43815_n680_1_bF_buf2), .Y(_abc_43815_n4075_1) );
  AND2X2 AND2X2_1817 ( .A(state_q_3_bF_buf0), .B(pc_q_7_), .Y(_abc_43815_n4076) );
  AND2X2 AND2X2_1818 ( .A(_abc_43815_n3985_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47730_7_), .Y(_abc_43815_n4077) );
  AND2X2 AND2X2_1819 ( .A(_abc_43815_n1198), .B(_abc_43815_n1108_1), .Y(_abc_43815_n4080) );
  AND2X2 AND2X2_182 ( .A(_abc_43815_n943), .B(_abc_43815_n944), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_) );
  AND2X2 AND2X2_1820 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_8_), .B(alu_op_r_6_), .Y(_abc_43815_n4081) );
  AND2X2 AND2X2_1821 ( .A(_abc_43815_n4053), .B(_abc_43815_n4068_1), .Y(_abc_43815_n4084) );
  AND2X2 AND2X2_1822 ( .A(_abc_43815_n4086), .B(_abc_43815_n1230_1), .Y(_abc_43815_n4087) );
  AND2X2 AND2X2_1823 ( .A(_abc_43815_n4087), .B(_abc_43815_n4083), .Y(_abc_43815_n4089_1) );
  AND2X2 AND2X2_1824 ( .A(_abc_43815_n4090), .B(_abc_43815_n4088), .Y(_abc_43815_n4091) );
  AND2X2 AND2X2_1825 ( .A(_abc_43815_n4091), .B(_abc_43815_n680_1_bF_buf1), .Y(_abc_43815_n4092) );
  AND2X2 AND2X2_1826 ( .A(state_q_3_bF_buf5), .B(pc_q_8_), .Y(_abc_43815_n4093) );
  AND2X2 AND2X2_1827 ( .A(_abc_43815_n3985_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47730_8_), .Y(_abc_43815_n4094_1) );
  AND2X2 AND2X2_1828 ( .A(_abc_43815_n4090), .B(_abc_43815_n4097), .Y(_abc_43815_n4098) );
  AND2X2 AND2X2_1829 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_9_), .B(alu_op_r_7_), .Y(_abc_43815_n4099) );
  AND2X2 AND2X2_183 ( .A(_abc_43815_n692_bF_buf1), .B(\mem_dat_i[26] ), .Y(_abc_43815_n946) );
  AND2X2 AND2X2_1830 ( .A(_abc_43815_n4100), .B(_abc_43815_n1212), .Y(_abc_43815_n4101_1) );
  AND2X2 AND2X2_1831 ( .A(_abc_43815_n4105), .B(_abc_43815_n4103), .Y(_abc_43815_n4106) );
  AND2X2 AND2X2_1832 ( .A(_abc_43815_n4106), .B(_abc_43815_n680_1_bF_buf0), .Y(_abc_43815_n4107) );
  AND2X2 AND2X2_1833 ( .A(state_q_3_bF_buf4), .B(pc_q_9_), .Y(_abc_43815_n4108) );
  AND2X2 AND2X2_1834 ( .A(_abc_43815_n3985_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47730_9_), .Y(_abc_43815_n4109) );
  AND2X2 AND2X2_1835 ( .A(_abc_43815_n4083), .B(_abc_43815_n4101_1), .Y(_abc_43815_n4112_1) );
  AND2X2 AND2X2_1836 ( .A(_abc_43815_n4087), .B(_abc_43815_n4112_1), .Y(_abc_43815_n4113) );
  AND2X2 AND2X2_1837 ( .A(_abc_43815_n4097), .B(_abc_43815_n4100), .Y(_abc_43815_n4114) );
  AND2X2 AND2X2_1838 ( .A(_abc_43815_n1201), .B(_abc_43815_n1199), .Y(_abc_43815_n4118) );
  AND2X2 AND2X2_1839 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_10_), .B(int32_r_10_), .Y(_abc_43815_n4119_1) );
  AND2X2 AND2X2_184 ( .A(_abc_43815_n947), .B(_abc_43815_n686_1_bF_buf3), .Y(_abc_43815_n948) );
  AND2X2 AND2X2_1840 ( .A(_abc_43815_n4117), .B(_abc_43815_n4121), .Y(_abc_43815_n4123) );
  AND2X2 AND2X2_1841 ( .A(_abc_43815_n4124_1), .B(_abc_43815_n4122), .Y(_abc_43815_n4125) );
  AND2X2 AND2X2_1842 ( .A(_abc_43815_n4125), .B(_abc_43815_n680_1_bF_buf4), .Y(_abc_43815_n4126) );
  AND2X2 AND2X2_1843 ( .A(state_q_3_bF_buf3), .B(pc_q_10_), .Y(_abc_43815_n4127) );
  AND2X2 AND2X2_1844 ( .A(_abc_43815_n3985_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47730_10_), .Y(_abc_43815_n4128) );
  AND2X2 AND2X2_1845 ( .A(_abc_43815_n4124_1), .B(_abc_43815_n4131_1), .Y(_abc_43815_n4132) );
  AND2X2 AND2X2_1846 ( .A(_abc_43815_n652), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_43815_n4133) );
  AND2X2 AND2X2_1847 ( .A(_abc_43815_n3509), .B(opcode_q_21_), .Y(_abc_43815_n4134) );
  AND2X2 AND2X2_1848 ( .A(_abc_43815_n4135), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_43815_n4136) );
  AND2X2 AND2X2_1849 ( .A(_abc_43815_n4137), .B(_abc_43815_n4138_1), .Y(_abc_43815_n4139) );
  AND2X2 AND2X2_185 ( .A(_abc_43815_n949), .B(_abc_43815_n950), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_) );
  AND2X2 AND2X2_1850 ( .A(_abc_43815_n4143), .B(_abc_43815_n4141), .Y(_abc_43815_n4144) );
  AND2X2 AND2X2_1851 ( .A(_abc_43815_n4144), .B(_abc_43815_n680_1_bF_buf3), .Y(_abc_43815_n4145_1) );
  AND2X2 AND2X2_1852 ( .A(state_q_3_bF_buf2), .B(pc_q_11_), .Y(_abc_43815_n4146) );
  AND2X2 AND2X2_1853 ( .A(_abc_43815_n3985_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47730_11_), .Y(_abc_43815_n4147) );
  AND2X2 AND2X2_1854 ( .A(_abc_43815_n652), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_43815_n4150_1) );
  AND2X2 AND2X2_1855 ( .A(_abc_43815_n3509), .B(opcode_q_22_), .Y(_abc_43815_n4151) );
  AND2X2 AND2X2_1856 ( .A(_abc_43815_n4152), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_43815_n4153) );
  AND2X2 AND2X2_1857 ( .A(_abc_43815_n4154), .B(_abc_43815_n4155), .Y(_abc_43815_n4156) );
  AND2X2 AND2X2_1858 ( .A(_abc_43815_n4139), .B(_abc_43815_n4121), .Y(_abc_43815_n4157_1) );
  AND2X2 AND2X2_1859 ( .A(_abc_43815_n4157_1), .B(_abc_43815_n4112_1), .Y(_abc_43815_n4158_1) );
  AND2X2 AND2X2_186 ( .A(_abc_43815_n692_bF_buf0), .B(\mem_dat_i[27] ), .Y(_abc_43815_n952) );
  AND2X2 AND2X2_1860 ( .A(_abc_43815_n4087), .B(_abc_43815_n4158_1), .Y(_abc_43815_n4159) );
  AND2X2 AND2X2_1861 ( .A(_abc_43815_n4138_1), .B(_abc_43815_n4119_1), .Y(_abc_43815_n4160) );
  AND2X2 AND2X2_1862 ( .A(_abc_43815_n4157_1), .B(_abc_43815_n4116), .Y(_abc_43815_n4162_1) );
  AND2X2 AND2X2_1863 ( .A(_abc_43815_n4164_1), .B(_abc_43815_n4156), .Y(_abc_43815_n4166_1) );
  AND2X2 AND2X2_1864 ( .A(_abc_43815_n4167_1), .B(_abc_43815_n4165_1), .Y(_abc_43815_n4168) );
  AND2X2 AND2X2_1865 ( .A(_abc_43815_n4168), .B(_abc_43815_n680_1_bF_buf2), .Y(_abc_43815_n4169) );
  AND2X2 AND2X2_1866 ( .A(state_q_3_bF_buf1), .B(pc_q_12_), .Y(_abc_43815_n4170) );
  AND2X2 AND2X2_1867 ( .A(_abc_43815_n3985_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47730_12_), .Y(_abc_43815_n4171) );
  AND2X2 AND2X2_1868 ( .A(_abc_43815_n652), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_43815_n4174) );
  AND2X2 AND2X2_1869 ( .A(_abc_43815_n3509), .B(opcode_q_23_), .Y(_abc_43815_n4175) );
  AND2X2 AND2X2_187 ( .A(_abc_43815_n953), .B(_abc_43815_n686_1_bF_buf2), .Y(_abc_43815_n954) );
  AND2X2 AND2X2_1870 ( .A(_abc_43815_n4176), .B(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_43815_n4177) );
  AND2X2 AND2X2_1871 ( .A(_abc_43815_n4178), .B(_abc_43815_n4179), .Y(_abc_43815_n4180) );
  AND2X2 AND2X2_1872 ( .A(_abc_43815_n4156), .B(_abc_43815_n4180), .Y(_abc_43815_n4183) );
  AND2X2 AND2X2_1873 ( .A(_abc_43815_n4164_1), .B(_abc_43815_n4183), .Y(_abc_43815_n4184) );
  AND2X2 AND2X2_1874 ( .A(_abc_43815_n4180), .B(_abc_43815_n4153), .Y(_abc_43815_n4186) );
  AND2X2 AND2X2_1875 ( .A(_abc_43815_n4187), .B(_abc_43815_n680_1_bF_buf1), .Y(_abc_43815_n4188) );
  AND2X2 AND2X2_1876 ( .A(_abc_43815_n4185), .B(_abc_43815_n4188), .Y(_abc_43815_n4189) );
  AND2X2 AND2X2_1877 ( .A(_abc_43815_n4189), .B(_abc_43815_n4182), .Y(_abc_43815_n4190) );
  AND2X2 AND2X2_1878 ( .A(state_q_3_bF_buf0), .B(pc_q_13_), .Y(_abc_43815_n4191) );
  AND2X2 AND2X2_1879 ( .A(_abc_43815_n3985_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47730_13_), .Y(_abc_43815_n4192) );
  AND2X2 AND2X2_188 ( .A(_abc_43815_n955_1), .B(_abc_43815_n956_1), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_) );
  AND2X2 AND2X2_1880 ( .A(_abc_43815_n4187), .B(_abc_43815_n4178), .Y(_abc_43815_n4195) );
  AND2X2 AND2X2_1881 ( .A(_abc_43815_n4185), .B(_abc_43815_n4195), .Y(_abc_43815_n4196) );
  AND2X2 AND2X2_1882 ( .A(_abc_43815_n652), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_43815_n4198) );
  AND2X2 AND2X2_1883 ( .A(_abc_43815_n3509), .B(opcode_q_24_), .Y(_abc_43815_n4199) );
  AND2X2 AND2X2_1884 ( .A(_abc_43815_n4200), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_43815_n4201) );
  AND2X2 AND2X2_1885 ( .A(_abc_43815_n4202), .B(_abc_43815_n4203), .Y(_abc_43815_n4204) );
  AND2X2 AND2X2_1886 ( .A(_abc_43815_n4197), .B(_abc_43815_n4204), .Y(_abc_43815_n4205) );
  AND2X2 AND2X2_1887 ( .A(_abc_43815_n4207), .B(_abc_43815_n680_1_bF_buf0), .Y(_abc_43815_n4208) );
  AND2X2 AND2X2_1888 ( .A(_abc_43815_n4208), .B(_abc_43815_n4206), .Y(_abc_43815_n4209) );
  AND2X2 AND2X2_1889 ( .A(state_q_3_bF_buf5), .B(pc_q_14_), .Y(_abc_43815_n4210) );
  AND2X2 AND2X2_189 ( .A(_abc_43815_n692_bF_buf3), .B(\mem_dat_i[28] ), .Y(_abc_43815_n958) );
  AND2X2 AND2X2_1890 ( .A(_abc_43815_n3985_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47730_14_), .Y(_abc_43815_n4211) );
  AND2X2 AND2X2_1891 ( .A(_abc_43815_n4206), .B(_abc_43815_n4202), .Y(_abc_43815_n4214) );
  AND2X2 AND2X2_1892 ( .A(_abc_43815_n652), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3), .Y(_abc_43815_n4215) );
  AND2X2 AND2X2_1893 ( .A(_abc_43815_n3509), .B(opcode_q_25_), .Y(_abc_43815_n4216) );
  AND2X2 AND2X2_1894 ( .A(_abc_43815_n4217_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_43815_n4218) );
  AND2X2 AND2X2_1895 ( .A(_abc_43815_n4220), .B(_abc_43815_n1205_1), .Y(_abc_43815_n4221) );
  AND2X2 AND2X2_1896 ( .A(_abc_43815_n4222), .B(_abc_43815_n4219), .Y(_abc_43815_n4223) );
  AND2X2 AND2X2_1897 ( .A(_abc_43815_n4227), .B(_abc_43815_n4225), .Y(_abc_43815_n4228) );
  AND2X2 AND2X2_1898 ( .A(_abc_43815_n4228), .B(_abc_43815_n680_1_bF_buf4), .Y(_abc_43815_n4229) );
  AND2X2 AND2X2_1899 ( .A(state_q_3_bF_buf4), .B(pc_q_15_), .Y(_abc_43815_n4230) );
  AND2X2 AND2X2_19 ( .A(inst_r_1_), .B(inst_r_0_), .Y(_abc_43815_n647_1) );
  AND2X2 AND2X2_190 ( .A(_abc_43815_n959), .B(_abc_43815_n686_1_bF_buf1), .Y(_abc_43815_n960) );
  AND2X2 AND2X2_1900 ( .A(_abc_43815_n3985_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47730_15_), .Y(_abc_43815_n4231) );
  AND2X2 AND2X2_1901 ( .A(_abc_43815_n4223), .B(_abc_43815_n4204), .Y(_abc_43815_n4234) );
  AND2X2 AND2X2_1902 ( .A(_abc_43815_n4222), .B(_abc_43815_n4201), .Y(_abc_43815_n4237) );
  AND2X2 AND2X2_1903 ( .A(_abc_43815_n4236), .B(_abc_43815_n4239), .Y(_abc_43815_n4240) );
  AND2X2 AND2X2_1904 ( .A(_abc_43815_n4234), .B(_abc_43815_n4183), .Y(_abc_43815_n4242) );
  AND2X2 AND2X2_1905 ( .A(_abc_43815_n4164_1), .B(_abc_43815_n4242), .Y(_abc_43815_n4243) );
  AND2X2 AND2X2_1906 ( .A(_abc_43815_n4217_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_43815_n4245) );
  AND2X2 AND2X2_1907 ( .A(_abc_43815_n4246), .B(_abc_43815_n4247), .Y(_abc_43815_n4248) );
  AND2X2 AND2X2_1908 ( .A(_abc_43815_n4244), .B(_abc_43815_n4248), .Y(_abc_43815_n4250) );
  AND2X2 AND2X2_1909 ( .A(_abc_43815_n4251), .B(_abc_43815_n4249), .Y(_abc_43815_n4252) );
  AND2X2 AND2X2_191 ( .A(_abc_43815_n961), .B(_abc_43815_n962), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_) );
  AND2X2 AND2X2_1910 ( .A(_abc_43815_n4252), .B(_abc_43815_n680_1_bF_buf3), .Y(_abc_43815_n4253) );
  AND2X2 AND2X2_1911 ( .A(state_q_3_bF_buf3), .B(pc_q_16_), .Y(_abc_43815_n4254) );
  AND2X2 AND2X2_1912 ( .A(_abc_43815_n3985_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47730_16_), .Y(_abc_43815_n4255) );
  AND2X2 AND2X2_1913 ( .A(_abc_43815_n4251), .B(_abc_43815_n4246), .Y(_abc_43815_n4258) );
  AND2X2 AND2X2_1914 ( .A(_abc_43815_n4217_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_43815_n4259) );
  AND2X2 AND2X2_1915 ( .A(_abc_43815_n4260), .B(_abc_43815_n4261), .Y(_abc_43815_n4262) );
  AND2X2 AND2X2_1916 ( .A(_abc_43815_n4266), .B(_abc_43815_n4264), .Y(_abc_43815_n4267) );
  AND2X2 AND2X2_1917 ( .A(_abc_43815_n4267), .B(_abc_43815_n680_1_bF_buf2), .Y(_abc_43815_n4268) );
  AND2X2 AND2X2_1918 ( .A(state_q_3_bF_buf2), .B(pc_q_17_), .Y(_abc_43815_n4269) );
  AND2X2 AND2X2_1919 ( .A(_abc_43815_n3985_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47730_17_), .Y(_abc_43815_n4270) );
  AND2X2 AND2X2_192 ( .A(_abc_43815_n692_bF_buf2), .B(\mem_dat_i[29] ), .Y(_abc_43815_n964_1) );
  AND2X2 AND2X2_1920 ( .A(_abc_43815_n4217_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_43815_n4273) );
  AND2X2 AND2X2_1921 ( .A(_abc_43815_n4274), .B(_abc_43815_n4275), .Y(_abc_43815_n4276) );
  AND2X2 AND2X2_1922 ( .A(_abc_43815_n4246), .B(_abc_43815_n4260), .Y(_abc_43815_n4277) );
  AND2X2 AND2X2_1923 ( .A(_abc_43815_n4248), .B(_abc_43815_n4262), .Y(_abc_43815_n4279) );
  AND2X2 AND2X2_1924 ( .A(_abc_43815_n4244), .B(_abc_43815_n4279), .Y(_abc_43815_n4280) );
  AND2X2 AND2X2_1925 ( .A(_abc_43815_n4281), .B(_abc_43815_n4276), .Y(_abc_43815_n4283) );
  AND2X2 AND2X2_1926 ( .A(_abc_43815_n4284), .B(_abc_43815_n4282), .Y(_abc_43815_n4285) );
  AND2X2 AND2X2_1927 ( .A(_abc_43815_n4285), .B(_abc_43815_n680_1_bF_buf1), .Y(_abc_43815_n4286) );
  AND2X2 AND2X2_1928 ( .A(state_q_3_bF_buf1), .B(pc_q_18_), .Y(_abc_43815_n4287) );
  AND2X2 AND2X2_1929 ( .A(_abc_43815_n3985_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47730_18_), .Y(_abc_43815_n4288) );
  AND2X2 AND2X2_193 ( .A(_abc_43815_n965), .B(_abc_43815_n686_1_bF_buf0), .Y(_abc_43815_n966) );
  AND2X2 AND2X2_1930 ( .A(_abc_43815_n4284), .B(_abc_43815_n4274), .Y(_abc_43815_n4291) );
  AND2X2 AND2X2_1931 ( .A(_abc_43815_n4217_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_43815_n4292) );
  AND2X2 AND2X2_1932 ( .A(_abc_43815_n4293), .B(_abc_43815_n4294), .Y(_abc_43815_n4295) );
  AND2X2 AND2X2_1933 ( .A(_abc_43815_n4299), .B(_abc_43815_n4297), .Y(_abc_43815_n4300) );
  AND2X2 AND2X2_1934 ( .A(_abc_43815_n4300), .B(_abc_43815_n680_1_bF_buf0), .Y(_abc_43815_n4301) );
  AND2X2 AND2X2_1935 ( .A(state_q_3_bF_buf0), .B(pc_q_19_), .Y(_abc_43815_n4302) );
  AND2X2 AND2X2_1936 ( .A(_abc_43815_n3985_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47730_19_), .Y(_abc_43815_n4303) );
  AND2X2 AND2X2_1937 ( .A(_abc_43815_n4276), .B(_abc_43815_n4295), .Y(_abc_43815_n4306) );
  AND2X2 AND2X2_1938 ( .A(_abc_43815_n4279), .B(_abc_43815_n4306), .Y(_abc_43815_n4307) );
  AND2X2 AND2X2_1939 ( .A(_abc_43815_n4244), .B(_abc_43815_n4307), .Y(_abc_43815_n4308) );
  AND2X2 AND2X2_194 ( .A(_abc_43815_n967), .B(_abc_43815_n968), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_) );
  AND2X2 AND2X2_1940 ( .A(_abc_43815_n4306), .B(_abc_43815_n4278), .Y(_abc_43815_n4309) );
  AND2X2 AND2X2_1941 ( .A(_abc_43815_n4274), .B(_abc_43815_n4293), .Y(_abc_43815_n4311) );
  AND2X2 AND2X2_1942 ( .A(_abc_43815_n4310), .B(_abc_43815_n4311), .Y(_abc_43815_n4312) );
  AND2X2 AND2X2_1943 ( .A(_abc_43815_n4217_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_43815_n4315) );
  AND2X2 AND2X2_1944 ( .A(_abc_43815_n4316), .B(_abc_43815_n4317), .Y(_abc_43815_n4318) );
  AND2X2 AND2X2_1945 ( .A(_abc_43815_n4314), .B(_abc_43815_n4318), .Y(_abc_43815_n4320) );
  AND2X2 AND2X2_1946 ( .A(_abc_43815_n4321), .B(_abc_43815_n4319), .Y(_abc_43815_n4322) );
  AND2X2 AND2X2_1947 ( .A(_abc_43815_n4322), .B(_abc_43815_n680_1_bF_buf4), .Y(_abc_43815_n4323) );
  AND2X2 AND2X2_1948 ( .A(state_q_3_bF_buf5), .B(pc_q_20_), .Y(_abc_43815_n4324) );
  AND2X2 AND2X2_1949 ( .A(_abc_43815_n3985_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47730_20_), .Y(_abc_43815_n4325) );
  AND2X2 AND2X2_195 ( .A(_abc_43815_n692_bF_buf1), .B(\mem_dat_i[30] ), .Y(_abc_43815_n970) );
  AND2X2 AND2X2_1950 ( .A(_abc_43815_n4321), .B(_abc_43815_n4316), .Y(_abc_43815_n4328) );
  AND2X2 AND2X2_1951 ( .A(_abc_43815_n4217_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_43815_n4329) );
  AND2X2 AND2X2_1952 ( .A(_abc_43815_n4330), .B(_abc_43815_n4331), .Y(_abc_43815_n4332) );
  AND2X2 AND2X2_1953 ( .A(_abc_43815_n4336), .B(_abc_43815_n4334), .Y(_abc_43815_n4337) );
  AND2X2 AND2X2_1954 ( .A(_abc_43815_n4337), .B(_abc_43815_n680_1_bF_buf3), .Y(_abc_43815_n4338) );
  AND2X2 AND2X2_1955 ( .A(state_q_3_bF_buf4), .B(pc_q_21_), .Y(_abc_43815_n4339) );
  AND2X2 AND2X2_1956 ( .A(_abc_43815_n3985_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47730_21_), .Y(_abc_43815_n4340) );
  AND2X2 AND2X2_1957 ( .A(_abc_43815_n4318), .B(_abc_43815_n4332), .Y(_abc_43815_n4344) );
  AND2X2 AND2X2_1958 ( .A(_abc_43815_n4314), .B(_abc_43815_n4344), .Y(_abc_43815_n4345) );
  AND2X2 AND2X2_1959 ( .A(_abc_43815_n4217_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_43815_n4347) );
  AND2X2 AND2X2_196 ( .A(_abc_43815_n971), .B(_abc_43815_n686_1_bF_buf4), .Y(_abc_43815_n972) );
  AND2X2 AND2X2_1960 ( .A(_abc_43815_n4348), .B(_abc_43815_n4349), .Y(_abc_43815_n4350) );
  AND2X2 AND2X2_1961 ( .A(_abc_43815_n4346), .B(_abc_43815_n4350), .Y(_abc_43815_n4352) );
  AND2X2 AND2X2_1962 ( .A(_abc_43815_n4353), .B(_abc_43815_n4351), .Y(_abc_43815_n4354) );
  AND2X2 AND2X2_1963 ( .A(_abc_43815_n4354), .B(_abc_43815_n680_1_bF_buf2), .Y(_abc_43815_n4355) );
  AND2X2 AND2X2_1964 ( .A(state_q_3_bF_buf3), .B(pc_q_22_), .Y(_abc_43815_n4356) );
  AND2X2 AND2X2_1965 ( .A(_abc_43815_n3985_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47730_22_), .Y(_abc_43815_n4357) );
  AND2X2 AND2X2_1966 ( .A(_abc_43815_n4353), .B(_abc_43815_n4348), .Y(_abc_43815_n4360) );
  AND2X2 AND2X2_1967 ( .A(_abc_43815_n4217_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_43815_n4362) );
  AND2X2 AND2X2_1968 ( .A(_abc_43815_n4363), .B(_abc_43815_n4364), .Y(_abc_43815_n4365) );
  AND2X2 AND2X2_1969 ( .A(_abc_43815_n4368), .B(_abc_43815_n680_1_bF_buf1), .Y(_abc_43815_n4369) );
  AND2X2 AND2X2_197 ( .A(_abc_43815_n973), .B(_abc_43815_n974), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_) );
  AND2X2 AND2X2_1970 ( .A(_abc_43815_n4369), .B(_abc_43815_n4366), .Y(_abc_43815_n4370) );
  AND2X2 AND2X2_1971 ( .A(state_q_3_bF_buf2), .B(pc_q_23_), .Y(_abc_43815_n4371) );
  AND2X2 AND2X2_1972 ( .A(_abc_43815_n3985_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47730_23_), .Y(_abc_43815_n4372) );
  AND2X2 AND2X2_1973 ( .A(_abc_43815_n4350), .B(_abc_43815_n4365), .Y(_abc_43815_n4375) );
  AND2X2 AND2X2_1974 ( .A(_abc_43815_n4375), .B(_abc_43815_n4343), .Y(_abc_43815_n4376) );
  AND2X2 AND2X2_1975 ( .A(_abc_43815_n4348), .B(_abc_43815_n4363), .Y(_abc_43815_n4378) );
  AND2X2 AND2X2_1976 ( .A(_abc_43815_n4377), .B(_abc_43815_n4378), .Y(_abc_43815_n4379) );
  AND2X2 AND2X2_1977 ( .A(_abc_43815_n4344), .B(_abc_43815_n4375), .Y(_abc_43815_n4381) );
  AND2X2 AND2X2_1978 ( .A(_abc_43815_n4314), .B(_abc_43815_n4381), .Y(_abc_43815_n4382) );
  AND2X2 AND2X2_1979 ( .A(_abc_43815_n4217_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_43815_n4384) );
  AND2X2 AND2X2_198 ( .A(_abc_43815_n692_bF_buf0), .B(\mem_dat_i[31] ), .Y(_abc_43815_n976) );
  AND2X2 AND2X2_1980 ( .A(_abc_43815_n4385), .B(_abc_43815_n4386), .Y(_abc_43815_n4387) );
  AND2X2 AND2X2_1981 ( .A(_abc_43815_n4383), .B(_abc_43815_n4387), .Y(_abc_43815_n4389) );
  AND2X2 AND2X2_1982 ( .A(_abc_43815_n4390), .B(_abc_43815_n4388), .Y(_abc_43815_n4391) );
  AND2X2 AND2X2_1983 ( .A(_abc_43815_n4391), .B(_abc_43815_n680_1_bF_buf0), .Y(_abc_43815_n4392) );
  AND2X2 AND2X2_1984 ( .A(state_q_3_bF_buf1), .B(pc_q_24_), .Y(_abc_43815_n4393) );
  AND2X2 AND2X2_1985 ( .A(_abc_43815_n3985_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47730_24_), .Y(_abc_43815_n4394) );
  AND2X2 AND2X2_1986 ( .A(_abc_43815_n4390), .B(_abc_43815_n4385), .Y(_abc_43815_n4397) );
  AND2X2 AND2X2_1987 ( .A(_abc_43815_n4217_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_43815_n4398) );
  AND2X2 AND2X2_1988 ( .A(_abc_43815_n4399), .B(_abc_43815_n4400), .Y(_abc_43815_n4401) );
  AND2X2 AND2X2_1989 ( .A(_abc_43815_n4405), .B(_abc_43815_n4403), .Y(_abc_43815_n4406) );
  AND2X2 AND2X2_199 ( .A(_abc_43815_n977), .B(_abc_43815_n686_1_bF_buf3), .Y(_abc_43815_n978) );
  AND2X2 AND2X2_1990 ( .A(_abc_43815_n4406), .B(_abc_43815_n680_1_bF_buf4), .Y(_abc_43815_n4407) );
  AND2X2 AND2X2_1991 ( .A(state_q_3_bF_buf0), .B(pc_q_25_), .Y(_abc_43815_n4408) );
  AND2X2 AND2X2_1992 ( .A(_abc_43815_n3985_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47730_25_), .Y(_abc_43815_n4409) );
  AND2X2 AND2X2_1993 ( .A(_abc_43815_n4387), .B(_abc_43815_n4401), .Y(_abc_43815_n4412) );
  AND2X2 AND2X2_1994 ( .A(_abc_43815_n4383), .B(_abc_43815_n4412), .Y(_abc_43815_n4413) );
  AND2X2 AND2X2_1995 ( .A(_abc_43815_n4385), .B(_abc_43815_n4399), .Y(_abc_43815_n4414) );
  AND2X2 AND2X2_1996 ( .A(_abc_43815_n4217_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_43815_n4417) );
  AND2X2 AND2X2_1997 ( .A(_abc_43815_n4418), .B(_abc_43815_n4419), .Y(_abc_43815_n4420) );
  AND2X2 AND2X2_1998 ( .A(_abc_43815_n4416), .B(_abc_43815_n4420), .Y(_abc_43815_n4422) );
  AND2X2 AND2X2_1999 ( .A(_abc_43815_n4423), .B(_abc_43815_n4421), .Y(_abc_43815_n4424) );
  AND2X2 AND2X2_2 ( .A(_abc_43815_n618), .B(enable_i_bF_buf7), .Y(_abc_43815_n619) );
  AND2X2 AND2X2_20 ( .A(_abc_43815_n638), .B(_abc_43815_n647_1), .Y(_abc_43815_n648) );
  AND2X2 AND2X2_200 ( .A(_abc_43815_n979), .B(_abc_43815_n980), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_) );
  AND2X2 AND2X2_2000 ( .A(_abc_43815_n4424), .B(_abc_43815_n680_1_bF_buf3), .Y(_abc_43815_n4425) );
  AND2X2 AND2X2_2001 ( .A(state_q_3_bF_buf5), .B(pc_q_26_), .Y(_abc_43815_n4426) );
  AND2X2 AND2X2_2002 ( .A(_abc_43815_n3985_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47730_26_), .Y(_abc_43815_n4427) );
  AND2X2 AND2X2_2003 ( .A(_abc_43815_n4423), .B(_abc_43815_n4418), .Y(_abc_43815_n4430) );
  AND2X2 AND2X2_2004 ( .A(_abc_43815_n4217_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_43815_n4431) );
  AND2X2 AND2X2_2005 ( .A(_abc_43815_n4432), .B(_abc_43815_n4433), .Y(_abc_43815_n4434) );
  AND2X2 AND2X2_2006 ( .A(_abc_43815_n4438), .B(_abc_43815_n4436), .Y(_abc_43815_n4439) );
  AND2X2 AND2X2_2007 ( .A(_abc_43815_n4439), .B(_abc_43815_n680_1_bF_buf2), .Y(_abc_43815_n4440) );
  AND2X2 AND2X2_2008 ( .A(state_q_3_bF_buf4), .B(pc_q_27_), .Y(_abc_43815_n4441) );
  AND2X2 AND2X2_2009 ( .A(_abc_43815_n3985_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_47730_27_), .Y(_abc_43815_n4442) );
  AND2X2 AND2X2_201 ( .A(inst_r_3_), .B(inst_r_2_), .Y(_abc_43815_n983) );
  AND2X2 AND2X2_2010 ( .A(_abc_43815_n4420), .B(_abc_43815_n4434), .Y(_abc_43815_n4447) );
  AND2X2 AND2X2_2011 ( .A(_abc_43815_n4447), .B(_abc_43815_n4415), .Y(_abc_43815_n4451) );
  AND2X2 AND2X2_2012 ( .A(_abc_43815_n4418), .B(_abc_43815_n4432), .Y(_abc_43815_n4453) );
  AND2X2 AND2X2_2013 ( .A(_abc_43815_n4452), .B(_abc_43815_n4453), .Y(_abc_43815_n4454) );
  AND2X2 AND2X2_2014 ( .A(_abc_43815_n4450), .B(_abc_43815_n4454), .Y(_abc_43815_n4455) );
  AND2X2 AND2X2_2015 ( .A(_abc_43815_n4217_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_43815_n4457) );
  AND2X2 AND2X2_2016 ( .A(_abc_43815_n4220), .B(_abc_43815_n4458), .Y(_abc_43815_n4459) );
  AND2X2 AND2X2_2017 ( .A(_abc_43815_n4456), .B(_abc_43815_n4461), .Y(_abc_43815_n4463) );
  AND2X2 AND2X2_2018 ( .A(_abc_43815_n4464), .B(_abc_43815_n4462), .Y(_abc_43815_n4465) );
  AND2X2 AND2X2_2019 ( .A(_abc_43815_n4465), .B(_abc_43815_n680_1_bF_buf1), .Y(_abc_43815_n4466) );
  AND2X2 AND2X2_202 ( .A(_abc_43815_n659), .B(_abc_43815_n983), .Y(_abc_43815_n984) );
  AND2X2 AND2X2_2020 ( .A(state_q_3_bF_buf3), .B(pc_q_28_), .Y(_abc_43815_n4467) );
  AND2X2 AND2X2_2021 ( .A(_abc_43815_n3985_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_47730_28_), .Y(_abc_43815_n4468) );
  AND2X2 AND2X2_2022 ( .A(_abc_43815_n4217_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_43815_n4473) );
  AND2X2 AND2X2_2023 ( .A(_abc_43815_n4220), .B(_abc_43815_n4474), .Y(_abc_43815_n4475) );
  AND2X2 AND2X2_2024 ( .A(_abc_43815_n4479), .B(_abc_43815_n680_1_bF_buf0), .Y(_abc_43815_n4480) );
  AND2X2 AND2X2_2025 ( .A(_abc_43815_n4480), .B(_abc_43815_n4477), .Y(_abc_43815_n4481) );
  AND2X2 AND2X2_2026 ( .A(state_q_3_bF_buf2), .B(pc_q_29_), .Y(_abc_43815_n4482) );
  AND2X2 AND2X2_2027 ( .A(_abc_43815_n3985_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_47730_29_), .Y(_abc_43815_n4483) );
  AND2X2 AND2X2_2028 ( .A(_abc_43815_n4217_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_43815_n4486) );
  AND2X2 AND2X2_2029 ( .A(_abc_43815_n4487), .B(_abc_43815_n4488), .Y(_abc_43815_n4489) );
  AND2X2 AND2X2_203 ( .A(_abc_43815_n626), .B(_abc_43815_n636), .Y(_abc_43815_n985) );
  AND2X2 AND2X2_2030 ( .A(_abc_43815_n4458), .B(_abc_43815_n4474), .Y(_abc_43815_n4490) );
  AND2X2 AND2X2_2031 ( .A(_abc_43815_n4461), .B(_abc_43815_n4478), .Y(_abc_43815_n4492) );
  AND2X2 AND2X2_2032 ( .A(_abc_43815_n4494), .B(_abc_43815_n4491), .Y(_abc_43815_n4495) );
  AND2X2 AND2X2_2033 ( .A(_abc_43815_n4499), .B(_abc_43815_n680_1_bF_buf4), .Y(_abc_43815_n4500) );
  AND2X2 AND2X2_2034 ( .A(_abc_43815_n4500), .B(_abc_43815_n4497), .Y(_abc_43815_n4501) );
  AND2X2 AND2X2_2035 ( .A(state_q_3_bF_buf1), .B(pc_q_30_), .Y(_abc_43815_n4502) );
  AND2X2 AND2X2_2036 ( .A(_abc_43815_n3985_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_47730_30_), .Y(_abc_43815_n4503) );
  AND2X2 AND2X2_2037 ( .A(_abc_43815_n4499), .B(_abc_43815_n4487), .Y(_abc_43815_n4506) );
  AND2X2 AND2X2_2038 ( .A(_abc_43815_n4508), .B(_abc_43815_n4509), .Y(_abc_43815_n4510) );
  AND2X2 AND2X2_2039 ( .A(_abc_43815_n4514), .B(_abc_43815_n4512), .Y(_abc_43815_n4515) );
  AND2X2 AND2X2_204 ( .A(_abc_43815_n985), .B(_abc_43815_n643_1), .Y(_abc_43815_n986) );
  AND2X2 AND2X2_2040 ( .A(_abc_43815_n4515), .B(_abc_43815_n680_1_bF_buf3), .Y(_abc_43815_n4516) );
  AND2X2 AND2X2_2041 ( .A(state_q_3_bF_buf0), .B(pc_q_31_), .Y(_abc_43815_n4517) );
  AND2X2 AND2X2_2042 ( .A(_abc_43815_n3985_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_47730_31_), .Y(_abc_43815_n4518) );
  AND2X2 AND2X2_2043 ( .A(_abc_43815_n634), .B(state_q_0_), .Y(_abc_27555_n4360) );
  AND2X2 AND2X2_2044 ( .A(_abc_43815_n1195), .B(enable_i_bF_buf0), .Y(_abc_43815_n4522) );
  AND2X2 AND2X2_2045 ( .A(_abc_43815_n1692), .B(_abc_43815_n4522), .Y(nmi_q_FF_INPUT) );
  AND2X2 AND2X2_2046 ( .A(_abc_43815_n4524), .B(enable_i_bF_buf7), .Y(fault_o_FF_INPUT) );
  AND2X2 AND2X2_2047 ( .A(REGFILE_SIM_reg_bank_rd_i_3_), .B(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2099_1) );
  AND2X2 AND2X2_2048 ( .A(REGFILE_SIM_reg_bank_rd_i_1_), .B(REGFILE_SIM_reg_bank_rd_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2100) );
  AND2X2 AND2X2_2049 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2099_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2100), .Y(REGFILE_SIM_reg_bank__abc_33898_n2101_1) );
  AND2X2 AND2X2_205 ( .A(_abc_43815_n988), .B(opcode_q_22_), .Y(_abc_43815_n989) );
  AND2X2 AND2X2_2050 ( .A(REGFILE_SIM_reg_bank_rd_i_4_), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2102) );
  AND2X2 AND2X2_2051 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2101_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1) );
  AND2X2 AND2X2_2052 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2106_1) );
  AND2X2 AND2X2_2053 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2107), .B(REGFILE_SIM_reg_bank__abc_33898_n2104), .Y(REGFILE_SIM_reg_bank_reg_r31_0__FF_INPUT) );
  AND2X2 AND2X2_2054 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n2111_1) );
  AND2X2 AND2X2_2055 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2112_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2109_1), .Y(REGFILE_SIM_reg_bank_reg_r31_1__FF_INPUT) );
  AND2X2 AND2X2_2056 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2116) );
  AND2X2 AND2X2_2057 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2117_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2114_1), .Y(REGFILE_SIM_reg_bank_reg_r31_2__FF_INPUT) );
  AND2X2 AND2X2_2058 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2121_1) );
  AND2X2 AND2X2_2059 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2122), .B(REGFILE_SIM_reg_bank__abc_33898_n2119), .Y(REGFILE_SIM_reg_bank_reg_r31_3__FF_INPUT) );
  AND2X2 AND2X2_206 ( .A(inst_r_0_), .B(inst_r_3_), .Y(_abc_43815_n990) );
  AND2X2 AND2X2_2060 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n2126_1) );
  AND2X2 AND2X2_2061 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2127_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2124_1), .Y(REGFILE_SIM_reg_bank_reg_r31_4__FF_INPUT) );
  AND2X2 AND2X2_2062 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2131) );
  AND2X2 AND2X2_2063 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2132_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2129_1), .Y(REGFILE_SIM_reg_bank_reg_r31_5__FF_INPUT) );
  AND2X2 AND2X2_2064 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2136_1) );
  AND2X2 AND2X2_2065 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2137), .B(REGFILE_SIM_reg_bank__abc_33898_n2134), .Y(REGFILE_SIM_reg_bank_reg_r31_6__FF_INPUT) );
  AND2X2 AND2X2_2066 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n2141_1) );
  AND2X2 AND2X2_2067 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2142_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2139_1), .Y(REGFILE_SIM_reg_bank_reg_r31_7__FF_INPUT) );
  AND2X2 AND2X2_2068 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2146) );
  AND2X2 AND2X2_2069 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2147_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2144_1), .Y(REGFILE_SIM_reg_bank_reg_r31_8__FF_INPUT) );
  AND2X2 AND2X2_207 ( .A(_abc_43815_n621), .B(inst_r_5_), .Y(_abc_43815_n991) );
  AND2X2 AND2X2_2070 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2151_1) );
  AND2X2 AND2X2_2071 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2152), .B(REGFILE_SIM_reg_bank__abc_33898_n2149), .Y(REGFILE_SIM_reg_bank_reg_r31_9__FF_INPUT) );
  AND2X2 AND2X2_2072 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n2156_1) );
  AND2X2 AND2X2_2073 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2157_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2154_1), .Y(REGFILE_SIM_reg_bank_reg_r31_10__FF_INPUT) );
  AND2X2 AND2X2_2074 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2161) );
  AND2X2 AND2X2_2075 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2162_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2159_1), .Y(REGFILE_SIM_reg_bank_reg_r31_11__FF_INPUT) );
  AND2X2 AND2X2_2076 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2166_1) );
  AND2X2 AND2X2_2077 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2167), .B(REGFILE_SIM_reg_bank__abc_33898_n2164), .Y(REGFILE_SIM_reg_bank_reg_r31_12__FF_INPUT) );
  AND2X2 AND2X2_2078 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n2171_1) );
  AND2X2 AND2X2_2079 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2172_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2169_1), .Y(REGFILE_SIM_reg_bank_reg_r31_13__FF_INPUT) );
  AND2X2 AND2X2_208 ( .A(_abc_43815_n991), .B(_abc_43815_n990), .Y(_abc_43815_n992) );
  AND2X2 AND2X2_2080 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2176) );
  AND2X2 AND2X2_2081 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2177_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2174_1), .Y(REGFILE_SIM_reg_bank_reg_r31_14__FF_INPUT) );
  AND2X2 AND2X2_2082 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2181_1) );
  AND2X2 AND2X2_2083 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2182), .B(REGFILE_SIM_reg_bank__abc_33898_n2179), .Y(REGFILE_SIM_reg_bank_reg_r31_15__FF_INPUT) );
  AND2X2 AND2X2_2084 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n2186_1) );
  AND2X2 AND2X2_2085 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2187_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2184_1), .Y(REGFILE_SIM_reg_bank_reg_r31_16__FF_INPUT) );
  AND2X2 AND2X2_2086 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2191) );
  AND2X2 AND2X2_2087 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2192_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2189_1), .Y(REGFILE_SIM_reg_bank_reg_r31_17__FF_INPUT) );
  AND2X2 AND2X2_2088 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2196_1) );
  AND2X2 AND2X2_2089 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2197), .B(REGFILE_SIM_reg_bank__abc_33898_n2194), .Y(REGFILE_SIM_reg_bank_reg_r31_18__FF_INPUT) );
  AND2X2 AND2X2_209 ( .A(_abc_43815_n992), .B(_abc_43815_n994_1), .Y(_abc_43815_n995) );
  AND2X2 AND2X2_2090 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2201) );
  AND2X2 AND2X2_2091 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2202_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2199), .Y(REGFILE_SIM_reg_bank_reg_r31_19__FF_INPUT) );
  AND2X2 AND2X2_2092 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2206_1) );
  AND2X2 AND2X2_2093 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2207), .B(REGFILE_SIM_reg_bank__abc_33898_n2204), .Y(REGFILE_SIM_reg_bank_reg_r31_20__FF_INPUT) );
  AND2X2 AND2X2_2094 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n2211_1) );
  AND2X2 AND2X2_2095 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2212_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2209_1), .Y(REGFILE_SIM_reg_bank_reg_r31_21__FF_INPUT) );
  AND2X2 AND2X2_2096 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2216) );
  AND2X2 AND2X2_2097 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2217_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2214_1), .Y(REGFILE_SIM_reg_bank_reg_r31_22__FF_INPUT) );
  AND2X2 AND2X2_2098 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2221_1) );
  AND2X2 AND2X2_2099 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2222), .B(REGFILE_SIM_reg_bank__abc_33898_n2219), .Y(REGFILE_SIM_reg_bank_reg_r31_23__FF_INPUT) );
  AND2X2 AND2X2_21 ( .A(_abc_43815_n648), .B(_abc_43815_n636), .Y(_abc_43815_n649) );
  AND2X2 AND2X2_210 ( .A(_abc_43815_n995), .B(_abc_43815_n989), .Y(_abc_43815_n996) );
  AND2X2 AND2X2_2100 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n2226_1) );
  AND2X2 AND2X2_2101 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2227_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2224_1), .Y(REGFILE_SIM_reg_bank_reg_r31_24__FF_INPUT) );
  AND2X2 AND2X2_2102 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2231) );
  AND2X2 AND2X2_2103 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2232_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2229_1), .Y(REGFILE_SIM_reg_bank_reg_r31_25__FF_INPUT) );
  AND2X2 AND2X2_2104 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2236_1) );
  AND2X2 AND2X2_2105 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2237), .B(REGFILE_SIM_reg_bank__abc_33898_n2234), .Y(REGFILE_SIM_reg_bank_reg_r31_26__FF_INPUT) );
  AND2X2 AND2X2_2106 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n2241_1) );
  AND2X2 AND2X2_2107 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2242_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2239_1), .Y(REGFILE_SIM_reg_bank_reg_r31_27__FF_INPUT) );
  AND2X2 AND2X2_2108 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2246) );
  AND2X2 AND2X2_2109 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2247_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2244_1), .Y(REGFILE_SIM_reg_bank_reg_r31_28__FF_INPUT) );
  AND2X2 AND2X2_211 ( .A(_abc_43815_n987), .B(_abc_43815_n996), .Y(_abc_43815_n997) );
  AND2X2 AND2X2_2110 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2251_1) );
  AND2X2 AND2X2_2111 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2252), .B(REGFILE_SIM_reg_bank__abc_33898_n2249), .Y(REGFILE_SIM_reg_bank_reg_r31_29__FF_INPUT) );
  AND2X2 AND2X2_2112 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n2256_1) );
  AND2X2 AND2X2_2113 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2257_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2254_1), .Y(REGFILE_SIM_reg_bank_reg_r31_30__FF_INPUT) );
  AND2X2 AND2X2_2114 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2261) );
  AND2X2 AND2X2_2115 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2262_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2259_1), .Y(REGFILE_SIM_reg_bank_reg_r31_31__FF_INPUT) );
  AND2X2 AND2X2_2116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2264), .B(REGFILE_SIM_reg_bank_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2265_1) );
  AND2X2 AND2X2_2117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2265_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2099_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2266_1) );
  AND2X2 AND2X2_2118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2266_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n2267) );
  AND2X2 AND2X2_2119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2270), .B(REGFILE_SIM_reg_bank__abc_33898_n2268_1), .Y(REGFILE_SIM_reg_bank_reg_r30_0__FF_INPUT) );
  AND2X2 AND2X2_212 ( .A(_abc_43815_n1002), .B(opcode_q_24_), .Y(_abc_43815_n1003) );
  AND2X2 AND2X2_2120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2273), .B(REGFILE_SIM_reg_bank__abc_33898_n2272_1), .Y(REGFILE_SIM_reg_bank_reg_r30_1__FF_INPUT) );
  AND2X2 AND2X2_2121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2276), .B(REGFILE_SIM_reg_bank__abc_33898_n2275_1), .Y(REGFILE_SIM_reg_bank_reg_r30_2__FF_INPUT) );
  AND2X2 AND2X2_2122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2279), .B(REGFILE_SIM_reg_bank__abc_33898_n2278_1), .Y(REGFILE_SIM_reg_bank_reg_r30_3__FF_INPUT) );
  AND2X2 AND2X2_2123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2282), .B(REGFILE_SIM_reg_bank__abc_33898_n2281_1), .Y(REGFILE_SIM_reg_bank_reg_r30_4__FF_INPUT) );
  AND2X2 AND2X2_2124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2285), .B(REGFILE_SIM_reg_bank__abc_33898_n2284_1), .Y(REGFILE_SIM_reg_bank_reg_r30_5__FF_INPUT) );
  AND2X2 AND2X2_2125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2288), .B(REGFILE_SIM_reg_bank__abc_33898_n2287_1), .Y(REGFILE_SIM_reg_bank_reg_r30_6__FF_INPUT) );
  AND2X2 AND2X2_2126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2291), .B(REGFILE_SIM_reg_bank__abc_33898_n2290_1), .Y(REGFILE_SIM_reg_bank_reg_r30_7__FF_INPUT) );
  AND2X2 AND2X2_2127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2294), .B(REGFILE_SIM_reg_bank__abc_33898_n2293_1), .Y(REGFILE_SIM_reg_bank_reg_r30_8__FF_INPUT) );
  AND2X2 AND2X2_2128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2297_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2296), .Y(REGFILE_SIM_reg_bank_reg_r30_9__FF_INPUT) );
  AND2X2 AND2X2_2129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2300_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2299_1), .Y(REGFILE_SIM_reg_bank_reg_r30_10__FF_INPUT) );
  AND2X2 AND2X2_213 ( .A(_abc_43815_n1007), .B(_abc_43815_n998), .Y(_abc_43815_n1008) );
  AND2X2 AND2X2_2130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2303_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2302_1), .Y(REGFILE_SIM_reg_bank_reg_r30_11__FF_INPUT) );
  AND2X2 AND2X2_2131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2306_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2305_1), .Y(REGFILE_SIM_reg_bank_reg_r30_12__FF_INPUT) );
  AND2X2 AND2X2_2132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2309_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2308_1), .Y(REGFILE_SIM_reg_bank_reg_r30_13__FF_INPUT) );
  AND2X2 AND2X2_2133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2312_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2311_1), .Y(REGFILE_SIM_reg_bank_reg_r30_14__FF_INPUT) );
  AND2X2 AND2X2_2134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2315_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2314_1), .Y(REGFILE_SIM_reg_bank_reg_r30_15__FF_INPUT) );
  AND2X2 AND2X2_2135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2318_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2317_1), .Y(REGFILE_SIM_reg_bank_reg_r30_16__FF_INPUT) );
  AND2X2 AND2X2_2136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2321_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2320_1), .Y(REGFILE_SIM_reg_bank_reg_r30_17__FF_INPUT) );
  AND2X2 AND2X2_2137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2324_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2323_1), .Y(REGFILE_SIM_reg_bank_reg_r30_18__FF_INPUT) );
  AND2X2 AND2X2_2138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2327_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2326_1), .Y(REGFILE_SIM_reg_bank_reg_r30_19__FF_INPUT) );
  AND2X2 AND2X2_2139 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2330_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2329_1), .Y(REGFILE_SIM_reg_bank_reg_r30_20__FF_INPUT) );
  AND2X2 AND2X2_214 ( .A(opcode_q_24_), .B(opcode_q_23_), .Y(_abc_43815_n1011) );
  AND2X2 AND2X2_2140 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2333_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2332_1), .Y(REGFILE_SIM_reg_bank_reg_r30_21__FF_INPUT) );
  AND2X2 AND2X2_2141 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2336_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2335_1), .Y(REGFILE_SIM_reg_bank_reg_r30_22__FF_INPUT) );
  AND2X2 AND2X2_2142 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2339_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2338_1), .Y(REGFILE_SIM_reg_bank_reg_r30_23__FF_INPUT) );
  AND2X2 AND2X2_2143 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2342_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2341_1), .Y(REGFILE_SIM_reg_bank_reg_r30_24__FF_INPUT) );
  AND2X2 AND2X2_2144 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2345_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2344_1), .Y(REGFILE_SIM_reg_bank_reg_r30_25__FF_INPUT) );
  AND2X2 AND2X2_2145 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2348_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2347_1), .Y(REGFILE_SIM_reg_bank_reg_r30_26__FF_INPUT) );
  AND2X2 AND2X2_2146 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2351_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2350_1), .Y(REGFILE_SIM_reg_bank_reg_r30_27__FF_INPUT) );
  AND2X2 AND2X2_2147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2354_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2353_1), .Y(REGFILE_SIM_reg_bank_reg_r30_28__FF_INPUT) );
  AND2X2 AND2X2_2148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2357_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2356_1), .Y(REGFILE_SIM_reg_bank_reg_r30_29__FF_INPUT) );
  AND2X2 AND2X2_2149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2360_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2359_1), .Y(REGFILE_SIM_reg_bank_reg_r30_30__FF_INPUT) );
  AND2X2 AND2X2_215 ( .A(_abc_43815_n1010), .B(_abc_43815_n1011), .Y(_abc_43815_n1012) );
  AND2X2 AND2X2_2150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2363_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2362_1), .Y(REGFILE_SIM_reg_bank_reg_r30_31__FF_INPUT) );
  AND2X2 AND2X2_2151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2365_1), .B(REGFILE_SIM_reg_bank_rd_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2366_1) );
  AND2X2 AND2X2_2152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2366_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2099_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2367) );
  AND2X2 AND2X2_2153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2367), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n2368_1) );
  AND2X2 AND2X2_2154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2371_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2369_1), .Y(REGFILE_SIM_reg_bank_reg_r29_0__FF_INPUT) );
  AND2X2 AND2X2_2155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2374_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2373), .Y(REGFILE_SIM_reg_bank_reg_r29_1__FF_INPUT) );
  AND2X2 AND2X2_2156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2377_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2376), .Y(REGFILE_SIM_reg_bank_reg_r29_2__FF_INPUT) );
  AND2X2 AND2X2_2157 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2380_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2379), .Y(REGFILE_SIM_reg_bank_reg_r29_3__FF_INPUT) );
  AND2X2 AND2X2_2158 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2383_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2382), .Y(REGFILE_SIM_reg_bank_reg_r29_4__FF_INPUT) );
  AND2X2 AND2X2_2159 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2386_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2385), .Y(REGFILE_SIM_reg_bank_reg_r29_5__FF_INPUT) );
  AND2X2 AND2X2_216 ( .A(_abc_43815_n1012), .B(_abc_43815_n992), .Y(_abc_43815_n1013) );
  AND2X2 AND2X2_2160 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2389_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2388), .Y(REGFILE_SIM_reg_bank_reg_r29_6__FF_INPUT) );
  AND2X2 AND2X2_2161 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2392_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2391), .Y(REGFILE_SIM_reg_bank_reg_r29_7__FF_INPUT) );
  AND2X2 AND2X2_2162 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2395), .B(REGFILE_SIM_reg_bank__abc_33898_n2394_1), .Y(REGFILE_SIM_reg_bank_reg_r29_8__FF_INPUT) );
  AND2X2 AND2X2_2163 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2398), .B(REGFILE_SIM_reg_bank__abc_33898_n2397_1), .Y(REGFILE_SIM_reg_bank_reg_r29_9__FF_INPUT) );
  AND2X2 AND2X2_2164 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2401), .B(REGFILE_SIM_reg_bank__abc_33898_n2400_1), .Y(REGFILE_SIM_reg_bank_reg_r29_10__FF_INPUT) );
  AND2X2 AND2X2_2165 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2404), .B(REGFILE_SIM_reg_bank__abc_33898_n2403_1), .Y(REGFILE_SIM_reg_bank_reg_r29_11__FF_INPUT) );
  AND2X2 AND2X2_2166 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2407), .B(REGFILE_SIM_reg_bank__abc_33898_n2406_1), .Y(REGFILE_SIM_reg_bank_reg_r29_12__FF_INPUT) );
  AND2X2 AND2X2_2167 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2410), .B(REGFILE_SIM_reg_bank__abc_33898_n2409_1), .Y(REGFILE_SIM_reg_bank_reg_r29_13__FF_INPUT) );
  AND2X2 AND2X2_2168 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2413), .B(REGFILE_SIM_reg_bank__abc_33898_n2412_1), .Y(REGFILE_SIM_reg_bank_reg_r29_14__FF_INPUT) );
  AND2X2 AND2X2_2169 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2416), .B(REGFILE_SIM_reg_bank__abc_33898_n2415_1), .Y(REGFILE_SIM_reg_bank_reg_r29_15__FF_INPUT) );
  AND2X2 AND2X2_217 ( .A(_abc_43815_n987), .B(_abc_43815_n1013), .Y(_abc_43815_n1014) );
  AND2X2 AND2X2_2170 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2419), .B(REGFILE_SIM_reg_bank__abc_33898_n2418_1), .Y(REGFILE_SIM_reg_bank_reg_r29_16__FF_INPUT) );
  AND2X2 AND2X2_2171 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2422), .B(REGFILE_SIM_reg_bank__abc_33898_n2421_1), .Y(REGFILE_SIM_reg_bank_reg_r29_17__FF_INPUT) );
  AND2X2 AND2X2_2172 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2425), .B(REGFILE_SIM_reg_bank__abc_33898_n2424_1), .Y(REGFILE_SIM_reg_bank_reg_r29_18__FF_INPUT) );
  AND2X2 AND2X2_2173 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2428), .B(REGFILE_SIM_reg_bank__abc_33898_n2427_1), .Y(REGFILE_SIM_reg_bank_reg_r29_19__FF_INPUT) );
  AND2X2 AND2X2_2174 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2431), .B(REGFILE_SIM_reg_bank__abc_33898_n2430_1), .Y(REGFILE_SIM_reg_bank_reg_r29_20__FF_INPUT) );
  AND2X2 AND2X2_2175 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2434), .B(REGFILE_SIM_reg_bank__abc_33898_n2433_1), .Y(REGFILE_SIM_reg_bank_reg_r29_21__FF_INPUT) );
  AND2X2 AND2X2_2176 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2437), .B(REGFILE_SIM_reg_bank__abc_33898_n2436_1), .Y(REGFILE_SIM_reg_bank_reg_r29_22__FF_INPUT) );
  AND2X2 AND2X2_2177 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2440), .B(REGFILE_SIM_reg_bank__abc_33898_n2439_1), .Y(REGFILE_SIM_reg_bank_reg_r29_23__FF_INPUT) );
  AND2X2 AND2X2_2178 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2443), .B(REGFILE_SIM_reg_bank__abc_33898_n2442_1), .Y(REGFILE_SIM_reg_bank_reg_r29_24__FF_INPUT) );
  AND2X2 AND2X2_2179 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2446), .B(REGFILE_SIM_reg_bank__abc_33898_n2445_1), .Y(REGFILE_SIM_reg_bank_reg_r29_25__FF_INPUT) );
  AND2X2 AND2X2_218 ( .A(_abc_43815_n1016), .B(opcode_q_23_), .Y(_abc_43815_n1017) );
  AND2X2 AND2X2_2180 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2449), .B(REGFILE_SIM_reg_bank__abc_33898_n2448_1), .Y(REGFILE_SIM_reg_bank_reg_r29_26__FF_INPUT) );
  AND2X2 AND2X2_2181 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2452), .B(REGFILE_SIM_reg_bank__abc_33898_n2451_1), .Y(REGFILE_SIM_reg_bank_reg_r29_27__FF_INPUT) );
  AND2X2 AND2X2_2182 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2455), .B(REGFILE_SIM_reg_bank__abc_33898_n2454_1), .Y(REGFILE_SIM_reg_bank_reg_r29_28__FF_INPUT) );
  AND2X2 AND2X2_2183 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2458), .B(REGFILE_SIM_reg_bank__abc_33898_n2457_1), .Y(REGFILE_SIM_reg_bank_reg_r29_29__FF_INPUT) );
  AND2X2 AND2X2_2184 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2461), .B(REGFILE_SIM_reg_bank__abc_33898_n2460_1), .Y(REGFILE_SIM_reg_bank_reg_r29_30__FF_INPUT) );
  AND2X2 AND2X2_2185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2464), .B(REGFILE_SIM_reg_bank__abc_33898_n2463_1), .Y(REGFILE_SIM_reg_bank_reg_r29_31__FF_INPUT) );
  AND2X2 AND2X2_2186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2365_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2264), .Y(REGFILE_SIM_reg_bank__abc_33898_n2466_1) );
  AND2X2 AND2X2_2187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2466_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n2467) );
  AND2X2 AND2X2_2188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2467), .B(REGFILE_SIM_reg_bank__abc_33898_n2099_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1) );
  AND2X2 AND2X2_2189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2470) );
  AND2X2 AND2X2_219 ( .A(_abc_43815_n1010), .B(_abc_43815_n1017), .Y(_abc_43815_n1018) );
  AND2X2 AND2X2_2190 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2471_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2469_1), .Y(REGFILE_SIM_reg_bank_reg_r28_0__FF_INPUT) );
  AND2X2 AND2X2_2191 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n2474_1) );
  AND2X2 AND2X2_2192 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2475_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2473), .Y(REGFILE_SIM_reg_bank_reg_r28_1__FF_INPUT) );
  AND2X2 AND2X2_2193 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2478_1) );
  AND2X2 AND2X2_2194 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2479), .B(REGFILE_SIM_reg_bank__abc_33898_n2477_1), .Y(REGFILE_SIM_reg_bank_reg_r28_2__FF_INPUT) );
  AND2X2 AND2X2_2195 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2482) );
  AND2X2 AND2X2_2196 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2483_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2481_1), .Y(REGFILE_SIM_reg_bank_reg_r28_3__FF_INPUT) );
  AND2X2 AND2X2_2197 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n2486_1) );
  AND2X2 AND2X2_2198 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2487_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2485), .Y(REGFILE_SIM_reg_bank_reg_r28_4__FF_INPUT) );
  AND2X2 AND2X2_2199 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2490) );
  AND2X2 AND2X2_22 ( .A(_abc_43815_n646_1_bF_buf3), .B(_abc_43815_n650_bF_buf4), .Y(_abc_43815_n651_1) );
  AND2X2 AND2X2_220 ( .A(_abc_43815_n1018), .B(_abc_43815_n992), .Y(_abc_43815_n1019) );
  AND2X2 AND2X2_2200 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2491_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2489_1), .Y(REGFILE_SIM_reg_bank_reg_r28_5__FF_INPUT) );
  AND2X2 AND2X2_2201 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2494_1) );
  AND2X2 AND2X2_2202 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2495), .B(REGFILE_SIM_reg_bank__abc_33898_n2493_1), .Y(REGFILE_SIM_reg_bank_reg_r28_6__FF_INPUT) );
  AND2X2 AND2X2_2203 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n2498) );
  AND2X2 AND2X2_2204 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2499_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2497_1), .Y(REGFILE_SIM_reg_bank_reg_r28_7__FF_INPUT) );
  AND2X2 AND2X2_2205 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2502_1) );
  AND2X2 AND2X2_2206 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2503_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2501), .Y(REGFILE_SIM_reg_bank_reg_r28_8__FF_INPUT) );
  AND2X2 AND2X2_2207 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2506_1) );
  AND2X2 AND2X2_2208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2507), .B(REGFILE_SIM_reg_bank__abc_33898_n2505_1), .Y(REGFILE_SIM_reg_bank_reg_r28_9__FF_INPUT) );
  AND2X2 AND2X2_2209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n2510) );
  AND2X2 AND2X2_221 ( .A(_abc_43815_n987), .B(_abc_43815_n1019), .Y(_abc_43815_n1020) );
  AND2X2 AND2X2_2210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2511_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2509_1), .Y(REGFILE_SIM_reg_bank_reg_r28_10__FF_INPUT) );
  AND2X2 AND2X2_2211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2514_1) );
  AND2X2 AND2X2_2212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2515_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2513), .Y(REGFILE_SIM_reg_bank_reg_r28_11__FF_INPUT) );
  AND2X2 AND2X2_2213 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2518_1) );
  AND2X2 AND2X2_2214 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2519), .B(REGFILE_SIM_reg_bank__abc_33898_n2517_1), .Y(REGFILE_SIM_reg_bank_reg_r28_12__FF_INPUT) );
  AND2X2 AND2X2_2215 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n2522) );
  AND2X2 AND2X2_2216 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2523_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2521_1), .Y(REGFILE_SIM_reg_bank_reg_r28_13__FF_INPUT) );
  AND2X2 AND2X2_2217 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2526_1) );
  AND2X2 AND2X2_2218 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2527_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2525), .Y(REGFILE_SIM_reg_bank_reg_r28_14__FF_INPUT) );
  AND2X2 AND2X2_2219 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2530_1) );
  AND2X2 AND2X2_222 ( .A(_abc_43815_n1015), .B(_abc_43815_n1021), .Y(_abc_43815_n1022) );
  AND2X2 AND2X2_2220 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2531), .B(REGFILE_SIM_reg_bank__abc_33898_n2529_1), .Y(REGFILE_SIM_reg_bank_reg_r28_15__FF_INPUT) );
  AND2X2 AND2X2_2221 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n2534) );
  AND2X2 AND2X2_2222 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2535_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2533_1), .Y(REGFILE_SIM_reg_bank_reg_r28_16__FF_INPUT) );
  AND2X2 AND2X2_2223 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2538_1) );
  AND2X2 AND2X2_2224 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2539_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2537), .Y(REGFILE_SIM_reg_bank_reg_r28_17__FF_INPUT) );
  AND2X2 AND2X2_2225 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2542_1) );
  AND2X2 AND2X2_2226 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2543), .B(REGFILE_SIM_reg_bank__abc_33898_n2541_1), .Y(REGFILE_SIM_reg_bank_reg_r28_18__FF_INPUT) );
  AND2X2 AND2X2_2227 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2546) );
  AND2X2 AND2X2_2228 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2547_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2545_1), .Y(REGFILE_SIM_reg_bank_reg_r28_19__FF_INPUT) );
  AND2X2 AND2X2_2229 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2550_1) );
  AND2X2 AND2X2_223 ( .A(_abc_43815_n1008), .B(_abc_43815_n1022), .Y(_abc_43815_n1023) );
  AND2X2 AND2X2_2230 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2551_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2549), .Y(REGFILE_SIM_reg_bank_reg_r28_20__FF_INPUT) );
  AND2X2 AND2X2_2231 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n2554_1) );
  AND2X2 AND2X2_2232 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2555), .B(REGFILE_SIM_reg_bank__abc_33898_n2553_1), .Y(REGFILE_SIM_reg_bank_reg_r28_21__FF_INPUT) );
  AND2X2 AND2X2_2233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2558) );
  AND2X2 AND2X2_2234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2559_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2557_1), .Y(REGFILE_SIM_reg_bank_reg_r28_22__FF_INPUT) );
  AND2X2 AND2X2_2235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2562_1) );
  AND2X2 AND2X2_2236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2563_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2561), .Y(REGFILE_SIM_reg_bank_reg_r28_23__FF_INPUT) );
  AND2X2 AND2X2_2237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n2566_1) );
  AND2X2 AND2X2_2238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2567), .B(REGFILE_SIM_reg_bank__abc_33898_n2565_1), .Y(REGFILE_SIM_reg_bank_reg_r28_24__FF_INPUT) );
  AND2X2 AND2X2_2239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2570) );
  AND2X2 AND2X2_224 ( .A(opcode_q_21_), .B(opcode_q_22_), .Y(_abc_43815_n1024) );
  AND2X2 AND2X2_2240 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2571_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2569_1), .Y(REGFILE_SIM_reg_bank_reg_r28_25__FF_INPUT) );
  AND2X2 AND2X2_2241 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2574_1) );
  AND2X2 AND2X2_2242 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2575_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2573), .Y(REGFILE_SIM_reg_bank_reg_r28_26__FF_INPUT) );
  AND2X2 AND2X2_2243 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n2578_1) );
  AND2X2 AND2X2_2244 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2579), .B(REGFILE_SIM_reg_bank__abc_33898_n2577_1), .Y(REGFILE_SIM_reg_bank_reg_r28_27__FF_INPUT) );
  AND2X2 AND2X2_2245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2582) );
  AND2X2 AND2X2_2246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2583_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2581_1), .Y(REGFILE_SIM_reg_bank_reg_r28_28__FF_INPUT) );
  AND2X2 AND2X2_2247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2586_1) );
  AND2X2 AND2X2_2248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2587), .B(REGFILE_SIM_reg_bank__abc_33898_n2585), .Y(REGFILE_SIM_reg_bank_reg_r28_29__FF_INPUT) );
  AND2X2 AND2X2_2249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n2590_1) );
  AND2X2 AND2X2_225 ( .A(_abc_43815_n1028), .B(_abc_43815_n1031_1), .Y(_abc_43815_n1032_1) );
  AND2X2 AND2X2_2250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2591_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2589), .Y(REGFILE_SIM_reg_bank_reg_r28_30__FF_INPUT) );
  AND2X2 AND2X2_2251 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2594_1) );
  AND2X2 AND2X2_2252 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2595), .B(REGFILE_SIM_reg_bank__abc_33898_n2593_1), .Y(REGFILE_SIM_reg_bank_reg_r28_31__FF_INPUT) );
  AND2X2 AND2X2_2253 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2597_1), .B(REGFILE_SIM_reg_bank_rd_i_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2598) );
  AND2X2 AND2X2_2254 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2598), .B(REGFILE_SIM_reg_bank__abc_33898_n2100), .Y(REGFILE_SIM_reg_bank__abc_33898_n2599_1) );
  AND2X2 AND2X2_2255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2599_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n2600_1) );
  AND2X2 AND2X2_2256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2603_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2601), .Y(REGFILE_SIM_reg_bank_reg_r27_0__FF_INPUT) );
  AND2X2 AND2X2_2257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2606_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2605_1), .Y(REGFILE_SIM_reg_bank_reg_r27_1__FF_INPUT) );
  AND2X2 AND2X2_2258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2609_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2608_1), .Y(REGFILE_SIM_reg_bank_reg_r27_2__FF_INPUT) );
  AND2X2 AND2X2_2259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2612_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2611_1), .Y(REGFILE_SIM_reg_bank_reg_r27_3__FF_INPUT) );
  AND2X2 AND2X2_226 ( .A(_abc_43815_n988), .B(_abc_43815_n1033), .Y(_abc_43815_n1034) );
  AND2X2 AND2X2_2260 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2615_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2614_1), .Y(REGFILE_SIM_reg_bank_reg_r27_4__FF_INPUT) );
  AND2X2 AND2X2_2261 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2618_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2617_1), .Y(REGFILE_SIM_reg_bank_reg_r27_5__FF_INPUT) );
  AND2X2 AND2X2_2262 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2621_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2620_1), .Y(REGFILE_SIM_reg_bank_reg_r27_6__FF_INPUT) );
  AND2X2 AND2X2_2263 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2624_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2623_1), .Y(REGFILE_SIM_reg_bank_reg_r27_7__FF_INPUT) );
  AND2X2 AND2X2_2264 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2627_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2626_1), .Y(REGFILE_SIM_reg_bank_reg_r27_8__FF_INPUT) );
  AND2X2 AND2X2_2265 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2630_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2629_1), .Y(REGFILE_SIM_reg_bank_reg_r27_9__FF_INPUT) );
  AND2X2 AND2X2_2266 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2633_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2632_1), .Y(REGFILE_SIM_reg_bank_reg_r27_10__FF_INPUT) );
  AND2X2 AND2X2_2267 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2636_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2635_1), .Y(REGFILE_SIM_reg_bank_reg_r27_11__FF_INPUT) );
  AND2X2 AND2X2_2268 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2639_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2638_1), .Y(REGFILE_SIM_reg_bank_reg_r27_12__FF_INPUT) );
  AND2X2 AND2X2_2269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2642_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2641_1), .Y(REGFILE_SIM_reg_bank_reg_r27_13__FF_INPUT) );
  AND2X2 AND2X2_227 ( .A(_abc_43815_n1032_1), .B(_abc_43815_n1038), .Y(_abc_43815_n1039) );
  AND2X2 AND2X2_2270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2645_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2644_1), .Y(REGFILE_SIM_reg_bank_reg_r27_14__FF_INPUT) );
  AND2X2 AND2X2_2271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2648_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2647_1), .Y(REGFILE_SIM_reg_bank_reg_r27_15__FF_INPUT) );
  AND2X2 AND2X2_2272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2651_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2650_1), .Y(REGFILE_SIM_reg_bank_reg_r27_16__FF_INPUT) );
  AND2X2 AND2X2_2273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2654_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2653_1), .Y(REGFILE_SIM_reg_bank_reg_r27_17__FF_INPUT) );
  AND2X2 AND2X2_2274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2657_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2656_1), .Y(REGFILE_SIM_reg_bank_reg_r27_18__FF_INPUT) );
  AND2X2 AND2X2_2275 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2660_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2659_1), .Y(REGFILE_SIM_reg_bank_reg_r27_19__FF_INPUT) );
  AND2X2 AND2X2_2276 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2663_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2662_1), .Y(REGFILE_SIM_reg_bank_reg_r27_20__FF_INPUT) );
  AND2X2 AND2X2_2277 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2666_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2665_1), .Y(REGFILE_SIM_reg_bank_reg_r27_21__FF_INPUT) );
  AND2X2 AND2X2_2278 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2669_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2668_1), .Y(REGFILE_SIM_reg_bank_reg_r27_22__FF_INPUT) );
  AND2X2 AND2X2_2279 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2672_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2671_1), .Y(REGFILE_SIM_reg_bank_reg_r27_23__FF_INPUT) );
  AND2X2 AND2X2_228 ( .A(_abc_43815_n1039), .B(_abc_43815_n1023), .Y(_abc_43815_n1040) );
  AND2X2 AND2X2_2280 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2675_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2674_1), .Y(REGFILE_SIM_reg_bank_reg_r27_24__FF_INPUT) );
  AND2X2 AND2X2_2281 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2678_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2677_1), .Y(REGFILE_SIM_reg_bank_reg_r27_25__FF_INPUT) );
  AND2X2 AND2X2_2282 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2681_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2680_1), .Y(REGFILE_SIM_reg_bank_reg_r27_26__FF_INPUT) );
  AND2X2 AND2X2_2283 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2684), .B(REGFILE_SIM_reg_bank__abc_33898_n2683_1), .Y(REGFILE_SIM_reg_bank_reg_r27_27__FF_INPUT) );
  AND2X2 AND2X2_2284 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2687_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2686), .Y(REGFILE_SIM_reg_bank_reg_r27_28__FF_INPUT) );
  AND2X2 AND2X2_2285 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2690_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2689), .Y(REGFILE_SIM_reg_bank_reg_r27_29__FF_INPUT) );
  AND2X2 AND2X2_2286 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2693_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2692), .Y(REGFILE_SIM_reg_bank_reg_r27_30__FF_INPUT) );
  AND2X2 AND2X2_2287 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2696_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2695), .Y(REGFILE_SIM_reg_bank_reg_r27_31__FF_INPUT) );
  AND2X2 AND2X2_2288 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2265_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2598), .Y(REGFILE_SIM_reg_bank__abc_33898_n2698) );
  AND2X2 AND2X2_2289 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2698), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1) );
  AND2X2 AND2X2_229 ( .A(_abc_43815_n639), .B(_abc_43815_n653), .Y(_abc_43815_n1043_1) );
  AND2X2 AND2X2_2290 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2701) );
  AND2X2 AND2X2_2291 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2702_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2700_1), .Y(REGFILE_SIM_reg_bank_reg_r26_0__FF_INPUT) );
  AND2X2 AND2X2_2292 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n2705_1) );
  AND2X2 AND2X2_2293 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2706_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2704), .Y(REGFILE_SIM_reg_bank_reg_r26_1__FF_INPUT) );
  AND2X2 AND2X2_2294 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2709_1) );
  AND2X2 AND2X2_2295 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2710), .B(REGFILE_SIM_reg_bank__abc_33898_n2708_1), .Y(REGFILE_SIM_reg_bank_reg_r26_2__FF_INPUT) );
  AND2X2 AND2X2_2296 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2713) );
  AND2X2 AND2X2_2297 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2714_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2712_1), .Y(REGFILE_SIM_reg_bank_reg_r26_3__FF_INPUT) );
  AND2X2 AND2X2_2298 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n2717_1) );
  AND2X2 AND2X2_2299 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2718_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2716), .Y(REGFILE_SIM_reg_bank_reg_r26_4__FF_INPUT) );
  AND2X2 AND2X2_23 ( .A(_abc_43815_n651_1), .B(_abc_43815_n642_1_bF_buf5), .Y(_abc_43815_n652) );
  AND2X2 AND2X2_230 ( .A(_abc_43815_n1043_1), .B(_abc_43815_n626), .Y(_abc_43815_n1044) );
  AND2X2 AND2X2_2300 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2721_1) );
  AND2X2 AND2X2_2301 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2722), .B(REGFILE_SIM_reg_bank__abc_33898_n2720_1), .Y(REGFILE_SIM_reg_bank_reg_r26_5__FF_INPUT) );
  AND2X2 AND2X2_2302 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2725) );
  AND2X2 AND2X2_2303 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2726_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2724_1), .Y(REGFILE_SIM_reg_bank_reg_r26_6__FF_INPUT) );
  AND2X2 AND2X2_2304 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n2729_1) );
  AND2X2 AND2X2_2305 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2730_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2728), .Y(REGFILE_SIM_reg_bank_reg_r26_7__FF_INPUT) );
  AND2X2 AND2X2_2306 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2733_1) );
  AND2X2 AND2X2_2307 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2734), .B(REGFILE_SIM_reg_bank__abc_33898_n2732_1), .Y(REGFILE_SIM_reg_bank_reg_r26_8__FF_INPUT) );
  AND2X2 AND2X2_2308 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2737) );
  AND2X2 AND2X2_2309 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2738_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2736_1), .Y(REGFILE_SIM_reg_bank_reg_r26_9__FF_INPUT) );
  AND2X2 AND2X2_231 ( .A(_abc_43815_n1042), .B(_abc_43815_n1045), .Y(_abc_43815_n1046_1) );
  AND2X2 AND2X2_2310 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n2741_1) );
  AND2X2 AND2X2_2311 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2742_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2740), .Y(REGFILE_SIM_reg_bank_reg_r26_10__FF_INPUT) );
  AND2X2 AND2X2_2312 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2745_1) );
  AND2X2 AND2X2_2313 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2746), .B(REGFILE_SIM_reg_bank__abc_33898_n2744_1), .Y(REGFILE_SIM_reg_bank_reg_r26_11__FF_INPUT) );
  AND2X2 AND2X2_2314 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2749) );
  AND2X2 AND2X2_2315 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2750_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2748_1), .Y(REGFILE_SIM_reg_bank_reg_r26_12__FF_INPUT) );
  AND2X2 AND2X2_2316 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n2753_1) );
  AND2X2 AND2X2_2317 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2754_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2752), .Y(REGFILE_SIM_reg_bank_reg_r26_13__FF_INPUT) );
  AND2X2 AND2X2_2318 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2757_1) );
  AND2X2 AND2X2_2319 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2758), .B(REGFILE_SIM_reg_bank__abc_33898_n2756_1), .Y(REGFILE_SIM_reg_bank_reg_r26_14__FF_INPUT) );
  AND2X2 AND2X2_232 ( .A(_abc_43815_n631), .B(_abc_43815_n656), .Y(_abc_43815_n1047) );
  AND2X2 AND2X2_2320 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2761) );
  AND2X2 AND2X2_2321 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2762_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2760_1), .Y(REGFILE_SIM_reg_bank_reg_r26_15__FF_INPUT) );
  AND2X2 AND2X2_2322 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n2765_1) );
  AND2X2 AND2X2_2323 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2766_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2764), .Y(REGFILE_SIM_reg_bank_reg_r26_16__FF_INPUT) );
  AND2X2 AND2X2_2324 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2769_1) );
  AND2X2 AND2X2_2325 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2770), .B(REGFILE_SIM_reg_bank__abc_33898_n2768_1), .Y(REGFILE_SIM_reg_bank_reg_r26_17__FF_INPUT) );
  AND2X2 AND2X2_2326 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2773) );
  AND2X2 AND2X2_2327 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2774_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2772_1), .Y(REGFILE_SIM_reg_bank_reg_r26_18__FF_INPUT) );
  AND2X2 AND2X2_2328 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2777_1) );
  AND2X2 AND2X2_2329 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2778_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2776), .Y(REGFILE_SIM_reg_bank_reg_r26_19__FF_INPUT) );
  AND2X2 AND2X2_233 ( .A(_abc_43815_n1047), .B(_abc_43815_n624_1), .Y(_abc_43815_n1048) );
  AND2X2 AND2X2_2330 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2781) );
  AND2X2 AND2X2_2331 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2782_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2780_1), .Y(REGFILE_SIM_reg_bank_reg_r26_20__FF_INPUT) );
  AND2X2 AND2X2_2332 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n2785_1) );
  AND2X2 AND2X2_2333 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2786), .B(REGFILE_SIM_reg_bank__abc_33898_n2784_1), .Y(REGFILE_SIM_reg_bank_reg_r26_21__FF_INPUT) );
  AND2X2 AND2X2_2334 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2789) );
  AND2X2 AND2X2_2335 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2790_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2788_1), .Y(REGFILE_SIM_reg_bank_reg_r26_22__FF_INPUT) );
  AND2X2 AND2X2_2336 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2793_1) );
  AND2X2 AND2X2_2337 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2794_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2792), .Y(REGFILE_SIM_reg_bank_reg_r26_23__FF_INPUT) );
  AND2X2 AND2X2_2338 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n2797_1) );
  AND2X2 AND2X2_2339 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2798), .B(REGFILE_SIM_reg_bank__abc_33898_n2796_1), .Y(REGFILE_SIM_reg_bank_reg_r26_24__FF_INPUT) );
  AND2X2 AND2X2_234 ( .A(_abc_43815_n659), .B(_abc_43815_n626), .Y(_abc_43815_n1050) );
  AND2X2 AND2X2_2340 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2801) );
  AND2X2 AND2X2_2341 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2802_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2800_1), .Y(REGFILE_SIM_reg_bank_reg_r26_25__FF_INPUT) );
  AND2X2 AND2X2_2342 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2805_1) );
  AND2X2 AND2X2_2343 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2806_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2804), .Y(REGFILE_SIM_reg_bank_reg_r26_26__FF_INPUT) );
  AND2X2 AND2X2_2344 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n2809_1) );
  AND2X2 AND2X2_2345 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2810), .B(REGFILE_SIM_reg_bank__abc_33898_n2808_1), .Y(REGFILE_SIM_reg_bank_reg_r26_27__FF_INPUT) );
  AND2X2 AND2X2_2346 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2813) );
  AND2X2 AND2X2_2347 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2814_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2812_1), .Y(REGFILE_SIM_reg_bank_reg_r26_28__FF_INPUT) );
  AND2X2 AND2X2_2348 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2817_1) );
  AND2X2 AND2X2_2349 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2818_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2816), .Y(REGFILE_SIM_reg_bank_reg_r26_29__FF_INPUT) );
  AND2X2 AND2X2_235 ( .A(_abc_43815_n1049), .B(_abc_43815_n1051), .Y(_abc_43815_n1052) );
  AND2X2 AND2X2_2350 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n2821_1) );
  AND2X2 AND2X2_2351 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2822), .B(REGFILE_SIM_reg_bank__abc_33898_n2820_1), .Y(REGFILE_SIM_reg_bank_reg_r26_30__FF_INPUT) );
  AND2X2 AND2X2_2352 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2825) );
  AND2X2 AND2X2_2353 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2826_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2824_1), .Y(REGFILE_SIM_reg_bank_reg_r26_31__FF_INPUT) );
  AND2X2 AND2X2_2354 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2366_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2598), .Y(REGFILE_SIM_reg_bank__abc_33898_n2828) );
  AND2X2 AND2X2_2355 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2828), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1) );
  AND2X2 AND2X2_2356 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2831) );
  AND2X2 AND2X2_2357 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2832_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2830_1), .Y(REGFILE_SIM_reg_bank_reg_r25_0__FF_INPUT) );
  AND2X2 AND2X2_2358 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n2835_1) );
  AND2X2 AND2X2_2359 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2836_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2834), .Y(REGFILE_SIM_reg_bank_reg_r25_1__FF_INPUT) );
  AND2X2 AND2X2_236 ( .A(_abc_43815_n1046_1), .B(_abc_43815_n1052), .Y(_abc_43815_n1053) );
  AND2X2 AND2X2_2360 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2839_1) );
  AND2X2 AND2X2_2361 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2840), .B(REGFILE_SIM_reg_bank__abc_33898_n2838_1), .Y(REGFILE_SIM_reg_bank_reg_r25_2__FF_INPUT) );
  AND2X2 AND2X2_2362 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2843) );
  AND2X2 AND2X2_2363 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2844_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2842_1), .Y(REGFILE_SIM_reg_bank_reg_r25_3__FF_INPUT) );
  AND2X2 AND2X2_2364 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n2847_1) );
  AND2X2 AND2X2_2365 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2848_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2846), .Y(REGFILE_SIM_reg_bank_reg_r25_4__FF_INPUT) );
  AND2X2 AND2X2_2366 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2851_1) );
  AND2X2 AND2X2_2367 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2852), .B(REGFILE_SIM_reg_bank__abc_33898_n2850_1), .Y(REGFILE_SIM_reg_bank_reg_r25_5__FF_INPUT) );
  AND2X2 AND2X2_2368 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2855) );
  AND2X2 AND2X2_2369 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2856_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2854_1), .Y(REGFILE_SIM_reg_bank_reg_r25_6__FF_INPUT) );
  AND2X2 AND2X2_237 ( .A(_abc_43815_n659), .B(_abc_43815_n638), .Y(_abc_43815_n1054) );
  AND2X2 AND2X2_2370 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n2859_1) );
  AND2X2 AND2X2_2371 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2860_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2858), .Y(REGFILE_SIM_reg_bank_reg_r25_7__FF_INPUT) );
  AND2X2 AND2X2_2372 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2863_1) );
  AND2X2 AND2X2_2373 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2864), .B(REGFILE_SIM_reg_bank__abc_33898_n2862_1), .Y(REGFILE_SIM_reg_bank_reg_r25_8__FF_INPUT) );
  AND2X2 AND2X2_2374 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2867) );
  AND2X2 AND2X2_2375 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2868_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2866_1), .Y(REGFILE_SIM_reg_bank_reg_r25_9__FF_INPUT) );
  AND2X2 AND2X2_2376 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n2871_1) );
  AND2X2 AND2X2_2377 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2872_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2870), .Y(REGFILE_SIM_reg_bank_reg_r25_10__FF_INPUT) );
  AND2X2 AND2X2_2378 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2875_1) );
  AND2X2 AND2X2_2379 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2876), .B(REGFILE_SIM_reg_bank__abc_33898_n2874_1), .Y(REGFILE_SIM_reg_bank_reg_r25_11__FF_INPUT) );
  AND2X2 AND2X2_238 ( .A(_abc_43815_n654), .B(_abc_43815_n626), .Y(_abc_43815_n1055) );
  AND2X2 AND2X2_2380 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2879_1) );
  AND2X2 AND2X2_2381 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2880), .B(REGFILE_SIM_reg_bank__abc_33898_n2878), .Y(REGFILE_SIM_reg_bank_reg_r25_12__FF_INPUT) );
  AND2X2 AND2X2_2382 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n2883) );
  AND2X2 AND2X2_2383 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2884_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2882_1), .Y(REGFILE_SIM_reg_bank_reg_r25_13__FF_INPUT) );
  AND2X2 AND2X2_2384 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2887_1) );
  AND2X2 AND2X2_2385 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2888_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2886), .Y(REGFILE_SIM_reg_bank_reg_r25_14__FF_INPUT) );
  AND2X2 AND2X2_2386 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2891_1) );
  AND2X2 AND2X2_2387 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2892), .B(REGFILE_SIM_reg_bank__abc_33898_n2890_1), .Y(REGFILE_SIM_reg_bank_reg_r25_15__FF_INPUT) );
  AND2X2 AND2X2_2388 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n2895) );
  AND2X2 AND2X2_2389 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2896_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2894_1), .Y(REGFILE_SIM_reg_bank_reg_r25_16__FF_INPUT) );
  AND2X2 AND2X2_239 ( .A(_abc_43815_n654), .B(_abc_43815_n983), .Y(_abc_43815_n1058) );
  AND2X2 AND2X2_2390 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2899_1) );
  AND2X2 AND2X2_2391 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2900_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2898), .Y(REGFILE_SIM_reg_bank_reg_r25_17__FF_INPUT) );
  AND2X2 AND2X2_2392 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2903_1) );
  AND2X2 AND2X2_2393 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2904), .B(REGFILE_SIM_reg_bank__abc_33898_n2902_1), .Y(REGFILE_SIM_reg_bank_reg_r25_18__FF_INPUT) );
  AND2X2 AND2X2_2394 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2907) );
  AND2X2 AND2X2_2395 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2908_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2906_1), .Y(REGFILE_SIM_reg_bank_reg_r25_19__FF_INPUT) );
  AND2X2 AND2X2_2396 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2911_1) );
  AND2X2 AND2X2_2397 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2912_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2910), .Y(REGFILE_SIM_reg_bank_reg_r25_20__FF_INPUT) );
  AND2X2 AND2X2_2398 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n2915_1) );
  AND2X2 AND2X2_2399 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2916), .B(REGFILE_SIM_reg_bank__abc_33898_n2914_1), .Y(REGFILE_SIM_reg_bank_reg_r25_21__FF_INPUT) );
  AND2X2 AND2X2_24 ( .A(_abc_43815_n622), .B(inst_r_5_), .Y(_abc_43815_n653) );
  AND2X2 AND2X2_240 ( .A(_abc_43815_n640), .B(_abc_43815_n624_1), .Y(_abc_43815_n1060) );
  AND2X2 AND2X2_2400 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2919) );
  AND2X2 AND2X2_2401 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2920_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2918_1), .Y(REGFILE_SIM_reg_bank_reg_r25_22__FF_INPUT) );
  AND2X2 AND2X2_2402 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2923_1) );
  AND2X2 AND2X2_2403 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2924_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2922), .Y(REGFILE_SIM_reg_bank_reg_r25_23__FF_INPUT) );
  AND2X2 AND2X2_2404 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n2927_1) );
  AND2X2 AND2X2_2405 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2928), .B(REGFILE_SIM_reg_bank__abc_33898_n2926_1), .Y(REGFILE_SIM_reg_bank_reg_r25_24__FF_INPUT) );
  AND2X2 AND2X2_2406 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2931) );
  AND2X2 AND2X2_2407 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2932_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2930_1), .Y(REGFILE_SIM_reg_bank_reg_r25_25__FF_INPUT) );
  AND2X2 AND2X2_2408 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2935_1) );
  AND2X2 AND2X2_2409 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2936_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2934), .Y(REGFILE_SIM_reg_bank_reg_r25_26__FF_INPUT) );
  AND2X2 AND2X2_241 ( .A(_abc_43815_n1059), .B(_abc_43815_n1061), .Y(_abc_43815_n1062) );
  AND2X2 AND2X2_2410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n2939_1) );
  AND2X2 AND2X2_2411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2940), .B(REGFILE_SIM_reg_bank__abc_33898_n2938_1), .Y(REGFILE_SIM_reg_bank_reg_r25_27__FF_INPUT) );
  AND2X2 AND2X2_2412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2943) );
  AND2X2 AND2X2_2413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2944_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2942_1), .Y(REGFILE_SIM_reg_bank_reg_r25_28__FF_INPUT) );
  AND2X2 AND2X2_2414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2947_1) );
  AND2X2 AND2X2_2415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2948_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2946), .Y(REGFILE_SIM_reg_bank_reg_r25_29__FF_INPUT) );
  AND2X2 AND2X2_2416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n2951_1) );
  AND2X2 AND2X2_2417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2952), .B(REGFILE_SIM_reg_bank__abc_33898_n2950_1), .Y(REGFILE_SIM_reg_bank_reg_r25_30__FF_INPUT) );
  AND2X2 AND2X2_2418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2955) );
  AND2X2 AND2X2_2419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2956_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2954_1), .Y(REGFILE_SIM_reg_bank_reg_r25_31__FF_INPUT) );
  AND2X2 AND2X2_242 ( .A(_abc_43815_n1057), .B(_abc_43815_n1062), .Y(_abc_43815_n1063) );
  AND2X2 AND2X2_2420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2467), .B(REGFILE_SIM_reg_bank__abc_33898_n2598), .Y(REGFILE_SIM_reg_bank__abc_33898_n2958) );
  AND2X2 AND2X2_2421 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2961), .B(REGFILE_SIM_reg_bank__abc_33898_n2959_1), .Y(REGFILE_SIM_reg_bank_reg_r24_0__FF_INPUT) );
  AND2X2 AND2X2_2422 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2964), .B(REGFILE_SIM_reg_bank__abc_33898_n2963_1), .Y(REGFILE_SIM_reg_bank_reg_r24_1__FF_INPUT) );
  AND2X2 AND2X2_2423 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2967), .B(REGFILE_SIM_reg_bank__abc_33898_n2966_1), .Y(REGFILE_SIM_reg_bank_reg_r24_2__FF_INPUT) );
  AND2X2 AND2X2_2424 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2970), .B(REGFILE_SIM_reg_bank__abc_33898_n2969_1), .Y(REGFILE_SIM_reg_bank_reg_r24_3__FF_INPUT) );
  AND2X2 AND2X2_2425 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2973), .B(REGFILE_SIM_reg_bank__abc_33898_n2972_1), .Y(REGFILE_SIM_reg_bank_reg_r24_4__FF_INPUT) );
  AND2X2 AND2X2_2426 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2976_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2975), .Y(REGFILE_SIM_reg_bank_reg_r24_5__FF_INPUT) );
  AND2X2 AND2X2_2427 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2979_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2978_1), .Y(REGFILE_SIM_reg_bank_reg_r24_6__FF_INPUT) );
  AND2X2 AND2X2_2428 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2982_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2981_1), .Y(REGFILE_SIM_reg_bank_reg_r24_7__FF_INPUT) );
  AND2X2 AND2X2_2429 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2985_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2984_1), .Y(REGFILE_SIM_reg_bank_reg_r24_8__FF_INPUT) );
  AND2X2 AND2X2_243 ( .A(_abc_43815_n1063), .B(_abc_43815_n1053), .Y(_abc_43815_n1064_1) );
  AND2X2 AND2X2_2430 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2988_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2987_1), .Y(REGFILE_SIM_reg_bank_reg_r24_9__FF_INPUT) );
  AND2X2 AND2X2_2431 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2991_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2990_1), .Y(REGFILE_SIM_reg_bank_reg_r24_10__FF_INPUT) );
  AND2X2 AND2X2_2432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2994_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2993_1), .Y(REGFILE_SIM_reg_bank_reg_r24_11__FF_INPUT) );
  AND2X2 AND2X2_2433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2997_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2996_1), .Y(REGFILE_SIM_reg_bank_reg_r24_12__FF_INPUT) );
  AND2X2 AND2X2_2434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3000_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2999_1), .Y(REGFILE_SIM_reg_bank_reg_r24_13__FF_INPUT) );
  AND2X2 AND2X2_2435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3003_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3002_1), .Y(REGFILE_SIM_reg_bank_reg_r24_14__FF_INPUT) );
  AND2X2 AND2X2_2436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3006_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3005_1), .Y(REGFILE_SIM_reg_bank_reg_r24_15__FF_INPUT) );
  AND2X2 AND2X2_2437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3009_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3008_1), .Y(REGFILE_SIM_reg_bank_reg_r24_16__FF_INPUT) );
  AND2X2 AND2X2_2438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3012_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3011_1), .Y(REGFILE_SIM_reg_bank_reg_r24_17__FF_INPUT) );
  AND2X2 AND2X2_2439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3015_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3014_1), .Y(REGFILE_SIM_reg_bank_reg_r24_18__FF_INPUT) );
  AND2X2 AND2X2_244 ( .A(_abc_43815_n627_1), .B(_abc_43815_n643_1), .Y(_abc_43815_n1065_1) );
  AND2X2 AND2X2_2440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3018_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3017_1), .Y(REGFILE_SIM_reg_bank_reg_r24_19__FF_INPUT) );
  AND2X2 AND2X2_2441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3021_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3020_1), .Y(REGFILE_SIM_reg_bank_reg_r24_20__FF_INPUT) );
  AND2X2 AND2X2_2442 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3024_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3023_1), .Y(REGFILE_SIM_reg_bank_reg_r24_21__FF_INPUT) );
  AND2X2 AND2X2_2443 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3027_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3026_1), .Y(REGFILE_SIM_reg_bank_reg_r24_22__FF_INPUT) );
  AND2X2 AND2X2_2444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3030_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3029_1), .Y(REGFILE_SIM_reg_bank_reg_r24_23__FF_INPUT) );
  AND2X2 AND2X2_2445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3033_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3032_1), .Y(REGFILE_SIM_reg_bank_reg_r24_24__FF_INPUT) );
  AND2X2 AND2X2_2446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3036_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3035_1), .Y(REGFILE_SIM_reg_bank_reg_r24_25__FF_INPUT) );
  AND2X2 AND2X2_2447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3039_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3038_1), .Y(REGFILE_SIM_reg_bank_reg_r24_26__FF_INPUT) );
  AND2X2 AND2X2_2448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3042_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3041_1), .Y(REGFILE_SIM_reg_bank_reg_r24_27__FF_INPUT) );
  AND2X2 AND2X2_2449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3045_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3044_1), .Y(REGFILE_SIM_reg_bank_reg_r24_28__FF_INPUT) );
  AND2X2 AND2X2_245 ( .A(_abc_43815_n656), .B(_abc_43815_n643_1), .Y(_abc_43815_n1067) );
  AND2X2 AND2X2_2450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3048_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3047_1), .Y(REGFILE_SIM_reg_bank_reg_r24_29__FF_INPUT) );
  AND2X2 AND2X2_2451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3051_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3050_1), .Y(REGFILE_SIM_reg_bank_reg_r24_30__FF_INPUT) );
  AND2X2 AND2X2_2452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3054_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3053_1), .Y(REGFILE_SIM_reg_bank_reg_r24_31__FF_INPUT) );
  AND2X2 AND2X2_2453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3056_1), .B(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3057_1) );
  AND2X2 AND2X2_2454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3057_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2100), .Y(REGFILE_SIM_reg_bank__abc_33898_n3058) );
  AND2X2 AND2X2_2455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3058), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n3059_1) );
  AND2X2 AND2X2_2456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3062_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3060_1), .Y(REGFILE_SIM_reg_bank_reg_r23_0__FF_INPUT) );
  AND2X2 AND2X2_2457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3065_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3064), .Y(REGFILE_SIM_reg_bank_reg_r23_1__FF_INPUT) );
  AND2X2 AND2X2_2458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3068_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3067), .Y(REGFILE_SIM_reg_bank_reg_r23_2__FF_INPUT) );
  AND2X2 AND2X2_2459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3071_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3070), .Y(REGFILE_SIM_reg_bank_reg_r23_3__FF_INPUT) );
  AND2X2 AND2X2_246 ( .A(_abc_43815_n623), .B(inst_r_4_), .Y(_abc_43815_n1068) );
  AND2X2 AND2X2_2460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3074_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3073), .Y(REGFILE_SIM_reg_bank_reg_r23_4__FF_INPUT) );
  AND2X2 AND2X2_2461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3077_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3076), .Y(REGFILE_SIM_reg_bank_reg_r23_5__FF_INPUT) );
  AND2X2 AND2X2_2462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3080), .B(REGFILE_SIM_reg_bank__abc_33898_n3079_1), .Y(REGFILE_SIM_reg_bank_reg_r23_6__FF_INPUT) );
  AND2X2 AND2X2_2463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3083), .B(REGFILE_SIM_reg_bank__abc_33898_n3082), .Y(REGFILE_SIM_reg_bank_reg_r23_7__FF_INPUT) );
  AND2X2 AND2X2_2464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3086), .B(REGFILE_SIM_reg_bank__abc_33898_n3085), .Y(REGFILE_SIM_reg_bank_reg_r23_8__FF_INPUT) );
  AND2X2 AND2X2_2465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3089), .B(REGFILE_SIM_reg_bank__abc_33898_n3088), .Y(REGFILE_SIM_reg_bank_reg_r23_9__FF_INPUT) );
  AND2X2 AND2X2_2466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3092), .B(REGFILE_SIM_reg_bank__abc_33898_n3091), .Y(REGFILE_SIM_reg_bank_reg_r23_10__FF_INPUT) );
  AND2X2 AND2X2_2467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3095), .B(REGFILE_SIM_reg_bank__abc_33898_n3094), .Y(REGFILE_SIM_reg_bank_reg_r23_11__FF_INPUT) );
  AND2X2 AND2X2_2468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3098), .B(REGFILE_SIM_reg_bank__abc_33898_n3097), .Y(REGFILE_SIM_reg_bank_reg_r23_12__FF_INPUT) );
  AND2X2 AND2X2_2469 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3101), .B(REGFILE_SIM_reg_bank__abc_33898_n3100), .Y(REGFILE_SIM_reg_bank_reg_r23_13__FF_INPUT) );
  AND2X2 AND2X2_247 ( .A(_abc_43815_n1067), .B(_abc_43815_n1068), .Y(_abc_43815_n1069) );
  AND2X2 AND2X2_2470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3104), .B(REGFILE_SIM_reg_bank__abc_33898_n3103), .Y(REGFILE_SIM_reg_bank_reg_r23_14__FF_INPUT) );
  AND2X2 AND2X2_2471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3107), .B(REGFILE_SIM_reg_bank__abc_33898_n3106), .Y(REGFILE_SIM_reg_bank_reg_r23_15__FF_INPUT) );
  AND2X2 AND2X2_2472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3110), .B(REGFILE_SIM_reg_bank__abc_33898_n3109), .Y(REGFILE_SIM_reg_bank_reg_r23_16__FF_INPUT) );
  AND2X2 AND2X2_2473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3113), .B(REGFILE_SIM_reg_bank__abc_33898_n3112), .Y(REGFILE_SIM_reg_bank_reg_r23_17__FF_INPUT) );
  AND2X2 AND2X2_2474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3116), .B(REGFILE_SIM_reg_bank__abc_33898_n3115), .Y(REGFILE_SIM_reg_bank_reg_r23_18__FF_INPUT) );
  AND2X2 AND2X2_2475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3119), .B(REGFILE_SIM_reg_bank__abc_33898_n3118), .Y(REGFILE_SIM_reg_bank_reg_r23_19__FF_INPUT) );
  AND2X2 AND2X2_2476 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3122), .B(REGFILE_SIM_reg_bank__abc_33898_n3121), .Y(REGFILE_SIM_reg_bank_reg_r23_20__FF_INPUT) );
  AND2X2 AND2X2_2477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3125), .B(REGFILE_SIM_reg_bank__abc_33898_n3124), .Y(REGFILE_SIM_reg_bank_reg_r23_21__FF_INPUT) );
  AND2X2 AND2X2_2478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3128), .B(REGFILE_SIM_reg_bank__abc_33898_n3127), .Y(REGFILE_SIM_reg_bank_reg_r23_22__FF_INPUT) );
  AND2X2 AND2X2_2479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3131), .B(REGFILE_SIM_reg_bank__abc_33898_n3130), .Y(REGFILE_SIM_reg_bank_reg_r23_23__FF_INPUT) );
  AND2X2 AND2X2_248 ( .A(_abc_43815_n1066), .B(_abc_43815_n1070), .Y(_abc_43815_n1071) );
  AND2X2 AND2X2_2480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3134), .B(REGFILE_SIM_reg_bank__abc_33898_n3133), .Y(REGFILE_SIM_reg_bank_reg_r23_24__FF_INPUT) );
  AND2X2 AND2X2_2481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3137), .B(REGFILE_SIM_reg_bank__abc_33898_n3136), .Y(REGFILE_SIM_reg_bank_reg_r23_25__FF_INPUT) );
  AND2X2 AND2X2_2482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3140), .B(REGFILE_SIM_reg_bank__abc_33898_n3139), .Y(REGFILE_SIM_reg_bank_reg_r23_26__FF_INPUT) );
  AND2X2 AND2X2_2483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3143), .B(REGFILE_SIM_reg_bank__abc_33898_n3142), .Y(REGFILE_SIM_reg_bank_reg_r23_27__FF_INPUT) );
  AND2X2 AND2X2_2484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3146), .B(REGFILE_SIM_reg_bank__abc_33898_n3145), .Y(REGFILE_SIM_reg_bank_reg_r23_28__FF_INPUT) );
  AND2X2 AND2X2_2485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3149), .B(REGFILE_SIM_reg_bank__abc_33898_n3148), .Y(REGFILE_SIM_reg_bank_reg_r23_29__FF_INPUT) );
  AND2X2 AND2X2_2486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3152), .B(REGFILE_SIM_reg_bank__abc_33898_n3151), .Y(REGFILE_SIM_reg_bank_reg_r23_30__FF_INPUT) );
  AND2X2 AND2X2_2487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3155), .B(REGFILE_SIM_reg_bank__abc_33898_n3154), .Y(REGFILE_SIM_reg_bank_reg_r23_31__FF_INPUT) );
  AND2X2 AND2X2_2488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2265_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3057_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3157) );
  AND2X2 AND2X2_2489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3157), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158) );
  AND2X2 AND2X2_249 ( .A(_abc_43815_n656), .B(_abc_43815_n647_1), .Y(_abc_43815_n1072) );
  AND2X2 AND2X2_2490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3160) );
  AND2X2 AND2X2_2491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3161), .B(REGFILE_SIM_reg_bank__abc_33898_n3159), .Y(REGFILE_SIM_reg_bank_reg_r22_0__FF_INPUT) );
  AND2X2 AND2X2_2492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n3164) );
  AND2X2 AND2X2_2493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3165), .B(REGFILE_SIM_reg_bank__abc_33898_n3163), .Y(REGFILE_SIM_reg_bank_reg_r22_1__FF_INPUT) );
  AND2X2 AND2X2_2494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3168) );
  AND2X2 AND2X2_2495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3169), .B(REGFILE_SIM_reg_bank__abc_33898_n3167), .Y(REGFILE_SIM_reg_bank_reg_r22_2__FF_INPUT) );
  AND2X2 AND2X2_2496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3172) );
  AND2X2 AND2X2_2497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3173), .B(REGFILE_SIM_reg_bank__abc_33898_n3171), .Y(REGFILE_SIM_reg_bank_reg_r22_3__FF_INPUT) );
  AND2X2 AND2X2_2498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n3176) );
  AND2X2 AND2X2_2499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3177), .B(REGFILE_SIM_reg_bank__abc_33898_n3175), .Y(REGFILE_SIM_reg_bank_reg_r22_4__FF_INPUT) );
  AND2X2 AND2X2_25 ( .A(_abc_43815_n643_1), .B(_abc_43815_n653), .Y(_abc_43815_n654) );
  AND2X2 AND2X2_250 ( .A(_abc_43815_n1072), .B(_abc_43815_n624_1), .Y(_abc_43815_n1073) );
  AND2X2 AND2X2_2500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3180) );
  AND2X2 AND2X2_2501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3181), .B(REGFILE_SIM_reg_bank__abc_33898_n3179), .Y(REGFILE_SIM_reg_bank_reg_r22_5__FF_INPUT) );
  AND2X2 AND2X2_2502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3184) );
  AND2X2 AND2X2_2503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3185), .B(REGFILE_SIM_reg_bank__abc_33898_n3183), .Y(REGFILE_SIM_reg_bank_reg_r22_6__FF_INPUT) );
  AND2X2 AND2X2_2504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n3188) );
  AND2X2 AND2X2_2505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3189), .B(REGFILE_SIM_reg_bank__abc_33898_n3187), .Y(REGFILE_SIM_reg_bank_reg_r22_7__FF_INPUT) );
  AND2X2 AND2X2_2506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3192) );
  AND2X2 AND2X2_2507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3193), .B(REGFILE_SIM_reg_bank__abc_33898_n3191), .Y(REGFILE_SIM_reg_bank_reg_r22_8__FF_INPUT) );
  AND2X2 AND2X2_2508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3196) );
  AND2X2 AND2X2_2509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3197_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3195), .Y(REGFILE_SIM_reg_bank_reg_r22_9__FF_INPUT) );
  AND2X2 AND2X2_251 ( .A(_abc_43815_n666), .B(_abc_43815_n624_1), .Y(_abc_43815_n1075) );
  AND2X2 AND2X2_2510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n3200) );
  AND2X2 AND2X2_2511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3201), .B(REGFILE_SIM_reg_bank__abc_33898_n3199), .Y(REGFILE_SIM_reg_bank_reg_r22_10__FF_INPUT) );
  AND2X2 AND2X2_2512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3204) );
  AND2X2 AND2X2_2513 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3205), .B(REGFILE_SIM_reg_bank__abc_33898_n3203), .Y(REGFILE_SIM_reg_bank_reg_r22_11__FF_INPUT) );
  AND2X2 AND2X2_2514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3208) );
  AND2X2 AND2X2_2515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3209), .B(REGFILE_SIM_reg_bank__abc_33898_n3207), .Y(REGFILE_SIM_reg_bank_reg_r22_12__FF_INPUT) );
  AND2X2 AND2X2_2516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n3212) );
  AND2X2 AND2X2_2517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3213), .B(REGFILE_SIM_reg_bank__abc_33898_n3211), .Y(REGFILE_SIM_reg_bank_reg_r22_13__FF_INPUT) );
  AND2X2 AND2X2_2518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3216) );
  AND2X2 AND2X2_2519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3217), .B(REGFILE_SIM_reg_bank__abc_33898_n3215), .Y(REGFILE_SIM_reg_bank_reg_r22_14__FF_INPUT) );
  AND2X2 AND2X2_252 ( .A(_abc_43815_n1076), .B(_abc_43815_n1074), .Y(_abc_43815_n1077) );
  AND2X2 AND2X2_2520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3220) );
  AND2X2 AND2X2_2521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3221), .B(REGFILE_SIM_reg_bank__abc_33898_n3219), .Y(REGFILE_SIM_reg_bank_reg_r22_15__FF_INPUT) );
  AND2X2 AND2X2_2522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n3224) );
  AND2X2 AND2X2_2523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3225), .B(REGFILE_SIM_reg_bank__abc_33898_n3223), .Y(REGFILE_SIM_reg_bank_reg_r22_16__FF_INPUT) );
  AND2X2 AND2X2_2524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3228) );
  AND2X2 AND2X2_2525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3229_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3227), .Y(REGFILE_SIM_reg_bank_reg_r22_17__FF_INPUT) );
  AND2X2 AND2X2_2526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3232) );
  AND2X2 AND2X2_2527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3233), .B(REGFILE_SIM_reg_bank__abc_33898_n3231), .Y(REGFILE_SIM_reg_bank_reg_r22_18__FF_INPUT) );
  AND2X2 AND2X2_2528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3236) );
  AND2X2 AND2X2_2529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3237), .B(REGFILE_SIM_reg_bank__abc_33898_n3235), .Y(REGFILE_SIM_reg_bank_reg_r22_19__FF_INPUT) );
  AND2X2 AND2X2_253 ( .A(_abc_43815_n1071), .B(_abc_43815_n1077), .Y(_abc_43815_n1078) );
  AND2X2 AND2X2_2530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3240) );
  AND2X2 AND2X2_2531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3241), .B(REGFILE_SIM_reg_bank__abc_33898_n3239), .Y(REGFILE_SIM_reg_bank_reg_r22_20__FF_INPUT) );
  AND2X2 AND2X2_2532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n3244) );
  AND2X2 AND2X2_2533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3245), .B(REGFILE_SIM_reg_bank__abc_33898_n3243), .Y(REGFILE_SIM_reg_bank_reg_r22_21__FF_INPUT) );
  AND2X2 AND2X2_2534 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3248) );
  AND2X2 AND2X2_2535 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3249), .B(REGFILE_SIM_reg_bank__abc_33898_n3247), .Y(REGFILE_SIM_reg_bank_reg_r22_22__FF_INPUT) );
  AND2X2 AND2X2_2536 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3252) );
  AND2X2 AND2X2_2537 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3253), .B(REGFILE_SIM_reg_bank__abc_33898_n3251), .Y(REGFILE_SIM_reg_bank_reg_r22_23__FF_INPUT) );
  AND2X2 AND2X2_2538 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n3256) );
  AND2X2 AND2X2_2539 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3257), .B(REGFILE_SIM_reg_bank__abc_33898_n3255), .Y(REGFILE_SIM_reg_bank_reg_r22_24__FF_INPUT) );
  AND2X2 AND2X2_254 ( .A(_abc_43815_n642_1_bF_buf4), .B(_abc_43815_n650_bF_buf3), .Y(_abc_43815_n1079) );
  AND2X2 AND2X2_2540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3260) );
  AND2X2 AND2X2_2541 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3261_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3259), .Y(REGFILE_SIM_reg_bank_reg_r22_25__FF_INPUT) );
  AND2X2 AND2X2_2542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3264) );
  AND2X2 AND2X2_2543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3265), .B(REGFILE_SIM_reg_bank__abc_33898_n3263), .Y(REGFILE_SIM_reg_bank_reg_r22_26__FF_INPUT) );
  AND2X2 AND2X2_2544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n3268) );
  AND2X2 AND2X2_2545 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3269), .B(REGFILE_SIM_reg_bank__abc_33898_n3267), .Y(REGFILE_SIM_reg_bank_reg_r22_27__FF_INPUT) );
  AND2X2 AND2X2_2546 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3272) );
  AND2X2 AND2X2_2547 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3273), .B(REGFILE_SIM_reg_bank__abc_33898_n3271), .Y(REGFILE_SIM_reg_bank_reg_r22_28__FF_INPUT) );
  AND2X2 AND2X2_2548 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3276) );
  AND2X2 AND2X2_2549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3277), .B(REGFILE_SIM_reg_bank__abc_33898_n3275), .Y(REGFILE_SIM_reg_bank_reg_r22_29__FF_INPUT) );
  AND2X2 AND2X2_255 ( .A(_abc_43815_n1047), .B(_abc_43815_n636), .Y(_abc_43815_n1080) );
  AND2X2 AND2X2_2550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n3280) );
  AND2X2 AND2X2_2551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3281), .B(REGFILE_SIM_reg_bank__abc_33898_n3279), .Y(REGFILE_SIM_reg_bank_reg_r22_30__FF_INPUT) );
  AND2X2 AND2X2_2552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3284) );
  AND2X2 AND2X2_2553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3285), .B(REGFILE_SIM_reg_bank__abc_33898_n3283), .Y(REGFILE_SIM_reg_bank_reg_r22_31__FF_INPUT) );
  AND2X2 AND2X2_2554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2366_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3057_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3287) );
  AND2X2 AND2X2_2555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3287), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288) );
  AND2X2 AND2X2_2556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3290) );
  AND2X2 AND2X2_2557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3291), .B(REGFILE_SIM_reg_bank__abc_33898_n3289), .Y(REGFILE_SIM_reg_bank_reg_r21_0__FF_INPUT) );
  AND2X2 AND2X2_2558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n3294) );
  AND2X2 AND2X2_2559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3295), .B(REGFILE_SIM_reg_bank__abc_33898_n3293_1), .Y(REGFILE_SIM_reg_bank_reg_r21_1__FF_INPUT) );
  AND2X2 AND2X2_256 ( .A(_abc_43815_n1081), .B(_abc_43815_n646_1_bF_buf2), .Y(_abc_43815_n1082) );
  AND2X2 AND2X2_2560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3298) );
  AND2X2 AND2X2_2561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3299), .B(REGFILE_SIM_reg_bank__abc_33898_n3297), .Y(REGFILE_SIM_reg_bank_reg_r21_2__FF_INPUT) );
  AND2X2 AND2X2_2562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3302) );
  AND2X2 AND2X2_2563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3303), .B(REGFILE_SIM_reg_bank__abc_33898_n3301), .Y(REGFILE_SIM_reg_bank_reg_r21_3__FF_INPUT) );
  AND2X2 AND2X2_2564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n3306) );
  AND2X2 AND2X2_2565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3307), .B(REGFILE_SIM_reg_bank__abc_33898_n3305), .Y(REGFILE_SIM_reg_bank_reg_r21_4__FF_INPUT) );
  AND2X2 AND2X2_2566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3310) );
  AND2X2 AND2X2_2567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3311), .B(REGFILE_SIM_reg_bank__abc_33898_n3309), .Y(REGFILE_SIM_reg_bank_reg_r21_5__FF_INPUT) );
  AND2X2 AND2X2_2568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3314) );
  AND2X2 AND2X2_2569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3315), .B(REGFILE_SIM_reg_bank__abc_33898_n3313), .Y(REGFILE_SIM_reg_bank_reg_r21_6__FF_INPUT) );
  AND2X2 AND2X2_257 ( .A(_abc_43815_n1082), .B(_abc_43815_n1079), .Y(_abc_43815_n1083_1) );
  AND2X2 AND2X2_2570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n3318) );
  AND2X2 AND2X2_2571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3319), .B(REGFILE_SIM_reg_bank__abc_33898_n3317), .Y(REGFILE_SIM_reg_bank_reg_r21_7__FF_INPUT) );
  AND2X2 AND2X2_2572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3322) );
  AND2X2 AND2X2_2573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3323), .B(REGFILE_SIM_reg_bank__abc_33898_n3321), .Y(REGFILE_SIM_reg_bank_reg_r21_8__FF_INPUT) );
  AND2X2 AND2X2_2574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3326) );
  AND2X2 AND2X2_2575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3327), .B(REGFILE_SIM_reg_bank__abc_33898_n3325_1), .Y(REGFILE_SIM_reg_bank_reg_r21_9__FF_INPUT) );
  AND2X2 AND2X2_2576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n3330) );
  AND2X2 AND2X2_2577 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3331), .B(REGFILE_SIM_reg_bank__abc_33898_n3329), .Y(REGFILE_SIM_reg_bank_reg_r21_10__FF_INPUT) );
  AND2X2 AND2X2_2578 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3334) );
  AND2X2 AND2X2_2579 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3335), .B(REGFILE_SIM_reg_bank__abc_33898_n3333), .Y(REGFILE_SIM_reg_bank_reg_r21_11__FF_INPUT) );
  AND2X2 AND2X2_258 ( .A(_abc_43815_n1078), .B(_abc_43815_n1083_1), .Y(_abc_43815_n1084) );
  AND2X2 AND2X2_2580 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3338) );
  AND2X2 AND2X2_2581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3339), .B(REGFILE_SIM_reg_bank__abc_33898_n3337), .Y(REGFILE_SIM_reg_bank_reg_r21_12__FF_INPUT) );
  AND2X2 AND2X2_2582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n3342) );
  AND2X2 AND2X2_2583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3343), .B(REGFILE_SIM_reg_bank__abc_33898_n3341), .Y(REGFILE_SIM_reg_bank_reg_r21_13__FF_INPUT) );
  AND2X2 AND2X2_2584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3346) );
  AND2X2 AND2X2_2585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3347), .B(REGFILE_SIM_reg_bank__abc_33898_n3345), .Y(REGFILE_SIM_reg_bank_reg_r21_14__FF_INPUT) );
  AND2X2 AND2X2_2586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3350) );
  AND2X2 AND2X2_2587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3351), .B(REGFILE_SIM_reg_bank__abc_33898_n3349), .Y(REGFILE_SIM_reg_bank_reg_r21_15__FF_INPUT) );
  AND2X2 AND2X2_2588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n3354) );
  AND2X2 AND2X2_2589 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3355), .B(REGFILE_SIM_reg_bank__abc_33898_n3353), .Y(REGFILE_SIM_reg_bank_reg_r21_16__FF_INPUT) );
  AND2X2 AND2X2_259 ( .A(_abc_43815_n1064_1), .B(_abc_43815_n1084), .Y(_abc_43815_n1085) );
  AND2X2 AND2X2_2590 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3358) );
  AND2X2 AND2X2_2591 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3359), .B(REGFILE_SIM_reg_bank__abc_33898_n3357_1), .Y(REGFILE_SIM_reg_bank_reg_r21_17__FF_INPUT) );
  AND2X2 AND2X2_2592 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3362) );
  AND2X2 AND2X2_2593 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3363), .B(REGFILE_SIM_reg_bank__abc_33898_n3361), .Y(REGFILE_SIM_reg_bank_reg_r21_18__FF_INPUT) );
  AND2X2 AND2X2_2594 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3366) );
  AND2X2 AND2X2_2595 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3367), .B(REGFILE_SIM_reg_bank__abc_33898_n3365), .Y(REGFILE_SIM_reg_bank_reg_r21_19__FF_INPUT) );
  AND2X2 AND2X2_2596 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3370) );
  AND2X2 AND2X2_2597 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3371), .B(REGFILE_SIM_reg_bank__abc_33898_n3369), .Y(REGFILE_SIM_reg_bank_reg_r21_20__FF_INPUT) );
  AND2X2 AND2X2_2598 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n3374) );
  AND2X2 AND2X2_2599 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3375), .B(REGFILE_SIM_reg_bank__abc_33898_n3373), .Y(REGFILE_SIM_reg_bank_reg_r21_21__FF_INPUT) );
  AND2X2 AND2X2_26 ( .A(_abc_43815_n654), .B(_abc_43815_n637), .Y(_abc_43815_n655) );
  AND2X2 AND2X2_260 ( .A(_abc_43815_n1089), .B(_abc_43815_n1093), .Y(_abc_43815_n1094) );
  AND2X2 AND2X2_2600 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3378) );
  AND2X2 AND2X2_2601 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3379), .B(REGFILE_SIM_reg_bank__abc_33898_n3377), .Y(REGFILE_SIM_reg_bank_reg_r21_22__FF_INPUT) );
  AND2X2 AND2X2_2602 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3382) );
  AND2X2 AND2X2_2603 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3383), .B(REGFILE_SIM_reg_bank__abc_33898_n3381), .Y(REGFILE_SIM_reg_bank_reg_r21_23__FF_INPUT) );
  AND2X2 AND2X2_2604 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n3386) );
  AND2X2 AND2X2_2605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3387), .B(REGFILE_SIM_reg_bank__abc_33898_n3385), .Y(REGFILE_SIM_reg_bank_reg_r21_24__FF_INPUT) );
  AND2X2 AND2X2_2606 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3390) );
  AND2X2 AND2X2_2607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3391), .B(REGFILE_SIM_reg_bank__abc_33898_n3389_1), .Y(REGFILE_SIM_reg_bank_reg_r21_25__FF_INPUT) );
  AND2X2 AND2X2_2608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3394) );
  AND2X2 AND2X2_2609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3395), .B(REGFILE_SIM_reg_bank__abc_33898_n3393), .Y(REGFILE_SIM_reg_bank_reg_r21_26__FF_INPUT) );
  AND2X2 AND2X2_261 ( .A(_abc_43815_n631), .B(_abc_43815_n1016), .Y(_abc_43815_n1095) );
  AND2X2 AND2X2_2610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n3398) );
  AND2X2 AND2X2_2611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3399), .B(REGFILE_SIM_reg_bank__abc_33898_n3397), .Y(REGFILE_SIM_reg_bank_reg_r21_27__FF_INPUT) );
  AND2X2 AND2X2_2612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3402) );
  AND2X2 AND2X2_2613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3403), .B(REGFILE_SIM_reg_bank__abc_33898_n3401), .Y(REGFILE_SIM_reg_bank_reg_r21_28__FF_INPUT) );
  AND2X2 AND2X2_2614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3406) );
  AND2X2 AND2X2_2615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3407), .B(REGFILE_SIM_reg_bank__abc_33898_n3405), .Y(REGFILE_SIM_reg_bank_reg_r21_29__FF_INPUT) );
  AND2X2 AND2X2_2616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n3410) );
  AND2X2 AND2X2_2617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3411), .B(REGFILE_SIM_reg_bank__abc_33898_n3409), .Y(REGFILE_SIM_reg_bank_reg_r21_30__FF_INPUT) );
  AND2X2 AND2X2_2618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3414) );
  AND2X2 AND2X2_2619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3415), .B(REGFILE_SIM_reg_bank__abc_33898_n3413), .Y(REGFILE_SIM_reg_bank_reg_r21_31__FF_INPUT) );
  AND2X2 AND2X2_262 ( .A(_abc_43815_n628), .B(_abc_43815_n1095), .Y(_abc_43815_n1096) );
  AND2X2 AND2X2_2620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2467), .B(REGFILE_SIM_reg_bank__abc_33898_n3057_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3417) );
  AND2X2 AND2X2_2621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3420), .B(REGFILE_SIM_reg_bank__abc_33898_n3418), .Y(REGFILE_SIM_reg_bank_reg_r20_0__FF_INPUT) );
  AND2X2 AND2X2_2622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3423), .B(REGFILE_SIM_reg_bank__abc_33898_n3422), .Y(REGFILE_SIM_reg_bank_reg_r20_1__FF_INPUT) );
  AND2X2 AND2X2_2623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3426), .B(REGFILE_SIM_reg_bank__abc_33898_n3425), .Y(REGFILE_SIM_reg_bank_reg_r20_2__FF_INPUT) );
  AND2X2 AND2X2_2624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3429), .B(REGFILE_SIM_reg_bank__abc_33898_n3428), .Y(REGFILE_SIM_reg_bank_reg_r20_3__FF_INPUT) );
  AND2X2 AND2X2_2625 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3432), .B(REGFILE_SIM_reg_bank__abc_33898_n3431), .Y(REGFILE_SIM_reg_bank_reg_r20_4__FF_INPUT) );
  AND2X2 AND2X2_2626 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3435), .B(REGFILE_SIM_reg_bank__abc_33898_n3434), .Y(REGFILE_SIM_reg_bank_reg_r20_5__FF_INPUT) );
  AND2X2 AND2X2_2627 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3438), .B(REGFILE_SIM_reg_bank__abc_33898_n3437), .Y(REGFILE_SIM_reg_bank_reg_r20_6__FF_INPUT) );
  AND2X2 AND2X2_2628 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3441), .B(REGFILE_SIM_reg_bank__abc_33898_n3440), .Y(REGFILE_SIM_reg_bank_reg_r20_7__FF_INPUT) );
  AND2X2 AND2X2_2629 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3444), .B(REGFILE_SIM_reg_bank__abc_33898_n3443), .Y(REGFILE_SIM_reg_bank_reg_r20_8__FF_INPUT) );
  AND2X2 AND2X2_263 ( .A(_abc_43815_n1101), .B(_abc_43815_n1098), .Y(_abc_43815_n1102_1) );
  AND2X2 AND2X2_2630 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3447), .B(REGFILE_SIM_reg_bank__abc_33898_n3446), .Y(REGFILE_SIM_reg_bank_reg_r20_9__FF_INPUT) );
  AND2X2 AND2X2_2631 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3450), .B(REGFILE_SIM_reg_bank__abc_33898_n3449), .Y(REGFILE_SIM_reg_bank_reg_r20_10__FF_INPUT) );
  AND2X2 AND2X2_2632 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3453_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3452), .Y(REGFILE_SIM_reg_bank_reg_r20_11__FF_INPUT) );
  AND2X2 AND2X2_2633 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3456), .B(REGFILE_SIM_reg_bank__abc_33898_n3455), .Y(REGFILE_SIM_reg_bank_reg_r20_12__FF_INPUT) );
  AND2X2 AND2X2_2634 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3459), .B(REGFILE_SIM_reg_bank__abc_33898_n3458), .Y(REGFILE_SIM_reg_bank_reg_r20_13__FF_INPUT) );
  AND2X2 AND2X2_2635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3462), .B(REGFILE_SIM_reg_bank__abc_33898_n3461), .Y(REGFILE_SIM_reg_bank_reg_r20_14__FF_INPUT) );
  AND2X2 AND2X2_2636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3465), .B(REGFILE_SIM_reg_bank__abc_33898_n3464), .Y(REGFILE_SIM_reg_bank_reg_r20_15__FF_INPUT) );
  AND2X2 AND2X2_2637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3468), .B(REGFILE_SIM_reg_bank__abc_33898_n3467), .Y(REGFILE_SIM_reg_bank_reg_r20_16__FF_INPUT) );
  AND2X2 AND2X2_2638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3471), .B(REGFILE_SIM_reg_bank__abc_33898_n3470), .Y(REGFILE_SIM_reg_bank_reg_r20_17__FF_INPUT) );
  AND2X2 AND2X2_2639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3474), .B(REGFILE_SIM_reg_bank__abc_33898_n3473), .Y(REGFILE_SIM_reg_bank_reg_r20_18__FF_INPUT) );
  AND2X2 AND2X2_264 ( .A(_abc_43815_n1094), .B(_abc_43815_n1102_1), .Y(_abc_43815_n1103_1) );
  AND2X2 AND2X2_2640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3477), .B(REGFILE_SIM_reg_bank__abc_33898_n3476), .Y(REGFILE_SIM_reg_bank_reg_r20_19__FF_INPUT) );
  AND2X2 AND2X2_2641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3480), .B(REGFILE_SIM_reg_bank__abc_33898_n3479), .Y(REGFILE_SIM_reg_bank_reg_r20_20__FF_INPUT) );
  AND2X2 AND2X2_2642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3483), .B(REGFILE_SIM_reg_bank__abc_33898_n3482), .Y(REGFILE_SIM_reg_bank_reg_r20_21__FF_INPUT) );
  AND2X2 AND2X2_2643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3486), .B(REGFILE_SIM_reg_bank__abc_33898_n3485_1), .Y(REGFILE_SIM_reg_bank_reg_r20_22__FF_INPUT) );
  AND2X2 AND2X2_2644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3489), .B(REGFILE_SIM_reg_bank__abc_33898_n3488), .Y(REGFILE_SIM_reg_bank_reg_r20_23__FF_INPUT) );
  AND2X2 AND2X2_2645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3492), .B(REGFILE_SIM_reg_bank__abc_33898_n3491), .Y(REGFILE_SIM_reg_bank_reg_r20_24__FF_INPUT) );
  AND2X2 AND2X2_2646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3495), .B(REGFILE_SIM_reg_bank__abc_33898_n3494), .Y(REGFILE_SIM_reg_bank_reg_r20_25__FF_INPUT) );
  AND2X2 AND2X2_2647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3498), .B(REGFILE_SIM_reg_bank__abc_33898_n3497), .Y(REGFILE_SIM_reg_bank_reg_r20_26__FF_INPUT) );
  AND2X2 AND2X2_2648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3501), .B(REGFILE_SIM_reg_bank__abc_33898_n3500), .Y(REGFILE_SIM_reg_bank_reg_r20_27__FF_INPUT) );
  AND2X2 AND2X2_2649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3504), .B(REGFILE_SIM_reg_bank__abc_33898_n3503), .Y(REGFILE_SIM_reg_bank_reg_r20_28__FF_INPUT) );
  AND2X2 AND2X2_265 ( .A(_abc_43815_n1103_1), .B(_abc_43815_n1085), .Y(_abc_43815_n1104) );
  AND2X2 AND2X2_2650 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3507), .B(REGFILE_SIM_reg_bank__abc_33898_n3506), .Y(REGFILE_SIM_reg_bank_reg_r20_29__FF_INPUT) );
  AND2X2 AND2X2_2651 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3510), .B(REGFILE_SIM_reg_bank__abc_33898_n3509), .Y(REGFILE_SIM_reg_bank_reg_r20_30__FF_INPUT) );
  AND2X2 AND2X2_2652 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3513), .B(REGFILE_SIM_reg_bank__abc_33898_n3512), .Y(REGFILE_SIM_reg_bank_reg_r20_31__FF_INPUT) );
  AND2X2 AND2X2_2653 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3056_1), .B(REGFILE_SIM_reg_bank__abc_33898_n2597_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3515) );
  AND2X2 AND2X2_2654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3515), .B(REGFILE_SIM_reg_bank__abc_33898_n2100), .Y(REGFILE_SIM_reg_bank__abc_33898_n3516) );
  AND2X2 AND2X2_2655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3516), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n3517_1) );
  AND2X2 AND2X2_2656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3520), .B(REGFILE_SIM_reg_bank__abc_33898_n3518), .Y(REGFILE_SIM_reg_bank_reg_r19_0__FF_INPUT) );
  AND2X2 AND2X2_2657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3523), .B(REGFILE_SIM_reg_bank__abc_33898_n3522), .Y(REGFILE_SIM_reg_bank_reg_r19_1__FF_INPUT) );
  AND2X2 AND2X2_2658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3526), .B(REGFILE_SIM_reg_bank__abc_33898_n3525), .Y(REGFILE_SIM_reg_bank_reg_r19_2__FF_INPUT) );
  AND2X2 AND2X2_2659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3529), .B(REGFILE_SIM_reg_bank__abc_33898_n3528), .Y(REGFILE_SIM_reg_bank_reg_r19_3__FF_INPUT) );
  AND2X2 AND2X2_266 ( .A(_abc_43815_n1040), .B(_abc_43815_n1104), .Y(_abc_43815_n1105) );
  AND2X2 AND2X2_2660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3532), .B(REGFILE_SIM_reg_bank__abc_33898_n3531), .Y(REGFILE_SIM_reg_bank_reg_r19_4__FF_INPUT) );
  AND2X2 AND2X2_2661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3535), .B(REGFILE_SIM_reg_bank__abc_33898_n3534), .Y(REGFILE_SIM_reg_bank_reg_r19_5__FF_INPUT) );
  AND2X2 AND2X2_2662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3538), .B(REGFILE_SIM_reg_bank__abc_33898_n3537), .Y(REGFILE_SIM_reg_bank_reg_r19_6__FF_INPUT) );
  AND2X2 AND2X2_2663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3541), .B(REGFILE_SIM_reg_bank__abc_33898_n3540), .Y(REGFILE_SIM_reg_bank_reg_r19_7__FF_INPUT) );
  AND2X2 AND2X2_2664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3544), .B(REGFILE_SIM_reg_bank__abc_33898_n3543), .Y(REGFILE_SIM_reg_bank_reg_r19_8__FF_INPUT) );
  AND2X2 AND2X2_2665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3547), .B(REGFILE_SIM_reg_bank__abc_33898_n3546), .Y(REGFILE_SIM_reg_bank_reg_r19_9__FF_INPUT) );
  AND2X2 AND2X2_2666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3550), .B(REGFILE_SIM_reg_bank__abc_33898_n3549_1), .Y(REGFILE_SIM_reg_bank_reg_r19_10__FF_INPUT) );
  AND2X2 AND2X2_2667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3553), .B(REGFILE_SIM_reg_bank__abc_33898_n3552), .Y(REGFILE_SIM_reg_bank_reg_r19_11__FF_INPUT) );
  AND2X2 AND2X2_2668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3556), .B(REGFILE_SIM_reg_bank__abc_33898_n3555), .Y(REGFILE_SIM_reg_bank_reg_r19_12__FF_INPUT) );
  AND2X2 AND2X2_2669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3559), .B(REGFILE_SIM_reg_bank__abc_33898_n3558), .Y(REGFILE_SIM_reg_bank_reg_r19_13__FF_INPUT) );
  AND2X2 AND2X2_267 ( .A(_abc_43815_n985), .B(_abc_43815_n631), .Y(_abc_43815_n1106) );
  AND2X2 AND2X2_2670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3562), .B(REGFILE_SIM_reg_bank__abc_33898_n3561), .Y(REGFILE_SIM_reg_bank_reg_r19_14__FF_INPUT) );
  AND2X2 AND2X2_2671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3565), .B(REGFILE_SIM_reg_bank__abc_33898_n3564), .Y(REGFILE_SIM_reg_bank_reg_r19_15__FF_INPUT) );
  AND2X2 AND2X2_2672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3568), .B(REGFILE_SIM_reg_bank__abc_33898_n3567), .Y(REGFILE_SIM_reg_bank_reg_r19_16__FF_INPUT) );
  AND2X2 AND2X2_2673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3571), .B(REGFILE_SIM_reg_bank__abc_33898_n3570), .Y(REGFILE_SIM_reg_bank_reg_r19_17__FF_INPUT) );
  AND2X2 AND2X2_2674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3574), .B(REGFILE_SIM_reg_bank__abc_33898_n3573), .Y(REGFILE_SIM_reg_bank_reg_r19_18__FF_INPUT) );
  AND2X2 AND2X2_2675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3577), .B(REGFILE_SIM_reg_bank__abc_33898_n3576), .Y(REGFILE_SIM_reg_bank_reg_r19_19__FF_INPUT) );
  AND2X2 AND2X2_2676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3580), .B(REGFILE_SIM_reg_bank__abc_33898_n3579), .Y(REGFILE_SIM_reg_bank_reg_r19_20__FF_INPUT) );
  AND2X2 AND2X2_2677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3583), .B(REGFILE_SIM_reg_bank__abc_33898_n3582), .Y(REGFILE_SIM_reg_bank_reg_r19_21__FF_INPUT) );
  AND2X2 AND2X2_2678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3586), .B(REGFILE_SIM_reg_bank__abc_33898_n3585), .Y(REGFILE_SIM_reg_bank_reg_r19_22__FF_INPUT) );
  AND2X2 AND2X2_2679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3589), .B(REGFILE_SIM_reg_bank__abc_33898_n3588), .Y(REGFILE_SIM_reg_bank_reg_r19_23__FF_INPUT) );
  AND2X2 AND2X2_268 ( .A(_abc_43815_n1107), .B(_abc_43815_n1108_1), .Y(_abc_43815_n1109) );
  AND2X2 AND2X2_2680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3592), .B(REGFILE_SIM_reg_bank__abc_33898_n3591), .Y(REGFILE_SIM_reg_bank_reg_r19_24__FF_INPUT) );
  AND2X2 AND2X2_2681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3595), .B(REGFILE_SIM_reg_bank__abc_33898_n3594), .Y(REGFILE_SIM_reg_bank_reg_r19_25__FF_INPUT) );
  AND2X2 AND2X2_2682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3598), .B(REGFILE_SIM_reg_bank__abc_33898_n3597), .Y(REGFILE_SIM_reg_bank_reg_r19_26__FF_INPUT) );
  AND2X2 AND2X2_2683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3601), .B(REGFILE_SIM_reg_bank__abc_33898_n3600), .Y(REGFILE_SIM_reg_bank_reg_r19_27__FF_INPUT) );
  AND2X2 AND2X2_2684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3604), .B(REGFILE_SIM_reg_bank__abc_33898_n3603), .Y(REGFILE_SIM_reg_bank_reg_r19_28__FF_INPUT) );
  AND2X2 AND2X2_2685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3607), .B(REGFILE_SIM_reg_bank__abc_33898_n3606), .Y(REGFILE_SIM_reg_bank_reg_r19_29__FF_INPUT) );
  AND2X2 AND2X2_2686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3610), .B(REGFILE_SIM_reg_bank__abc_33898_n3609), .Y(REGFILE_SIM_reg_bank_reg_r19_30__FF_INPUT) );
  AND2X2 AND2X2_2687 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3613_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3612), .Y(REGFILE_SIM_reg_bank_reg_r19_31__FF_INPUT) );
  AND2X2 AND2X2_2688 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3515), .B(REGFILE_SIM_reg_bank__abc_33898_n2265_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3615) );
  AND2X2 AND2X2_2689 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3615), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n3616) );
  AND2X2 AND2X2_269 ( .A(_abc_43815_n1110), .B(_abc_43815_n1111), .Y(_abc_43815_n1112) );
  AND2X2 AND2X2_2690 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3619), .B(REGFILE_SIM_reg_bank__abc_33898_n3617), .Y(REGFILE_SIM_reg_bank_reg_r18_0__FF_INPUT) );
  AND2X2 AND2X2_2691 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3622), .B(REGFILE_SIM_reg_bank__abc_33898_n3621), .Y(REGFILE_SIM_reg_bank_reg_r18_1__FF_INPUT) );
  AND2X2 AND2X2_2692 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3625), .B(REGFILE_SIM_reg_bank__abc_33898_n3624), .Y(REGFILE_SIM_reg_bank_reg_r18_2__FF_INPUT) );
  AND2X2 AND2X2_2693 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3628), .B(REGFILE_SIM_reg_bank__abc_33898_n3627), .Y(REGFILE_SIM_reg_bank_reg_r18_3__FF_INPUT) );
  AND2X2 AND2X2_2694 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3631), .B(REGFILE_SIM_reg_bank__abc_33898_n3630), .Y(REGFILE_SIM_reg_bank_reg_r18_4__FF_INPUT) );
  AND2X2 AND2X2_2695 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3634), .B(REGFILE_SIM_reg_bank__abc_33898_n3633), .Y(REGFILE_SIM_reg_bank_reg_r18_5__FF_INPUT) );
  AND2X2 AND2X2_2696 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3637), .B(REGFILE_SIM_reg_bank__abc_33898_n3636), .Y(REGFILE_SIM_reg_bank_reg_r18_6__FF_INPUT) );
  AND2X2 AND2X2_2697 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3640), .B(REGFILE_SIM_reg_bank__abc_33898_n3639), .Y(REGFILE_SIM_reg_bank_reg_r18_7__FF_INPUT) );
  AND2X2 AND2X2_2698 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3643), .B(REGFILE_SIM_reg_bank__abc_33898_n3642), .Y(REGFILE_SIM_reg_bank_reg_r18_8__FF_INPUT) );
  AND2X2 AND2X2_2699 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3646), .B(REGFILE_SIM_reg_bank__abc_33898_n3645_1), .Y(REGFILE_SIM_reg_bank_reg_r18_9__FF_INPUT) );
  AND2X2 AND2X2_27 ( .A(_abc_43815_n637), .B(_abc_43815_n625), .Y(_abc_43815_n656) );
  AND2X2 AND2X2_270 ( .A(_abc_43815_n1109), .B(_abc_43815_n1112), .Y(_abc_43815_n1113) );
  AND2X2 AND2X2_2700 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3649), .B(REGFILE_SIM_reg_bank__abc_33898_n3648), .Y(REGFILE_SIM_reg_bank_reg_r18_10__FF_INPUT) );
  AND2X2 AND2X2_2701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3652), .B(REGFILE_SIM_reg_bank__abc_33898_n3651), .Y(REGFILE_SIM_reg_bank_reg_r18_11__FF_INPUT) );
  AND2X2 AND2X2_2702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3655), .B(REGFILE_SIM_reg_bank__abc_33898_n3654), .Y(REGFILE_SIM_reg_bank_reg_r18_12__FF_INPUT) );
  AND2X2 AND2X2_2703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3658), .B(REGFILE_SIM_reg_bank__abc_33898_n3657), .Y(REGFILE_SIM_reg_bank_reg_r18_13__FF_INPUT) );
  AND2X2 AND2X2_2704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3661), .B(REGFILE_SIM_reg_bank__abc_33898_n3660), .Y(REGFILE_SIM_reg_bank_reg_r18_14__FF_INPUT) );
  AND2X2 AND2X2_2705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3664), .B(REGFILE_SIM_reg_bank__abc_33898_n3663), .Y(REGFILE_SIM_reg_bank_reg_r18_15__FF_INPUT) );
  AND2X2 AND2X2_2706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3667), .B(REGFILE_SIM_reg_bank__abc_33898_n3666), .Y(REGFILE_SIM_reg_bank_reg_r18_16__FF_INPUT) );
  AND2X2 AND2X2_2707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3670), .B(REGFILE_SIM_reg_bank__abc_33898_n3669), .Y(REGFILE_SIM_reg_bank_reg_r18_17__FF_INPUT) );
  AND2X2 AND2X2_2708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3673), .B(REGFILE_SIM_reg_bank__abc_33898_n3672), .Y(REGFILE_SIM_reg_bank_reg_r18_18__FF_INPUT) );
  AND2X2 AND2X2_2709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3676), .B(REGFILE_SIM_reg_bank__abc_33898_n3675), .Y(REGFILE_SIM_reg_bank_reg_r18_19__FF_INPUT) );
  AND2X2 AND2X2_271 ( .A(_abc_43815_n1114), .B(alu_op_r_3_), .Y(_abc_43815_n1115) );
  AND2X2 AND2X2_2710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3679), .B(REGFILE_SIM_reg_bank__abc_33898_n3678), .Y(REGFILE_SIM_reg_bank_reg_r18_20__FF_INPUT) );
  AND2X2 AND2X2_2711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3682), .B(REGFILE_SIM_reg_bank__abc_33898_n3681), .Y(REGFILE_SIM_reg_bank_reg_r18_21__FF_INPUT) );
  AND2X2 AND2X2_2712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3685), .B(REGFILE_SIM_reg_bank__abc_33898_n3684), .Y(REGFILE_SIM_reg_bank_reg_r18_22__FF_INPUT) );
  AND2X2 AND2X2_2713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3688), .B(REGFILE_SIM_reg_bank__abc_33898_n3687), .Y(REGFILE_SIM_reg_bank_reg_r18_23__FF_INPUT) );
  AND2X2 AND2X2_2714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3691), .B(REGFILE_SIM_reg_bank__abc_33898_n3690), .Y(REGFILE_SIM_reg_bank_reg_r18_24__FF_INPUT) );
  AND2X2 AND2X2_2715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3694), .B(REGFILE_SIM_reg_bank__abc_33898_n3693), .Y(REGFILE_SIM_reg_bank_reg_r18_25__FF_INPUT) );
  AND2X2 AND2X2_2716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3697), .B(REGFILE_SIM_reg_bank__abc_33898_n3696), .Y(REGFILE_SIM_reg_bank_reg_r18_26__FF_INPUT) );
  AND2X2 AND2X2_2717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3700), .B(REGFILE_SIM_reg_bank__abc_33898_n3699), .Y(REGFILE_SIM_reg_bank_reg_r18_27__FF_INPUT) );
  AND2X2 AND2X2_2718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3703), .B(REGFILE_SIM_reg_bank__abc_33898_n3702), .Y(REGFILE_SIM_reg_bank_reg_r18_28__FF_INPUT) );
  AND2X2 AND2X2_2719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3706), .B(REGFILE_SIM_reg_bank__abc_33898_n3705), .Y(REGFILE_SIM_reg_bank_reg_r18_29__FF_INPUT) );
  AND2X2 AND2X2_272 ( .A(_abc_43815_n1116_1), .B(_abc_43815_n1117), .Y(_abc_43815_n1118) );
  AND2X2 AND2X2_2720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3709_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3708), .Y(REGFILE_SIM_reg_bank_reg_r18_30__FF_INPUT) );
  AND2X2 AND2X2_2721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3712), .B(REGFILE_SIM_reg_bank__abc_33898_n3711), .Y(REGFILE_SIM_reg_bank_reg_r18_31__FF_INPUT) );
  AND2X2 AND2X2_2722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3515), .B(REGFILE_SIM_reg_bank__abc_33898_n2366_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3714) );
  AND2X2 AND2X2_2723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3714), .B(REGFILE_SIM_reg_bank__abc_33898_n2102), .Y(REGFILE_SIM_reg_bank__abc_33898_n3715) );
  AND2X2 AND2X2_2724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3718), .B(REGFILE_SIM_reg_bank__abc_33898_n3716), .Y(REGFILE_SIM_reg_bank_reg_r17_0__FF_INPUT) );
  AND2X2 AND2X2_2725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3721), .B(REGFILE_SIM_reg_bank__abc_33898_n3720), .Y(REGFILE_SIM_reg_bank_reg_r17_1__FF_INPUT) );
  AND2X2 AND2X2_2726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3724), .B(REGFILE_SIM_reg_bank__abc_33898_n3723), .Y(REGFILE_SIM_reg_bank_reg_r17_2__FF_INPUT) );
  AND2X2 AND2X2_2727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3727), .B(REGFILE_SIM_reg_bank__abc_33898_n3726), .Y(REGFILE_SIM_reg_bank_reg_r17_3__FF_INPUT) );
  AND2X2 AND2X2_2728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3730), .B(REGFILE_SIM_reg_bank__abc_33898_n3729), .Y(REGFILE_SIM_reg_bank_reg_r17_4__FF_INPUT) );
  AND2X2 AND2X2_2729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3733), .B(REGFILE_SIM_reg_bank__abc_33898_n3732), .Y(REGFILE_SIM_reg_bank_reg_r17_5__FF_INPUT) );
  AND2X2 AND2X2_273 ( .A(_abc_43815_n1118), .B(_abc_43815_n1115), .Y(_abc_43815_n1119_1) );
  AND2X2 AND2X2_2730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3736), .B(REGFILE_SIM_reg_bank__abc_33898_n3735), .Y(REGFILE_SIM_reg_bank_reg_r17_6__FF_INPUT) );
  AND2X2 AND2X2_2731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3739), .B(REGFILE_SIM_reg_bank__abc_33898_n3738), .Y(REGFILE_SIM_reg_bank_reg_r17_7__FF_INPUT) );
  AND2X2 AND2X2_2732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3742), .B(REGFILE_SIM_reg_bank__abc_33898_n3741_1), .Y(REGFILE_SIM_reg_bank_reg_r17_8__FF_INPUT) );
  AND2X2 AND2X2_2733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3745), .B(REGFILE_SIM_reg_bank__abc_33898_n3744), .Y(REGFILE_SIM_reg_bank_reg_r17_9__FF_INPUT) );
  AND2X2 AND2X2_2734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3748), .B(REGFILE_SIM_reg_bank__abc_33898_n3747), .Y(REGFILE_SIM_reg_bank_reg_r17_10__FF_INPUT) );
  AND2X2 AND2X2_2735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3751), .B(REGFILE_SIM_reg_bank__abc_33898_n3750), .Y(REGFILE_SIM_reg_bank_reg_r17_11__FF_INPUT) );
  AND2X2 AND2X2_2736 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3754), .B(REGFILE_SIM_reg_bank__abc_33898_n3753), .Y(REGFILE_SIM_reg_bank_reg_r17_12__FF_INPUT) );
  AND2X2 AND2X2_2737 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3757), .B(REGFILE_SIM_reg_bank__abc_33898_n3756), .Y(REGFILE_SIM_reg_bank_reg_r17_13__FF_INPUT) );
  AND2X2 AND2X2_2738 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3760), .B(REGFILE_SIM_reg_bank__abc_33898_n3759), .Y(REGFILE_SIM_reg_bank_reg_r17_14__FF_INPUT) );
  AND2X2 AND2X2_2739 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3763), .B(REGFILE_SIM_reg_bank__abc_33898_n3762), .Y(REGFILE_SIM_reg_bank_reg_r17_15__FF_INPUT) );
  AND2X2 AND2X2_274 ( .A(_abc_43815_n1113), .B(_abc_43815_n1119_1), .Y(_abc_43815_n1120) );
  AND2X2 AND2X2_2740 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3766), .B(REGFILE_SIM_reg_bank__abc_33898_n3765), .Y(REGFILE_SIM_reg_bank_reg_r17_16__FF_INPUT) );
  AND2X2 AND2X2_2741 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3769), .B(REGFILE_SIM_reg_bank__abc_33898_n3768), .Y(REGFILE_SIM_reg_bank_reg_r17_17__FF_INPUT) );
  AND2X2 AND2X2_2742 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3772), .B(REGFILE_SIM_reg_bank__abc_33898_n3771), .Y(REGFILE_SIM_reg_bank_reg_r17_18__FF_INPUT) );
  AND2X2 AND2X2_2743 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3775), .B(REGFILE_SIM_reg_bank__abc_33898_n3774), .Y(REGFILE_SIM_reg_bank_reg_r17_19__FF_INPUT) );
  AND2X2 AND2X2_2744 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3778), .B(REGFILE_SIM_reg_bank__abc_33898_n3777), .Y(REGFILE_SIM_reg_bank_reg_r17_20__FF_INPUT) );
  AND2X2 AND2X2_2745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3781), .B(REGFILE_SIM_reg_bank__abc_33898_n3780), .Y(REGFILE_SIM_reg_bank_reg_r17_21__FF_INPUT) );
  AND2X2 AND2X2_2746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3784), .B(REGFILE_SIM_reg_bank__abc_33898_n3783), .Y(REGFILE_SIM_reg_bank_reg_r17_22__FF_INPUT) );
  AND2X2 AND2X2_2747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3787), .B(REGFILE_SIM_reg_bank__abc_33898_n3786), .Y(REGFILE_SIM_reg_bank_reg_r17_23__FF_INPUT) );
  AND2X2 AND2X2_2748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3790), .B(REGFILE_SIM_reg_bank__abc_33898_n3789), .Y(REGFILE_SIM_reg_bank_reg_r17_24__FF_INPUT) );
  AND2X2 AND2X2_2749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3793), .B(REGFILE_SIM_reg_bank__abc_33898_n3792), .Y(REGFILE_SIM_reg_bank_reg_r17_25__FF_INPUT) );
  AND2X2 AND2X2_275 ( .A(_abc_43815_n1120), .B(_abc_43815_n1106), .Y(_abc_43815_n1121) );
  AND2X2 AND2X2_2750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3796), .B(REGFILE_SIM_reg_bank__abc_33898_n3795), .Y(REGFILE_SIM_reg_bank_reg_r17_26__FF_INPUT) );
  AND2X2 AND2X2_2751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3799), .B(REGFILE_SIM_reg_bank__abc_33898_n3798), .Y(REGFILE_SIM_reg_bank_reg_r17_27__FF_INPUT) );
  AND2X2 AND2X2_2752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3802), .B(REGFILE_SIM_reg_bank__abc_33898_n3801), .Y(REGFILE_SIM_reg_bank_reg_r17_28__FF_INPUT) );
  AND2X2 AND2X2_2753 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3805_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3804), .Y(REGFILE_SIM_reg_bank_reg_r17_29__FF_INPUT) );
  AND2X2 AND2X2_2754 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3808), .B(REGFILE_SIM_reg_bank__abc_33898_n3807), .Y(REGFILE_SIM_reg_bank_reg_r17_30__FF_INPUT) );
  AND2X2 AND2X2_2755 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3811), .B(REGFILE_SIM_reg_bank__abc_33898_n3810), .Y(REGFILE_SIM_reg_bank_reg_r17_31__FF_INPUT) );
  AND2X2 AND2X2_2756 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2467), .B(REGFILE_SIM_reg_bank__abc_33898_n3515), .Y(REGFILE_SIM_reg_bank__abc_33898_n3813) );
  AND2X2 AND2X2_2757 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3816), .B(REGFILE_SIM_reg_bank__abc_33898_n3814), .Y(REGFILE_SIM_reg_bank_reg_r16_0__FF_INPUT) );
  AND2X2 AND2X2_2758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3819), .B(REGFILE_SIM_reg_bank__abc_33898_n3818), .Y(REGFILE_SIM_reg_bank_reg_r16_1__FF_INPUT) );
  AND2X2 AND2X2_2759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3822), .B(REGFILE_SIM_reg_bank__abc_33898_n3821), .Y(REGFILE_SIM_reg_bank_reg_r16_2__FF_INPUT) );
  AND2X2 AND2X2_276 ( .A(_abc_43815_n1110), .B(alu_op_r_5_), .Y(_abc_43815_n1123) );
  AND2X2 AND2X2_2760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3825), .B(REGFILE_SIM_reg_bank__abc_33898_n3824), .Y(REGFILE_SIM_reg_bank_reg_r16_3__FF_INPUT) );
  AND2X2 AND2X2_2761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3828), .B(REGFILE_SIM_reg_bank__abc_33898_n3827), .Y(REGFILE_SIM_reg_bank_reg_r16_4__FF_INPUT) );
  AND2X2 AND2X2_2762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3831), .B(REGFILE_SIM_reg_bank__abc_33898_n3830), .Y(REGFILE_SIM_reg_bank_reg_r16_5__FF_INPUT) );
  AND2X2 AND2X2_2763 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3834), .B(REGFILE_SIM_reg_bank__abc_33898_n3833), .Y(REGFILE_SIM_reg_bank_reg_r16_6__FF_INPUT) );
  AND2X2 AND2X2_2764 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3837_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3836), .Y(REGFILE_SIM_reg_bank_reg_r16_7__FF_INPUT) );
  AND2X2 AND2X2_2765 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3840), .B(REGFILE_SIM_reg_bank__abc_33898_n3839), .Y(REGFILE_SIM_reg_bank_reg_r16_8__FF_INPUT) );
  AND2X2 AND2X2_2766 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3843), .B(REGFILE_SIM_reg_bank__abc_33898_n3842), .Y(REGFILE_SIM_reg_bank_reg_r16_9__FF_INPUT) );
  AND2X2 AND2X2_2767 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3846), .B(REGFILE_SIM_reg_bank__abc_33898_n3845), .Y(REGFILE_SIM_reg_bank_reg_r16_10__FF_INPUT) );
  AND2X2 AND2X2_2768 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3849), .B(REGFILE_SIM_reg_bank__abc_33898_n3848), .Y(REGFILE_SIM_reg_bank_reg_r16_11__FF_INPUT) );
  AND2X2 AND2X2_2769 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3852), .B(REGFILE_SIM_reg_bank__abc_33898_n3851), .Y(REGFILE_SIM_reg_bank_reg_r16_12__FF_INPUT) );
  AND2X2 AND2X2_277 ( .A(_abc_43815_n1109), .B(_abc_43815_n1123), .Y(_abc_43815_n1124) );
  AND2X2 AND2X2_2770 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3855), .B(REGFILE_SIM_reg_bank__abc_33898_n3854), .Y(REGFILE_SIM_reg_bank_reg_r16_13__FF_INPUT) );
  AND2X2 AND2X2_2771 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3858), .B(REGFILE_SIM_reg_bank__abc_33898_n3857), .Y(REGFILE_SIM_reg_bank_reg_r16_14__FF_INPUT) );
  AND2X2 AND2X2_2772 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3861), .B(REGFILE_SIM_reg_bank__abc_33898_n3860), .Y(REGFILE_SIM_reg_bank_reg_r16_15__FF_INPUT) );
  AND2X2 AND2X2_2773 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3864), .B(REGFILE_SIM_reg_bank__abc_33898_n3863), .Y(REGFILE_SIM_reg_bank_reg_r16_16__FF_INPUT) );
  AND2X2 AND2X2_2774 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3867), .B(REGFILE_SIM_reg_bank__abc_33898_n3866), .Y(REGFILE_SIM_reg_bank_reg_r16_17__FF_INPUT) );
  AND2X2 AND2X2_2775 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3870), .B(REGFILE_SIM_reg_bank__abc_33898_n3869_1), .Y(REGFILE_SIM_reg_bank_reg_r16_18__FF_INPUT) );
  AND2X2 AND2X2_2776 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3873), .B(REGFILE_SIM_reg_bank__abc_33898_n3872), .Y(REGFILE_SIM_reg_bank_reg_r16_19__FF_INPUT) );
  AND2X2 AND2X2_2777 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3876), .B(REGFILE_SIM_reg_bank__abc_33898_n3875), .Y(REGFILE_SIM_reg_bank_reg_r16_20__FF_INPUT) );
  AND2X2 AND2X2_2778 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3879), .B(REGFILE_SIM_reg_bank__abc_33898_n3878), .Y(REGFILE_SIM_reg_bank_reg_r16_21__FF_INPUT) );
  AND2X2 AND2X2_2779 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3882), .B(REGFILE_SIM_reg_bank__abc_33898_n3881), .Y(REGFILE_SIM_reg_bank_reg_r16_22__FF_INPUT) );
  AND2X2 AND2X2_278 ( .A(_abc_43815_n1119_1), .B(_abc_43815_n1124), .Y(_abc_43815_n1125) );
  AND2X2 AND2X2_2780 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3885), .B(REGFILE_SIM_reg_bank__abc_33898_n3884), .Y(REGFILE_SIM_reg_bank_reg_r16_23__FF_INPUT) );
  AND2X2 AND2X2_2781 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3888), .B(REGFILE_SIM_reg_bank__abc_33898_n3887), .Y(REGFILE_SIM_reg_bank_reg_r16_24__FF_INPUT) );
  AND2X2 AND2X2_2782 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3891), .B(REGFILE_SIM_reg_bank__abc_33898_n3890), .Y(REGFILE_SIM_reg_bank_reg_r16_25__FF_INPUT) );
  AND2X2 AND2X2_2783 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3894), .B(REGFILE_SIM_reg_bank__abc_33898_n3893), .Y(REGFILE_SIM_reg_bank_reg_r16_26__FF_INPUT) );
  AND2X2 AND2X2_2784 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3897), .B(REGFILE_SIM_reg_bank__abc_33898_n3896), .Y(REGFILE_SIM_reg_bank_reg_r16_27__FF_INPUT) );
  AND2X2 AND2X2_2785 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3900), .B(REGFILE_SIM_reg_bank__abc_33898_n3899), .Y(REGFILE_SIM_reg_bank_reg_r16_28__FF_INPUT) );
  AND2X2 AND2X2_2786 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3903), .B(REGFILE_SIM_reg_bank__abc_33898_n3902), .Y(REGFILE_SIM_reg_bank_reg_r16_29__FF_INPUT) );
  AND2X2 AND2X2_2787 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3906), .B(REGFILE_SIM_reg_bank__abc_33898_n3905), .Y(REGFILE_SIM_reg_bank_reg_r16_30__FF_INPUT) );
  AND2X2 AND2X2_2788 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3909), .B(REGFILE_SIM_reg_bank__abc_33898_n3908), .Y(REGFILE_SIM_reg_bank_reg_r16_31__FF_INPUT) );
  AND2X2 AND2X2_2789 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3911), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3912) );
  AND2X2 AND2X2_279 ( .A(_abc_43815_n1125), .B(_abc_43815_n1106), .Y(_abc_43815_n1126) );
  AND2X2 AND2X2_2790 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2101_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913) );
  AND2X2 AND2X2_2791 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3915) );
  AND2X2 AND2X2_2792 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3916), .B(REGFILE_SIM_reg_bank__abc_33898_n3914), .Y(REGFILE_SIM_reg_bank_reg_r15_0__FF_INPUT) );
  AND2X2 AND2X2_2793 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n3919) );
  AND2X2 AND2X2_2794 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3920), .B(REGFILE_SIM_reg_bank__abc_33898_n3918), .Y(REGFILE_SIM_reg_bank_reg_r15_1__FF_INPUT) );
  AND2X2 AND2X2_2795 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3923) );
  AND2X2 AND2X2_2796 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3924), .B(REGFILE_SIM_reg_bank__abc_33898_n3922), .Y(REGFILE_SIM_reg_bank_reg_r15_2__FF_INPUT) );
  AND2X2 AND2X2_2797 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3927) );
  AND2X2 AND2X2_2798 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3928), .B(REGFILE_SIM_reg_bank__abc_33898_n3926), .Y(REGFILE_SIM_reg_bank_reg_r15_3__FF_INPUT) );
  AND2X2 AND2X2_2799 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n3931) );
  AND2X2 AND2X2_28 ( .A(_abc_43815_n656), .B(_abc_43815_n639), .Y(_abc_43815_n657) );
  AND2X2 AND2X2_280 ( .A(_abc_43815_n1127), .B(_abc_43815_n1122), .Y(_abc_43815_n1128) );
  AND2X2 AND2X2_2800 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3932), .B(REGFILE_SIM_reg_bank__abc_33898_n3930), .Y(REGFILE_SIM_reg_bank_reg_r15_4__FF_INPUT) );
  AND2X2 AND2X2_2801 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3935) );
  AND2X2 AND2X2_2802 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3936), .B(REGFILE_SIM_reg_bank__abc_33898_n3934), .Y(REGFILE_SIM_reg_bank_reg_r15_5__FF_INPUT) );
  AND2X2 AND2X2_2803 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3939) );
  AND2X2 AND2X2_2804 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3940), .B(REGFILE_SIM_reg_bank__abc_33898_n3938), .Y(REGFILE_SIM_reg_bank_reg_r15_6__FF_INPUT) );
  AND2X2 AND2X2_2805 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n3943) );
  AND2X2 AND2X2_2806 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3944), .B(REGFILE_SIM_reg_bank__abc_33898_n3942), .Y(REGFILE_SIM_reg_bank_reg_r15_7__FF_INPUT) );
  AND2X2 AND2X2_2807 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3947) );
  AND2X2 AND2X2_2808 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3948), .B(REGFILE_SIM_reg_bank__abc_33898_n3946), .Y(REGFILE_SIM_reg_bank_reg_r15_8__FF_INPUT) );
  AND2X2 AND2X2_2809 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3951) );
  AND2X2 AND2X2_281 ( .A(_abc_43815_n1129), .B(_abc_43815_n1114), .Y(_abc_43815_n1130) );
  AND2X2 AND2X2_2810 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3952), .B(REGFILE_SIM_reg_bank__abc_33898_n3950), .Y(REGFILE_SIM_reg_bank_reg_r15_9__FF_INPUT) );
  AND2X2 AND2X2_2811 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n3955) );
  AND2X2 AND2X2_2812 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3956), .B(REGFILE_SIM_reg_bank__abc_33898_n3954), .Y(REGFILE_SIM_reg_bank_reg_r15_10__FF_INPUT) );
  AND2X2 AND2X2_2813 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3959) );
  AND2X2 AND2X2_2814 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3960), .B(REGFILE_SIM_reg_bank__abc_33898_n3958), .Y(REGFILE_SIM_reg_bank_reg_r15_11__FF_INPUT) );
  AND2X2 AND2X2_2815 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3963) );
  AND2X2 AND2X2_2816 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3964), .B(REGFILE_SIM_reg_bank__abc_33898_n3962), .Y(REGFILE_SIM_reg_bank_reg_r15_12__FF_INPUT) );
  AND2X2 AND2X2_2817 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n3967) );
  AND2X2 AND2X2_2818 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3968), .B(REGFILE_SIM_reg_bank__abc_33898_n3966), .Y(REGFILE_SIM_reg_bank_reg_r15_13__FF_INPUT) );
  AND2X2 AND2X2_2819 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3971) );
  AND2X2 AND2X2_282 ( .A(_abc_43815_n1117), .B(alu_op_r_1_), .Y(_abc_43815_n1131) );
  AND2X2 AND2X2_2820 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3972), .B(REGFILE_SIM_reg_bank__abc_33898_n3970), .Y(REGFILE_SIM_reg_bank_reg_r15_14__FF_INPUT) );
  AND2X2 AND2X2_2821 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3975) );
  AND2X2 AND2X2_2822 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3976), .B(REGFILE_SIM_reg_bank__abc_33898_n3974), .Y(REGFILE_SIM_reg_bank_reg_r15_15__FF_INPUT) );
  AND2X2 AND2X2_2823 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n3979) );
  AND2X2 AND2X2_2824 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3980), .B(REGFILE_SIM_reg_bank__abc_33898_n3978), .Y(REGFILE_SIM_reg_bank_reg_r15_16__FF_INPUT) );
  AND2X2 AND2X2_2825 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3983) );
  AND2X2 AND2X2_2826 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3984), .B(REGFILE_SIM_reg_bank__abc_33898_n3982), .Y(REGFILE_SIM_reg_bank_reg_r15_17__FF_INPUT) );
  AND2X2 AND2X2_2827 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3987) );
  AND2X2 AND2X2_2828 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3988), .B(REGFILE_SIM_reg_bank__abc_33898_n3986), .Y(REGFILE_SIM_reg_bank_reg_r15_18__FF_INPUT) );
  AND2X2 AND2X2_2829 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3991) );
  AND2X2 AND2X2_283 ( .A(_abc_43815_n1130), .B(_abc_43815_n1131), .Y(_abc_43815_n1132) );
  AND2X2 AND2X2_2830 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3992), .B(REGFILE_SIM_reg_bank__abc_33898_n3990), .Y(REGFILE_SIM_reg_bank_reg_r15_19__FF_INPUT) );
  AND2X2 AND2X2_2831 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3995) );
  AND2X2 AND2X2_2832 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3996), .B(REGFILE_SIM_reg_bank__abc_33898_n3994), .Y(REGFILE_SIM_reg_bank_reg_r15_20__FF_INPUT) );
  AND2X2 AND2X2_2833 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n3999) );
  AND2X2 AND2X2_2834 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4000), .B(REGFILE_SIM_reg_bank__abc_33898_n3998), .Y(REGFILE_SIM_reg_bank_reg_r15_21__FF_INPUT) );
  AND2X2 AND2X2_2835 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4003) );
  AND2X2 AND2X2_2836 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4004), .B(REGFILE_SIM_reg_bank__abc_33898_n4002), .Y(REGFILE_SIM_reg_bank_reg_r15_22__FF_INPUT) );
  AND2X2 AND2X2_2837 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4007) );
  AND2X2 AND2X2_2838 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4008), .B(REGFILE_SIM_reg_bank__abc_33898_n4006), .Y(REGFILE_SIM_reg_bank_reg_r15_23__FF_INPUT) );
  AND2X2 AND2X2_2839 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n4011) );
  AND2X2 AND2X2_284 ( .A(_abc_43815_n1113), .B(_abc_43815_n1132), .Y(_abc_43815_n1133) );
  AND2X2 AND2X2_2840 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4012), .B(REGFILE_SIM_reg_bank__abc_33898_n4010), .Y(REGFILE_SIM_reg_bank_reg_r15_24__FF_INPUT) );
  AND2X2 AND2X2_2841 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4015) );
  AND2X2 AND2X2_2842 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4016), .B(REGFILE_SIM_reg_bank__abc_33898_n4014), .Y(REGFILE_SIM_reg_bank_reg_r15_25__FF_INPUT) );
  AND2X2 AND2X2_2843 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4019) );
  AND2X2 AND2X2_2844 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4020), .B(REGFILE_SIM_reg_bank__abc_33898_n4018), .Y(REGFILE_SIM_reg_bank_reg_r15_26__FF_INPUT) );
  AND2X2 AND2X2_2845 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n4023) );
  AND2X2 AND2X2_2846 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4024), .B(REGFILE_SIM_reg_bank__abc_33898_n4022), .Y(REGFILE_SIM_reg_bank_reg_r15_27__FF_INPUT) );
  AND2X2 AND2X2_2847 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4027) );
  AND2X2 AND2X2_2848 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4028), .B(REGFILE_SIM_reg_bank__abc_33898_n4026), .Y(REGFILE_SIM_reg_bank_reg_r15_28__FF_INPUT) );
  AND2X2 AND2X2_2849 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4031) );
  AND2X2 AND2X2_285 ( .A(_abc_43815_n1133), .B(_abc_43815_n1106), .Y(_abc_43815_n1134) );
  AND2X2 AND2X2_2850 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4032), .B(REGFILE_SIM_reg_bank__abc_33898_n4030), .Y(REGFILE_SIM_reg_bank_reg_r15_29__FF_INPUT) );
  AND2X2 AND2X2_2851 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n4035) );
  AND2X2 AND2X2_2852 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4036), .B(REGFILE_SIM_reg_bank__abc_33898_n4034), .Y(REGFILE_SIM_reg_bank_reg_r15_30__FF_INPUT) );
  AND2X2 AND2X2_2853 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4039) );
  AND2X2 AND2X2_2854 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4040), .B(REGFILE_SIM_reg_bank__abc_33898_n4038), .Y(REGFILE_SIM_reg_bank_reg_r15_31__FF_INPUT) );
  AND2X2 AND2X2_2855 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2266_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n4042) );
  AND2X2 AND2X2_2856 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4045), .B(REGFILE_SIM_reg_bank__abc_33898_n4043), .Y(REGFILE_SIM_reg_bank_reg_r14_0__FF_INPUT) );
  AND2X2 AND2X2_2857 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4048), .B(REGFILE_SIM_reg_bank__abc_33898_n4047), .Y(REGFILE_SIM_reg_bank_reg_r14_1__FF_INPUT) );
  AND2X2 AND2X2_2858 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4051), .B(REGFILE_SIM_reg_bank__abc_33898_n4050), .Y(REGFILE_SIM_reg_bank_reg_r14_2__FF_INPUT) );
  AND2X2 AND2X2_2859 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4054), .B(REGFILE_SIM_reg_bank__abc_33898_n4053), .Y(REGFILE_SIM_reg_bank_reg_r14_3__FF_INPUT) );
  AND2X2 AND2X2_286 ( .A(_abc_43815_n1111), .B(alu_op_r_4_), .Y(_abc_43815_n1137) );
  AND2X2 AND2X2_2860 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4057), .B(REGFILE_SIM_reg_bank__abc_33898_n4056), .Y(REGFILE_SIM_reg_bank_reg_r14_4__FF_INPUT) );
  AND2X2 AND2X2_2861 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4060), .B(REGFILE_SIM_reg_bank__abc_33898_n4059), .Y(REGFILE_SIM_reg_bank_reg_r14_5__FF_INPUT) );
  AND2X2 AND2X2_2862 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4063), .B(REGFILE_SIM_reg_bank__abc_33898_n4062), .Y(REGFILE_SIM_reg_bank_reg_r14_6__FF_INPUT) );
  AND2X2 AND2X2_2863 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4066), .B(REGFILE_SIM_reg_bank__abc_33898_n4065), .Y(REGFILE_SIM_reg_bank_reg_r14_7__FF_INPUT) );
  AND2X2 AND2X2_2864 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4069), .B(REGFILE_SIM_reg_bank__abc_33898_n4068), .Y(REGFILE_SIM_reg_bank_reg_r14_8__FF_INPUT) );
  AND2X2 AND2X2_2865 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4072), .B(REGFILE_SIM_reg_bank__abc_33898_n4071), .Y(REGFILE_SIM_reg_bank_reg_r14_9__FF_INPUT) );
  AND2X2 AND2X2_2866 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4075), .B(REGFILE_SIM_reg_bank__abc_33898_n4074), .Y(REGFILE_SIM_reg_bank_reg_r14_10__FF_INPUT) );
  AND2X2 AND2X2_2867 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4078), .B(REGFILE_SIM_reg_bank__abc_33898_n4077), .Y(REGFILE_SIM_reg_bank_reg_r14_11__FF_INPUT) );
  AND2X2 AND2X2_2868 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4081), .B(REGFILE_SIM_reg_bank__abc_33898_n4080), .Y(REGFILE_SIM_reg_bank_reg_r14_12__FF_INPUT) );
  AND2X2 AND2X2_2869 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4084), .B(REGFILE_SIM_reg_bank__abc_33898_n4083), .Y(REGFILE_SIM_reg_bank_reg_r14_13__FF_INPUT) );
  AND2X2 AND2X2_287 ( .A(_abc_43815_n1109), .B(_abc_43815_n1137), .Y(_abc_43815_n1138) );
  AND2X2 AND2X2_2870 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4087), .B(REGFILE_SIM_reg_bank__abc_33898_n4086), .Y(REGFILE_SIM_reg_bank_reg_r14_14__FF_INPUT) );
  AND2X2 AND2X2_2871 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4090), .B(REGFILE_SIM_reg_bank__abc_33898_n4089), .Y(REGFILE_SIM_reg_bank_reg_r14_15__FF_INPUT) );
  AND2X2 AND2X2_2872 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4093_1), .B(REGFILE_SIM_reg_bank__abc_33898_n4092), .Y(REGFILE_SIM_reg_bank_reg_r14_16__FF_INPUT) );
  AND2X2 AND2X2_2873 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4096), .B(REGFILE_SIM_reg_bank__abc_33898_n4095), .Y(REGFILE_SIM_reg_bank_reg_r14_17__FF_INPUT) );
  AND2X2 AND2X2_2874 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4099), .B(REGFILE_SIM_reg_bank__abc_33898_n4098), .Y(REGFILE_SIM_reg_bank_reg_r14_18__FF_INPUT) );
  AND2X2 AND2X2_2875 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4102), .B(REGFILE_SIM_reg_bank__abc_33898_n4101), .Y(REGFILE_SIM_reg_bank_reg_r14_19__FF_INPUT) );
  AND2X2 AND2X2_2876 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4105), .B(REGFILE_SIM_reg_bank__abc_33898_n4104), .Y(REGFILE_SIM_reg_bank_reg_r14_20__FF_INPUT) );
  AND2X2 AND2X2_2877 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4108), .B(REGFILE_SIM_reg_bank__abc_33898_n4107), .Y(REGFILE_SIM_reg_bank_reg_r14_21__FF_INPUT) );
  AND2X2 AND2X2_2878 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4111), .B(REGFILE_SIM_reg_bank__abc_33898_n4110), .Y(REGFILE_SIM_reg_bank_reg_r14_22__FF_INPUT) );
  AND2X2 AND2X2_2879 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4114), .B(REGFILE_SIM_reg_bank__abc_33898_n4113), .Y(REGFILE_SIM_reg_bank_reg_r14_23__FF_INPUT) );
  AND2X2 AND2X2_288 ( .A(_abc_43815_n1119_1), .B(_abc_43815_n1138), .Y(_abc_43815_n1139) );
  AND2X2 AND2X2_2880 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4117), .B(REGFILE_SIM_reg_bank__abc_33898_n4116), .Y(REGFILE_SIM_reg_bank_reg_r14_24__FF_INPUT) );
  AND2X2 AND2X2_2881 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4120), .B(REGFILE_SIM_reg_bank__abc_33898_n4119), .Y(REGFILE_SIM_reg_bank_reg_r14_25__FF_INPUT) );
  AND2X2 AND2X2_2882 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4123), .B(REGFILE_SIM_reg_bank__abc_33898_n4122), .Y(REGFILE_SIM_reg_bank_reg_r14_26__FF_INPUT) );
  AND2X2 AND2X2_2883 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4126), .B(REGFILE_SIM_reg_bank__abc_33898_n4125_1), .Y(REGFILE_SIM_reg_bank_reg_r14_27__FF_INPUT) );
  AND2X2 AND2X2_2884 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4129), .B(REGFILE_SIM_reg_bank__abc_33898_n4128), .Y(REGFILE_SIM_reg_bank_reg_r14_28__FF_INPUT) );
  AND2X2 AND2X2_2885 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4132), .B(REGFILE_SIM_reg_bank__abc_33898_n4131), .Y(REGFILE_SIM_reg_bank_reg_r14_29__FF_INPUT) );
  AND2X2 AND2X2_2886 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4135), .B(REGFILE_SIM_reg_bank__abc_33898_n4134), .Y(REGFILE_SIM_reg_bank_reg_r14_30__FF_INPUT) );
  AND2X2 AND2X2_2887 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4138), .B(REGFILE_SIM_reg_bank__abc_33898_n4137), .Y(REGFILE_SIM_reg_bank_reg_r14_31__FF_INPUT) );
  AND2X2 AND2X2_2888 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2367), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n4140) );
  AND2X2 AND2X2_2889 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4143), .B(REGFILE_SIM_reg_bank__abc_33898_n4141), .Y(REGFILE_SIM_reg_bank_reg_r13_0__FF_INPUT) );
  AND2X2 AND2X2_289 ( .A(_abc_43815_n1141), .B(_abc_43815_n1135_1), .Y(_abc_43815_n1142_1) );
  AND2X2 AND2X2_2890 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4146), .B(REGFILE_SIM_reg_bank__abc_33898_n4145), .Y(REGFILE_SIM_reg_bank_reg_r13_1__FF_INPUT) );
  AND2X2 AND2X2_2891 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4149), .B(REGFILE_SIM_reg_bank__abc_33898_n4148), .Y(REGFILE_SIM_reg_bank_reg_r13_2__FF_INPUT) );
  AND2X2 AND2X2_2892 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4152), .B(REGFILE_SIM_reg_bank__abc_33898_n4151), .Y(REGFILE_SIM_reg_bank_reg_r13_3__FF_INPUT) );
  AND2X2 AND2X2_2893 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4155), .B(REGFILE_SIM_reg_bank__abc_33898_n4154), .Y(REGFILE_SIM_reg_bank_reg_r13_4__FF_INPUT) );
  AND2X2 AND2X2_2894 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4158), .B(REGFILE_SIM_reg_bank__abc_33898_n4157_1), .Y(REGFILE_SIM_reg_bank_reg_r13_5__FF_INPUT) );
  AND2X2 AND2X2_2895 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4161), .B(REGFILE_SIM_reg_bank__abc_33898_n4160), .Y(REGFILE_SIM_reg_bank_reg_r13_6__FF_INPUT) );
  AND2X2 AND2X2_2896 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4164), .B(REGFILE_SIM_reg_bank__abc_33898_n4163), .Y(REGFILE_SIM_reg_bank_reg_r13_7__FF_INPUT) );
  AND2X2 AND2X2_2897 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4167), .B(REGFILE_SIM_reg_bank__abc_33898_n4166), .Y(REGFILE_SIM_reg_bank_reg_r13_8__FF_INPUT) );
  AND2X2 AND2X2_2898 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4170), .B(REGFILE_SIM_reg_bank__abc_33898_n4169), .Y(REGFILE_SIM_reg_bank_reg_r13_9__FF_INPUT) );
  AND2X2 AND2X2_2899 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4173), .B(REGFILE_SIM_reg_bank__abc_33898_n4172), .Y(REGFILE_SIM_reg_bank_reg_r13_10__FF_INPUT) );
  AND2X2 AND2X2_29 ( .A(_abc_43815_n657), .B(_abc_43815_n653), .Y(_abc_43815_n658) );
  AND2X2 AND2X2_290 ( .A(_abc_43815_n1142_1), .B(_abc_43815_n1128), .Y(_abc_43815_n1143) );
  AND2X2 AND2X2_2900 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4176), .B(REGFILE_SIM_reg_bank__abc_33898_n4175), .Y(REGFILE_SIM_reg_bank_reg_r13_11__FF_INPUT) );
  AND2X2 AND2X2_2901 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4179), .B(REGFILE_SIM_reg_bank__abc_33898_n4178), .Y(REGFILE_SIM_reg_bank_reg_r13_12__FF_INPUT) );
  AND2X2 AND2X2_2902 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4182), .B(REGFILE_SIM_reg_bank__abc_33898_n4181), .Y(REGFILE_SIM_reg_bank_reg_r13_13__FF_INPUT) );
  AND2X2 AND2X2_2903 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4185), .B(REGFILE_SIM_reg_bank__abc_33898_n4184), .Y(REGFILE_SIM_reg_bank_reg_r13_14__FF_INPUT) );
  AND2X2 AND2X2_2904 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4188), .B(REGFILE_SIM_reg_bank__abc_33898_n4187), .Y(REGFILE_SIM_reg_bank_reg_r13_15__FF_INPUT) );
  AND2X2 AND2X2_2905 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4191), .B(REGFILE_SIM_reg_bank__abc_33898_n4190_1), .Y(REGFILE_SIM_reg_bank_reg_r13_16__FF_INPUT) );
  AND2X2 AND2X2_2906 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4194), .B(REGFILE_SIM_reg_bank__abc_33898_n4193_1), .Y(REGFILE_SIM_reg_bank_reg_r13_17__FF_INPUT) );
  AND2X2 AND2X2_2907 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4197_1), .B(REGFILE_SIM_reg_bank__abc_33898_n4196), .Y(REGFILE_SIM_reg_bank_reg_r13_18__FF_INPUT) );
  AND2X2 AND2X2_2908 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4200), .B(REGFILE_SIM_reg_bank__abc_33898_n4199), .Y(REGFILE_SIM_reg_bank_reg_r13_19__FF_INPUT) );
  AND2X2 AND2X2_2909 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4203), .B(REGFILE_SIM_reg_bank__abc_33898_n4202), .Y(REGFILE_SIM_reg_bank_reg_r13_20__FF_INPUT) );
  AND2X2 AND2X2_291 ( .A(_abc_43815_n1116_1), .B(alu_op_r_0_), .Y(_abc_43815_n1150) );
  AND2X2 AND2X2_2910 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4206), .B(REGFILE_SIM_reg_bank__abc_33898_n4205), .Y(REGFILE_SIM_reg_bank_reg_r13_21__FF_INPUT) );
  AND2X2 AND2X2_2911 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4209), .B(REGFILE_SIM_reg_bank__abc_33898_n4208), .Y(REGFILE_SIM_reg_bank_reg_r13_22__FF_INPUT) );
  AND2X2 AND2X2_2912 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4212), .B(REGFILE_SIM_reg_bank__abc_33898_n4211), .Y(REGFILE_SIM_reg_bank_reg_r13_23__FF_INPUT) );
  AND2X2 AND2X2_2913 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4215), .B(REGFILE_SIM_reg_bank__abc_33898_n4214), .Y(REGFILE_SIM_reg_bank_reg_r13_24__FF_INPUT) );
  AND2X2 AND2X2_2914 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4218), .B(REGFILE_SIM_reg_bank__abc_33898_n4217), .Y(REGFILE_SIM_reg_bank_reg_r13_25__FF_INPUT) );
  AND2X2 AND2X2_2915 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4221), .B(REGFILE_SIM_reg_bank__abc_33898_n4220), .Y(REGFILE_SIM_reg_bank_reg_r13_26__FF_INPUT) );
  AND2X2 AND2X2_2916 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4224), .B(REGFILE_SIM_reg_bank__abc_33898_n4223), .Y(REGFILE_SIM_reg_bank_reg_r13_27__FF_INPUT) );
  AND2X2 AND2X2_2917 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4227), .B(REGFILE_SIM_reg_bank__abc_33898_n4226), .Y(REGFILE_SIM_reg_bank_reg_r13_28__FF_INPUT) );
  AND2X2 AND2X2_2918 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4230), .B(REGFILE_SIM_reg_bank__abc_33898_n4229), .Y(REGFILE_SIM_reg_bank_reg_r13_29__FF_INPUT) );
  AND2X2 AND2X2_2919 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4233), .B(REGFILE_SIM_reg_bank__abc_33898_n4232), .Y(REGFILE_SIM_reg_bank_reg_r13_30__FF_INPUT) );
  AND2X2 AND2X2_292 ( .A(_abc_43815_n1130), .B(_abc_43815_n1150), .Y(_abc_43815_n1151) );
  AND2X2 AND2X2_2920 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4236), .B(REGFILE_SIM_reg_bank__abc_33898_n4235), .Y(REGFILE_SIM_reg_bank_reg_r13_31__FF_INPUT) );
  AND2X2 AND2X2_2921 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2466_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n4238) );
  AND2X2 AND2X2_2922 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4238), .B(REGFILE_SIM_reg_bank__abc_33898_n2099_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4239) );
  AND2X2 AND2X2_2923 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4242), .B(REGFILE_SIM_reg_bank__abc_33898_n4240), .Y(REGFILE_SIM_reg_bank_reg_r12_0__FF_INPUT) );
  AND2X2 AND2X2_2924 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4245), .B(REGFILE_SIM_reg_bank__abc_33898_n4244), .Y(REGFILE_SIM_reg_bank_reg_r12_1__FF_INPUT) );
  AND2X2 AND2X2_2925 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4248), .B(REGFILE_SIM_reg_bank__abc_33898_n4247), .Y(REGFILE_SIM_reg_bank_reg_r12_2__FF_INPUT) );
  AND2X2 AND2X2_2926 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4251), .B(REGFILE_SIM_reg_bank__abc_33898_n4250), .Y(REGFILE_SIM_reg_bank_reg_r12_3__FF_INPUT) );
  AND2X2 AND2X2_2927 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4254), .B(REGFILE_SIM_reg_bank__abc_33898_n4253), .Y(REGFILE_SIM_reg_bank_reg_r12_4__FF_INPUT) );
  AND2X2 AND2X2_2928 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4257), .B(REGFILE_SIM_reg_bank__abc_33898_n4256), .Y(REGFILE_SIM_reg_bank_reg_r12_5__FF_INPUT) );
  AND2X2 AND2X2_2929 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4260), .B(REGFILE_SIM_reg_bank__abc_33898_n4259), .Y(REGFILE_SIM_reg_bank_reg_r12_6__FF_INPUT) );
  AND2X2 AND2X2_293 ( .A(_abc_43815_n1113), .B(_abc_43815_n1151), .Y(_abc_43815_n1152) );
  AND2X2 AND2X2_2930 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4263), .B(REGFILE_SIM_reg_bank__abc_33898_n4262), .Y(REGFILE_SIM_reg_bank_reg_r12_7__FF_INPUT) );
  AND2X2 AND2X2_2931 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4266), .B(REGFILE_SIM_reg_bank__abc_33898_n4265), .Y(REGFILE_SIM_reg_bank_reg_r12_8__FF_INPUT) );
  AND2X2 AND2X2_2932 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4269), .B(REGFILE_SIM_reg_bank__abc_33898_n4268), .Y(REGFILE_SIM_reg_bank_reg_r12_9__FF_INPUT) );
  AND2X2 AND2X2_2933 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4272), .B(REGFILE_SIM_reg_bank__abc_33898_n4271), .Y(REGFILE_SIM_reg_bank_reg_r12_10__FF_INPUT) );
  AND2X2 AND2X2_2934 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4275), .B(REGFILE_SIM_reg_bank__abc_33898_n4274), .Y(REGFILE_SIM_reg_bank_reg_r12_11__FF_INPUT) );
  AND2X2 AND2X2_2935 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4278), .B(REGFILE_SIM_reg_bank__abc_33898_n4277), .Y(REGFILE_SIM_reg_bank_reg_r12_12__FF_INPUT) );
  AND2X2 AND2X2_2936 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4281), .B(REGFILE_SIM_reg_bank__abc_33898_n4280), .Y(REGFILE_SIM_reg_bank_reg_r12_13__FF_INPUT) );
  AND2X2 AND2X2_2937 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4284), .B(REGFILE_SIM_reg_bank__abc_33898_n4283), .Y(REGFILE_SIM_reg_bank_reg_r12_14__FF_INPUT) );
  AND2X2 AND2X2_2938 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4287), .B(REGFILE_SIM_reg_bank__abc_33898_n4286), .Y(REGFILE_SIM_reg_bank_reg_r12_15__FF_INPUT) );
  AND2X2 AND2X2_2939 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4290), .B(REGFILE_SIM_reg_bank__abc_33898_n4289), .Y(REGFILE_SIM_reg_bank_reg_r12_16__FF_INPUT) );
  AND2X2 AND2X2_294 ( .A(_abc_43815_n1152), .B(_abc_43815_n1106), .Y(_abc_43815_n1153_1) );
  AND2X2 AND2X2_2940 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4293), .B(REGFILE_SIM_reg_bank__abc_33898_n4292), .Y(REGFILE_SIM_reg_bank_reg_r12_17__FF_INPUT) );
  AND2X2 AND2X2_2941 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4296), .B(REGFILE_SIM_reg_bank__abc_33898_n4295), .Y(REGFILE_SIM_reg_bank_reg_r12_18__FF_INPUT) );
  AND2X2 AND2X2_2942 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4299), .B(REGFILE_SIM_reg_bank__abc_33898_n4298), .Y(REGFILE_SIM_reg_bank_reg_r12_19__FF_INPUT) );
  AND2X2 AND2X2_2943 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4302), .B(REGFILE_SIM_reg_bank__abc_33898_n4301), .Y(REGFILE_SIM_reg_bank_reg_r12_20__FF_INPUT) );
  AND2X2 AND2X2_2944 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4305), .B(REGFILE_SIM_reg_bank__abc_33898_n4304), .Y(REGFILE_SIM_reg_bank_reg_r12_21__FF_INPUT) );
  AND2X2 AND2X2_2945 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4308), .B(REGFILE_SIM_reg_bank__abc_33898_n4307), .Y(REGFILE_SIM_reg_bank_reg_r12_22__FF_INPUT) );
  AND2X2 AND2X2_2946 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4311), .B(REGFILE_SIM_reg_bank__abc_33898_n4310), .Y(REGFILE_SIM_reg_bank_reg_r12_23__FF_INPUT) );
  AND2X2 AND2X2_2947 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4314), .B(REGFILE_SIM_reg_bank__abc_33898_n4313_1), .Y(REGFILE_SIM_reg_bank_reg_r12_24__FF_INPUT) );
  AND2X2 AND2X2_2948 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4317), .B(REGFILE_SIM_reg_bank__abc_33898_n4316), .Y(REGFILE_SIM_reg_bank_reg_r12_25__FF_INPUT) );
  AND2X2 AND2X2_2949 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4320), .B(REGFILE_SIM_reg_bank__abc_33898_n4319), .Y(REGFILE_SIM_reg_bank_reg_r12_26__FF_INPUT) );
  AND2X2 AND2X2_295 ( .A(_abc_43815_n1149), .B(_abc_43815_n1154), .Y(_abc_43815_n1155) );
  AND2X2 AND2X2_2950 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4323), .B(REGFILE_SIM_reg_bank__abc_33898_n4322), .Y(REGFILE_SIM_reg_bank_reg_r12_27__FF_INPUT) );
  AND2X2 AND2X2_2951 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4326), .B(REGFILE_SIM_reg_bank__abc_33898_n4325), .Y(REGFILE_SIM_reg_bank_reg_r12_28__FF_INPUT) );
  AND2X2 AND2X2_2952 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4329), .B(REGFILE_SIM_reg_bank__abc_33898_n4328), .Y(REGFILE_SIM_reg_bank_reg_r12_29__FF_INPUT) );
  AND2X2 AND2X2_2953 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4332), .B(REGFILE_SIM_reg_bank__abc_33898_n4331), .Y(REGFILE_SIM_reg_bank_reg_r12_30__FF_INPUT) );
  AND2X2 AND2X2_2954 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4335), .B(REGFILE_SIM_reg_bank__abc_33898_n4334), .Y(REGFILE_SIM_reg_bank_reg_r12_31__FF_INPUT) );
  AND2X2 AND2X2_2955 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2599_1), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n4337) );
  AND2X2 AND2X2_2956 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4340), .B(REGFILE_SIM_reg_bank__abc_33898_n4338), .Y(REGFILE_SIM_reg_bank_reg_r11_0__FF_INPUT) );
  AND2X2 AND2X2_2957 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4343_1), .B(REGFILE_SIM_reg_bank__abc_33898_n4342), .Y(REGFILE_SIM_reg_bank_reg_r11_1__FF_INPUT) );
  AND2X2 AND2X2_2958 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4346), .B(REGFILE_SIM_reg_bank__abc_33898_n4345), .Y(REGFILE_SIM_reg_bank_reg_r11_2__FF_INPUT) );
  AND2X2 AND2X2_2959 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4349), .B(REGFILE_SIM_reg_bank__abc_33898_n4348), .Y(REGFILE_SIM_reg_bank_reg_r11_3__FF_INPUT) );
  AND2X2 AND2X2_296 ( .A(_abc_43815_n1129), .B(alu_op_r_2_), .Y(_abc_43815_n1156_1) );
  AND2X2 AND2X2_2960 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4352), .B(REGFILE_SIM_reg_bank__abc_33898_n4351), .Y(REGFILE_SIM_reg_bank_reg_r11_4__FF_INPUT) );
  AND2X2 AND2X2_2961 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4355), .B(REGFILE_SIM_reg_bank__abc_33898_n4354), .Y(REGFILE_SIM_reg_bank_reg_r11_5__FF_INPUT) );
  AND2X2 AND2X2_2962 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4358), .B(REGFILE_SIM_reg_bank__abc_33898_n4357), .Y(REGFILE_SIM_reg_bank_reg_r11_6__FF_INPUT) );
  AND2X2 AND2X2_2963 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4361), .B(REGFILE_SIM_reg_bank__abc_33898_n4360), .Y(REGFILE_SIM_reg_bank_reg_r11_7__FF_INPUT) );
  AND2X2 AND2X2_2964 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4364), .B(REGFILE_SIM_reg_bank__abc_33898_n4363), .Y(REGFILE_SIM_reg_bank_reg_r11_8__FF_INPUT) );
  AND2X2 AND2X2_2965 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4367), .B(REGFILE_SIM_reg_bank__abc_33898_n4366), .Y(REGFILE_SIM_reg_bank_reg_r11_9__FF_INPUT) );
  AND2X2 AND2X2_2966 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4370), .B(REGFILE_SIM_reg_bank__abc_33898_n4369), .Y(REGFILE_SIM_reg_bank_reg_r11_10__FF_INPUT) );
  AND2X2 AND2X2_2967 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4373_1), .B(REGFILE_SIM_reg_bank__abc_33898_n4372), .Y(REGFILE_SIM_reg_bank_reg_r11_11__FF_INPUT) );
  AND2X2 AND2X2_2968 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4376), .B(REGFILE_SIM_reg_bank__abc_33898_n4375), .Y(REGFILE_SIM_reg_bank_reg_r11_12__FF_INPUT) );
  AND2X2 AND2X2_2969 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4379), .B(REGFILE_SIM_reg_bank__abc_33898_n4378), .Y(REGFILE_SIM_reg_bank_reg_r11_13__FF_INPUT) );
  AND2X2 AND2X2_297 ( .A(_abc_43815_n1118), .B(_abc_43815_n1156_1), .Y(_abc_43815_n1157) );
  AND2X2 AND2X2_2970 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4382), .B(REGFILE_SIM_reg_bank__abc_33898_n4381), .Y(REGFILE_SIM_reg_bank_reg_r11_14__FF_INPUT) );
  AND2X2 AND2X2_2971 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4385), .B(REGFILE_SIM_reg_bank__abc_33898_n4384), .Y(REGFILE_SIM_reg_bank_reg_r11_15__FF_INPUT) );
  AND2X2 AND2X2_2972 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4388), .B(REGFILE_SIM_reg_bank__abc_33898_n4387), .Y(REGFILE_SIM_reg_bank_reg_r11_16__FF_INPUT) );
  AND2X2 AND2X2_2973 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4391), .B(REGFILE_SIM_reg_bank__abc_33898_n4390), .Y(REGFILE_SIM_reg_bank_reg_r11_17__FF_INPUT) );
  AND2X2 AND2X2_2974 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4394), .B(REGFILE_SIM_reg_bank__abc_33898_n4393), .Y(REGFILE_SIM_reg_bank_reg_r11_18__FF_INPUT) );
  AND2X2 AND2X2_2975 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4397), .B(REGFILE_SIM_reg_bank__abc_33898_n4396), .Y(REGFILE_SIM_reg_bank_reg_r11_19__FF_INPUT) );
  AND2X2 AND2X2_2976 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4400), .B(REGFILE_SIM_reg_bank__abc_33898_n4399), .Y(REGFILE_SIM_reg_bank_reg_r11_20__FF_INPUT) );
  AND2X2 AND2X2_2977 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4403_1), .B(REGFILE_SIM_reg_bank__abc_33898_n4402), .Y(REGFILE_SIM_reg_bank_reg_r11_21__FF_INPUT) );
  AND2X2 AND2X2_2978 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4406), .B(REGFILE_SIM_reg_bank__abc_33898_n4405), .Y(REGFILE_SIM_reg_bank_reg_r11_22__FF_INPUT) );
  AND2X2 AND2X2_2979 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4409), .B(REGFILE_SIM_reg_bank__abc_33898_n4408), .Y(REGFILE_SIM_reg_bank_reg_r11_23__FF_INPUT) );
  AND2X2 AND2X2_298 ( .A(_abc_43815_n1113), .B(_abc_43815_n1157), .Y(_abc_43815_n1158) );
  AND2X2 AND2X2_2980 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4412), .B(REGFILE_SIM_reg_bank__abc_33898_n4411), .Y(REGFILE_SIM_reg_bank_reg_r11_24__FF_INPUT) );
  AND2X2 AND2X2_2981 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4415), .B(REGFILE_SIM_reg_bank__abc_33898_n4414), .Y(REGFILE_SIM_reg_bank_reg_r11_25__FF_INPUT) );
  AND2X2 AND2X2_2982 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4418), .B(REGFILE_SIM_reg_bank__abc_33898_n4417), .Y(REGFILE_SIM_reg_bank_reg_r11_26__FF_INPUT) );
  AND2X2 AND2X2_2983 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4421), .B(REGFILE_SIM_reg_bank__abc_33898_n4420), .Y(REGFILE_SIM_reg_bank_reg_r11_27__FF_INPUT) );
  AND2X2 AND2X2_2984 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4424), .B(REGFILE_SIM_reg_bank__abc_33898_n4423), .Y(REGFILE_SIM_reg_bank_reg_r11_28__FF_INPUT) );
  AND2X2 AND2X2_2985 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4427), .B(REGFILE_SIM_reg_bank__abc_33898_n4426), .Y(REGFILE_SIM_reg_bank_reg_r11_29__FF_INPUT) );
  AND2X2 AND2X2_2986 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4430), .B(REGFILE_SIM_reg_bank__abc_33898_n4429), .Y(REGFILE_SIM_reg_bank_reg_r11_30__FF_INPUT) );
  AND2X2 AND2X2_2987 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4433_1), .B(REGFILE_SIM_reg_bank__abc_33898_n4432), .Y(REGFILE_SIM_reg_bank_reg_r11_31__FF_INPUT) );
  AND2X2 AND2X2_2988 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2698), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435) );
  AND2X2 AND2X2_2989 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4437) );
  AND2X2 AND2X2_299 ( .A(_abc_43815_n1158), .B(_abc_43815_n1106), .Y(_abc_43815_n1159) );
  AND2X2 AND2X2_2990 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4438), .B(REGFILE_SIM_reg_bank__abc_33898_n4436), .Y(REGFILE_SIM_reg_bank_reg_r10_0__FF_INPUT) );
  AND2X2 AND2X2_2991 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n4441) );
  AND2X2 AND2X2_2992 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4442), .B(REGFILE_SIM_reg_bank__abc_33898_n4440), .Y(REGFILE_SIM_reg_bank_reg_r10_1__FF_INPUT) );
  AND2X2 AND2X2_2993 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4445) );
  AND2X2 AND2X2_2994 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4446), .B(REGFILE_SIM_reg_bank__abc_33898_n4444), .Y(REGFILE_SIM_reg_bank_reg_r10_2__FF_INPUT) );
  AND2X2 AND2X2_2995 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4449) );
  AND2X2 AND2X2_2996 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4450), .B(REGFILE_SIM_reg_bank__abc_33898_n4448), .Y(REGFILE_SIM_reg_bank_reg_r10_3__FF_INPUT) );
  AND2X2 AND2X2_2997 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n4453) );
  AND2X2 AND2X2_2998 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4454), .B(REGFILE_SIM_reg_bank__abc_33898_n4452), .Y(REGFILE_SIM_reg_bank_reg_r10_4__FF_INPUT) );
  AND2X2 AND2X2_2999 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4457) );
  AND2X2 AND2X2_3 ( .A(_abc_43815_n622), .B(_abc_43815_n623), .Y(_abc_43815_n624_1) );
  AND2X2 AND2X2_30 ( .A(_abc_43815_n653), .B(_abc_43815_n647_1), .Y(_abc_43815_n659) );
  AND2X2 AND2X2_300 ( .A(alu_op_r_1_), .B(alu_op_r_0_), .Y(_abc_43815_n1161) );
  AND2X2 AND2X2_3000 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4458), .B(REGFILE_SIM_reg_bank__abc_33898_n4456), .Y(REGFILE_SIM_reg_bank_reg_r10_5__FF_INPUT) );
  AND2X2 AND2X2_3001 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4461) );
  AND2X2 AND2X2_3002 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4462), .B(REGFILE_SIM_reg_bank__abc_33898_n4460), .Y(REGFILE_SIM_reg_bank_reg_r10_6__FF_INPUT) );
  AND2X2 AND2X2_3003 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n4465) );
  AND2X2 AND2X2_3004 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4466), .B(REGFILE_SIM_reg_bank__abc_33898_n4464), .Y(REGFILE_SIM_reg_bank_reg_r10_7__FF_INPUT) );
  AND2X2 AND2X2_3005 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4469) );
  AND2X2 AND2X2_3006 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4470), .B(REGFILE_SIM_reg_bank__abc_33898_n4468), .Y(REGFILE_SIM_reg_bank_reg_r10_8__FF_INPUT) );
  AND2X2 AND2X2_3007 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4473) );
  AND2X2 AND2X2_3008 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4474), .B(REGFILE_SIM_reg_bank__abc_33898_n4472), .Y(REGFILE_SIM_reg_bank_reg_r10_9__FF_INPUT) );
  AND2X2 AND2X2_3009 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n4477) );
  AND2X2 AND2X2_301 ( .A(_abc_43815_n1130), .B(_abc_43815_n1161), .Y(_abc_43815_n1162) );
  AND2X2 AND2X2_3010 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4478), .B(REGFILE_SIM_reg_bank__abc_33898_n4476), .Y(REGFILE_SIM_reg_bank_reg_r10_10__FF_INPUT) );
  AND2X2 AND2X2_3011 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4481) );
  AND2X2 AND2X2_3012 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4482), .B(REGFILE_SIM_reg_bank__abc_33898_n4480), .Y(REGFILE_SIM_reg_bank_reg_r10_11__FF_INPUT) );
  AND2X2 AND2X2_3013 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4485) );
  AND2X2 AND2X2_3014 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4486), .B(REGFILE_SIM_reg_bank__abc_33898_n4484), .Y(REGFILE_SIM_reg_bank_reg_r10_12__FF_INPUT) );
  AND2X2 AND2X2_3015 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n4489) );
  AND2X2 AND2X2_3016 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4490), .B(REGFILE_SIM_reg_bank__abc_33898_n4488), .Y(REGFILE_SIM_reg_bank_reg_r10_13__FF_INPUT) );
  AND2X2 AND2X2_3017 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4493_1) );
  AND2X2 AND2X2_3018 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4494), .B(REGFILE_SIM_reg_bank__abc_33898_n4492), .Y(REGFILE_SIM_reg_bank_reg_r10_14__FF_INPUT) );
  AND2X2 AND2X2_3019 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4497) );
  AND2X2 AND2X2_302 ( .A(_abc_43815_n1113), .B(_abc_43815_n1162), .Y(_abc_43815_n1163) );
  AND2X2 AND2X2_3020 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4498), .B(REGFILE_SIM_reg_bank__abc_33898_n4496), .Y(REGFILE_SIM_reg_bank_reg_r10_15__FF_INPUT) );
  AND2X2 AND2X2_3021 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n4501) );
  AND2X2 AND2X2_3022 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4502), .B(REGFILE_SIM_reg_bank__abc_33898_n4500), .Y(REGFILE_SIM_reg_bank_reg_r10_16__FF_INPUT) );
  AND2X2 AND2X2_3023 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4505) );
  AND2X2 AND2X2_3024 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4506), .B(REGFILE_SIM_reg_bank__abc_33898_n4504), .Y(REGFILE_SIM_reg_bank_reg_r10_17__FF_INPUT) );
  AND2X2 AND2X2_3025 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4509) );
  AND2X2 AND2X2_3026 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4510), .B(REGFILE_SIM_reg_bank__abc_33898_n4508), .Y(REGFILE_SIM_reg_bank_reg_r10_18__FF_INPUT) );
  AND2X2 AND2X2_3027 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4513) );
  AND2X2 AND2X2_3028 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4514), .B(REGFILE_SIM_reg_bank__abc_33898_n4512), .Y(REGFILE_SIM_reg_bank_reg_r10_19__FF_INPUT) );
  AND2X2 AND2X2_3029 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4517) );
  AND2X2 AND2X2_303 ( .A(_abc_43815_n1163), .B(_abc_43815_n1106), .Y(_abc_43815_n1164) );
  AND2X2 AND2X2_3030 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4518), .B(REGFILE_SIM_reg_bank__abc_33898_n4516), .Y(REGFILE_SIM_reg_bank_reg_r10_20__FF_INPUT) );
  AND2X2 AND2X2_3031 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n4521) );
  AND2X2 AND2X2_3032 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4522), .B(REGFILE_SIM_reg_bank__abc_33898_n4520), .Y(REGFILE_SIM_reg_bank_reg_r10_21__FF_INPUT) );
  AND2X2 AND2X2_3033 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4525) );
  AND2X2 AND2X2_3034 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4526), .B(REGFILE_SIM_reg_bank__abc_33898_n4524), .Y(REGFILE_SIM_reg_bank_reg_r10_22__FF_INPUT) );
  AND2X2 AND2X2_3035 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4529) );
  AND2X2 AND2X2_3036 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4530), .B(REGFILE_SIM_reg_bank__abc_33898_n4528), .Y(REGFILE_SIM_reg_bank_reg_r10_23__FF_INPUT) );
  AND2X2 AND2X2_3037 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n4533) );
  AND2X2 AND2X2_3038 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4534), .B(REGFILE_SIM_reg_bank__abc_33898_n4532), .Y(REGFILE_SIM_reg_bank_reg_r10_24__FF_INPUT) );
  AND2X2 AND2X2_3039 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4537) );
  AND2X2 AND2X2_304 ( .A(_abc_43815_n1160), .B(_abc_43815_n1165), .Y(_abc_43815_n1166) );
  AND2X2 AND2X2_3040 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4538), .B(REGFILE_SIM_reg_bank__abc_33898_n4536), .Y(REGFILE_SIM_reg_bank_reg_r10_25__FF_INPUT) );
  AND2X2 AND2X2_3041 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4541) );
  AND2X2 AND2X2_3042 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4542), .B(REGFILE_SIM_reg_bank__abc_33898_n4540), .Y(REGFILE_SIM_reg_bank_reg_r10_26__FF_INPUT) );
  AND2X2 AND2X2_3043 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n4545) );
  AND2X2 AND2X2_3044 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4546), .B(REGFILE_SIM_reg_bank__abc_33898_n4544), .Y(REGFILE_SIM_reg_bank_reg_r10_27__FF_INPUT) );
  AND2X2 AND2X2_3045 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4549) );
  AND2X2 AND2X2_3046 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4550), .B(REGFILE_SIM_reg_bank__abc_33898_n4548), .Y(REGFILE_SIM_reg_bank_reg_r10_28__FF_INPUT) );
  AND2X2 AND2X2_3047 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4553_1) );
  AND2X2 AND2X2_3048 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4554), .B(REGFILE_SIM_reg_bank__abc_33898_n4552), .Y(REGFILE_SIM_reg_bank_reg_r10_29__FF_INPUT) );
  AND2X2 AND2X2_3049 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n4557) );
  AND2X2 AND2X2_305 ( .A(_abc_43815_n1155), .B(_abc_43815_n1166), .Y(_abc_43815_n1167) );
  AND2X2 AND2X2_3050 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4558), .B(REGFILE_SIM_reg_bank__abc_33898_n4556), .Y(REGFILE_SIM_reg_bank_reg_r10_30__FF_INPUT) );
  AND2X2 AND2X2_3051 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4561) );
  AND2X2 AND2X2_3052 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4562), .B(REGFILE_SIM_reg_bank__abc_33898_n4560), .Y(REGFILE_SIM_reg_bank_reg_r10_31__FF_INPUT) );
  AND2X2 AND2X2_3053 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2828), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564) );
  AND2X2 AND2X2_3054 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4566) );
  AND2X2 AND2X2_3055 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4567), .B(REGFILE_SIM_reg_bank__abc_33898_n4565), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_0__FF_INPUT) );
  AND2X2 AND2X2_3056 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n4570) );
  AND2X2 AND2X2_3057 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4571), .B(REGFILE_SIM_reg_bank__abc_33898_n4569), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_1__FF_INPUT) );
  AND2X2 AND2X2_3058 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4574) );
  AND2X2 AND2X2_3059 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4575), .B(REGFILE_SIM_reg_bank__abc_33898_n4573), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_2__FF_INPUT) );
  AND2X2 AND2X2_306 ( .A(_abc_43815_n1167), .B(_abc_43815_n1143), .Y(_abc_43815_n1168) );
  AND2X2 AND2X2_3060 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4578) );
  AND2X2 AND2X2_3061 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4579), .B(REGFILE_SIM_reg_bank__abc_33898_n4577), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_3__FF_INPUT) );
  AND2X2 AND2X2_3062 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n4582) );
  AND2X2 AND2X2_3063 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4583_1), .B(REGFILE_SIM_reg_bank__abc_33898_n4581), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_4__FF_INPUT) );
  AND2X2 AND2X2_3064 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4586) );
  AND2X2 AND2X2_3065 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4587), .B(REGFILE_SIM_reg_bank__abc_33898_n4585), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_5__FF_INPUT) );
  AND2X2 AND2X2_3066 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4590) );
  AND2X2 AND2X2_3067 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4591), .B(REGFILE_SIM_reg_bank__abc_33898_n4589), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_6__FF_INPUT) );
  AND2X2 AND2X2_3068 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n4594) );
  AND2X2 AND2X2_3069 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4595), .B(REGFILE_SIM_reg_bank__abc_33898_n4593), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_7__FF_INPUT) );
  AND2X2 AND2X2_307 ( .A(_abc_43815_n657), .B(_abc_43815_n1068), .Y(_abc_43815_n1169) );
  AND2X2 AND2X2_3070 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4598) );
  AND2X2 AND2X2_3071 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4599), .B(REGFILE_SIM_reg_bank__abc_33898_n4597), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_8__FF_INPUT) );
  AND2X2 AND2X2_3072 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4602) );
  AND2X2 AND2X2_3073 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4603), .B(REGFILE_SIM_reg_bank__abc_33898_n4601), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_9__FF_INPUT) );
  AND2X2 AND2X2_3074 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n4606) );
  AND2X2 AND2X2_3075 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4607), .B(REGFILE_SIM_reg_bank__abc_33898_n4605), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_10__FF_INPUT) );
  AND2X2 AND2X2_3076 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4610) );
  AND2X2 AND2X2_3077 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4611), .B(REGFILE_SIM_reg_bank__abc_33898_n4609), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_11__FF_INPUT) );
  AND2X2 AND2X2_3078 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4614) );
  AND2X2 AND2X2_3079 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4615), .B(REGFILE_SIM_reg_bank__abc_33898_n4613_1), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_12__FF_INPUT) );
  AND2X2 AND2X2_308 ( .A(_abc_43815_n1067), .B(_abc_43815_n624_1), .Y(_abc_43815_n1170) );
  AND2X2 AND2X2_3080 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n4618) );
  AND2X2 AND2X2_3081 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4619), .B(REGFILE_SIM_reg_bank__abc_33898_n4617), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_13__FF_INPUT) );
  AND2X2 AND2X2_3082 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4622) );
  AND2X2 AND2X2_3083 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4623), .B(REGFILE_SIM_reg_bank__abc_33898_n4621), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_14__FF_INPUT) );
  AND2X2 AND2X2_3084 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4626) );
  AND2X2 AND2X2_3085 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4627), .B(REGFILE_SIM_reg_bank__abc_33898_n4625), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_15__FF_INPUT) );
  AND2X2 AND2X2_3086 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n4630) );
  AND2X2 AND2X2_3087 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4631), .B(REGFILE_SIM_reg_bank__abc_33898_n4629), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_16__FF_INPUT) );
  AND2X2 AND2X2_3088 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4634) );
  AND2X2 AND2X2_3089 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4635), .B(REGFILE_SIM_reg_bank__abc_33898_n4633), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_17__FF_INPUT) );
  AND2X2 AND2X2_309 ( .A(_abc_43815_n1172_1_bF_buf4), .B(_abc_43815_n669), .Y(_abc_43815_n1173_1) );
  AND2X2 AND2X2_3090 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4638) );
  AND2X2 AND2X2_3091 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4639), .B(REGFILE_SIM_reg_bank__abc_33898_n4637), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_18__FF_INPUT) );
  AND2X2 AND2X2_3092 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4642) );
  AND2X2 AND2X2_3093 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4643_1), .B(REGFILE_SIM_reg_bank__abc_33898_n4641), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_19__FF_INPUT) );
  AND2X2 AND2X2_3094 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4646) );
  AND2X2 AND2X2_3095 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4647), .B(REGFILE_SIM_reg_bank__abc_33898_n4645), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_20__FF_INPUT) );
  AND2X2 AND2X2_3096 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n4650) );
  AND2X2 AND2X2_3097 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4651), .B(REGFILE_SIM_reg_bank__abc_33898_n4649), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_21__FF_INPUT) );
  AND2X2 AND2X2_3098 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4654) );
  AND2X2 AND2X2_3099 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4655), .B(REGFILE_SIM_reg_bank__abc_33898_n4653), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_22__FF_INPUT) );
  AND2X2 AND2X2_31 ( .A(_abc_43815_n659), .B(_abc_43815_n656), .Y(_abc_43815_n660) );
  AND2X2 AND2X2_310 ( .A(_abc_43815_n663), .B(_abc_43815_n1173_1), .Y(_abc_43815_n1174) );
  AND2X2 AND2X2_3100 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4658) );
  AND2X2 AND2X2_3101 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4659), .B(REGFILE_SIM_reg_bank__abc_33898_n4657), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_23__FF_INPUT) );
  AND2X2 AND2X2_3102 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n4662) );
  AND2X2 AND2X2_3103 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4663), .B(REGFILE_SIM_reg_bank__abc_33898_n4661), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_24__FF_INPUT) );
  AND2X2 AND2X2_3104 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4666) );
  AND2X2 AND2X2_3105 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4667), .B(REGFILE_SIM_reg_bank__abc_33898_n4665), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_25__FF_INPUT) );
  AND2X2 AND2X2_3106 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4670) );
  AND2X2 AND2X2_3107 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4671), .B(REGFILE_SIM_reg_bank__abc_33898_n4669), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_26__FF_INPUT) );
  AND2X2 AND2X2_3108 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n4674) );
  AND2X2 AND2X2_3109 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4675), .B(REGFILE_SIM_reg_bank__abc_33898_n4673_1), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_27__FF_INPUT) );
  AND2X2 AND2X2_311 ( .A(_abc_43815_n1150), .B(_abc_43815_n1156_1), .Y(_abc_43815_n1175) );
  AND2X2 AND2X2_3110 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4678) );
  AND2X2 AND2X2_3111 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4679), .B(REGFILE_SIM_reg_bank__abc_33898_n4677), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_28__FF_INPUT) );
  AND2X2 AND2X2_3112 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4682) );
  AND2X2 AND2X2_3113 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4683), .B(REGFILE_SIM_reg_bank__abc_33898_n4681), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_29__FF_INPUT) );
  AND2X2 AND2X2_3114 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n4686) );
  AND2X2 AND2X2_3115 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4687), .B(REGFILE_SIM_reg_bank__abc_33898_n4685), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_30__FF_INPUT) );
  AND2X2 AND2X2_3116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4690) );
  AND2X2 AND2X2_3117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4691), .B(REGFILE_SIM_reg_bank__abc_33898_n4689), .Y(REGFILE_SIM_reg_bank_reg_r9_lr_31__FF_INPUT) );
  AND2X2 AND2X2_3118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4238), .B(REGFILE_SIM_reg_bank__abc_33898_n2598), .Y(REGFILE_SIM_reg_bank__abc_33898_n4693) );
  AND2X2 AND2X2_3119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4696), .B(REGFILE_SIM_reg_bank__abc_33898_n4694), .Y(REGFILE_SIM_reg_bank_reg_r8_0__FF_INPUT) );
  AND2X2 AND2X2_312 ( .A(_abc_43815_n1113), .B(_abc_43815_n1175), .Y(_abc_43815_n1176) );
  AND2X2 AND2X2_3120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4699), .B(REGFILE_SIM_reg_bank__abc_33898_n4698), .Y(REGFILE_SIM_reg_bank_reg_r8_1__FF_INPUT) );
  AND2X2 AND2X2_3121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4702), .B(REGFILE_SIM_reg_bank__abc_33898_n4701), .Y(REGFILE_SIM_reg_bank_reg_r8_2__FF_INPUT) );
  AND2X2 AND2X2_3122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4705), .B(REGFILE_SIM_reg_bank__abc_33898_n4704), .Y(REGFILE_SIM_reg_bank_reg_r8_3__FF_INPUT) );
  AND2X2 AND2X2_3123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4708), .B(REGFILE_SIM_reg_bank__abc_33898_n4707), .Y(REGFILE_SIM_reg_bank_reg_r8_4__FF_INPUT) );
  AND2X2 AND2X2_3124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4711), .B(REGFILE_SIM_reg_bank__abc_33898_n4710), .Y(REGFILE_SIM_reg_bank_reg_r8_5__FF_INPUT) );
  AND2X2 AND2X2_3125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4714), .B(REGFILE_SIM_reg_bank__abc_33898_n4713), .Y(REGFILE_SIM_reg_bank_reg_r8_6__FF_INPUT) );
  AND2X2 AND2X2_3126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4717), .B(REGFILE_SIM_reg_bank__abc_33898_n4716), .Y(REGFILE_SIM_reg_bank_reg_r8_7__FF_INPUT) );
  AND2X2 AND2X2_3127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4720), .B(REGFILE_SIM_reg_bank__abc_33898_n4719), .Y(REGFILE_SIM_reg_bank_reg_r8_8__FF_INPUT) );
  AND2X2 AND2X2_3128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4723), .B(REGFILE_SIM_reg_bank__abc_33898_n4722), .Y(REGFILE_SIM_reg_bank_reg_r8_9__FF_INPUT) );
  AND2X2 AND2X2_3129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4726), .B(REGFILE_SIM_reg_bank__abc_33898_n4725), .Y(REGFILE_SIM_reg_bank_reg_r8_10__FF_INPUT) );
  AND2X2 AND2X2_313 ( .A(_abc_43815_n1176), .B(_abc_43815_n1106), .Y(_abc_43815_n1177) );
  AND2X2 AND2X2_3130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4729), .B(REGFILE_SIM_reg_bank__abc_33898_n4728), .Y(REGFILE_SIM_reg_bank_reg_r8_11__FF_INPUT) );
  AND2X2 AND2X2_3131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4732), .B(REGFILE_SIM_reg_bank__abc_33898_n4731), .Y(REGFILE_SIM_reg_bank_reg_r8_12__FF_INPUT) );
  AND2X2 AND2X2_3132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4735), .B(REGFILE_SIM_reg_bank__abc_33898_n4734), .Y(REGFILE_SIM_reg_bank_reg_r8_13__FF_INPUT) );
  AND2X2 AND2X2_3133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4738), .B(REGFILE_SIM_reg_bank__abc_33898_n4737), .Y(REGFILE_SIM_reg_bank_reg_r8_14__FF_INPUT) );
  AND2X2 AND2X2_3134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4741), .B(REGFILE_SIM_reg_bank__abc_33898_n4740), .Y(REGFILE_SIM_reg_bank_reg_r8_15__FF_INPUT) );
  AND2X2 AND2X2_3135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4744), .B(REGFILE_SIM_reg_bank__abc_33898_n4743), .Y(REGFILE_SIM_reg_bank_reg_r8_16__FF_INPUT) );
  AND2X2 AND2X2_3136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4747), .B(REGFILE_SIM_reg_bank__abc_33898_n4746), .Y(REGFILE_SIM_reg_bank_reg_r8_17__FF_INPUT) );
  AND2X2 AND2X2_3137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4750), .B(REGFILE_SIM_reg_bank__abc_33898_n4749), .Y(REGFILE_SIM_reg_bank_reg_r8_18__FF_INPUT) );
  AND2X2 AND2X2_3138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4753), .B(REGFILE_SIM_reg_bank__abc_33898_n4752), .Y(REGFILE_SIM_reg_bank_reg_r8_19__FF_INPUT) );
  AND2X2 AND2X2_3139 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4756), .B(REGFILE_SIM_reg_bank__abc_33898_n4755), .Y(REGFILE_SIM_reg_bank_reg_r8_20__FF_INPUT) );
  AND2X2 AND2X2_314 ( .A(_abc_43815_n1043_1), .B(_abc_43815_n983), .Y(_abc_43815_n1179) );
  AND2X2 AND2X2_3140 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4759), .B(REGFILE_SIM_reg_bank__abc_33898_n4758), .Y(REGFILE_SIM_reg_bank_reg_r8_21__FF_INPUT) );
  AND2X2 AND2X2_3141 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4762), .B(REGFILE_SIM_reg_bank__abc_33898_n4761), .Y(REGFILE_SIM_reg_bank_reg_r8_22__FF_INPUT) );
  AND2X2 AND2X2_3142 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4765), .B(REGFILE_SIM_reg_bank__abc_33898_n4764), .Y(REGFILE_SIM_reg_bank_reg_r8_23__FF_INPUT) );
  AND2X2 AND2X2_3143 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4768), .B(REGFILE_SIM_reg_bank__abc_33898_n4767), .Y(REGFILE_SIM_reg_bank_reg_r8_24__FF_INPUT) );
  AND2X2 AND2X2_3144 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4771), .B(REGFILE_SIM_reg_bank__abc_33898_n4770), .Y(REGFILE_SIM_reg_bank_reg_r8_25__FF_INPUT) );
  AND2X2 AND2X2_3145 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4774), .B(REGFILE_SIM_reg_bank__abc_33898_n4773), .Y(REGFILE_SIM_reg_bank_reg_r8_26__FF_INPUT) );
  AND2X2 AND2X2_3146 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4777), .B(REGFILE_SIM_reg_bank__abc_33898_n4776), .Y(REGFILE_SIM_reg_bank_reg_r8_27__FF_INPUT) );
  AND2X2 AND2X2_3147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4780), .B(REGFILE_SIM_reg_bank__abc_33898_n4779), .Y(REGFILE_SIM_reg_bank_reg_r8_28__FF_INPUT) );
  AND2X2 AND2X2_3148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4783), .B(REGFILE_SIM_reg_bank__abc_33898_n4782), .Y(REGFILE_SIM_reg_bank_reg_r8_29__FF_INPUT) );
  AND2X2 AND2X2_3149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4786), .B(REGFILE_SIM_reg_bank__abc_33898_n4785), .Y(REGFILE_SIM_reg_bank_reg_r8_30__FF_INPUT) );
  AND2X2 AND2X2_315 ( .A(_abc_43815_n1179), .B(_abc_43815_n1112), .Y(_abc_43815_n1180) );
  AND2X2 AND2X2_3150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4789), .B(REGFILE_SIM_reg_bank__abc_33898_n4788), .Y(REGFILE_SIM_reg_bank_reg_r8_31__FF_INPUT) );
  AND2X2 AND2X2_3151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3058), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n4791) );
  AND2X2 AND2X2_3152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4794), .B(REGFILE_SIM_reg_bank__abc_33898_n4792), .Y(REGFILE_SIM_reg_bank_reg_r7_0__FF_INPUT) );
  AND2X2 AND2X2_3153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4797), .B(REGFILE_SIM_reg_bank__abc_33898_n4796), .Y(REGFILE_SIM_reg_bank_reg_r7_1__FF_INPUT) );
  AND2X2 AND2X2_3154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4800), .B(REGFILE_SIM_reg_bank__abc_33898_n4799), .Y(REGFILE_SIM_reg_bank_reg_r7_2__FF_INPUT) );
  AND2X2 AND2X2_3155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4803), .B(REGFILE_SIM_reg_bank__abc_33898_n4802), .Y(REGFILE_SIM_reg_bank_reg_r7_3__FF_INPUT) );
  AND2X2 AND2X2_3156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4806), .B(REGFILE_SIM_reg_bank__abc_33898_n4805), .Y(REGFILE_SIM_reg_bank_reg_r7_4__FF_INPUT) );
  AND2X2 AND2X2_3157 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4809), .B(REGFILE_SIM_reg_bank__abc_33898_n4808), .Y(REGFILE_SIM_reg_bank_reg_r7_5__FF_INPUT) );
  AND2X2 AND2X2_3158 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4812), .B(REGFILE_SIM_reg_bank__abc_33898_n4811), .Y(REGFILE_SIM_reg_bank_reg_r7_6__FF_INPUT) );
  AND2X2 AND2X2_3159 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4815), .B(REGFILE_SIM_reg_bank__abc_33898_n4814), .Y(REGFILE_SIM_reg_bank_reg_r7_7__FF_INPUT) );
  AND2X2 AND2X2_316 ( .A(_abc_43815_n1178_1), .B(_abc_43815_n1181), .Y(_abc_43815_n1182) );
  AND2X2 AND2X2_3160 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4818), .B(REGFILE_SIM_reg_bank__abc_33898_n4817), .Y(REGFILE_SIM_reg_bank_reg_r7_8__FF_INPUT) );
  AND2X2 AND2X2_3161 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4821), .B(REGFILE_SIM_reg_bank__abc_33898_n4820), .Y(REGFILE_SIM_reg_bank_reg_r7_9__FF_INPUT) );
  AND2X2 AND2X2_3162 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4824), .B(REGFILE_SIM_reg_bank__abc_33898_n4823_1), .Y(REGFILE_SIM_reg_bank_reg_r7_10__FF_INPUT) );
  AND2X2 AND2X2_3163 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4827), .B(REGFILE_SIM_reg_bank__abc_33898_n4826), .Y(REGFILE_SIM_reg_bank_reg_r7_11__FF_INPUT) );
  AND2X2 AND2X2_3164 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4830), .B(REGFILE_SIM_reg_bank__abc_33898_n4829), .Y(REGFILE_SIM_reg_bank_reg_r7_12__FF_INPUT) );
  AND2X2 AND2X2_3165 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4833), .B(REGFILE_SIM_reg_bank__abc_33898_n4832), .Y(REGFILE_SIM_reg_bank_reg_r7_13__FF_INPUT) );
  AND2X2 AND2X2_3166 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4836), .B(REGFILE_SIM_reg_bank__abc_33898_n4835), .Y(REGFILE_SIM_reg_bank_reg_r7_14__FF_INPUT) );
  AND2X2 AND2X2_3167 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4839), .B(REGFILE_SIM_reg_bank__abc_33898_n4838), .Y(REGFILE_SIM_reg_bank_reg_r7_15__FF_INPUT) );
  AND2X2 AND2X2_3168 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4842), .B(REGFILE_SIM_reg_bank__abc_33898_n4841), .Y(REGFILE_SIM_reg_bank_reg_r7_16__FF_INPUT) );
  AND2X2 AND2X2_3169 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4845), .B(REGFILE_SIM_reg_bank__abc_33898_n4844), .Y(REGFILE_SIM_reg_bank_reg_r7_17__FF_INPUT) );
  AND2X2 AND2X2_317 ( .A(_abc_43815_n1179), .B(_abc_43815_n1137), .Y(_abc_43815_n1183) );
  AND2X2 AND2X2_3170 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4848), .B(REGFILE_SIM_reg_bank__abc_33898_n4847), .Y(REGFILE_SIM_reg_bank_reg_r7_18__FF_INPUT) );
  AND2X2 AND2X2_3171 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4851), .B(REGFILE_SIM_reg_bank__abc_33898_n4850), .Y(REGFILE_SIM_reg_bank_reg_r7_19__FF_INPUT) );
  AND2X2 AND2X2_3172 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4854), .B(REGFILE_SIM_reg_bank__abc_33898_n4853_1), .Y(REGFILE_SIM_reg_bank_reg_r7_20__FF_INPUT) );
  AND2X2 AND2X2_3173 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4857), .B(REGFILE_SIM_reg_bank__abc_33898_n4856), .Y(REGFILE_SIM_reg_bank_reg_r7_21__FF_INPUT) );
  AND2X2 AND2X2_3174 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4860), .B(REGFILE_SIM_reg_bank__abc_33898_n4859), .Y(REGFILE_SIM_reg_bank_reg_r7_22__FF_INPUT) );
  AND2X2 AND2X2_3175 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4863), .B(REGFILE_SIM_reg_bank__abc_33898_n4862), .Y(REGFILE_SIM_reg_bank_reg_r7_23__FF_INPUT) );
  AND2X2 AND2X2_3176 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4866), .B(REGFILE_SIM_reg_bank__abc_33898_n4865), .Y(REGFILE_SIM_reg_bank_reg_r7_24__FF_INPUT) );
  AND2X2 AND2X2_3177 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4869), .B(REGFILE_SIM_reg_bank__abc_33898_n4868), .Y(REGFILE_SIM_reg_bank_reg_r7_25__FF_INPUT) );
  AND2X2 AND2X2_3178 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4872), .B(REGFILE_SIM_reg_bank__abc_33898_n4871), .Y(REGFILE_SIM_reg_bank_reg_r7_26__FF_INPUT) );
  AND2X2 AND2X2_3179 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4875), .B(REGFILE_SIM_reg_bank__abc_33898_n4874), .Y(REGFILE_SIM_reg_bank_reg_r7_27__FF_INPUT) );
  AND2X2 AND2X2_318 ( .A(_abc_43815_n1179), .B(_abc_43815_n1123), .Y(_abc_43815_n1184) );
  AND2X2 AND2X2_3180 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4878), .B(REGFILE_SIM_reg_bank__abc_33898_n4877), .Y(REGFILE_SIM_reg_bank_reg_r7_28__FF_INPUT) );
  AND2X2 AND2X2_3181 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4881), .B(REGFILE_SIM_reg_bank__abc_33898_n4880), .Y(REGFILE_SIM_reg_bank_reg_r7_29__FF_INPUT) );
  AND2X2 AND2X2_3182 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4884), .B(REGFILE_SIM_reg_bank__abc_33898_n4883_1), .Y(REGFILE_SIM_reg_bank_reg_r7_30__FF_INPUT) );
  AND2X2 AND2X2_3183 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4887), .B(REGFILE_SIM_reg_bank__abc_33898_n4886), .Y(REGFILE_SIM_reg_bank_reg_r7_31__FF_INPUT) );
  AND2X2 AND2X2_3184 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3157), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889) );
  AND2X2 AND2X2_3185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4891) );
  AND2X2 AND2X2_3186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4892), .B(REGFILE_SIM_reg_bank__abc_33898_n4890), .Y(REGFILE_SIM_reg_bank_reg_r6_0__FF_INPUT) );
  AND2X2 AND2X2_3187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n4895) );
  AND2X2 AND2X2_3188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4896), .B(REGFILE_SIM_reg_bank__abc_33898_n4894), .Y(REGFILE_SIM_reg_bank_reg_r6_1__FF_INPUT) );
  AND2X2 AND2X2_3189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4899) );
  AND2X2 AND2X2_319 ( .A(_abc_43815_n1186_1), .B(_abc_43815_n1182), .Y(_abc_43815_n1187) );
  AND2X2 AND2X2_3190 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4900), .B(REGFILE_SIM_reg_bank__abc_33898_n4898), .Y(REGFILE_SIM_reg_bank_reg_r6_2__FF_INPUT) );
  AND2X2 AND2X2_3191 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4903) );
  AND2X2 AND2X2_3192 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4904), .B(REGFILE_SIM_reg_bank__abc_33898_n4902), .Y(REGFILE_SIM_reg_bank_reg_r6_3__FF_INPUT) );
  AND2X2 AND2X2_3193 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n4907) );
  AND2X2 AND2X2_3194 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4908), .B(REGFILE_SIM_reg_bank__abc_33898_n4906), .Y(REGFILE_SIM_reg_bank_reg_r6_4__FF_INPUT) );
  AND2X2 AND2X2_3195 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4911) );
  AND2X2 AND2X2_3196 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4912), .B(REGFILE_SIM_reg_bank__abc_33898_n4910), .Y(REGFILE_SIM_reg_bank_reg_r6_5__FF_INPUT) );
  AND2X2 AND2X2_3197 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4915) );
  AND2X2 AND2X2_3198 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4916), .B(REGFILE_SIM_reg_bank__abc_33898_n4914), .Y(REGFILE_SIM_reg_bank_reg_r6_6__FF_INPUT) );
  AND2X2 AND2X2_3199 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n4919) );
  AND2X2 AND2X2_32 ( .A(_abc_43815_n631), .B(_abc_43815_n638), .Y(_abc_43815_n666) );
  AND2X2 AND2X2_320 ( .A(_abc_43815_n1174), .B(_abc_43815_n1187), .Y(_abc_43815_n1188) );
  AND2X2 AND2X2_3200 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4920), .B(REGFILE_SIM_reg_bank__abc_33898_n4918), .Y(REGFILE_SIM_reg_bank_reg_r6_7__FF_INPUT) );
  AND2X2 AND2X2_3201 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4923) );
  AND2X2 AND2X2_3202 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4924), .B(REGFILE_SIM_reg_bank__abc_33898_n4922), .Y(REGFILE_SIM_reg_bank_reg_r6_8__FF_INPUT) );
  AND2X2 AND2X2_3203 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4927) );
  AND2X2 AND2X2_3204 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4928), .B(REGFILE_SIM_reg_bank__abc_33898_n4926), .Y(REGFILE_SIM_reg_bank_reg_r6_9__FF_INPUT) );
  AND2X2 AND2X2_3205 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n4931) );
  AND2X2 AND2X2_3206 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4932), .B(REGFILE_SIM_reg_bank__abc_33898_n4930), .Y(REGFILE_SIM_reg_bank_reg_r6_10__FF_INPUT) );
  AND2X2 AND2X2_3207 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4935) );
  AND2X2 AND2X2_3208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4936), .B(REGFILE_SIM_reg_bank__abc_33898_n4934), .Y(REGFILE_SIM_reg_bank_reg_r6_11__FF_INPUT) );
  AND2X2 AND2X2_3209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4939) );
  AND2X2 AND2X2_321 ( .A(_abc_43815_n1168), .B(_abc_43815_n1188), .Y(_abc_43815_n1189_1) );
  AND2X2 AND2X2_3210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4940), .B(REGFILE_SIM_reg_bank__abc_33898_n4938), .Y(REGFILE_SIM_reg_bank_reg_r6_12__FF_INPUT) );
  AND2X2 AND2X2_3211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n4943_1) );
  AND2X2 AND2X2_3212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4944), .B(REGFILE_SIM_reg_bank__abc_33898_n4942), .Y(REGFILE_SIM_reg_bank_reg_r6_13__FF_INPUT) );
  AND2X2 AND2X2_3213 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4947) );
  AND2X2 AND2X2_3214 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4948), .B(REGFILE_SIM_reg_bank__abc_33898_n4946), .Y(REGFILE_SIM_reg_bank_reg_r6_14__FF_INPUT) );
  AND2X2 AND2X2_3215 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4951) );
  AND2X2 AND2X2_3216 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4952), .B(REGFILE_SIM_reg_bank__abc_33898_n4950), .Y(REGFILE_SIM_reg_bank_reg_r6_15__FF_INPUT) );
  AND2X2 AND2X2_3217 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n4955) );
  AND2X2 AND2X2_3218 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4956), .B(REGFILE_SIM_reg_bank__abc_33898_n4954), .Y(REGFILE_SIM_reg_bank_reg_r6_16__FF_INPUT) );
  AND2X2 AND2X2_3219 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4959) );
  AND2X2 AND2X2_322 ( .A(_abc_43815_n1105), .B(_abc_43815_n1189_1), .Y(_abc_43815_n1190) );
  AND2X2 AND2X2_3220 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4960), .B(REGFILE_SIM_reg_bank__abc_33898_n4958), .Y(REGFILE_SIM_reg_bank_reg_r6_17__FF_INPUT) );
  AND2X2 AND2X2_3221 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4963) );
  AND2X2 AND2X2_3222 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4964), .B(REGFILE_SIM_reg_bank__abc_33898_n4962), .Y(REGFILE_SIM_reg_bank_reg_r6_18__FF_INPUT) );
  AND2X2 AND2X2_3223 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4967) );
  AND2X2 AND2X2_3224 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4968), .B(REGFILE_SIM_reg_bank__abc_33898_n4966), .Y(REGFILE_SIM_reg_bank_reg_r6_19__FF_INPUT) );
  AND2X2 AND2X2_3225 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4971) );
  AND2X2 AND2X2_3226 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4972), .B(REGFILE_SIM_reg_bank__abc_33898_n4970), .Y(REGFILE_SIM_reg_bank_reg_r6_20__FF_INPUT) );
  AND2X2 AND2X2_3227 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n4975) );
  AND2X2 AND2X2_3228 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4976), .B(REGFILE_SIM_reg_bank__abc_33898_n4974), .Y(REGFILE_SIM_reg_bank_reg_r6_21__FF_INPUT) );
  AND2X2 AND2X2_3229 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4979) );
  AND2X2 AND2X2_323 ( .A(_abc_43815_n1193), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .Y(_abc_43815_n1194) );
  AND2X2 AND2X2_3230 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4980), .B(REGFILE_SIM_reg_bank__abc_33898_n4978), .Y(REGFILE_SIM_reg_bank_reg_r6_22__FF_INPUT) );
  AND2X2 AND2X2_3231 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4983) );
  AND2X2 AND2X2_3232 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4984), .B(REGFILE_SIM_reg_bank__abc_33898_n4982), .Y(REGFILE_SIM_reg_bank_reg_r6_23__FF_INPUT) );
  AND2X2 AND2X2_3233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n4987) );
  AND2X2 AND2X2_3234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4988), .B(REGFILE_SIM_reg_bank__abc_33898_n4986), .Y(REGFILE_SIM_reg_bank_reg_r6_24__FF_INPUT) );
  AND2X2 AND2X2_3235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4991) );
  AND2X2 AND2X2_3236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4992), .B(REGFILE_SIM_reg_bank__abc_33898_n4990), .Y(REGFILE_SIM_reg_bank_reg_r6_25__FF_INPUT) );
  AND2X2 AND2X2_3237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4995) );
  AND2X2 AND2X2_3238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4996), .B(REGFILE_SIM_reg_bank__abc_33898_n4994), .Y(REGFILE_SIM_reg_bank_reg_r6_26__FF_INPUT) );
  AND2X2 AND2X2_3239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n4999) );
  AND2X2 AND2X2_324 ( .A(_abc_43815_n1098), .B(_abc_43815_n1196), .Y(_abc_43815_n1197) );
  AND2X2 AND2X2_3240 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5000), .B(REGFILE_SIM_reg_bank__abc_33898_n4998), .Y(REGFILE_SIM_reg_bank_reg_r6_27__FF_INPUT) );
  AND2X2 AND2X2_3241 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5003_1) );
  AND2X2 AND2X2_3242 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5004), .B(REGFILE_SIM_reg_bank__abc_33898_n5002), .Y(REGFILE_SIM_reg_bank_reg_r6_28__FF_INPUT) );
  AND2X2 AND2X2_3243 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5007) );
  AND2X2 AND2X2_3244 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5008), .B(REGFILE_SIM_reg_bank__abc_33898_n5006), .Y(REGFILE_SIM_reg_bank_reg_r6_29__FF_INPUT) );
  AND2X2 AND2X2_3245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n5011) );
  AND2X2 AND2X2_3246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5012), .B(REGFILE_SIM_reg_bank__abc_33898_n5010), .Y(REGFILE_SIM_reg_bank_reg_r6_30__FF_INPUT) );
  AND2X2 AND2X2_3247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5015) );
  AND2X2 AND2X2_3248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5016), .B(REGFILE_SIM_reg_bank__abc_33898_n5014), .Y(REGFILE_SIM_reg_bank_reg_r6_31__FF_INPUT) );
  AND2X2 AND2X2_3249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3287), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018) );
  AND2X2 AND2X2_325 ( .A(_abc_43815_n1198), .B(_abc_43815_n1199), .Y(_abc_43815_n1200) );
  AND2X2 AND2X2_3250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2105_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5020) );
  AND2X2 AND2X2_3251 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5021), .B(REGFILE_SIM_reg_bank__abc_33898_n5019), .Y(REGFILE_SIM_reg_bank_reg_r5_0__FF_INPUT) );
  AND2X2 AND2X2_3252 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2110), .Y(REGFILE_SIM_reg_bank__abc_33898_n5024) );
  AND2X2 AND2X2_3253 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5025), .B(REGFILE_SIM_reg_bank__abc_33898_n5023), .Y(REGFILE_SIM_reg_bank_reg_r5_1__FF_INPUT) );
  AND2X2 AND2X2_3254 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2115_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5028) );
  AND2X2 AND2X2_3255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5029), .B(REGFILE_SIM_reg_bank__abc_33898_n5027), .Y(REGFILE_SIM_reg_bank_reg_r5_2__FF_INPUT) );
  AND2X2 AND2X2_3256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2120_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5032) );
  AND2X2 AND2X2_3257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5033_1), .B(REGFILE_SIM_reg_bank__abc_33898_n5031), .Y(REGFILE_SIM_reg_bank_reg_r5_3__FF_INPUT) );
  AND2X2 AND2X2_3258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2125), .Y(REGFILE_SIM_reg_bank__abc_33898_n5036) );
  AND2X2 AND2X2_3259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5037), .B(REGFILE_SIM_reg_bank__abc_33898_n5035), .Y(REGFILE_SIM_reg_bank_reg_r5_4__FF_INPUT) );
  AND2X2 AND2X2_326 ( .A(_abc_43815_n1201), .B(_abc_43815_n1108_1), .Y(_abc_43815_n1202) );
  AND2X2 AND2X2_3260 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2130_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5040) );
  AND2X2 AND2X2_3261 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5041), .B(REGFILE_SIM_reg_bank__abc_33898_n5039), .Y(REGFILE_SIM_reg_bank_reg_r5_5__FF_INPUT) );
  AND2X2 AND2X2_3262 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2135_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5044) );
  AND2X2 AND2X2_3263 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5045), .B(REGFILE_SIM_reg_bank__abc_33898_n5043), .Y(REGFILE_SIM_reg_bank_reg_r5_6__FF_INPUT) );
  AND2X2 AND2X2_3264 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2140), .Y(REGFILE_SIM_reg_bank__abc_33898_n5048) );
  AND2X2 AND2X2_3265 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5049), .B(REGFILE_SIM_reg_bank__abc_33898_n5047), .Y(REGFILE_SIM_reg_bank_reg_r5_7__FF_INPUT) );
  AND2X2 AND2X2_3266 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2145_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5052) );
  AND2X2 AND2X2_3267 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5053), .B(REGFILE_SIM_reg_bank__abc_33898_n5051), .Y(REGFILE_SIM_reg_bank_reg_r5_8__FF_INPUT) );
  AND2X2 AND2X2_3268 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2150_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5056) );
  AND2X2 AND2X2_3269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5057), .B(REGFILE_SIM_reg_bank__abc_33898_n5055), .Y(REGFILE_SIM_reg_bank_reg_r5_9__FF_INPUT) );
  AND2X2 AND2X2_327 ( .A(_abc_43815_n1200), .B(_abc_43815_n1202), .Y(_abc_43815_n1203) );
  AND2X2 AND2X2_3270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2155), .Y(REGFILE_SIM_reg_bank__abc_33898_n5060) );
  AND2X2 AND2X2_3271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5061), .B(REGFILE_SIM_reg_bank__abc_33898_n5059), .Y(REGFILE_SIM_reg_bank_reg_r5_10__FF_INPUT) );
  AND2X2 AND2X2_3272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2160_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5064) );
  AND2X2 AND2X2_3273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5065), .B(REGFILE_SIM_reg_bank__abc_33898_n5063_1), .Y(REGFILE_SIM_reg_bank_reg_r5_11__FF_INPUT) );
  AND2X2 AND2X2_3274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2165_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5068) );
  AND2X2 AND2X2_3275 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5069), .B(REGFILE_SIM_reg_bank__abc_33898_n5067), .Y(REGFILE_SIM_reg_bank_reg_r5_12__FF_INPUT) );
  AND2X2 AND2X2_3276 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2170), .Y(REGFILE_SIM_reg_bank__abc_33898_n5072) );
  AND2X2 AND2X2_3277 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5073), .B(REGFILE_SIM_reg_bank__abc_33898_n5071), .Y(REGFILE_SIM_reg_bank_reg_r5_13__FF_INPUT) );
  AND2X2 AND2X2_3278 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2175_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5076) );
  AND2X2 AND2X2_3279 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5077), .B(REGFILE_SIM_reg_bank__abc_33898_n5075), .Y(REGFILE_SIM_reg_bank_reg_r5_14__FF_INPUT) );
  AND2X2 AND2X2_328 ( .A(_abc_43815_n1205_1), .B(_abc_43815_n1206_1), .Y(_abc_43815_n1207) );
  AND2X2 AND2X2_3280 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2180_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5080) );
  AND2X2 AND2X2_3281 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5081), .B(REGFILE_SIM_reg_bank__abc_33898_n5079), .Y(REGFILE_SIM_reg_bank_reg_r5_15__FF_INPUT) );
  AND2X2 AND2X2_3282 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2185), .Y(REGFILE_SIM_reg_bank__abc_33898_n5084) );
  AND2X2 AND2X2_3283 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5085), .B(REGFILE_SIM_reg_bank__abc_33898_n5083), .Y(REGFILE_SIM_reg_bank_reg_r5_16__FF_INPUT) );
  AND2X2 AND2X2_3284 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2190_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5088) );
  AND2X2 AND2X2_3285 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5089), .B(REGFILE_SIM_reg_bank__abc_33898_n5087), .Y(REGFILE_SIM_reg_bank_reg_r5_17__FF_INPUT) );
  AND2X2 AND2X2_3286 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2195_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5092) );
  AND2X2 AND2X2_3287 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5093_1), .B(REGFILE_SIM_reg_bank__abc_33898_n5091), .Y(REGFILE_SIM_reg_bank_reg_r5_18__FF_INPUT) );
  AND2X2 AND2X2_3288 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2200_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5096) );
  AND2X2 AND2X2_3289 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5097), .B(REGFILE_SIM_reg_bank__abc_33898_n5095), .Y(REGFILE_SIM_reg_bank_reg_r5_19__FF_INPUT) );
  AND2X2 AND2X2_329 ( .A(_abc_43815_n1207), .B(_abc_43815_n1204), .Y(_abc_43815_n1208) );
  AND2X2 AND2X2_3290 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2205_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5100) );
  AND2X2 AND2X2_3291 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5101), .B(REGFILE_SIM_reg_bank__abc_33898_n5099), .Y(REGFILE_SIM_reg_bank_reg_r5_20__FF_INPUT) );
  AND2X2 AND2X2_3292 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2210), .Y(REGFILE_SIM_reg_bank__abc_33898_n5104) );
  AND2X2 AND2X2_3293 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5105), .B(REGFILE_SIM_reg_bank__abc_33898_n5103), .Y(REGFILE_SIM_reg_bank_reg_r5_21__FF_INPUT) );
  AND2X2 AND2X2_3294 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2215_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5108) );
  AND2X2 AND2X2_3295 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5109), .B(REGFILE_SIM_reg_bank__abc_33898_n5107), .Y(REGFILE_SIM_reg_bank_reg_r5_22__FF_INPUT) );
  AND2X2 AND2X2_3296 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2220_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5112) );
  AND2X2 AND2X2_3297 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5113), .B(REGFILE_SIM_reg_bank__abc_33898_n5111), .Y(REGFILE_SIM_reg_bank_reg_r5_23__FF_INPUT) );
  AND2X2 AND2X2_3298 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2225), .Y(REGFILE_SIM_reg_bank__abc_33898_n5116) );
  AND2X2 AND2X2_3299 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5117), .B(REGFILE_SIM_reg_bank__abc_33898_n5115), .Y(REGFILE_SIM_reg_bank_reg_r5_24__FF_INPUT) );
  AND2X2 AND2X2_33 ( .A(_abc_43815_n665), .B(_abc_43815_n667), .Y(_abc_43815_n668) );
  AND2X2 AND2X2_330 ( .A(_abc_43815_n1209), .B(_abc_43815_n1210), .Y(_abc_43815_n1211) );
  AND2X2 AND2X2_3300 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2230_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5120) );
  AND2X2 AND2X2_3301 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5121), .B(REGFILE_SIM_reg_bank__abc_33898_n5119), .Y(REGFILE_SIM_reg_bank_reg_r5_25__FF_INPUT) );
  AND2X2 AND2X2_3302 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2235_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5124) );
  AND2X2 AND2X2_3303 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5125), .B(REGFILE_SIM_reg_bank__abc_33898_n5123_1), .Y(REGFILE_SIM_reg_bank_reg_r5_26__FF_INPUT) );
  AND2X2 AND2X2_3304 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2240), .Y(REGFILE_SIM_reg_bank__abc_33898_n5128) );
  AND2X2 AND2X2_3305 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5129), .B(REGFILE_SIM_reg_bank__abc_33898_n5127), .Y(REGFILE_SIM_reg_bank_reg_r5_27__FF_INPUT) );
  AND2X2 AND2X2_3306 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6), .B(REGFILE_SIM_reg_bank__abc_33898_n2245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5132) );
  AND2X2 AND2X2_3307 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5133), .B(REGFILE_SIM_reg_bank__abc_33898_n5131), .Y(REGFILE_SIM_reg_bank_reg_r5_28__FF_INPUT) );
  AND2X2 AND2X2_3308 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4), .B(REGFILE_SIM_reg_bank__abc_33898_n2250_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5136) );
  AND2X2 AND2X2_3309 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5137), .B(REGFILE_SIM_reg_bank__abc_33898_n5135), .Y(REGFILE_SIM_reg_bank_reg_r5_29__FF_INPUT) );
  AND2X2 AND2X2_331 ( .A(_abc_43815_n1213), .B(_abc_43815_n1211), .Y(_abc_43815_n1214_1) );
  AND2X2 AND2X2_3310 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2), .B(REGFILE_SIM_reg_bank__abc_33898_n2255), .Y(REGFILE_SIM_reg_bank__abc_33898_n5140) );
  AND2X2 AND2X2_3311 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5141), .B(REGFILE_SIM_reg_bank__abc_33898_n5139), .Y(REGFILE_SIM_reg_bank_reg_r5_30__FF_INPUT) );
  AND2X2 AND2X2_3312 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0), .B(REGFILE_SIM_reg_bank__abc_33898_n2260_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5144) );
  AND2X2 AND2X2_3313 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5145), .B(REGFILE_SIM_reg_bank__abc_33898_n5143), .Y(REGFILE_SIM_reg_bank_reg_r5_31__FF_INPUT) );
  AND2X2 AND2X2_3314 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4238), .B(REGFILE_SIM_reg_bank__abc_33898_n3057_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5147) );
  AND2X2 AND2X2_3315 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5150), .B(REGFILE_SIM_reg_bank__abc_33898_n5148), .Y(REGFILE_SIM_reg_bank_reg_r4_0__FF_INPUT) );
  AND2X2 AND2X2_3316 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5153_1), .B(REGFILE_SIM_reg_bank__abc_33898_n5152), .Y(REGFILE_SIM_reg_bank_reg_r4_1__FF_INPUT) );
  AND2X2 AND2X2_3317 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5156), .B(REGFILE_SIM_reg_bank__abc_33898_n5155), .Y(REGFILE_SIM_reg_bank_reg_r4_2__FF_INPUT) );
  AND2X2 AND2X2_3318 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5159), .B(REGFILE_SIM_reg_bank__abc_33898_n5158), .Y(REGFILE_SIM_reg_bank_reg_r4_3__FF_INPUT) );
  AND2X2 AND2X2_3319 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5162), .B(REGFILE_SIM_reg_bank__abc_33898_n5161), .Y(REGFILE_SIM_reg_bank_reg_r4_4__FF_INPUT) );
  AND2X2 AND2X2_332 ( .A(_abc_43815_n1214_1), .B(_abc_43815_n1208), .Y(_abc_43815_n1215) );
  AND2X2 AND2X2_3320 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5165), .B(REGFILE_SIM_reg_bank__abc_33898_n5164), .Y(REGFILE_SIM_reg_bank_reg_r4_5__FF_INPUT) );
  AND2X2 AND2X2_3321 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5168), .B(REGFILE_SIM_reg_bank__abc_33898_n5167), .Y(REGFILE_SIM_reg_bank_reg_r4_6__FF_INPUT) );
  AND2X2 AND2X2_3322 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5171), .B(REGFILE_SIM_reg_bank__abc_33898_n5170), .Y(REGFILE_SIM_reg_bank_reg_r4_7__FF_INPUT) );
  AND2X2 AND2X2_3323 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5174), .B(REGFILE_SIM_reg_bank__abc_33898_n5173), .Y(REGFILE_SIM_reg_bank_reg_r4_8__FF_INPUT) );
  AND2X2 AND2X2_3324 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5177), .B(REGFILE_SIM_reg_bank__abc_33898_n5176), .Y(REGFILE_SIM_reg_bank_reg_r4_9__FF_INPUT) );
  AND2X2 AND2X2_3325 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5180), .B(REGFILE_SIM_reg_bank__abc_33898_n5179), .Y(REGFILE_SIM_reg_bank_reg_r4_10__FF_INPUT) );
  AND2X2 AND2X2_3326 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5183_1), .B(REGFILE_SIM_reg_bank__abc_33898_n5182), .Y(REGFILE_SIM_reg_bank_reg_r4_11__FF_INPUT) );
  AND2X2 AND2X2_3327 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5186), .B(REGFILE_SIM_reg_bank__abc_33898_n5185), .Y(REGFILE_SIM_reg_bank_reg_r4_12__FF_INPUT) );
  AND2X2 AND2X2_3328 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5189), .B(REGFILE_SIM_reg_bank__abc_33898_n5188), .Y(REGFILE_SIM_reg_bank_reg_r4_13__FF_INPUT) );
  AND2X2 AND2X2_3329 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5192), .B(REGFILE_SIM_reg_bank__abc_33898_n5191), .Y(REGFILE_SIM_reg_bank_reg_r4_14__FF_INPUT) );
  AND2X2 AND2X2_333 ( .A(_abc_43815_n1215), .B(_abc_43815_n1203), .Y(_abc_43815_n1216) );
  AND2X2 AND2X2_3330 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5195), .B(REGFILE_SIM_reg_bank__abc_33898_n5194), .Y(REGFILE_SIM_reg_bank_reg_r4_15__FF_INPUT) );
  AND2X2 AND2X2_3331 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5198), .B(REGFILE_SIM_reg_bank__abc_33898_n5197), .Y(REGFILE_SIM_reg_bank_reg_r4_16__FF_INPUT) );
  AND2X2 AND2X2_3332 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5201), .B(REGFILE_SIM_reg_bank__abc_33898_n5200), .Y(REGFILE_SIM_reg_bank_reg_r4_17__FF_INPUT) );
  AND2X2 AND2X2_3333 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5204), .B(REGFILE_SIM_reg_bank__abc_33898_n5203), .Y(REGFILE_SIM_reg_bank_reg_r4_18__FF_INPUT) );
  AND2X2 AND2X2_3334 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5207), .B(REGFILE_SIM_reg_bank__abc_33898_n5206), .Y(REGFILE_SIM_reg_bank_reg_r4_19__FF_INPUT) );
  AND2X2 AND2X2_3335 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5210), .B(REGFILE_SIM_reg_bank__abc_33898_n5209), .Y(REGFILE_SIM_reg_bank_reg_r4_20__FF_INPUT) );
  AND2X2 AND2X2_3336 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5213_1), .B(REGFILE_SIM_reg_bank__abc_33898_n5212), .Y(REGFILE_SIM_reg_bank_reg_r4_21__FF_INPUT) );
  AND2X2 AND2X2_3337 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5216), .B(REGFILE_SIM_reg_bank__abc_33898_n5215), .Y(REGFILE_SIM_reg_bank_reg_r4_22__FF_INPUT) );
  AND2X2 AND2X2_3338 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5219), .B(REGFILE_SIM_reg_bank__abc_33898_n5218), .Y(REGFILE_SIM_reg_bank_reg_r4_23__FF_INPUT) );
  AND2X2 AND2X2_3339 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5222), .B(REGFILE_SIM_reg_bank__abc_33898_n5221), .Y(REGFILE_SIM_reg_bank_reg_r4_24__FF_INPUT) );
  AND2X2 AND2X2_334 ( .A(_abc_43815_n1218), .B(_abc_43815_n1220), .Y(_abc_43815_n1221) );
  AND2X2 AND2X2_3340 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5225), .B(REGFILE_SIM_reg_bank__abc_33898_n5224), .Y(REGFILE_SIM_reg_bank_reg_r4_25__FF_INPUT) );
  AND2X2 AND2X2_3341 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5228), .B(REGFILE_SIM_reg_bank__abc_33898_n5227), .Y(REGFILE_SIM_reg_bank_reg_r4_26__FF_INPUT) );
  AND2X2 AND2X2_3342 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5231), .B(REGFILE_SIM_reg_bank__abc_33898_n5230), .Y(REGFILE_SIM_reg_bank_reg_r4_27__FF_INPUT) );
  AND2X2 AND2X2_3343 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5234), .B(REGFILE_SIM_reg_bank__abc_33898_n5233), .Y(REGFILE_SIM_reg_bank_reg_r4_28__FF_INPUT) );
  AND2X2 AND2X2_3344 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5237), .B(REGFILE_SIM_reg_bank__abc_33898_n5236), .Y(REGFILE_SIM_reg_bank_reg_r4_29__FF_INPUT) );
  AND2X2 AND2X2_3345 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5240), .B(REGFILE_SIM_reg_bank__abc_33898_n5239), .Y(REGFILE_SIM_reg_bank_reg_r4_30__FF_INPUT) );
  AND2X2 AND2X2_3346 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5243_1), .B(REGFILE_SIM_reg_bank__abc_33898_n5242), .Y(REGFILE_SIM_reg_bank_reg_r4_31__FF_INPUT) );
  AND2X2 AND2X2_3347 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3516), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_1) );
  AND2X2 AND2X2_3348 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5248), .B(REGFILE_SIM_reg_bank__abc_33898_n5246), .Y(REGFILE_SIM_reg_bank_reg_r3_0__FF_INPUT) );
  AND2X2 AND2X2_3349 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5251), .B(REGFILE_SIM_reg_bank__abc_33898_n5250), .Y(REGFILE_SIM_reg_bank_reg_r3_1__FF_INPUT) );
  AND2X2 AND2X2_335 ( .A(_abc_43815_n1223), .B(_abc_43815_n1225), .Y(_abc_43815_n1226) );
  AND2X2 AND2X2_3350 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5254), .B(REGFILE_SIM_reg_bank__abc_33898_n5253), .Y(REGFILE_SIM_reg_bank_reg_r3_2__FF_INPUT) );
  AND2X2 AND2X2_3351 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5257), .B(REGFILE_SIM_reg_bank__abc_33898_n5256), .Y(REGFILE_SIM_reg_bank_reg_r3_3__FF_INPUT) );
  AND2X2 AND2X2_3352 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5260), .B(REGFILE_SIM_reg_bank__abc_33898_n5259), .Y(REGFILE_SIM_reg_bank_reg_r3_4__FF_INPUT) );
  AND2X2 AND2X2_3353 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5263), .B(REGFILE_SIM_reg_bank__abc_33898_n5262), .Y(REGFILE_SIM_reg_bank_reg_r3_5__FF_INPUT) );
  AND2X2 AND2X2_3354 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5266), .B(REGFILE_SIM_reg_bank__abc_33898_n5265), .Y(REGFILE_SIM_reg_bank_reg_r3_6__FF_INPUT) );
  AND2X2 AND2X2_3355 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5269), .B(REGFILE_SIM_reg_bank__abc_33898_n5268), .Y(REGFILE_SIM_reg_bank_reg_r3_7__FF_INPUT) );
  AND2X2 AND2X2_3356 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5272), .B(REGFILE_SIM_reg_bank__abc_33898_n5271), .Y(REGFILE_SIM_reg_bank_reg_r3_8__FF_INPUT) );
  AND2X2 AND2X2_3357 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5275), .B(REGFILE_SIM_reg_bank__abc_33898_n5274), .Y(REGFILE_SIM_reg_bank_reg_r3_9__FF_INPUT) );
  AND2X2 AND2X2_3358 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5278), .B(REGFILE_SIM_reg_bank__abc_33898_n5277), .Y(REGFILE_SIM_reg_bank_reg_r3_10__FF_INPUT) );
  AND2X2 AND2X2_3359 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5281), .B(REGFILE_SIM_reg_bank__abc_33898_n5280), .Y(REGFILE_SIM_reg_bank_reg_r3_11__FF_INPUT) );
  AND2X2 AND2X2_336 ( .A(_abc_43815_n1221), .B(_abc_43815_n1226), .Y(_abc_43815_n1227) );
  AND2X2 AND2X2_3360 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5284), .B(REGFILE_SIM_reg_bank__abc_33898_n5283), .Y(REGFILE_SIM_reg_bank_reg_r3_12__FF_INPUT) );
  AND2X2 AND2X2_3361 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5287), .B(REGFILE_SIM_reg_bank__abc_33898_n5286), .Y(REGFILE_SIM_reg_bank_reg_r3_13__FF_INPUT) );
  AND2X2 AND2X2_3362 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5290), .B(REGFILE_SIM_reg_bank__abc_33898_n5289), .Y(REGFILE_SIM_reg_bank_reg_r3_14__FF_INPUT) );
  AND2X2 AND2X2_3363 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5293), .B(REGFILE_SIM_reg_bank__abc_33898_n5292), .Y(REGFILE_SIM_reg_bank_reg_r3_15__FF_INPUT) );
  AND2X2 AND2X2_3364 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5296), .B(REGFILE_SIM_reg_bank__abc_33898_n5295), .Y(REGFILE_SIM_reg_bank_reg_r3_16__FF_INPUT) );
  AND2X2 AND2X2_3365 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5299), .B(REGFILE_SIM_reg_bank__abc_33898_n5298), .Y(REGFILE_SIM_reg_bank_reg_r3_17__FF_INPUT) );
  AND2X2 AND2X2_3366 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5302), .B(REGFILE_SIM_reg_bank__abc_33898_n5301), .Y(REGFILE_SIM_reg_bank_reg_r3_18__FF_INPUT) );
  AND2X2 AND2X2_3367 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5305), .B(REGFILE_SIM_reg_bank__abc_33898_n5304), .Y(REGFILE_SIM_reg_bank_reg_r3_19__FF_INPUT) );
  AND2X2 AND2X2_3368 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5308), .B(REGFILE_SIM_reg_bank__abc_33898_n5307), .Y(REGFILE_SIM_reg_bank_reg_r3_20__FF_INPUT) );
  AND2X2 AND2X2_3369 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5311), .B(REGFILE_SIM_reg_bank__abc_33898_n5310), .Y(REGFILE_SIM_reg_bank_reg_r3_21__FF_INPUT) );
  AND2X2 AND2X2_337 ( .A(_abc_43815_n1229), .B(_abc_43815_n1231), .Y(_abc_43815_n1232) );
  AND2X2 AND2X2_3370 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5314), .B(REGFILE_SIM_reg_bank__abc_33898_n5313), .Y(REGFILE_SIM_reg_bank_reg_r3_22__FF_INPUT) );
  AND2X2 AND2X2_3371 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5317), .B(REGFILE_SIM_reg_bank__abc_33898_n5316), .Y(REGFILE_SIM_reg_bank_reg_r3_23__FF_INPUT) );
  AND2X2 AND2X2_3372 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5320), .B(REGFILE_SIM_reg_bank__abc_33898_n5319), .Y(REGFILE_SIM_reg_bank_reg_r3_24__FF_INPUT) );
  AND2X2 AND2X2_3373 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5323), .B(REGFILE_SIM_reg_bank__abc_33898_n5322), .Y(REGFILE_SIM_reg_bank_reg_r3_25__FF_INPUT) );
  AND2X2 AND2X2_3374 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5326), .B(REGFILE_SIM_reg_bank__abc_33898_n5325), .Y(REGFILE_SIM_reg_bank_reg_r3_26__FF_INPUT) );
  AND2X2 AND2X2_3375 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5329), .B(REGFILE_SIM_reg_bank__abc_33898_n5328), .Y(REGFILE_SIM_reg_bank_reg_r3_27__FF_INPUT) );
  AND2X2 AND2X2_3376 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5332), .B(REGFILE_SIM_reg_bank__abc_33898_n5331), .Y(REGFILE_SIM_reg_bank_reg_r3_28__FF_INPUT) );
  AND2X2 AND2X2_3377 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5335), .B(REGFILE_SIM_reg_bank__abc_33898_n5334), .Y(REGFILE_SIM_reg_bank_reg_r3_29__FF_INPUT) );
  AND2X2 AND2X2_3378 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5338), .B(REGFILE_SIM_reg_bank__abc_33898_n5337), .Y(REGFILE_SIM_reg_bank_reg_r3_30__FF_INPUT) );
  AND2X2 AND2X2_3379 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5341), .B(REGFILE_SIM_reg_bank__abc_33898_n5340), .Y(REGFILE_SIM_reg_bank_reg_r3_31__FF_INPUT) );
  AND2X2 AND2X2_338 ( .A(_abc_43815_n1235), .B(_abc_43815_n1233_1), .Y(_abc_43815_n1236) );
  AND2X2 AND2X2_3380 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3615), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n5343) );
  AND2X2 AND2X2_3381 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5346), .B(REGFILE_SIM_reg_bank__abc_33898_n5344), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_0__FF_INPUT) );
  AND2X2 AND2X2_3382 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5349), .B(REGFILE_SIM_reg_bank__abc_33898_n5348), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_1__FF_INPUT) );
  AND2X2 AND2X2_3383 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5352), .B(REGFILE_SIM_reg_bank__abc_33898_n5351), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_2__FF_INPUT) );
  AND2X2 AND2X2_3384 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5355), .B(REGFILE_SIM_reg_bank__abc_33898_n5354), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_3__FF_INPUT) );
  AND2X2 AND2X2_3385 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5358), .B(REGFILE_SIM_reg_bank__abc_33898_n5357), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_4__FF_INPUT) );
  AND2X2 AND2X2_3386 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5361), .B(REGFILE_SIM_reg_bank__abc_33898_n5360), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_5__FF_INPUT) );
  AND2X2 AND2X2_3387 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5364), .B(REGFILE_SIM_reg_bank__abc_33898_n5363), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_6__FF_INPUT) );
  AND2X2 AND2X2_3388 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5367), .B(REGFILE_SIM_reg_bank__abc_33898_n5366), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_7__FF_INPUT) );
  AND2X2 AND2X2_3389 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5370), .B(REGFILE_SIM_reg_bank__abc_33898_n5369), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_8__FF_INPUT) );
  AND2X2 AND2X2_339 ( .A(_abc_43815_n1232), .B(_abc_43815_n1236), .Y(_abc_43815_n1237) );
  AND2X2 AND2X2_3390 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5373), .B(REGFILE_SIM_reg_bank__abc_33898_n5372), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_9__FF_INPUT) );
  AND2X2 AND2X2_3391 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5376), .B(REGFILE_SIM_reg_bank__abc_33898_n5375), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_10__FF_INPUT) );
  AND2X2 AND2X2_3392 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5379), .B(REGFILE_SIM_reg_bank__abc_33898_n5378), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_11__FF_INPUT) );
  AND2X2 AND2X2_3393 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5382), .B(REGFILE_SIM_reg_bank__abc_33898_n5381), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_12__FF_INPUT) );
  AND2X2 AND2X2_3394 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5385), .B(REGFILE_SIM_reg_bank__abc_33898_n5384), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_13__FF_INPUT) );
  AND2X2 AND2X2_3395 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5388), .B(REGFILE_SIM_reg_bank__abc_33898_n5387), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_14__FF_INPUT) );
  AND2X2 AND2X2_3396 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5391), .B(REGFILE_SIM_reg_bank__abc_33898_n5390), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_15__FF_INPUT) );
  AND2X2 AND2X2_3397 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5394), .B(REGFILE_SIM_reg_bank__abc_33898_n5393), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_16__FF_INPUT) );
  AND2X2 AND2X2_3398 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5397), .B(REGFILE_SIM_reg_bank__abc_33898_n5396), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_17__FF_INPUT) );
  AND2X2 AND2X2_3399 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5400), .B(REGFILE_SIM_reg_bank__abc_33898_n5399), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_18__FF_INPUT) );
  AND2X2 AND2X2_34 ( .A(_abc_43815_n663), .B(_abc_43815_n669), .Y(_abc_43815_n670_1) );
  AND2X2 AND2X2_340 ( .A(_abc_43815_n1227), .B(_abc_43815_n1237), .Y(_abc_43815_n1238) );
  AND2X2 AND2X2_3400 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5403), .B(REGFILE_SIM_reg_bank__abc_33898_n5402), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_19__FF_INPUT) );
  AND2X2 AND2X2_3401 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5406), .B(REGFILE_SIM_reg_bank__abc_33898_n5405), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_20__FF_INPUT) );
  AND2X2 AND2X2_3402 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5409), .B(REGFILE_SIM_reg_bank__abc_33898_n5408), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_21__FF_INPUT) );
  AND2X2 AND2X2_3403 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5412), .B(REGFILE_SIM_reg_bank__abc_33898_n5411), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_22__FF_INPUT) );
  AND2X2 AND2X2_3404 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5415), .B(REGFILE_SIM_reg_bank__abc_33898_n5414), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_23__FF_INPUT) );
  AND2X2 AND2X2_3405 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5418), .B(REGFILE_SIM_reg_bank__abc_33898_n5417), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_24__FF_INPUT) );
  AND2X2 AND2X2_3406 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5421), .B(REGFILE_SIM_reg_bank__abc_33898_n5420), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_25__FF_INPUT) );
  AND2X2 AND2X2_3407 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5424), .B(REGFILE_SIM_reg_bank__abc_33898_n5423), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_26__FF_INPUT) );
  AND2X2 AND2X2_3408 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5427), .B(REGFILE_SIM_reg_bank__abc_33898_n5426), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_27__FF_INPUT) );
  AND2X2 AND2X2_3409 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5430), .B(REGFILE_SIM_reg_bank__abc_33898_n5429), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_28__FF_INPUT) );
  AND2X2 AND2X2_341 ( .A(_abc_43815_n1238), .B(_abc_43815_n1216), .Y(_abc_43815_n1239) );
  AND2X2 AND2X2_3410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5433), .B(REGFILE_SIM_reg_bank__abc_33898_n5432), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_29__FF_INPUT) );
  AND2X2 AND2X2_3411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5436), .B(REGFILE_SIM_reg_bank__abc_33898_n5435), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_30__FF_INPUT) );
  AND2X2 AND2X2_3412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5439), .B(REGFILE_SIM_reg_bank__abc_33898_n5438), .Y(REGFILE_SIM_reg_bank_reg_r2_fp_31__FF_INPUT) );
  AND2X2 AND2X2_3413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3714), .B(REGFILE_SIM_reg_bank__abc_33898_n3912), .Y(REGFILE_SIM_reg_bank__abc_33898_n5441) );
  AND2X2 AND2X2_3414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5444), .B(REGFILE_SIM_reg_bank__abc_33898_n5442), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_0__FF_INPUT) );
  AND2X2 AND2X2_3415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5447), .B(REGFILE_SIM_reg_bank__abc_33898_n5446), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_1__FF_INPUT) );
  AND2X2 AND2X2_3416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5450), .B(REGFILE_SIM_reg_bank__abc_33898_n5449), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_2__FF_INPUT) );
  AND2X2 AND2X2_3417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5453), .B(REGFILE_SIM_reg_bank__abc_33898_n5452), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_3__FF_INPUT) );
  AND2X2 AND2X2_3418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5456), .B(REGFILE_SIM_reg_bank__abc_33898_n5455), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_4__FF_INPUT) );
  AND2X2 AND2X2_3419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5459), .B(REGFILE_SIM_reg_bank__abc_33898_n5458), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_5__FF_INPUT) );
  AND2X2 AND2X2_342 ( .A(_abc_43815_n1239), .B(_abc_43815_n1080), .Y(_abc_43815_n1240) );
  AND2X2 AND2X2_3420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5462), .B(REGFILE_SIM_reg_bank__abc_33898_n5461), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_6__FF_INPUT) );
  AND2X2 AND2X2_3421 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5465), .B(REGFILE_SIM_reg_bank__abc_33898_n5464), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_7__FF_INPUT) );
  AND2X2 AND2X2_3422 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5468), .B(REGFILE_SIM_reg_bank__abc_33898_n5467), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_8__FF_INPUT) );
  AND2X2 AND2X2_3423 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5471), .B(REGFILE_SIM_reg_bank__abc_33898_n5470), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_9__FF_INPUT) );
  AND2X2 AND2X2_3424 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5474), .B(REGFILE_SIM_reg_bank__abc_33898_n5473), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_10__FF_INPUT) );
  AND2X2 AND2X2_3425 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5477), .B(REGFILE_SIM_reg_bank__abc_33898_n5476), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_11__FF_INPUT) );
  AND2X2 AND2X2_3426 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5480), .B(REGFILE_SIM_reg_bank__abc_33898_n5479), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_12__FF_INPUT) );
  AND2X2 AND2X2_3427 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5483), .B(REGFILE_SIM_reg_bank__abc_33898_n5482), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_13__FF_INPUT) );
  AND2X2 AND2X2_3428 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5486), .B(REGFILE_SIM_reg_bank__abc_33898_n5485), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_14__FF_INPUT) );
  AND2X2 AND2X2_3429 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5489), .B(REGFILE_SIM_reg_bank__abc_33898_n5488), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_15__FF_INPUT) );
  AND2X2 AND2X2_343 ( .A(_abc_43815_n1241), .B(esr_q_2_), .Y(_abc_43815_n1242) );
  AND2X2 AND2X2_3430 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5492), .B(REGFILE_SIM_reg_bank__abc_33898_n5491), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_16__FF_INPUT) );
  AND2X2 AND2X2_3431 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5495), .B(REGFILE_SIM_reg_bank__abc_33898_n5494), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_17__FF_INPUT) );
  AND2X2 AND2X2_3432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5498), .B(REGFILE_SIM_reg_bank__abc_33898_n5497), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_18__FF_INPUT) );
  AND2X2 AND2X2_3433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5501), .B(REGFILE_SIM_reg_bank__abc_33898_n5500), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_19__FF_INPUT) );
  AND2X2 AND2X2_3434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5504), .B(REGFILE_SIM_reg_bank__abc_33898_n5503), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_20__FF_INPUT) );
  AND2X2 AND2X2_3435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5507), .B(REGFILE_SIM_reg_bank__abc_33898_n5506), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_21__FF_INPUT) );
  AND2X2 AND2X2_3436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5510), .B(REGFILE_SIM_reg_bank__abc_33898_n5509), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_22__FF_INPUT) );
  AND2X2 AND2X2_3437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5513), .B(REGFILE_SIM_reg_bank__abc_33898_n5512), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_23__FF_INPUT) );
  AND2X2 AND2X2_3438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5516), .B(REGFILE_SIM_reg_bank__abc_33898_n5515), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_24__FF_INPUT) );
  AND2X2 AND2X2_3439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5519), .B(REGFILE_SIM_reg_bank__abc_33898_n5518), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_25__FF_INPUT) );
  AND2X2 AND2X2_344 ( .A(_abc_43815_n1240), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n1243) );
  AND2X2 AND2X2_3440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5522), .B(REGFILE_SIM_reg_bank__abc_33898_n5521), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_26__FF_INPUT) );
  AND2X2 AND2X2_3441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5525), .B(REGFILE_SIM_reg_bank__abc_33898_n5524), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_27__FF_INPUT) );
  AND2X2 AND2X2_3442 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5528), .B(REGFILE_SIM_reg_bank__abc_33898_n5527), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_28__FF_INPUT) );
  AND2X2 AND2X2_3443 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5531), .B(REGFILE_SIM_reg_bank__abc_33898_n5530), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_29__FF_INPUT) );
  AND2X2 AND2X2_3444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5534), .B(REGFILE_SIM_reg_bank__abc_33898_n5533), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_30__FF_INPUT) );
  AND2X2 AND2X2_3445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5537), .B(REGFILE_SIM_reg_bank__abc_33898_n5536), .Y(REGFILE_SIM_reg_bank_reg_r1_sp_31__FF_INPUT) );
  AND2X2 AND2X2_3446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5540), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5541) );
  AND2X2 AND2X2_3447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5541), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5542) );
  AND2X2 AND2X2_3448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5543), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5544) );
  AND2X2 AND2X2_3449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5542), .B(REGFILE_SIM_reg_bank__abc_33898_n5544), .Y(REGFILE_SIM_reg_bank__abc_33898_n5545) );
  AND2X2 AND2X2_345 ( .A(_abc_43815_n1244), .B(_abc_43815_n1197), .Y(_abc_43815_n1245) );
  AND2X2 AND2X2_3450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5546) );
  AND2X2 AND2X2_3451 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5547) );
  AND2X2 AND2X2_3452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5542), .B(REGFILE_SIM_reg_bank__abc_33898_n5547), .Y(REGFILE_SIM_reg_bank__abc_33898_n5548) );
  AND2X2 AND2X2_3453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5549) );
  AND2X2 AND2X2_3454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5540), .B(REGFILE_SIM_reg_bank__abc_33898_n5551), .Y(REGFILE_SIM_reg_bank__abc_33898_n5552) );
  AND2X2 AND2X2_3455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5552), .B(REGFILE_SIM_reg_bank__abc_33898_n5544), .Y(REGFILE_SIM_reg_bank__abc_33898_n5553) );
  AND2X2 AND2X2_3456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5553), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5554) );
  AND2X2 AND2X2_3457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5555) );
  AND2X2 AND2X2_3458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5552), .B(REGFILE_SIM_reg_bank__abc_33898_n5547), .Y(REGFILE_SIM_reg_bank__abc_33898_n5556) );
  AND2X2 AND2X2_3459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5556), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5557) );
  AND2X2 AND2X2_346 ( .A(_abc_43815_n1228), .B(_abc_43815_n1222), .Y(_abc_43815_n1246) );
  AND2X2 AND2X2_3460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5558) );
  AND2X2 AND2X2_3461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5561), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5562) );
  AND2X2 AND2X2_3462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5551), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5563) );
  AND2X2 AND2X2_3463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5562), .B(REGFILE_SIM_reg_bank__abc_33898_n5563), .Y(REGFILE_SIM_reg_bank__abc_33898_n5564) );
  AND2X2 AND2X2_3464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5564), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5565) );
  AND2X2 AND2X2_3465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5566) );
  AND2X2 AND2X2_3466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5563), .B(REGFILE_SIM_reg_bank__abc_33898_n5547), .Y(REGFILE_SIM_reg_bank__abc_33898_n5567) );
  AND2X2 AND2X2_3467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5567), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5568) );
  AND2X2 AND2X2_3468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5569) );
  AND2X2 AND2X2_3469 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5571) );
  AND2X2 AND2X2_347 ( .A(_abc_43815_n1231), .B(_abc_43815_n1251), .Y(_abc_43815_n1252) );
  AND2X2 AND2X2_3470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5562), .B(REGFILE_SIM_reg_bank__abc_33898_n5571), .Y(REGFILE_SIM_reg_bank__abc_33898_n5572) );
  AND2X2 AND2X2_3471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5572), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5573) );
  AND2X2 AND2X2_3472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5574) );
  AND2X2 AND2X2_3473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5544), .B(REGFILE_SIM_reg_bank__abc_33898_n5571), .Y(REGFILE_SIM_reg_bank__abc_33898_n5575) );
  AND2X2 AND2X2_3474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5575), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5576) );
  AND2X2 AND2X2_3475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5577) );
  AND2X2 AND2X2_3476 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5553), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5581) );
  AND2X2 AND2X2_3477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5582) );
  AND2X2 AND2X2_3478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5556), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5583) );
  AND2X2 AND2X2_3479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5584) );
  AND2X2 AND2X2_348 ( .A(_abc_43815_n1257), .B(sr_q_2_), .Y(_abc_43815_n1258) );
  AND2X2 AND2X2_3480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5541), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5586) );
  AND2X2 AND2X2_3481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5586), .B(REGFILE_SIM_reg_bank__abc_33898_n5562), .Y(REGFILE_SIM_reg_bank__abc_33898_n5587) );
  AND2X2 AND2X2_3482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5588) );
  AND2X2 AND2X2_3483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5561), .B(REGFILE_SIM_reg_bank__abc_33898_n5543), .Y(REGFILE_SIM_reg_bank__abc_33898_n5589) );
  AND2X2 AND2X2_3484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5586), .B(REGFILE_SIM_reg_bank__abc_33898_n5589), .Y(REGFILE_SIM_reg_bank__abc_33898_n5590) );
  AND2X2 AND2X2_3485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5591) );
  AND2X2 AND2X2_3486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5575), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5594) );
  AND2X2 AND2X2_3487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5595) );
  AND2X2 AND2X2_3488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5571), .B(REGFILE_SIM_reg_bank__abc_33898_n5547), .Y(REGFILE_SIM_reg_bank__abc_33898_n5596) );
  AND2X2 AND2X2_3489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5596), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5597) );
  AND2X2 AND2X2_349 ( .A(_abc_43815_n1231), .B(_abc_43815_n1225), .Y(_abc_43815_n1259) );
  AND2X2 AND2X2_3490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5598) );
  AND2X2 AND2X2_3491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5564), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5600) );
  AND2X2 AND2X2_3492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5601) );
  AND2X2 AND2X2_3493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5589), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5602) );
  AND2X2 AND2X2_3494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5602), .B(REGFILE_SIM_reg_bank__abc_33898_n5563), .Y(REGFILE_SIM_reg_bank__abc_33898_n5603) );
  AND2X2 AND2X2_3495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5604) );
  AND2X2 AND2X2_3496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5552), .B(REGFILE_SIM_reg_bank__abc_33898_n5562), .Y(REGFILE_SIM_reg_bank__abc_33898_n5609) );
  AND2X2 AND2X2_3497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5609), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5610) );
  AND2X2 AND2X2_3498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5611) );
  AND2X2 AND2X2_3499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5589), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5612) );
  AND2X2 AND2X2_35 ( .A(_abc_43815_n670_1), .B(state_q_5_), .Y(_abc_43815_n671) );
  AND2X2 AND2X2_350 ( .A(_abc_43815_n1259), .B(_abc_43815_n1246), .Y(_abc_43815_n1260) );
  AND2X2 AND2X2_3500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5612), .B(REGFILE_SIM_reg_bank__abc_33898_n5571), .Y(REGFILE_SIM_reg_bank__abc_33898_n5613) );
  AND2X2 AND2X2_3501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5614) );
  AND2X2 AND2X2_3502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5542), .B(REGFILE_SIM_reg_bank__abc_33898_n5589), .Y(REGFILE_SIM_reg_bank__abc_33898_n5616) );
  AND2X2 AND2X2_3503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5617) );
  AND2X2 AND2X2_3504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5542), .B(REGFILE_SIM_reg_bank__abc_33898_n5562), .Y(REGFILE_SIM_reg_bank__abc_33898_n5618) );
  AND2X2 AND2X2_3505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5619) );
  AND2X2 AND2X2_3506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5544), .B(REGFILE_SIM_reg_bank__abc_33898_n5563), .Y(REGFILE_SIM_reg_bank__abc_33898_n5622) );
  AND2X2 AND2X2_3507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5622), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5623) );
  AND2X2 AND2X2_3508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5624) );
  AND2X2 AND2X2_3509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5612), .B(REGFILE_SIM_reg_bank__abc_33898_n5563), .Y(REGFILE_SIM_reg_bank__abc_33898_n5625) );
  AND2X2 AND2X2_351 ( .A(_abc_43815_n1251), .B(_abc_43815_n1235), .Y(_abc_43815_n1261) );
  AND2X2 AND2X2_3510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5626) );
  AND2X2 AND2X2_3511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5596), .B(REGFILE_SIM_reg_bank__abc_33898_n5539), .Y(REGFILE_SIM_reg_bank__abc_33898_n5627) );
  AND2X2 AND2X2_3512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5628) );
  AND2X2 AND2X2_3513 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5586), .B(REGFILE_SIM_reg_bank__abc_33898_n5544), .Y(REGFILE_SIM_reg_bank__abc_33898_n5632) );
  AND2X2 AND2X2_3514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5633) );
  AND2X2 AND2X2_3515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5586), .B(REGFILE_SIM_reg_bank__abc_33898_n5547), .Y(REGFILE_SIM_reg_bank__abc_33898_n5634) );
  AND2X2 AND2X2_3516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5635) );
  AND2X2 AND2X2_3517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5609), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5637) );
  AND2X2 AND2X2_3518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5638) );
  AND2X2 AND2X2_3519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5602), .B(REGFILE_SIM_reg_bank__abc_33898_n5552), .Y(REGFILE_SIM_reg_bank__abc_33898_n5639) );
  AND2X2 AND2X2_352 ( .A(_abc_43815_n1221), .B(_abc_43815_n1261), .Y(_abc_43815_n1262) );
  AND2X2 AND2X2_3520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5640) );
  AND2X2 AND2X2_3521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5602), .B(REGFILE_SIM_reg_bank__abc_33898_n5571), .Y(REGFILE_SIM_reg_bank__abc_33898_n5643) );
  AND2X2 AND2X2_3522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5644) );
  AND2X2 AND2X2_3523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5572), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5645) );
  AND2X2 AND2X2_3524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5646) );
  AND2X2 AND2X2_3525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5622), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5648) );
  AND2X2 AND2X2_3526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5649) );
  AND2X2 AND2X2_3527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5567), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5650) );
  AND2X2 AND2X2_3528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5651) );
  AND2X2 AND2X2_3529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5657) );
  AND2X2 AND2X2_353 ( .A(_abc_43815_n1262), .B(_abc_43815_n1260), .Y(_abc_43815_n1263_1) );
  AND2X2 AND2X2_3530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5658) );
  AND2X2 AND2X2_3531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5660) );
  AND2X2 AND2X2_3532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5661) );
  AND2X2 AND2X2_3533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5664) );
  AND2X2 AND2X2_3534 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5665) );
  AND2X2 AND2X2_3535 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5667) );
  AND2X2 AND2X2_3536 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5668) );
  AND2X2 AND2X2_3537 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5672) );
  AND2X2 AND2X2_3538 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5673) );
  AND2X2 AND2X2_3539 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5675) );
  AND2X2 AND2X2_354 ( .A(_abc_43815_n1263_1), .B(_abc_43815_n1216), .Y(_abc_43815_n1264) );
  AND2X2 AND2X2_3540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5676) );
  AND2X2 AND2X2_3541 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5679) );
  AND2X2 AND2X2_3542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5680) );
  AND2X2 AND2X2_3543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5682) );
  AND2X2 AND2X2_3544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5683) );
  AND2X2 AND2X2_3545 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5688) );
  AND2X2 AND2X2_3546 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5689) );
  AND2X2 AND2X2_3547 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5691) );
  AND2X2 AND2X2_3548 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5692) );
  AND2X2 AND2X2_3549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5695) );
  AND2X2 AND2X2_355 ( .A(_abc_43815_n1264), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n1265) );
  AND2X2 AND2X2_3550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5696) );
  AND2X2 AND2X2_3551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5697) );
  AND2X2 AND2X2_3552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5701) );
  AND2X2 AND2X2_3553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5702) );
  AND2X2 AND2X2_3554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5704) );
  AND2X2 AND2X2_3555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5705) );
  AND2X2 AND2X2_3556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5708) );
  AND2X2 AND2X2_3557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5709) );
  AND2X2 AND2X2_3558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5711) );
  AND2X2 AND2X2_3559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5712) );
  AND2X2 AND2X2_356 ( .A(_abc_43815_n1266_1), .B(_abc_43815_n1080), .Y(_abc_43815_n1267) );
  AND2X2 AND2X2_3560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5718) );
  AND2X2 AND2X2_3561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5719) );
  AND2X2 AND2X2_3562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5721) );
  AND2X2 AND2X2_3563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5722) );
  AND2X2 AND2X2_3564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5725) );
  AND2X2 AND2X2_3565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5726) );
  AND2X2 AND2X2_3566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5728) );
  AND2X2 AND2X2_3567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5729) );
  AND2X2 AND2X2_3568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5733) );
  AND2X2 AND2X2_3569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5734) );
  AND2X2 AND2X2_357 ( .A(_abc_43815_n1066), .B(sr_q_2_), .Y(_abc_43815_n1268) );
  AND2X2 AND2X2_3570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5736) );
  AND2X2 AND2X2_3571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5737) );
  AND2X2 AND2X2_3572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5740) );
  AND2X2 AND2X2_3573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5741) );
  AND2X2 AND2X2_3574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5743) );
  AND2X2 AND2X2_3575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5744) );
  AND2X2 AND2X2_3576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5749) );
  AND2X2 AND2X2_3577 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5750) );
  AND2X2 AND2X2_3578 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5752) );
  AND2X2 AND2X2_3579 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5753) );
  AND2X2 AND2X2_358 ( .A(_abc_43815_n1065_1_bF_buf3), .B(esr_q_2_), .Y(_abc_43815_n1269) );
  AND2X2 AND2X2_3580 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5756) );
  AND2X2 AND2X2_3581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5757) );
  AND2X2 AND2X2_3582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5758) );
  AND2X2 AND2X2_3583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5762) );
  AND2X2 AND2X2_3584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5763) );
  AND2X2 AND2X2_3585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5765) );
  AND2X2 AND2X2_3586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5766) );
  AND2X2 AND2X2_3587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5769) );
  AND2X2 AND2X2_3588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5770) );
  AND2X2 AND2X2_3589 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5772) );
  AND2X2 AND2X2_359 ( .A(_abc_43815_n1270), .B(_abc_43815_n1081), .Y(_abc_43815_n1271) );
  AND2X2 AND2X2_3590 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5773) );
  AND2X2 AND2X2_3591 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5779) );
  AND2X2 AND2X2_3592 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5780) );
  AND2X2 AND2X2_3593 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5782) );
  AND2X2 AND2X2_3594 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5783) );
  AND2X2 AND2X2_3595 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5786) );
  AND2X2 AND2X2_3596 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5787) );
  AND2X2 AND2X2_3597 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5789) );
  AND2X2 AND2X2_3598 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5790) );
  AND2X2 AND2X2_3599 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5794) );
  AND2X2 AND2X2_36 ( .A(_abc_43815_n671_bF_buf4), .B(_abc_43815_n652), .Y(_abc_43815_n672) );
  AND2X2 AND2X2_360 ( .A(_abc_43815_n1272), .B(_abc_43815_n1274), .Y(_abc_43815_n1275) );
  AND2X2 AND2X2_3600 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5795) );
  AND2X2 AND2X2_3601 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5797) );
  AND2X2 AND2X2_3602 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5798) );
  AND2X2 AND2X2_3603 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5801) );
  AND2X2 AND2X2_3604 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5802) );
  AND2X2 AND2X2_3605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5804) );
  AND2X2 AND2X2_3606 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5805) );
  AND2X2 AND2X2_3607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5810) );
  AND2X2 AND2X2_3608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5811) );
  AND2X2 AND2X2_3609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5813) );
  AND2X2 AND2X2_361 ( .A(_abc_43815_n1194), .B(_abc_43815_n1276), .Y(_abc_43815_n1277) );
  AND2X2 AND2X2_3610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5814) );
  AND2X2 AND2X2_3611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5817) );
  AND2X2 AND2X2_3612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5818) );
  AND2X2 AND2X2_3613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5819) );
  AND2X2 AND2X2_3614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5823) );
  AND2X2 AND2X2_3615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5824) );
  AND2X2 AND2X2_3616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5826) );
  AND2X2 AND2X2_3617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5827) );
  AND2X2 AND2X2_3618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5830) );
  AND2X2 AND2X2_3619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5831) );
  AND2X2 AND2X2_362 ( .A(_abc_43815_n1278_bF_buf7), .B(esr_q_2_), .Y(_abc_43815_n1279) );
  AND2X2 AND2X2_3620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5833) );
  AND2X2 AND2X2_3621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5834) );
  AND2X2 AND2X2_3622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5840) );
  AND2X2 AND2X2_3623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5841) );
  AND2X2 AND2X2_3624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5843) );
  AND2X2 AND2X2_3625 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5844) );
  AND2X2 AND2X2_3626 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5847) );
  AND2X2 AND2X2_3627 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5848) );
  AND2X2 AND2X2_3628 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5850) );
  AND2X2 AND2X2_3629 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5851) );
  AND2X2 AND2X2_363 ( .A(_abc_43815_n1192), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .Y(_abc_43815_n1280) );
  AND2X2 AND2X2_3630 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5855) );
  AND2X2 AND2X2_3631 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5856) );
  AND2X2 AND2X2_3632 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5858) );
  AND2X2 AND2X2_3633 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5859) );
  AND2X2 AND2X2_3634 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5862) );
  AND2X2 AND2X2_3635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5863) );
  AND2X2 AND2X2_3636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5865) );
  AND2X2 AND2X2_3637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5866) );
  AND2X2 AND2X2_3638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5871) );
  AND2X2 AND2X2_3639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5872) );
  AND2X2 AND2X2_364 ( .A(_abc_43815_n1280), .B(_abc_43815_n1272), .Y(_abc_43815_n1281) );
  AND2X2 AND2X2_3640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5874) );
  AND2X2 AND2X2_3641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5875) );
  AND2X2 AND2X2_3642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5878) );
  AND2X2 AND2X2_3643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5879) );
  AND2X2 AND2X2_3644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5880) );
  AND2X2 AND2X2_3645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5884) );
  AND2X2 AND2X2_3646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5885) );
  AND2X2 AND2X2_3647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5887) );
  AND2X2 AND2X2_3648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5888) );
  AND2X2 AND2X2_3649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5891) );
  AND2X2 AND2X2_365 ( .A(_abc_43815_n1283_1), .B(enable_i_bF_buf5), .Y(esr_q_2__FF_INPUT) );
  AND2X2 AND2X2_3650 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5892) );
  AND2X2 AND2X2_3651 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5894) );
  AND2X2 AND2X2_3652 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5895) );
  AND2X2 AND2X2_3653 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5901) );
  AND2X2 AND2X2_3654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5902) );
  AND2X2 AND2X2_3655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5904) );
  AND2X2 AND2X2_3656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5905) );
  AND2X2 AND2X2_3657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5908) );
  AND2X2 AND2X2_3658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5909) );
  AND2X2 AND2X2_3659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5911) );
  AND2X2 AND2X2_366 ( .A(_abc_43815_n992), .B(_abc_43815_n1003), .Y(_abc_43815_n1287) );
  AND2X2 AND2X2_3660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5912) );
  AND2X2 AND2X2_3661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5916) );
  AND2X2 AND2X2_3662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5917) );
  AND2X2 AND2X2_3663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5919) );
  AND2X2 AND2X2_3664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5920) );
  AND2X2 AND2X2_3665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5923) );
  AND2X2 AND2X2_3666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5924) );
  AND2X2 AND2X2_3667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5926) );
  AND2X2 AND2X2_3668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5927) );
  AND2X2 AND2X2_3669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5932) );
  AND2X2 AND2X2_367 ( .A(_abc_43815_n987), .B(_abc_43815_n1024), .Y(_abc_43815_n1288) );
  AND2X2 AND2X2_3670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5933) );
  AND2X2 AND2X2_3671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5935) );
  AND2X2 AND2X2_3672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5936) );
  AND2X2 AND2X2_3673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5939) );
  AND2X2 AND2X2_3674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5940) );
  AND2X2 AND2X2_3675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5941) );
  AND2X2 AND2X2_3676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5945) );
  AND2X2 AND2X2_3677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5946) );
  AND2X2 AND2X2_3678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5948) );
  AND2X2 AND2X2_3679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5949) );
  AND2X2 AND2X2_368 ( .A(_abc_43815_n1288), .B(_abc_43815_n1287), .Y(_abc_43815_n1289_1) );
  AND2X2 AND2X2_3680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5952) );
  AND2X2 AND2X2_3681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5953) );
  AND2X2 AND2X2_3682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5955) );
  AND2X2 AND2X2_3683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5956) );
  AND2X2 AND2X2_3684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5962) );
  AND2X2 AND2X2_3685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5963) );
  AND2X2 AND2X2_3686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5965) );
  AND2X2 AND2X2_3687 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5966) );
  AND2X2 AND2X2_3688 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5969) );
  AND2X2 AND2X2_3689 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5970) );
  AND2X2 AND2X2_369 ( .A(_abc_43815_n987), .B(_abc_43815_n989), .Y(_abc_43815_n1290) );
  AND2X2 AND2X2_3690 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5972) );
  AND2X2 AND2X2_3691 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5973) );
  AND2X2 AND2X2_3692 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5977) );
  AND2X2 AND2X2_3693 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5978) );
  AND2X2 AND2X2_3694 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5980) );
  AND2X2 AND2X2_3695 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5981) );
  AND2X2 AND2X2_3696 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5984) );
  AND2X2 AND2X2_3697 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5985) );
  AND2X2 AND2X2_3698 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5987) );
  AND2X2 AND2X2_3699 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5988) );
  AND2X2 AND2X2_37 ( .A(_abc_43815_n674_1), .B(state_q_2_), .Y(_abc_43815_n675) );
  AND2X2 AND2X2_370 ( .A(_abc_43815_n1290), .B(_abc_43815_n1287), .Y(_abc_43815_n1291) );
  AND2X2 AND2X2_3700 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5993) );
  AND2X2 AND2X2_3701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5994) );
  AND2X2 AND2X2_3702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5996) );
  AND2X2 AND2X2_3703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5997) );
  AND2X2 AND2X2_3704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6000) );
  AND2X2 AND2X2_3705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6001) );
  AND2X2 AND2X2_3706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6002) );
  AND2X2 AND2X2_3707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6006) );
  AND2X2 AND2X2_3708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6007) );
  AND2X2 AND2X2_3709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6009) );
  AND2X2 AND2X2_371 ( .A(_abc_43815_n987), .B(_abc_43815_n1034), .Y(_abc_43815_n1293) );
  AND2X2 AND2X2_3710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6010) );
  AND2X2 AND2X2_3711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6013) );
  AND2X2 AND2X2_3712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6014) );
  AND2X2 AND2X2_3713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6016) );
  AND2X2 AND2X2_3714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6017) );
  AND2X2 AND2X2_3715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6023) );
  AND2X2 AND2X2_3716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6024) );
  AND2X2 AND2X2_3717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6026) );
  AND2X2 AND2X2_3718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6027) );
  AND2X2 AND2X2_3719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6030) );
  AND2X2 AND2X2_372 ( .A(_abc_43815_n992), .B(_abc_43815_n1017), .Y(_abc_43815_n1294) );
  AND2X2 AND2X2_3720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6031) );
  AND2X2 AND2X2_3721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6033) );
  AND2X2 AND2X2_3722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6034) );
  AND2X2 AND2X2_3723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6038) );
  AND2X2 AND2X2_3724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6039) );
  AND2X2 AND2X2_3725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6041) );
  AND2X2 AND2X2_3726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6042) );
  AND2X2 AND2X2_3727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6045) );
  AND2X2 AND2X2_3728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6046) );
  AND2X2 AND2X2_3729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6048) );
  AND2X2 AND2X2_373 ( .A(_abc_43815_n1293), .B(_abc_43815_n1294), .Y(_abc_43815_n1295) );
  AND2X2 AND2X2_3730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6049) );
  AND2X2 AND2X2_3731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6054) );
  AND2X2 AND2X2_3732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6055) );
  AND2X2 AND2X2_3733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6057) );
  AND2X2 AND2X2_3734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6058) );
  AND2X2 AND2X2_3735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6061) );
  AND2X2 AND2X2_3736 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6062) );
  AND2X2 AND2X2_3737 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6063) );
  AND2X2 AND2X2_3738 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6067) );
  AND2X2 AND2X2_3739 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6068) );
  AND2X2 AND2X2_374 ( .A(_abc_43815_n995), .B(_abc_43815_n1010), .Y(_abc_43815_n1297) );
  AND2X2 AND2X2_3740 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6070) );
  AND2X2 AND2X2_3741 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6071) );
  AND2X2 AND2X2_3742 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6074) );
  AND2X2 AND2X2_3743 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6075) );
  AND2X2 AND2X2_3744 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6077) );
  AND2X2 AND2X2_3745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6078) );
  AND2X2 AND2X2_3746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6084) );
  AND2X2 AND2X2_3747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6085) );
  AND2X2 AND2X2_3748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6087) );
  AND2X2 AND2X2_3749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6088) );
  AND2X2 AND2X2_375 ( .A(_abc_43815_n987), .B(_abc_43815_n1297), .Y(_abc_43815_n1298) );
  AND2X2 AND2X2_3750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6091) );
  AND2X2 AND2X2_3751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6092) );
  AND2X2 AND2X2_3752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6094) );
  AND2X2 AND2X2_3753 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6095) );
  AND2X2 AND2X2_3754 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6099) );
  AND2X2 AND2X2_3755 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6100) );
  AND2X2 AND2X2_3756 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6102) );
  AND2X2 AND2X2_3757 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6103) );
  AND2X2 AND2X2_3758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6106) );
  AND2X2 AND2X2_3759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6107) );
  AND2X2 AND2X2_376 ( .A(_abc_43815_n1301), .B(_abc_43815_n1299), .Y(_abc_43815_n1302) );
  AND2X2 AND2X2_3760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6109) );
  AND2X2 AND2X2_3761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6110) );
  AND2X2 AND2X2_3762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6115) );
  AND2X2 AND2X2_3763 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6116) );
  AND2X2 AND2X2_3764 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6118) );
  AND2X2 AND2X2_3765 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6119) );
  AND2X2 AND2X2_3766 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6122) );
  AND2X2 AND2X2_3767 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6123) );
  AND2X2 AND2X2_3768 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6124) );
  AND2X2 AND2X2_3769 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6128) );
  AND2X2 AND2X2_377 ( .A(_abc_43815_n1302), .B(_abc_43815_n1296), .Y(_abc_43815_n1303_1) );
  AND2X2 AND2X2_3770 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6129) );
  AND2X2 AND2X2_3771 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6131) );
  AND2X2 AND2X2_3772 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6132) );
  AND2X2 AND2X2_3773 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6135) );
  AND2X2 AND2X2_3774 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6136) );
  AND2X2 AND2X2_3775 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6138) );
  AND2X2 AND2X2_3776 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6139) );
  AND2X2 AND2X2_3777 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6145) );
  AND2X2 AND2X2_3778 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6146) );
  AND2X2 AND2X2_3779 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6148) );
  AND2X2 AND2X2_378 ( .A(_abc_43815_n992), .B(_abc_43815_n1011), .Y(_abc_43815_n1304) );
  AND2X2 AND2X2_3780 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6149) );
  AND2X2 AND2X2_3781 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6152) );
  AND2X2 AND2X2_3782 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6153) );
  AND2X2 AND2X2_3783 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6155) );
  AND2X2 AND2X2_3784 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6156) );
  AND2X2 AND2X2_3785 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6160) );
  AND2X2 AND2X2_3786 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6161) );
  AND2X2 AND2X2_3787 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6163) );
  AND2X2 AND2X2_3788 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6164) );
  AND2X2 AND2X2_3789 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6167) );
  AND2X2 AND2X2_379 ( .A(_abc_43815_n1293), .B(_abc_43815_n1304), .Y(_abc_43815_n1305) );
  AND2X2 AND2X2_3790 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6168) );
  AND2X2 AND2X2_3791 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6170) );
  AND2X2 AND2X2_3792 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6171) );
  AND2X2 AND2X2_3793 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6176) );
  AND2X2 AND2X2_3794 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6177) );
  AND2X2 AND2X2_3795 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6179) );
  AND2X2 AND2X2_3796 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6180) );
  AND2X2 AND2X2_3797 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6183) );
  AND2X2 AND2X2_3798 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6184) );
  AND2X2 AND2X2_3799 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6185) );
  AND2X2 AND2X2_38 ( .A(_abc_43815_n674_1), .B(state_q_1_bF_buf3), .Y(_abc_43815_n677) );
  AND2X2 AND2X2_380 ( .A(_abc_43815_n1295), .B(alu_less_than_o), .Y(_abc_43815_n1306) );
  AND2X2 AND2X2_3800 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6189) );
  AND2X2 AND2X2_3801 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6190) );
  AND2X2 AND2X2_3802 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6192) );
  AND2X2 AND2X2_3803 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6193) );
  AND2X2 AND2X2_3804 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6196) );
  AND2X2 AND2X2_3805 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6197) );
  AND2X2 AND2X2_3806 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6199) );
  AND2X2 AND2X2_3807 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6200) );
  AND2X2 AND2X2_3808 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6206) );
  AND2X2 AND2X2_3809 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6207) );
  AND2X2 AND2X2_381 ( .A(_abc_43815_n1308), .B(_abc_43815_n1309), .Y(_abc_43815_n1310) );
  AND2X2 AND2X2_3810 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6209) );
  AND2X2 AND2X2_3811 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6210) );
  AND2X2 AND2X2_3812 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6213) );
  AND2X2 AND2X2_3813 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6214) );
  AND2X2 AND2X2_3814 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6216) );
  AND2X2 AND2X2_3815 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6217) );
  AND2X2 AND2X2_3816 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6221) );
  AND2X2 AND2X2_3817 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6222) );
  AND2X2 AND2X2_3818 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6224) );
  AND2X2 AND2X2_3819 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6225) );
  AND2X2 AND2X2_382 ( .A(_abc_43815_n1311), .B(_abc_43815_n1313), .Y(_abc_43815_n1314) );
  AND2X2 AND2X2_3820 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6228) );
  AND2X2 AND2X2_3821 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6229) );
  AND2X2 AND2X2_3822 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6231) );
  AND2X2 AND2X2_3823 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6232) );
  AND2X2 AND2X2_3824 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6237) );
  AND2X2 AND2X2_3825 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6238) );
  AND2X2 AND2X2_3826 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6240) );
  AND2X2 AND2X2_3827 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6241) );
  AND2X2 AND2X2_3828 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6244) );
  AND2X2 AND2X2_3829 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6245) );
  AND2X2 AND2X2_383 ( .A(_abc_43815_n1315), .B(_abc_43815_n1317), .Y(_abc_43815_n1318) );
  AND2X2 AND2X2_3830 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6246) );
  AND2X2 AND2X2_3831 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6250) );
  AND2X2 AND2X2_3832 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6251) );
  AND2X2 AND2X2_3833 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6253) );
  AND2X2 AND2X2_3834 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6254) );
  AND2X2 AND2X2_3835 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6257) );
  AND2X2 AND2X2_3836 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6258) );
  AND2X2 AND2X2_3837 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6260) );
  AND2X2 AND2X2_3838 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6261) );
  AND2X2 AND2X2_3839 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6267) );
  AND2X2 AND2X2_384 ( .A(_abc_43815_n1319_1), .B(_abc_43815_n1320_1), .Y(_abc_43815_n1321) );
  AND2X2 AND2X2_3840 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6268) );
  AND2X2 AND2X2_3841 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6270) );
  AND2X2 AND2X2_3842 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6271) );
  AND2X2 AND2X2_3843 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6274) );
  AND2X2 AND2X2_3844 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6275) );
  AND2X2 AND2X2_3845 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6277) );
  AND2X2 AND2X2_3846 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6278) );
  AND2X2 AND2X2_3847 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6282) );
  AND2X2 AND2X2_3848 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6283) );
  AND2X2 AND2X2_3849 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6285) );
  AND2X2 AND2X2_385 ( .A(_abc_43815_n1321), .B(_abc_43815_n1292), .Y(_abc_43815_n1322) );
  AND2X2 AND2X2_3850 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6286) );
  AND2X2 AND2X2_3851 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6289) );
  AND2X2 AND2X2_3852 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6290) );
  AND2X2 AND2X2_3853 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6292) );
  AND2X2 AND2X2_3854 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6293) );
  AND2X2 AND2X2_3855 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6298) );
  AND2X2 AND2X2_3856 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6299) );
  AND2X2 AND2X2_3857 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6301) );
  AND2X2 AND2X2_3858 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6302) );
  AND2X2 AND2X2_3859 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6305) );
  AND2X2 AND2X2_386 ( .A(_abc_43815_n1288), .B(_abc_43815_n995), .Y(_abc_43815_n1323) );
  AND2X2 AND2X2_3860 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6306) );
  AND2X2 AND2X2_3861 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6307) );
  AND2X2 AND2X2_3862 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6311) );
  AND2X2 AND2X2_3863 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6312) );
  AND2X2 AND2X2_3864 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6314) );
  AND2X2 AND2X2_3865 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6315) );
  AND2X2 AND2X2_3866 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6318) );
  AND2X2 AND2X2_3867 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6319) );
  AND2X2 AND2X2_3868 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6321) );
  AND2X2 AND2X2_3869 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6322) );
  AND2X2 AND2X2_387 ( .A(_abc_43815_n1291), .B(alu_greater_than_signed_o), .Y(_abc_43815_n1324) );
  AND2X2 AND2X2_3870 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6328) );
  AND2X2 AND2X2_3871 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6329) );
  AND2X2 AND2X2_3872 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6331) );
  AND2X2 AND2X2_3873 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6332) );
  AND2X2 AND2X2_3874 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6335) );
  AND2X2 AND2X2_3875 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6336) );
  AND2X2 AND2X2_3876 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6338) );
  AND2X2 AND2X2_3877 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6339) );
  AND2X2 AND2X2_3878 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6343) );
  AND2X2 AND2X2_3879 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6344) );
  AND2X2 AND2X2_388 ( .A(_abc_43815_n1326), .B(_abc_43815_n1328), .Y(_abc_43815_n1329) );
  AND2X2 AND2X2_3880 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6346) );
  AND2X2 AND2X2_3881 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6347) );
  AND2X2 AND2X2_3882 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6350) );
  AND2X2 AND2X2_3883 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6351) );
  AND2X2 AND2X2_3884 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6353) );
  AND2X2 AND2X2_3885 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6354) );
  AND2X2 AND2X2_3886 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6359) );
  AND2X2 AND2X2_3887 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6360) );
  AND2X2 AND2X2_3888 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6362) );
  AND2X2 AND2X2_3889 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6363) );
  AND2X2 AND2X2_389 ( .A(_abc_43815_n1330), .B(_abc_43815_n1332), .Y(_abc_43815_n1333_1) );
  AND2X2 AND2X2_3890 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6366) );
  AND2X2 AND2X2_3891 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6367) );
  AND2X2 AND2X2_3892 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6368) );
  AND2X2 AND2X2_3893 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6372) );
  AND2X2 AND2X2_3894 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6373) );
  AND2X2 AND2X2_3895 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6375) );
  AND2X2 AND2X2_3896 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6376) );
  AND2X2 AND2X2_3897 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6379) );
  AND2X2 AND2X2_3898 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6380) );
  AND2X2 AND2X2_3899 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6382) );
  AND2X2 AND2X2_39 ( .A(_abc_43815_n670_1), .B(_abc_43815_n652), .Y(_abc_43815_n678) );
  AND2X2 AND2X2_390 ( .A(_abc_43815_n1334), .B(_abc_43815_n1285), .Y(_abc_43815_n1335) );
  AND2X2 AND2X2_3900 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6383) );
  AND2X2 AND2X2_3901 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6389) );
  AND2X2 AND2X2_3902 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6390) );
  AND2X2 AND2X2_3903 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6392) );
  AND2X2 AND2X2_3904 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6393) );
  AND2X2 AND2X2_3905 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6396) );
  AND2X2 AND2X2_3906 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6397) );
  AND2X2 AND2X2_3907 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6399) );
  AND2X2 AND2X2_3908 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6400) );
  AND2X2 AND2X2_3909 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6404) );
  AND2X2 AND2X2_391 ( .A(_abc_43815_n1335), .B(_abc_43815_n1257), .Y(_abc_43815_n1336_1) );
  AND2X2 AND2X2_3910 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6405) );
  AND2X2 AND2X2_3911 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6407) );
  AND2X2 AND2X2_3912 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6408) );
  AND2X2 AND2X2_3913 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6411) );
  AND2X2 AND2X2_3914 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6412) );
  AND2X2 AND2X2_3915 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6414) );
  AND2X2 AND2X2_3916 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6415) );
  AND2X2 AND2X2_3917 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6420) );
  AND2X2 AND2X2_3918 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6421) );
  AND2X2 AND2X2_3919 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6423) );
  AND2X2 AND2X2_392 ( .A(_abc_43815_n1264), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n1337) );
  AND2X2 AND2X2_3920 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6424) );
  AND2X2 AND2X2_3921 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6427) );
  AND2X2 AND2X2_3922 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6428) );
  AND2X2 AND2X2_3923 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6429) );
  AND2X2 AND2X2_3924 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6433) );
  AND2X2 AND2X2_3925 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6434) );
  AND2X2 AND2X2_3926 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6436) );
  AND2X2 AND2X2_3927 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6437) );
  AND2X2 AND2X2_3928 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6440) );
  AND2X2 AND2X2_3929 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6441) );
  AND2X2 AND2X2_393 ( .A(_abc_43815_n1341), .B(_abc_43815_n1066), .Y(_abc_43815_n1342) );
  AND2X2 AND2X2_3930 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6443) );
  AND2X2 AND2X2_3931 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6444) );
  AND2X2 AND2X2_3932 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6450) );
  AND2X2 AND2X2_3933 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6451) );
  AND2X2 AND2X2_3934 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6453) );
  AND2X2 AND2X2_3935 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6454) );
  AND2X2 AND2X2_3936 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6457) );
  AND2X2 AND2X2_3937 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6458) );
  AND2X2 AND2X2_3938 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6460) );
  AND2X2 AND2X2_3939 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6461) );
  AND2X2 AND2X2_394 ( .A(_abc_43815_n1340), .B(_abc_43815_n1342), .Y(_abc_43815_n1343) );
  AND2X2 AND2X2_3940 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6465) );
  AND2X2 AND2X2_3941 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6466) );
  AND2X2 AND2X2_3942 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6468) );
  AND2X2 AND2X2_3943 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6469) );
  AND2X2 AND2X2_3944 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6472) );
  AND2X2 AND2X2_3945 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6473) );
  AND2X2 AND2X2_3946 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6475) );
  AND2X2 AND2X2_3947 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6476) );
  AND2X2 AND2X2_3948 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6481) );
  AND2X2 AND2X2_3949 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6482) );
  AND2X2 AND2X2_395 ( .A(_abc_43815_n1065_1_bF_buf2), .B(esr_q_9_), .Y(_abc_43815_n1344) );
  AND2X2 AND2X2_3950 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6484) );
  AND2X2 AND2X2_3951 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6485) );
  AND2X2 AND2X2_3952 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6488) );
  AND2X2 AND2X2_3953 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6489) );
  AND2X2 AND2X2_3954 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6490) );
  AND2X2 AND2X2_3955 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6494) );
  AND2X2 AND2X2_3956 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6495) );
  AND2X2 AND2X2_3957 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6497) );
  AND2X2 AND2X2_3958 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6498) );
  AND2X2 AND2X2_3959 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6501) );
  AND2X2 AND2X2_396 ( .A(_abc_43815_n1346), .B(_abc_43815_n1339), .Y(_abc_43815_n1347) );
  AND2X2 AND2X2_3960 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6502) );
  AND2X2 AND2X2_3961 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6504) );
  AND2X2 AND2X2_3962 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6505) );
  AND2X2 AND2X2_3963 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6511) );
  AND2X2 AND2X2_3964 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6512) );
  AND2X2 AND2X2_3965 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6514) );
  AND2X2 AND2X2_3966 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6515) );
  AND2X2 AND2X2_3967 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6518) );
  AND2X2 AND2X2_3968 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6519) );
  AND2X2 AND2X2_3969 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6521) );
  AND2X2 AND2X2_397 ( .A(_abc_43815_n1272), .B(intr_i), .Y(_abc_43815_n1348) );
  AND2X2 AND2X2_3970 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6522) );
  AND2X2 AND2X2_3971 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6526) );
  AND2X2 AND2X2_3972 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6527) );
  AND2X2 AND2X2_3973 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6529) );
  AND2X2 AND2X2_3974 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6530) );
  AND2X2 AND2X2_3975 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6533) );
  AND2X2 AND2X2_3976 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6534) );
  AND2X2 AND2X2_3977 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6536) );
  AND2X2 AND2X2_3978 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6537) );
  AND2X2 AND2X2_3979 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6542) );
  AND2X2 AND2X2_398 ( .A(_abc_43815_n1349), .B(_abc_43815_n1196), .Y(_abc_43815_n1350) );
  AND2X2 AND2X2_3980 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6543) );
  AND2X2 AND2X2_3981 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6545) );
  AND2X2 AND2X2_3982 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6546) );
  AND2X2 AND2X2_3983 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6549) );
  AND2X2 AND2X2_3984 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6550) );
  AND2X2 AND2X2_3985 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6551) );
  AND2X2 AND2X2_3986 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6555) );
  AND2X2 AND2X2_3987 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6556) );
  AND2X2 AND2X2_3988 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6558) );
  AND2X2 AND2X2_3989 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6559) );
  AND2X2 AND2X2_399 ( .A(_abc_43815_n1193), .B(_abc_43815_n1098), .Y(_abc_43815_n1351) );
  AND2X2 AND2X2_3990 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6562) );
  AND2X2 AND2X2_3991 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6563) );
  AND2X2 AND2X2_3992 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6565) );
  AND2X2 AND2X2_3993 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6566) );
  AND2X2 AND2X2_3994 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6572) );
  AND2X2 AND2X2_3995 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6573) );
  AND2X2 AND2X2_3996 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6575) );
  AND2X2 AND2X2_3997 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6576) );
  AND2X2 AND2X2_3998 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6579) );
  AND2X2 AND2X2_3999 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6580) );
  AND2X2 AND2X2_4 ( .A(_abc_43815_n625), .B(inst_r_3_), .Y(_abc_43815_n626) );
  AND2X2 AND2X2_40 ( .A(_abc_43815_n679_1), .B(state_q_5_), .Y(_abc_43815_n680_1) );
  AND2X2 AND2X2_400 ( .A(_abc_43815_n1351_bF_buf4), .B(_abc_43815_n1350_bF_buf4), .Y(_abc_43815_n1352_1) );
  AND2X2 AND2X2_4000 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6582) );
  AND2X2 AND2X2_4001 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6583) );
  AND2X2 AND2X2_4002 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6587) );
  AND2X2 AND2X2_4003 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6588) );
  AND2X2 AND2X2_4004 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6590) );
  AND2X2 AND2X2_4005 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6591) );
  AND2X2 AND2X2_4006 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6594) );
  AND2X2 AND2X2_4007 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6595) );
  AND2X2 AND2X2_4008 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6597) );
  AND2X2 AND2X2_4009 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6598) );
  AND2X2 AND2X2_401 ( .A(_abc_43815_n1347), .B(_abc_43815_n1353_1), .Y(_abc_43815_n1354) );
  AND2X2 AND2X2_4010 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6603) );
  AND2X2 AND2X2_4011 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6604) );
  AND2X2 AND2X2_4012 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6606) );
  AND2X2 AND2X2_4013 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6607) );
  AND2X2 AND2X2_4014 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6610) );
  AND2X2 AND2X2_4015 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6611) );
  AND2X2 AND2X2_4016 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6612) );
  AND2X2 AND2X2_4017 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6616) );
  AND2X2 AND2X2_4018 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6617) );
  AND2X2 AND2X2_4019 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6619) );
  AND2X2 AND2X2_402 ( .A(_abc_43815_n1240), .B(_abc_43815_n1356), .Y(_abc_43815_n1357) );
  AND2X2 AND2X2_4020 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6620) );
  AND2X2 AND2X2_4021 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6623) );
  AND2X2 AND2X2_4022 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6624) );
  AND2X2 AND2X2_4023 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6626) );
  AND2X2 AND2X2_4024 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6627) );
  AND2X2 AND2X2_4025 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6633) );
  AND2X2 AND2X2_4026 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6634) );
  AND2X2 AND2X2_4027 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6636) );
  AND2X2 AND2X2_4028 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6637) );
  AND2X2 AND2X2_4029 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6640) );
  AND2X2 AND2X2_403 ( .A(_abc_43815_n1358), .B(_abc_43815_n1355), .Y(_abc_43815_n1359) );
  AND2X2 AND2X2_4030 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6641) );
  AND2X2 AND2X2_4031 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6643) );
  AND2X2 AND2X2_4032 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6644) );
  AND2X2 AND2X2_4033 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6648) );
  AND2X2 AND2X2_4034 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6649) );
  AND2X2 AND2X2_4035 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6651) );
  AND2X2 AND2X2_4036 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6652) );
  AND2X2 AND2X2_4037 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6655) );
  AND2X2 AND2X2_4038 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6656) );
  AND2X2 AND2X2_4039 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6658) );
  AND2X2 AND2X2_404 ( .A(_abc_43815_n1352_1), .B(_abc_43815_n1359), .Y(_abc_43815_n1360_1) );
  AND2X2 AND2X2_4040 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6659) );
  AND2X2 AND2X2_4041 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6664) );
  AND2X2 AND2X2_4042 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6665) );
  AND2X2 AND2X2_4043 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6667) );
  AND2X2 AND2X2_4044 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6668) );
  AND2X2 AND2X2_4045 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6671) );
  AND2X2 AND2X2_4046 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6672) );
  AND2X2 AND2X2_4047 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6673) );
  AND2X2 AND2X2_4048 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6677) );
  AND2X2 AND2X2_4049 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6678) );
  AND2X2 AND2X2_405 ( .A(_abc_43815_n1363), .B(enable_i_bF_buf4), .Y(_abc_43815_n1364) );
  AND2X2 AND2X2_4050 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6680) );
  AND2X2 AND2X2_4051 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6681) );
  AND2X2 AND2X2_4052 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6684) );
  AND2X2 AND2X2_4053 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6685) );
  AND2X2 AND2X2_4054 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6687) );
  AND2X2 AND2X2_4055 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6688) );
  AND2X2 AND2X2_4056 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6694) );
  AND2X2 AND2X2_4057 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6695) );
  AND2X2 AND2X2_4058 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6697) );
  AND2X2 AND2X2_4059 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6698) );
  AND2X2 AND2X2_406 ( .A(_abc_43815_n1362), .B(_abc_43815_n1364), .Y(esr_q_9__FF_INPUT) );
  AND2X2 AND2X2_4060 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6701) );
  AND2X2 AND2X2_4061 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6702) );
  AND2X2 AND2X2_4062 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6704) );
  AND2X2 AND2X2_4063 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6705) );
  AND2X2 AND2X2_4064 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6709) );
  AND2X2 AND2X2_4065 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6710) );
  AND2X2 AND2X2_4066 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6712) );
  AND2X2 AND2X2_4067 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6713) );
  AND2X2 AND2X2_4068 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6716) );
  AND2X2 AND2X2_4069 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6717) );
  AND2X2 AND2X2_407 ( .A(_abc_43815_n1368), .B(_abc_43815_n1366), .Y(_abc_43815_n1369) );
  AND2X2 AND2X2_4070 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6719) );
  AND2X2 AND2X2_4071 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6720) );
  AND2X2 AND2X2_4072 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6725) );
  AND2X2 AND2X2_4073 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6726) );
  AND2X2 AND2X2_4074 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6728) );
  AND2X2 AND2X2_4075 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6729) );
  AND2X2 AND2X2_4076 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6732) );
  AND2X2 AND2X2_4077 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6733) );
  AND2X2 AND2X2_4078 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6734) );
  AND2X2 AND2X2_4079 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6738) );
  AND2X2 AND2X2_408 ( .A(_abc_43815_n1066), .B(_abc_43815_n1369), .Y(_abc_43815_n1370) );
  AND2X2 AND2X2_4080 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6739) );
  AND2X2 AND2X2_4081 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6741) );
  AND2X2 AND2X2_4082 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6742) );
  AND2X2 AND2X2_4083 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6745) );
  AND2X2 AND2X2_4084 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6746) );
  AND2X2 AND2X2_4085 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6748) );
  AND2X2 AND2X2_4086 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6749) );
  AND2X2 AND2X2_4087 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6755) );
  AND2X2 AND2X2_4088 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6756) );
  AND2X2 AND2X2_4089 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6758) );
  AND2X2 AND2X2_409 ( .A(_abc_43815_n1065_1_bF_buf1), .B(esr_q_10_), .Y(_abc_43815_n1371) );
  AND2X2 AND2X2_4090 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6759) );
  AND2X2 AND2X2_4091 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6762) );
  AND2X2 AND2X2_4092 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6763) );
  AND2X2 AND2X2_4093 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6765) );
  AND2X2 AND2X2_4094 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6766) );
  AND2X2 AND2X2_4095 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6770) );
  AND2X2 AND2X2_4096 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6771) );
  AND2X2 AND2X2_4097 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6773) );
  AND2X2 AND2X2_4098 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6774) );
  AND2X2 AND2X2_4099 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6777) );
  AND2X2 AND2X2_41 ( .A(_abc_43815_n682), .B(alu_p_o_0_), .Y(_abc_43815_n683) );
  AND2X2 AND2X2_410 ( .A(_abc_43815_n1221), .B(_abc_43815_n1252), .Y(_abc_43815_n1374) );
  AND2X2 AND2X2_4100 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6778) );
  AND2X2 AND2X2_4101 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6780) );
  AND2X2 AND2X2_4102 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6781) );
  AND2X2 AND2X2_4103 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6786) );
  AND2X2 AND2X2_4104 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6787) );
  AND2X2 AND2X2_4105 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6789) );
  AND2X2 AND2X2_4106 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6790) );
  AND2X2 AND2X2_4107 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6793) );
  AND2X2 AND2X2_4108 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6794) );
  AND2X2 AND2X2_4109 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6795) );
  AND2X2 AND2X2_411 ( .A(_abc_43815_n1235), .B(_abc_43815_n1228), .Y(_abc_43815_n1375_1) );
  AND2X2 AND2X2_4110 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6799) );
  AND2X2 AND2X2_4111 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6800) );
  AND2X2 AND2X2_4112 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6802) );
  AND2X2 AND2X2_4113 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6803) );
  AND2X2 AND2X2_4114 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6806) );
  AND2X2 AND2X2_4115 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6807) );
  AND2X2 AND2X2_4116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6809) );
  AND2X2 AND2X2_4117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6810) );
  AND2X2 AND2X2_4118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6816) );
  AND2X2 AND2X2_4119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6817) );
  AND2X2 AND2X2_412 ( .A(_abc_43815_n1225), .B(_abc_43815_n1222), .Y(_abc_43815_n1376) );
  AND2X2 AND2X2_4120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6819) );
  AND2X2 AND2X2_4121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6820) );
  AND2X2 AND2X2_4122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6823) );
  AND2X2 AND2X2_4123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6824) );
  AND2X2 AND2X2_4124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6826) );
  AND2X2 AND2X2_4125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6827) );
  AND2X2 AND2X2_4126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6831) );
  AND2X2 AND2X2_4127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6832) );
  AND2X2 AND2X2_4128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6834) );
  AND2X2 AND2X2_4129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6835) );
  AND2X2 AND2X2_413 ( .A(_abc_43815_n1375_1), .B(_abc_43815_n1376), .Y(_abc_43815_n1377) );
  AND2X2 AND2X2_4130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6838) );
  AND2X2 AND2X2_4131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6839) );
  AND2X2 AND2X2_4132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6841) );
  AND2X2 AND2X2_4133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6842) );
  AND2X2 AND2X2_4134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6847) );
  AND2X2 AND2X2_4135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6848) );
  AND2X2 AND2X2_4136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6850) );
  AND2X2 AND2X2_4137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6851) );
  AND2X2 AND2X2_4138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6854) );
  AND2X2 AND2X2_4139 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6855) );
  AND2X2 AND2X2_414 ( .A(_abc_43815_n1374), .B(_abc_43815_n1377), .Y(_abc_43815_n1378) );
  AND2X2 AND2X2_4140 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6856) );
  AND2X2 AND2X2_4141 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6860) );
  AND2X2 AND2X2_4142 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6861) );
  AND2X2 AND2X2_4143 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6863) );
  AND2X2 AND2X2_4144 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6864) );
  AND2X2 AND2X2_4145 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6867) );
  AND2X2 AND2X2_4146 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6868) );
  AND2X2 AND2X2_4147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6870) );
  AND2X2 AND2X2_4148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6871) );
  AND2X2 AND2X2_4149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6877) );
  AND2X2 AND2X2_415 ( .A(_abc_43815_n1378), .B(_abc_43815_n1216), .Y(_abc_43815_n1379) );
  AND2X2 AND2X2_4150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6878) );
  AND2X2 AND2X2_4151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6880) );
  AND2X2 AND2X2_4152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6881) );
  AND2X2 AND2X2_4153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6884) );
  AND2X2 AND2X2_4154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6885) );
  AND2X2 AND2X2_4155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6887) );
  AND2X2 AND2X2_4156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6888) );
  AND2X2 AND2X2_4157 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6892) );
  AND2X2 AND2X2_4158 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6893) );
  AND2X2 AND2X2_4159 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6895) );
  AND2X2 AND2X2_416 ( .A(_abc_43815_n1379), .B(_abc_43815_n1381), .Y(_abc_43815_n1382) );
  AND2X2 AND2X2_4160 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6896) );
  AND2X2 AND2X2_4161 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6899) );
  AND2X2 AND2X2_4162 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6900) );
  AND2X2 AND2X2_4163 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6902) );
  AND2X2 AND2X2_4164 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6903) );
  AND2X2 AND2X2_4165 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6908) );
  AND2X2 AND2X2_4166 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6909) );
  AND2X2 AND2X2_4167 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6911) );
  AND2X2 AND2X2_4168 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6912) );
  AND2X2 AND2X2_4169 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6915) );
  AND2X2 AND2X2_417 ( .A(_abc_43815_n1383), .B(_abc_43815_n1380), .Y(_abc_43815_n1384) );
  AND2X2 AND2X2_4170 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6916) );
  AND2X2 AND2X2_4171 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6917) );
  AND2X2 AND2X2_4172 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6921) );
  AND2X2 AND2X2_4173 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6922) );
  AND2X2 AND2X2_4174 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6924) );
  AND2X2 AND2X2_4175 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6925) );
  AND2X2 AND2X2_4176 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6928) );
  AND2X2 AND2X2_4177 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6929) );
  AND2X2 AND2X2_4178 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6931) );
  AND2X2 AND2X2_4179 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6932) );
  AND2X2 AND2X2_418 ( .A(_abc_43815_n1385), .B(_abc_43815_n1373), .Y(_abc_43815_n1386) );
  AND2X2 AND2X2_4180 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6938) );
  AND2X2 AND2X2_4181 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6939) );
  AND2X2 AND2X2_4182 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6941) );
  AND2X2 AND2X2_4183 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6942) );
  AND2X2 AND2X2_4184 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6945) );
  AND2X2 AND2X2_4185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6946) );
  AND2X2 AND2X2_4186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6948) );
  AND2X2 AND2X2_4187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6949) );
  AND2X2 AND2X2_4188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6953) );
  AND2X2 AND2X2_4189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6954) );
  AND2X2 AND2X2_419 ( .A(_abc_43815_n1353_1), .B(_abc_43815_n1386), .Y(_abc_43815_n1387) );
  AND2X2 AND2X2_4190 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6956) );
  AND2X2 AND2X2_4191 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6957) );
  AND2X2 AND2X2_4192 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6960) );
  AND2X2 AND2X2_4193 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6961) );
  AND2X2 AND2X2_4194 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6963) );
  AND2X2 AND2X2_4195 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6964) );
  AND2X2 AND2X2_4196 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6969) );
  AND2X2 AND2X2_4197 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6970) );
  AND2X2 AND2X2_4198 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6972) );
  AND2X2 AND2X2_4199 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6973) );
  AND2X2 AND2X2_42 ( .A(_abc_43815_n666), .B(_abc_43815_n653), .Y(_abc_43815_n684) );
  AND2X2 AND2X2_420 ( .A(_abc_43815_n1240), .B(_abc_43815_n1381), .Y(_abc_43815_n1389) );
  AND2X2 AND2X2_4200 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6976) );
  AND2X2 AND2X2_4201 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6977) );
  AND2X2 AND2X2_4202 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6978) );
  AND2X2 AND2X2_4203 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6982) );
  AND2X2 AND2X2_4204 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6983) );
  AND2X2 AND2X2_4205 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6985) );
  AND2X2 AND2X2_4206 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6986) );
  AND2X2 AND2X2_4207 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6989) );
  AND2X2 AND2X2_4208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6990) );
  AND2X2 AND2X2_4209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6992) );
  AND2X2 AND2X2_421 ( .A(_abc_43815_n1390), .B(_abc_43815_n1388), .Y(_abc_43815_n1391_1) );
  AND2X2 AND2X2_4210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6993) );
  AND2X2 AND2X2_4211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n6999) );
  AND2X2 AND2X2_4212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7000) );
  AND2X2 AND2X2_4213 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7002) );
  AND2X2 AND2X2_4214 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7003) );
  AND2X2 AND2X2_4215 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7006) );
  AND2X2 AND2X2_4216 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7007) );
  AND2X2 AND2X2_4217 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7009) );
  AND2X2 AND2X2_4218 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7010) );
  AND2X2 AND2X2_4219 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7014) );
  AND2X2 AND2X2_422 ( .A(_abc_43815_n1352_1), .B(_abc_43815_n1391_1), .Y(_abc_43815_n1392_1) );
  AND2X2 AND2X2_4220 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7015) );
  AND2X2 AND2X2_4221 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7017) );
  AND2X2 AND2X2_4222 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7018) );
  AND2X2 AND2X2_4223 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7021) );
  AND2X2 AND2X2_4224 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7022) );
  AND2X2 AND2X2_4225 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7024) );
  AND2X2 AND2X2_4226 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7025) );
  AND2X2 AND2X2_4227 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7030) );
  AND2X2 AND2X2_4228 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7031) );
  AND2X2 AND2X2_4229 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7033) );
  AND2X2 AND2X2_423 ( .A(_abc_43815_n1395), .B(enable_i_bF_buf3), .Y(_abc_43815_n1396) );
  AND2X2 AND2X2_4230 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7034) );
  AND2X2 AND2X2_4231 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7037) );
  AND2X2 AND2X2_4232 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7038) );
  AND2X2 AND2X2_4233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7039) );
  AND2X2 AND2X2_4234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7043) );
  AND2X2 AND2X2_4235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7044) );
  AND2X2 AND2X2_4236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7046) );
  AND2X2 AND2X2_4237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7047) );
  AND2X2 AND2X2_4238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7050) );
  AND2X2 AND2X2_4239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7051) );
  AND2X2 AND2X2_424 ( .A(_abc_43815_n1394), .B(_abc_43815_n1396), .Y(esr_q_10__FF_INPUT) );
  AND2X2 AND2X2_4240 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7053) );
  AND2X2 AND2X2_4241 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7054) );
  AND2X2 AND2X2_4242 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7060) );
  AND2X2 AND2X2_4243 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7061) );
  AND2X2 AND2X2_4244 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7063) );
  AND2X2 AND2X2_4245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7064) );
  AND2X2 AND2X2_4246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7067) );
  AND2X2 AND2X2_4247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7068) );
  AND2X2 AND2X2_4248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7070) );
  AND2X2 AND2X2_4249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7071) );
  AND2X2 AND2X2_425 ( .A(_abc_43815_n1351_bF_buf3), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .Y(_abc_43815_n1398) );
  AND2X2 AND2X2_4250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7075) );
  AND2X2 AND2X2_4251 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7076) );
  AND2X2 AND2X2_4252 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7078) );
  AND2X2 AND2X2_4253 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7079) );
  AND2X2 AND2X2_4254 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7082) );
  AND2X2 AND2X2_4255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7083) );
  AND2X2 AND2X2_4256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7085) );
  AND2X2 AND2X2_4257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7086) );
  AND2X2 AND2X2_4258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7091) );
  AND2X2 AND2X2_4259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7092) );
  AND2X2 AND2X2_426 ( .A(_abc_43815_n1398), .B(_abc_43815_n1350_bF_buf3), .Y(_abc_43815_n1399) );
  AND2X2 AND2X2_4260 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7094) );
  AND2X2 AND2X2_4261 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7095) );
  AND2X2 AND2X2_4262 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7098) );
  AND2X2 AND2X2_4263 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7099) );
  AND2X2 AND2X2_4264 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7100) );
  AND2X2 AND2X2_4265 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7104) );
  AND2X2 AND2X2_4266 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7105) );
  AND2X2 AND2X2_4267 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7107) );
  AND2X2 AND2X2_4268 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7108) );
  AND2X2 AND2X2_4269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7111) );
  AND2X2 AND2X2_427 ( .A(_abc_43815_n1399_bF_buf4), .B(_abc_43815_n1272), .Y(_abc_43815_n1400) );
  AND2X2 AND2X2_4270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7112) );
  AND2X2 AND2X2_4271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7114) );
  AND2X2 AND2X2_4272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7115) );
  AND2X2 AND2X2_4273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7121) );
  AND2X2 AND2X2_4274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7122) );
  AND2X2 AND2X2_4275 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7124) );
  AND2X2 AND2X2_4276 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7125) );
  AND2X2 AND2X2_4277 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7128) );
  AND2X2 AND2X2_4278 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7129) );
  AND2X2 AND2X2_4279 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7131) );
  AND2X2 AND2X2_428 ( .A(_abc_43815_n1278_bF_buf4), .B(sr_q_2_), .Y(_abc_43815_n1401) );
  AND2X2 AND2X2_4280 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7132) );
  AND2X2 AND2X2_4281 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7136) );
  AND2X2 AND2X2_4282 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7137) );
  AND2X2 AND2X2_4283 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7139) );
  AND2X2 AND2X2_4284 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7140) );
  AND2X2 AND2X2_4285 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7143) );
  AND2X2 AND2X2_4286 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7144) );
  AND2X2 AND2X2_4287 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7146) );
  AND2X2 AND2X2_4288 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7147) );
  AND2X2 AND2X2_4289 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7152) );
  AND2X2 AND2X2_429 ( .A(_abc_43815_n1402), .B(enable_i_bF_buf2), .Y(sr_q_2__FF_INPUT) );
  AND2X2 AND2X2_4290 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7153) );
  AND2X2 AND2X2_4291 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7155) );
  AND2X2 AND2X2_4292 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7156) );
  AND2X2 AND2X2_4293 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7159) );
  AND2X2 AND2X2_4294 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7160) );
  AND2X2 AND2X2_4295 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7161) );
  AND2X2 AND2X2_4296 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7165) );
  AND2X2 AND2X2_4297 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7166) );
  AND2X2 AND2X2_4298 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7168) );
  AND2X2 AND2X2_4299 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7169) );
  AND2X2 AND2X2_43 ( .A(_abc_43815_n687), .B(_abc_43815_n688), .Y(_abc_43815_n689) );
  AND2X2 AND2X2_430 ( .A(_abc_43815_n1347), .B(_abc_43815_n1399_bF_buf3), .Y(_abc_43815_n1404) );
  AND2X2 AND2X2_4300 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7172) );
  AND2X2 AND2X2_4301 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7173) );
  AND2X2 AND2X2_4302 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7175) );
  AND2X2 AND2X2_4303 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7176) );
  AND2X2 AND2X2_4304 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7182) );
  AND2X2 AND2X2_4305 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7183) );
  AND2X2 AND2X2_4306 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7185) );
  AND2X2 AND2X2_4307 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7186) );
  AND2X2 AND2X2_4308 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7189) );
  AND2X2 AND2X2_4309 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7190) );
  AND2X2 AND2X2_431 ( .A(_abc_43815_n1278_bF_buf3), .B(sr_q_9_), .Y(_abc_43815_n1405_1) );
  AND2X2 AND2X2_4310 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7192) );
  AND2X2 AND2X2_4311 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7193) );
  AND2X2 AND2X2_4312 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7197) );
  AND2X2 AND2X2_4313 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7198) );
  AND2X2 AND2X2_4314 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7200) );
  AND2X2 AND2X2_4315 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7201) );
  AND2X2 AND2X2_4316 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7204) );
  AND2X2 AND2X2_4317 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7205) );
  AND2X2 AND2X2_4318 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7207) );
  AND2X2 AND2X2_4319 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7208) );
  AND2X2 AND2X2_432 ( .A(_abc_43815_n1406), .B(enable_i_bF_buf1), .Y(sr_q_9__FF_INPUT) );
  AND2X2 AND2X2_4320 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7213) );
  AND2X2 AND2X2_4321 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7214) );
  AND2X2 AND2X2_4322 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7216) );
  AND2X2 AND2X2_4323 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7217) );
  AND2X2 AND2X2_4324 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7220) );
  AND2X2 AND2X2_4325 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7221) );
  AND2X2 AND2X2_4326 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7222) );
  AND2X2 AND2X2_4327 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7226) );
  AND2X2 AND2X2_4328 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7227) );
  AND2X2 AND2X2_4329 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7229) );
  AND2X2 AND2X2_433 ( .A(_abc_43815_n1278_bF_buf2), .B(alu_c_i), .Y(_abc_43815_n1408_1) );
  AND2X2 AND2X2_4330 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7230) );
  AND2X2 AND2X2_4331 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7233) );
  AND2X2 AND2X2_4332 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7234) );
  AND2X2 AND2X2_4333 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7236) );
  AND2X2 AND2X2_4334 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7237) );
  AND2X2 AND2X2_4335 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7243) );
  AND2X2 AND2X2_4336 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7244) );
  AND2X2 AND2X2_4337 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7246) );
  AND2X2 AND2X2_4338 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7247) );
  AND2X2 AND2X2_4339 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7250) );
  AND2X2 AND2X2_434 ( .A(_abc_43815_n1399_bF_buf2), .B(_abc_43815_n1386), .Y(_abc_43815_n1409) );
  AND2X2 AND2X2_4340 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7251) );
  AND2X2 AND2X2_4341 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7253) );
  AND2X2 AND2X2_4342 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7254) );
  AND2X2 AND2X2_4343 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7258) );
  AND2X2 AND2X2_4344 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7259) );
  AND2X2 AND2X2_4345 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7261) );
  AND2X2 AND2X2_4346 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7262) );
  AND2X2 AND2X2_4347 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7265) );
  AND2X2 AND2X2_4348 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7266) );
  AND2X2 AND2X2_4349 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7268) );
  AND2X2 AND2X2_435 ( .A(_abc_43815_n1410), .B(enable_i_bF_buf0), .Y(sr_q_10__FF_INPUT) );
  AND2X2 AND2X2_4350 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7269) );
  AND2X2 AND2X2_4351 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7274) );
  AND2X2 AND2X2_4352 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7275) );
  AND2X2 AND2X2_4353 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7277) );
  AND2X2 AND2X2_4354 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7278) );
  AND2X2 AND2X2_4355 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7281) );
  AND2X2 AND2X2_4356 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7282) );
  AND2X2 AND2X2_4357 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7283) );
  AND2X2 AND2X2_4358 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7287) );
  AND2X2 AND2X2_4359 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7288) );
  AND2X2 AND2X2_436 ( .A(_abc_43815_n1251), .B(_abc_43815_n1234), .Y(_abc_43815_n1414) );
  AND2X2 AND2X2_4360 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7290) );
  AND2X2 AND2X2_4361 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7291) );
  AND2X2 AND2X2_4362 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7294) );
  AND2X2 AND2X2_4363 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7295) );
  AND2X2 AND2X2_4364 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7297) );
  AND2X2 AND2X2_4365 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7298) );
  AND2X2 AND2X2_4366 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7304) );
  AND2X2 AND2X2_4367 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7305) );
  AND2X2 AND2X2_4368 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7307) );
  AND2X2 AND2X2_4369 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7308) );
  AND2X2 AND2X2_437 ( .A(_abc_43815_n1232), .B(_abc_43815_n1414), .Y(_abc_43815_n1415) );
  AND2X2 AND2X2_4370 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7311) );
  AND2X2 AND2X2_4371 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7312) );
  AND2X2 AND2X2_4372 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7314) );
  AND2X2 AND2X2_4373 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7315) );
  AND2X2 AND2X2_4374 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7319) );
  AND2X2 AND2X2_4375 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7320) );
  AND2X2 AND2X2_4376 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7322) );
  AND2X2 AND2X2_4377 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7323) );
  AND2X2 AND2X2_4378 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7326) );
  AND2X2 AND2X2_4379 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7327) );
  AND2X2 AND2X2_438 ( .A(_abc_43815_n1227), .B(_abc_43815_n1415), .Y(_abc_43815_n1416) );
  AND2X2 AND2X2_4380 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7329) );
  AND2X2 AND2X2_4381 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7330) );
  AND2X2 AND2X2_4382 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7335) );
  AND2X2 AND2X2_4383 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7336) );
  AND2X2 AND2X2_4384 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7338) );
  AND2X2 AND2X2_4385 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7339) );
  AND2X2 AND2X2_4386 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7342) );
  AND2X2 AND2X2_4387 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7343) );
  AND2X2 AND2X2_4388 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7344) );
  AND2X2 AND2X2_4389 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7348) );
  AND2X2 AND2X2_439 ( .A(_abc_43815_n1416), .B(_abc_43815_n1216), .Y(_abc_43815_n1417) );
  AND2X2 AND2X2_4390 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7349) );
  AND2X2 AND2X2_4391 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7351) );
  AND2X2 AND2X2_4392 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7352) );
  AND2X2 AND2X2_4393 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7355) );
  AND2X2 AND2X2_4394 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7356) );
  AND2X2 AND2X2_4395 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7358) );
  AND2X2 AND2X2_4396 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7359) );
  AND2X2 AND2X2_4397 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7365) );
  AND2X2 AND2X2_4398 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7366) );
  AND2X2 AND2X2_4399 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7368) );
  AND2X2 AND2X2_44 ( .A(_abc_43815_n665), .B(_abc_43815_n690), .Y(_abc_43815_n691) );
  AND2X2 AND2X2_440 ( .A(_abc_43815_n1417), .B(_abc_43815_n1080), .Y(_abc_43815_n1418) );
  AND2X2 AND2X2_4400 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7369) );
  AND2X2 AND2X2_4401 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7372) );
  AND2X2 AND2X2_4402 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7373) );
  AND2X2 AND2X2_4403 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7375) );
  AND2X2 AND2X2_4404 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7376) );
  AND2X2 AND2X2_4405 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7380) );
  AND2X2 AND2X2_4406 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7381) );
  AND2X2 AND2X2_4407 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7383) );
  AND2X2 AND2X2_4408 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7384) );
  AND2X2 AND2X2_4409 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7387) );
  AND2X2 AND2X2_441 ( .A(_abc_43815_n1418_bF_buf4), .B(_abc_43815_n1420), .Y(_abc_43815_n1421) );
  AND2X2 AND2X2_4410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7388) );
  AND2X2 AND2X2_4411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7390) );
  AND2X2 AND2X2_4412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7391) );
  AND2X2 AND2X2_4413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7396) );
  AND2X2 AND2X2_4414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7397) );
  AND2X2 AND2X2_4415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7399) );
  AND2X2 AND2X2_4416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7400) );
  AND2X2 AND2X2_4417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7403) );
  AND2X2 AND2X2_4418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7404) );
  AND2X2 AND2X2_4419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7405) );
  AND2X2 AND2X2_442 ( .A(_abc_43815_n1422), .B(_abc_43815_n1419), .Y(_abc_43815_n1423) );
  AND2X2 AND2X2_4420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7409) );
  AND2X2 AND2X2_4421 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7410) );
  AND2X2 AND2X2_4422 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7412) );
  AND2X2 AND2X2_4423 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7413) );
  AND2X2 AND2X2_4424 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7416) );
  AND2X2 AND2X2_4425 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7417) );
  AND2X2 AND2X2_4426 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7419) );
  AND2X2 AND2X2_4427 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7420) );
  AND2X2 AND2X2_4428 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7426) );
  AND2X2 AND2X2_4429 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7427) );
  AND2X2 AND2X2_443 ( .A(_abc_43815_n1098), .B(_abc_43815_n1066), .Y(_abc_43815_n1425_1) );
  AND2X2 AND2X2_4430 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7429) );
  AND2X2 AND2X2_4431 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7430) );
  AND2X2 AND2X2_4432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7433) );
  AND2X2 AND2X2_4433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7434) );
  AND2X2 AND2X2_4434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7436) );
  AND2X2 AND2X2_4435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7437) );
  AND2X2 AND2X2_4436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7441) );
  AND2X2 AND2X2_4437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7442) );
  AND2X2 AND2X2_4438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7444) );
  AND2X2 AND2X2_4439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7445) );
  AND2X2 AND2X2_444 ( .A(_abc_43815_n1425_1_bF_buf4), .B(next_pc_r_0_), .Y(_abc_43815_n1426) );
  AND2X2 AND2X2_4440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7448) );
  AND2X2 AND2X2_4441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7449) );
  AND2X2 AND2X2_4442 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7451) );
  AND2X2 AND2X2_4443 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7452) );
  AND2X2 AND2X2_4444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7457) );
  AND2X2 AND2X2_4445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7458) );
  AND2X2 AND2X2_4446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7460) );
  AND2X2 AND2X2_4447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7461) );
  AND2X2 AND2X2_4448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7464) );
  AND2X2 AND2X2_4449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7465) );
  AND2X2 AND2X2_445 ( .A(_abc_43815_n1065_1_bF_buf0), .B(epc_q_0_), .Y(_abc_43815_n1427) );
  AND2X2 AND2X2_4450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7466) );
  AND2X2 AND2X2_4451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7470) );
  AND2X2 AND2X2_4452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7471) );
  AND2X2 AND2X2_4453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7473) );
  AND2X2 AND2X2_4454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7474) );
  AND2X2 AND2X2_4455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7477) );
  AND2X2 AND2X2_4456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7478) );
  AND2X2 AND2X2_4457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7480) );
  AND2X2 AND2X2_4458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7481) );
  AND2X2 AND2X2_4459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7487) );
  AND2X2 AND2X2_446 ( .A(_abc_43815_n1430), .B(_abc_43815_n1432), .Y(_abc_43815_n1433) );
  AND2X2 AND2X2_4460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7488) );
  AND2X2 AND2X2_4461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7490) );
  AND2X2 AND2X2_4462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7491) );
  AND2X2 AND2X2_4463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7494) );
  AND2X2 AND2X2_4464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7495) );
  AND2X2 AND2X2_4465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7497) );
  AND2X2 AND2X2_4466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7498) );
  AND2X2 AND2X2_4467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7502) );
  AND2X2 AND2X2_4468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7503) );
  AND2X2 AND2X2_4469 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7505) );
  AND2X2 AND2X2_447 ( .A(_abc_43815_n1424_1), .B(_abc_43815_n1434), .Y(_abc_43815_n1435) );
  AND2X2 AND2X2_4470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7506) );
  AND2X2 AND2X2_4471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7509) );
  AND2X2 AND2X2_4472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7510) );
  AND2X2 AND2X2_4473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7512) );
  AND2X2 AND2X2_4474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7513) );
  AND2X2 AND2X2_4475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7518) );
  AND2X2 AND2X2_4476 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7519) );
  AND2X2 AND2X2_4477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7521) );
  AND2X2 AND2X2_4478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7522) );
  AND2X2 AND2X2_4479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7525) );
  AND2X2 AND2X2_448 ( .A(_abc_43815_n1435), .B(_abc_43815_n1351_bF_buf2), .Y(_abc_43815_n1436) );
  AND2X2 AND2X2_4480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7526) );
  AND2X2 AND2X2_4481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7527) );
  AND2X2 AND2X2_4482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7531) );
  AND2X2 AND2X2_4483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7532) );
  AND2X2 AND2X2_4484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7534) );
  AND2X2 AND2X2_4485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7535) );
  AND2X2 AND2X2_4486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7538) );
  AND2X2 AND2X2_4487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7539) );
  AND2X2 AND2X2_4488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7541) );
  AND2X2 AND2X2_4489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7542) );
  AND2X2 AND2X2_449 ( .A(_abc_43815_n1438), .B(enable_i_bF_buf7), .Y(_abc_43815_n1439) );
  AND2X2 AND2X2_4490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7549), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7550) );
  AND2X2 AND2X2_4491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7550), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7551) );
  AND2X2 AND2X2_4492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7552), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7553) );
  AND2X2 AND2X2_4493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7551), .B(REGFILE_SIM_reg_bank__abc_33898_n7553), .Y(REGFILE_SIM_reg_bank__abc_33898_n7554) );
  AND2X2 AND2X2_4494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7555) );
  AND2X2 AND2X2_4495 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7556) );
  AND2X2 AND2X2_4496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7551), .B(REGFILE_SIM_reg_bank__abc_33898_n7556), .Y(REGFILE_SIM_reg_bank__abc_33898_n7557) );
  AND2X2 AND2X2_4497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7558) );
  AND2X2 AND2X2_4498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7549), .B(REGFILE_SIM_reg_bank__abc_33898_n7560), .Y(REGFILE_SIM_reg_bank__abc_33898_n7561) );
  AND2X2 AND2X2_4499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7561), .B(REGFILE_SIM_reg_bank__abc_33898_n7553), .Y(REGFILE_SIM_reg_bank__abc_33898_n7562) );
  AND2X2 AND2X2_45 ( .A(_abc_43815_n693), .B(_abc_43815_n689), .Y(_abc_43815_n694) );
  AND2X2 AND2X2_450 ( .A(_abc_43815_n1437), .B(_abc_43815_n1439), .Y(epc_q_0__FF_INPUT) );
  AND2X2 AND2X2_4500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7562), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7563) );
  AND2X2 AND2X2_4501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7564) );
  AND2X2 AND2X2_4502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7561), .B(REGFILE_SIM_reg_bank__abc_33898_n7556), .Y(REGFILE_SIM_reg_bank__abc_33898_n7565) );
  AND2X2 AND2X2_4503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7565), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7566) );
  AND2X2 AND2X2_4504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7567) );
  AND2X2 AND2X2_4505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7570), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7571) );
  AND2X2 AND2X2_4506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7560), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7572) );
  AND2X2 AND2X2_4507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7571), .B(REGFILE_SIM_reg_bank__abc_33898_n7572), .Y(REGFILE_SIM_reg_bank__abc_33898_n7573) );
  AND2X2 AND2X2_4508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7573), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7574) );
  AND2X2 AND2X2_4509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7575) );
  AND2X2 AND2X2_451 ( .A(_abc_43815_n1418_bF_buf2), .B(_abc_43815_n1442), .Y(_abc_43815_n1443_1) );
  AND2X2 AND2X2_4510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7572), .B(REGFILE_SIM_reg_bank__abc_33898_n7556), .Y(REGFILE_SIM_reg_bank__abc_33898_n7576) );
  AND2X2 AND2X2_4511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7576), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7577) );
  AND2X2 AND2X2_4512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7578) );
  AND2X2 AND2X2_4513 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7580) );
  AND2X2 AND2X2_4514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7571), .B(REGFILE_SIM_reg_bank__abc_33898_n7580), .Y(REGFILE_SIM_reg_bank__abc_33898_n7581) );
  AND2X2 AND2X2_4515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7581), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7582) );
  AND2X2 AND2X2_4516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7583) );
  AND2X2 AND2X2_4517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7553), .B(REGFILE_SIM_reg_bank__abc_33898_n7580), .Y(REGFILE_SIM_reg_bank__abc_33898_n7584) );
  AND2X2 AND2X2_4518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7584), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7585) );
  AND2X2 AND2X2_4519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7586) );
  AND2X2 AND2X2_452 ( .A(_abc_43815_n1444), .B(_abc_43815_n1441), .Y(_abc_43815_n1445) );
  AND2X2 AND2X2_4520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7562), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7590) );
  AND2X2 AND2X2_4521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7591) );
  AND2X2 AND2X2_4522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7565), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7592) );
  AND2X2 AND2X2_4523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7593) );
  AND2X2 AND2X2_4524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7550), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7595) );
  AND2X2 AND2X2_4525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7595), .B(REGFILE_SIM_reg_bank__abc_33898_n7571), .Y(REGFILE_SIM_reg_bank__abc_33898_n7596) );
  AND2X2 AND2X2_4526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7597) );
  AND2X2 AND2X2_4527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7570), .B(REGFILE_SIM_reg_bank__abc_33898_n7552), .Y(REGFILE_SIM_reg_bank__abc_33898_n7598) );
  AND2X2 AND2X2_4528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7595), .B(REGFILE_SIM_reg_bank__abc_33898_n7598), .Y(REGFILE_SIM_reg_bank__abc_33898_n7599) );
  AND2X2 AND2X2_4529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7600) );
  AND2X2 AND2X2_453 ( .A(_abc_43815_n1425_1_bF_buf3), .B(next_pc_r_1_), .Y(_abc_43815_n1447) );
  AND2X2 AND2X2_4530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7584), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7603) );
  AND2X2 AND2X2_4531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7604) );
  AND2X2 AND2X2_4532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7580), .B(REGFILE_SIM_reg_bank__abc_33898_n7556), .Y(REGFILE_SIM_reg_bank__abc_33898_n7605) );
  AND2X2 AND2X2_4533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7605), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7606) );
  AND2X2 AND2X2_4534 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7607) );
  AND2X2 AND2X2_4535 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7573), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7609) );
  AND2X2 AND2X2_4536 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7610) );
  AND2X2 AND2X2_4537 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7598), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7611) );
  AND2X2 AND2X2_4538 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7611), .B(REGFILE_SIM_reg_bank__abc_33898_n7572), .Y(REGFILE_SIM_reg_bank__abc_33898_n7612) );
  AND2X2 AND2X2_4539 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7613) );
  AND2X2 AND2X2_454 ( .A(_abc_43815_n1065_1_bF_buf4), .B(epc_q_1_), .Y(_abc_43815_n1448) );
  AND2X2 AND2X2_4540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7561), .B(REGFILE_SIM_reg_bank__abc_33898_n7571), .Y(REGFILE_SIM_reg_bank__abc_33898_n7618) );
  AND2X2 AND2X2_4541 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7618), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7619) );
  AND2X2 AND2X2_4542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7620) );
  AND2X2 AND2X2_4543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7598), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7621) );
  AND2X2 AND2X2_4544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7621), .B(REGFILE_SIM_reg_bank__abc_33898_n7580), .Y(REGFILE_SIM_reg_bank__abc_33898_n7622) );
  AND2X2 AND2X2_4545 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7623) );
  AND2X2 AND2X2_4546 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7551), .B(REGFILE_SIM_reg_bank__abc_33898_n7598), .Y(REGFILE_SIM_reg_bank__abc_33898_n7625) );
  AND2X2 AND2X2_4547 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7626) );
  AND2X2 AND2X2_4548 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7551), .B(REGFILE_SIM_reg_bank__abc_33898_n7571), .Y(REGFILE_SIM_reg_bank__abc_33898_n7627) );
  AND2X2 AND2X2_4549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7628) );
  AND2X2 AND2X2_455 ( .A(_abc_43815_n1450), .B(_abc_43815_n1451), .Y(_abc_43815_n1452) );
  AND2X2 AND2X2_4550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7553), .B(REGFILE_SIM_reg_bank__abc_33898_n7572), .Y(REGFILE_SIM_reg_bank__abc_33898_n7631) );
  AND2X2 AND2X2_4551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7631), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7632) );
  AND2X2 AND2X2_4552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7633) );
  AND2X2 AND2X2_4553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7621), .B(REGFILE_SIM_reg_bank__abc_33898_n7572), .Y(REGFILE_SIM_reg_bank__abc_33898_n7634) );
  AND2X2 AND2X2_4554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7635) );
  AND2X2 AND2X2_4555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7605), .B(REGFILE_SIM_reg_bank__abc_33898_n7548), .Y(REGFILE_SIM_reg_bank__abc_33898_n7636) );
  AND2X2 AND2X2_4556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7637) );
  AND2X2 AND2X2_4557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7595), .B(REGFILE_SIM_reg_bank__abc_33898_n7553), .Y(REGFILE_SIM_reg_bank__abc_33898_n7641) );
  AND2X2 AND2X2_4558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7642) );
  AND2X2 AND2X2_4559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7595), .B(REGFILE_SIM_reg_bank__abc_33898_n7556), .Y(REGFILE_SIM_reg_bank__abc_33898_n7643) );
  AND2X2 AND2X2_456 ( .A(_abc_43815_n1446), .B(_abc_43815_n1453), .Y(_abc_43815_n1454) );
  AND2X2 AND2X2_4560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7644) );
  AND2X2 AND2X2_4561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7618), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7646) );
  AND2X2 AND2X2_4562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7647) );
  AND2X2 AND2X2_4563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7611), .B(REGFILE_SIM_reg_bank__abc_33898_n7561), .Y(REGFILE_SIM_reg_bank__abc_33898_n7648) );
  AND2X2 AND2X2_4564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7649) );
  AND2X2 AND2X2_4565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7611), .B(REGFILE_SIM_reg_bank__abc_33898_n7580), .Y(REGFILE_SIM_reg_bank__abc_33898_n7652) );
  AND2X2 AND2X2_4566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7653) );
  AND2X2 AND2X2_4567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7581), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7654) );
  AND2X2 AND2X2_4568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7655) );
  AND2X2 AND2X2_4569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7631), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7657) );
  AND2X2 AND2X2_457 ( .A(_abc_43815_n1454), .B(_abc_43815_n1351_bF_buf1), .Y(_abc_43815_n1455) );
  AND2X2 AND2X2_4570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7658) );
  AND2X2 AND2X2_4571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7576), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7659) );
  AND2X2 AND2X2_4572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7660) );
  AND2X2 AND2X2_4573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7666) );
  AND2X2 AND2X2_4574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7667) );
  AND2X2 AND2X2_4575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7669) );
  AND2X2 AND2X2_4576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7670) );
  AND2X2 AND2X2_4577 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7673) );
  AND2X2 AND2X2_4578 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7674) );
  AND2X2 AND2X2_4579 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7676) );
  AND2X2 AND2X2_458 ( .A(_abc_43815_n1458), .B(enable_i_bF_buf6), .Y(_abc_43815_n1459_1) );
  AND2X2 AND2X2_4580 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7677) );
  AND2X2 AND2X2_4581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7681) );
  AND2X2 AND2X2_4582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7682) );
  AND2X2 AND2X2_4583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7684) );
  AND2X2 AND2X2_4584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7685) );
  AND2X2 AND2X2_4585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7688) );
  AND2X2 AND2X2_4586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7689) );
  AND2X2 AND2X2_4587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7691) );
  AND2X2 AND2X2_4588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7692) );
  AND2X2 AND2X2_4589 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7697) );
  AND2X2 AND2X2_459 ( .A(_abc_43815_n1457), .B(_abc_43815_n1459_1), .Y(epc_q_1__FF_INPUT) );
  AND2X2 AND2X2_4590 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7698) );
  AND2X2 AND2X2_4591 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7700) );
  AND2X2 AND2X2_4592 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7701) );
  AND2X2 AND2X2_4593 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7704) );
  AND2X2 AND2X2_4594 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7705) );
  AND2X2 AND2X2_4595 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7706) );
  AND2X2 AND2X2_4596 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7710) );
  AND2X2 AND2X2_4597 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7711) );
  AND2X2 AND2X2_4598 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7713) );
  AND2X2 AND2X2_4599 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7714) );
  AND2X2 AND2X2_46 ( .A(_abc_43815_n694), .B(\mem_dat_i[16] ), .Y(_abc_43815_n695) );
  AND2X2 AND2X2_460 ( .A(_abc_43815_n1075), .B(_abc_43815_n1462), .Y(_abc_43815_n1463) );
  AND2X2 AND2X2_4600 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7717) );
  AND2X2 AND2X2_4601 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7718) );
  AND2X2 AND2X2_4602 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7720) );
  AND2X2 AND2X2_4603 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7721) );
  AND2X2 AND2X2_4604 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7727) );
  AND2X2 AND2X2_4605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7728) );
  AND2X2 AND2X2_4606 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7730) );
  AND2X2 AND2X2_4607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7731) );
  AND2X2 AND2X2_4608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7734) );
  AND2X2 AND2X2_4609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7735) );
  AND2X2 AND2X2_461 ( .A(_abc_43815_n1172_1_bF_buf3), .B(_abc_43815_n1049), .Y(_abc_43815_n1465) );
  AND2X2 AND2X2_4610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7737) );
  AND2X2 AND2X2_4611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7738) );
  AND2X2 AND2X2_4612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7742) );
  AND2X2 AND2X2_4613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7743) );
  AND2X2 AND2X2_4614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7745) );
  AND2X2 AND2X2_4615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7746) );
  AND2X2 AND2X2_4616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7749) );
  AND2X2 AND2X2_4617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7750) );
  AND2X2 AND2X2_4618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7752) );
  AND2X2 AND2X2_4619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7753) );
  AND2X2 AND2X2_462 ( .A(_abc_43815_n1465), .B(_abc_43815_n1071), .Y(_abc_43815_n1466) );
  AND2X2 AND2X2_4620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7758) );
  AND2X2 AND2X2_4621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7759) );
  AND2X2 AND2X2_4622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7761) );
  AND2X2 AND2X2_4623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7762) );
  AND2X2 AND2X2_4624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7765) );
  AND2X2 AND2X2_4625 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7766) );
  AND2X2 AND2X2_4626 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7767) );
  AND2X2 AND2X2_4627 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7771) );
  AND2X2 AND2X2_4628 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7772) );
  AND2X2 AND2X2_4629 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7774) );
  AND2X2 AND2X2_463 ( .A(_abc_43815_n1466), .B(_abc_43815_n1098), .Y(_abc_43815_n1467) );
  AND2X2 AND2X2_4630 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7775) );
  AND2X2 AND2X2_4631 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7778) );
  AND2X2 AND2X2_4632 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7779) );
  AND2X2 AND2X2_4633 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7781) );
  AND2X2 AND2X2_4634 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7782) );
  AND2X2 AND2X2_4635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7788) );
  AND2X2 AND2X2_4636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7789) );
  AND2X2 AND2X2_4637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7791) );
  AND2X2 AND2X2_4638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7792) );
  AND2X2 AND2X2_4639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7795) );
  AND2X2 AND2X2_464 ( .A(_abc_43815_n1073), .B(_abc_43815_n1462), .Y(_abc_43815_n1469) );
  AND2X2 AND2X2_4640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7796) );
  AND2X2 AND2X2_4641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7798) );
  AND2X2 AND2X2_4642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7799) );
  AND2X2 AND2X2_4643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7803) );
  AND2X2 AND2X2_4644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7804) );
  AND2X2 AND2X2_4645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7806) );
  AND2X2 AND2X2_4646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7807) );
  AND2X2 AND2X2_4647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7810) );
  AND2X2 AND2X2_4648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7811) );
  AND2X2 AND2X2_4649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7813) );
  AND2X2 AND2X2_465 ( .A(_abc_43815_n1471), .B(_abc_43815_n1464), .Y(_abc_43815_n1472_1) );
  AND2X2 AND2X2_4650 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7814) );
  AND2X2 AND2X2_4651 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7819) );
  AND2X2 AND2X2_4652 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7820) );
  AND2X2 AND2X2_4653 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7822) );
  AND2X2 AND2X2_4654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7823) );
  AND2X2 AND2X2_4655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7826) );
  AND2X2 AND2X2_4656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7827) );
  AND2X2 AND2X2_4657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7828) );
  AND2X2 AND2X2_4658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7832) );
  AND2X2 AND2X2_4659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7833) );
  AND2X2 AND2X2_466 ( .A(alu_op_r_0_), .B(pc_q_2_), .Y(_abc_43815_n1474) );
  AND2X2 AND2X2_4660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7835) );
  AND2X2 AND2X2_4661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7836) );
  AND2X2 AND2X2_4662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7839) );
  AND2X2 AND2X2_4663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7840) );
  AND2X2 AND2X2_4664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7842) );
  AND2X2 AND2X2_4665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7843) );
  AND2X2 AND2X2_4666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7849) );
  AND2X2 AND2X2_4667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7850) );
  AND2X2 AND2X2_4668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7852) );
  AND2X2 AND2X2_4669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7853) );
  AND2X2 AND2X2_467 ( .A(_abc_43815_n1475_1), .B(_abc_43815_n1476), .Y(_abc_43815_n1477) );
  AND2X2 AND2X2_4670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7856) );
  AND2X2 AND2X2_4671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7857) );
  AND2X2 AND2X2_4672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7859) );
  AND2X2 AND2X2_4673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7860) );
  AND2X2 AND2X2_4674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7864) );
  AND2X2 AND2X2_4675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7865) );
  AND2X2 AND2X2_4676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7867) );
  AND2X2 AND2X2_4677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7868) );
  AND2X2 AND2X2_4678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7871) );
  AND2X2 AND2X2_4679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7872) );
  AND2X2 AND2X2_468 ( .A(_abc_43815_n1425_1_bF_buf2), .B(_abc_43815_n1477), .Y(_abc_43815_n1478) );
  AND2X2 AND2X2_4680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7874) );
  AND2X2 AND2X2_4681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7875) );
  AND2X2 AND2X2_4682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7880) );
  AND2X2 AND2X2_4683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7881) );
  AND2X2 AND2X2_4684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7883) );
  AND2X2 AND2X2_4685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7884) );
  AND2X2 AND2X2_4686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7887) );
  AND2X2 AND2X2_4687 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7888) );
  AND2X2 AND2X2_4688 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7889) );
  AND2X2 AND2X2_4689 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7893) );
  AND2X2 AND2X2_469 ( .A(_abc_43815_n1065_1_bF_buf3), .B(epc_q_2_), .Y(_abc_43815_n1479) );
  AND2X2 AND2X2_4690 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7894) );
  AND2X2 AND2X2_4691 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7896) );
  AND2X2 AND2X2_4692 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7897) );
  AND2X2 AND2X2_4693 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7900) );
  AND2X2 AND2X2_4694 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7901) );
  AND2X2 AND2X2_4695 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7903) );
  AND2X2 AND2X2_4696 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7904) );
  AND2X2 AND2X2_4697 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7910) );
  AND2X2 AND2X2_4698 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7911) );
  AND2X2 AND2X2_4699 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7913) );
  AND2X2 AND2X2_47 ( .A(_abc_43815_n687), .B(mem_offset_q_1_), .Y(_abc_43815_n696) );
  AND2X2 AND2X2_470 ( .A(_abc_43815_n1481), .B(_abc_43815_n1482), .Y(_abc_43815_n1483) );
  AND2X2 AND2X2_4700 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7914) );
  AND2X2 AND2X2_4701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7917) );
  AND2X2 AND2X2_4702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7918) );
  AND2X2 AND2X2_4703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7920) );
  AND2X2 AND2X2_4704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7921) );
  AND2X2 AND2X2_4705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7925) );
  AND2X2 AND2X2_4706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7926) );
  AND2X2 AND2X2_4707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7928) );
  AND2X2 AND2X2_4708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7929) );
  AND2X2 AND2X2_4709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7932) );
  AND2X2 AND2X2_471 ( .A(_abc_43815_n1484), .B(_abc_43815_n1486), .Y(_abc_43815_n1487) );
  AND2X2 AND2X2_4710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7933) );
  AND2X2 AND2X2_4711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7935) );
  AND2X2 AND2X2_4712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7936) );
  AND2X2 AND2X2_4713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7941) );
  AND2X2 AND2X2_4714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7942) );
  AND2X2 AND2X2_4715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7944) );
  AND2X2 AND2X2_4716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7945) );
  AND2X2 AND2X2_4717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7948) );
  AND2X2 AND2X2_4718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7949) );
  AND2X2 AND2X2_4719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7950) );
  AND2X2 AND2X2_472 ( .A(_abc_43815_n1489_bF_buf4), .B(epc_q_2_), .Y(_abc_43815_n1490) );
  AND2X2 AND2X2_4720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7954) );
  AND2X2 AND2X2_4721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7955) );
  AND2X2 AND2X2_4722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7957) );
  AND2X2 AND2X2_4723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7958) );
  AND2X2 AND2X2_4724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7961) );
  AND2X2 AND2X2_4725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7962) );
  AND2X2 AND2X2_4726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7964) );
  AND2X2 AND2X2_4727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7965) );
  AND2X2 AND2X2_4728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7971) );
  AND2X2 AND2X2_4729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7972) );
  AND2X2 AND2X2_473 ( .A(_abc_43815_n1418_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n1491_1) );
  AND2X2 AND2X2_4730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7974) );
  AND2X2 AND2X2_4731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7975) );
  AND2X2 AND2X2_4732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7978) );
  AND2X2 AND2X2_4733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7979) );
  AND2X2 AND2X2_4734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7981) );
  AND2X2 AND2X2_4735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7982) );
  AND2X2 AND2X2_4736 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7986) );
  AND2X2 AND2X2_4737 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7987) );
  AND2X2 AND2X2_4738 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7989) );
  AND2X2 AND2X2_4739 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7990) );
  AND2X2 AND2X2_474 ( .A(_abc_43815_n1493), .B(_abc_43815_n1488), .Y(_abc_43815_n1494) );
  AND2X2 AND2X2_4740 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7993) );
  AND2X2 AND2X2_4741 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7994) );
  AND2X2 AND2X2_4742 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7996) );
  AND2X2 AND2X2_4743 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7997) );
  AND2X2 AND2X2_4744 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8002) );
  AND2X2 AND2X2_4745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8003) );
  AND2X2 AND2X2_4746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8005) );
  AND2X2 AND2X2_4747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8006) );
  AND2X2 AND2X2_4748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8009) );
  AND2X2 AND2X2_4749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8010) );
  AND2X2 AND2X2_475 ( .A(_abc_43815_n1495), .B(_abc_43815_n1496), .Y(_abc_43815_n1497) );
  AND2X2 AND2X2_4750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8011) );
  AND2X2 AND2X2_4751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8015) );
  AND2X2 AND2X2_4752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8016) );
  AND2X2 AND2X2_4753 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8018) );
  AND2X2 AND2X2_4754 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8019) );
  AND2X2 AND2X2_4755 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8022) );
  AND2X2 AND2X2_4756 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8023) );
  AND2X2 AND2X2_4757 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8025) );
  AND2X2 AND2X2_4758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8026) );
  AND2X2 AND2X2_4759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8032) );
  AND2X2 AND2X2_476 ( .A(_abc_43815_n1499), .B(enable_i_bF_buf5), .Y(_abc_43815_n1500) );
  AND2X2 AND2X2_4760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8033) );
  AND2X2 AND2X2_4761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8035) );
  AND2X2 AND2X2_4762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8036) );
  AND2X2 AND2X2_4763 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8039) );
  AND2X2 AND2X2_4764 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8040) );
  AND2X2 AND2X2_4765 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8042) );
  AND2X2 AND2X2_4766 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8043) );
  AND2X2 AND2X2_4767 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8047) );
  AND2X2 AND2X2_4768 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8048) );
  AND2X2 AND2X2_4769 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8050) );
  AND2X2 AND2X2_477 ( .A(_abc_43815_n1498), .B(_abc_43815_n1500), .Y(epc_q_2__FF_INPUT) );
  AND2X2 AND2X2_4770 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8051) );
  AND2X2 AND2X2_4771 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8054) );
  AND2X2 AND2X2_4772 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8055) );
  AND2X2 AND2X2_4773 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8057) );
  AND2X2 AND2X2_4774 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8058) );
  AND2X2 AND2X2_4775 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8063) );
  AND2X2 AND2X2_4776 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8064) );
  AND2X2 AND2X2_4777 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8066) );
  AND2X2 AND2X2_4778 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8067) );
  AND2X2 AND2X2_4779 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8070) );
  AND2X2 AND2X2_478 ( .A(_abc_43815_n1418_bF_buf4), .B(_abc_43815_n1503), .Y(_abc_43815_n1504) );
  AND2X2 AND2X2_4780 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8071) );
  AND2X2 AND2X2_4781 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8072) );
  AND2X2 AND2X2_4782 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8076) );
  AND2X2 AND2X2_4783 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8077) );
  AND2X2 AND2X2_4784 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8079) );
  AND2X2 AND2X2_4785 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8080) );
  AND2X2 AND2X2_4786 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8083) );
  AND2X2 AND2X2_4787 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8084) );
  AND2X2 AND2X2_4788 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8086) );
  AND2X2 AND2X2_4789 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8087) );
  AND2X2 AND2X2_479 ( .A(_abc_43815_n1505), .B(_abc_43815_n1502), .Y(_abc_43815_n1506) );
  AND2X2 AND2X2_4790 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8093) );
  AND2X2 AND2X2_4791 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8094) );
  AND2X2 AND2X2_4792 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8096) );
  AND2X2 AND2X2_4793 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8097) );
  AND2X2 AND2X2_4794 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8100) );
  AND2X2 AND2X2_4795 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8101) );
  AND2X2 AND2X2_4796 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8103) );
  AND2X2 AND2X2_4797 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8104) );
  AND2X2 AND2X2_4798 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8108) );
  AND2X2 AND2X2_4799 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8109) );
  AND2X2 AND2X2_48 ( .A(_abc_43815_n697), .B(\mem_dat_i[0] ), .Y(_abc_43815_n698) );
  AND2X2 AND2X2_480 ( .A(alu_op_r_1_), .B(pc_q_3_), .Y(_abc_43815_n1510) );
  AND2X2 AND2X2_4800 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8111) );
  AND2X2 AND2X2_4801 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8112) );
  AND2X2 AND2X2_4802 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8115) );
  AND2X2 AND2X2_4803 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8116) );
  AND2X2 AND2X2_4804 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8118) );
  AND2X2 AND2X2_4805 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8119) );
  AND2X2 AND2X2_4806 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8124) );
  AND2X2 AND2X2_4807 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8125) );
  AND2X2 AND2X2_4808 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8127) );
  AND2X2 AND2X2_4809 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8128) );
  AND2X2 AND2X2_481 ( .A(_abc_43815_n1511), .B(_abc_43815_n1509), .Y(_abc_43815_n1512) );
  AND2X2 AND2X2_4810 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8131) );
  AND2X2 AND2X2_4811 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8132) );
  AND2X2 AND2X2_4812 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8133) );
  AND2X2 AND2X2_4813 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8137) );
  AND2X2 AND2X2_4814 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8138) );
  AND2X2 AND2X2_4815 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8140) );
  AND2X2 AND2X2_4816 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8141) );
  AND2X2 AND2X2_4817 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8144) );
  AND2X2 AND2X2_4818 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8145) );
  AND2X2 AND2X2_4819 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8147) );
  AND2X2 AND2X2_482 ( .A(_abc_43815_n1512), .B(_abc_43815_n1474), .Y(_abc_43815_n1513) );
  AND2X2 AND2X2_4820 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8148) );
  AND2X2 AND2X2_4821 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8154) );
  AND2X2 AND2X2_4822 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8155) );
  AND2X2 AND2X2_4823 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8157) );
  AND2X2 AND2X2_4824 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8158) );
  AND2X2 AND2X2_4825 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8161) );
  AND2X2 AND2X2_4826 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8162) );
  AND2X2 AND2X2_4827 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8164) );
  AND2X2 AND2X2_4828 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8165) );
  AND2X2 AND2X2_4829 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8169) );
  AND2X2 AND2X2_483 ( .A(_abc_43815_n1514), .B(_abc_43815_n1515_1), .Y(_abc_43815_n1516) );
  AND2X2 AND2X2_4830 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8170) );
  AND2X2 AND2X2_4831 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8172) );
  AND2X2 AND2X2_4832 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8173) );
  AND2X2 AND2X2_4833 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8176) );
  AND2X2 AND2X2_4834 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8177) );
  AND2X2 AND2X2_4835 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8179) );
  AND2X2 AND2X2_4836 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8180) );
  AND2X2 AND2X2_4837 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8185) );
  AND2X2 AND2X2_4838 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8186) );
  AND2X2 AND2X2_4839 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8188) );
  AND2X2 AND2X2_484 ( .A(_abc_43815_n1425_1_bF_buf1), .B(_abc_43815_n1516), .Y(_abc_43815_n1517) );
  AND2X2 AND2X2_4840 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8189) );
  AND2X2 AND2X2_4841 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8192) );
  AND2X2 AND2X2_4842 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8193) );
  AND2X2 AND2X2_4843 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8194) );
  AND2X2 AND2X2_4844 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8198) );
  AND2X2 AND2X2_4845 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8199) );
  AND2X2 AND2X2_4846 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8201) );
  AND2X2 AND2X2_4847 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8202) );
  AND2X2 AND2X2_4848 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8205) );
  AND2X2 AND2X2_4849 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8206) );
  AND2X2 AND2X2_485 ( .A(_abc_43815_n1065_1_bF_buf2), .B(epc_q_3_), .Y(_abc_43815_n1518_1) );
  AND2X2 AND2X2_4850 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8208) );
  AND2X2 AND2X2_4851 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8209) );
  AND2X2 AND2X2_4852 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8215) );
  AND2X2 AND2X2_4853 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8216) );
  AND2X2 AND2X2_4854 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8218) );
  AND2X2 AND2X2_4855 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8219) );
  AND2X2 AND2X2_4856 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8222) );
  AND2X2 AND2X2_4857 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8223) );
  AND2X2 AND2X2_4858 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8225) );
  AND2X2 AND2X2_4859 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8226) );
  AND2X2 AND2X2_486 ( .A(_abc_43815_n1520), .B(_abc_43815_n1508), .Y(_abc_43815_n1521) );
  AND2X2 AND2X2_4860 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8230) );
  AND2X2 AND2X2_4861 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8231) );
  AND2X2 AND2X2_4862 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8233) );
  AND2X2 AND2X2_4863 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8234) );
  AND2X2 AND2X2_4864 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8237) );
  AND2X2 AND2X2_4865 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8238) );
  AND2X2 AND2X2_4866 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8240) );
  AND2X2 AND2X2_4867 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8241) );
  AND2X2 AND2X2_4868 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8246) );
  AND2X2 AND2X2_4869 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8247) );
  AND2X2 AND2X2_487 ( .A(pc_q_2_), .B(pc_q_3_), .Y(_abc_43815_n1524) );
  AND2X2 AND2X2_4870 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8249) );
  AND2X2 AND2X2_4871 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8250) );
  AND2X2 AND2X2_4872 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8253) );
  AND2X2 AND2X2_4873 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8254) );
  AND2X2 AND2X2_4874 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8255) );
  AND2X2 AND2X2_4875 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8259) );
  AND2X2 AND2X2_4876 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8260) );
  AND2X2 AND2X2_4877 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8262) );
  AND2X2 AND2X2_4878 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8263) );
  AND2X2 AND2X2_4879 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8266) );
  AND2X2 AND2X2_488 ( .A(_abc_43815_n1525), .B(_abc_43815_n1523), .Y(_abc_43815_n1526) );
  AND2X2 AND2X2_4880 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8267) );
  AND2X2 AND2X2_4881 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8269) );
  AND2X2 AND2X2_4882 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8270) );
  AND2X2 AND2X2_4883 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8276) );
  AND2X2 AND2X2_4884 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8277) );
  AND2X2 AND2X2_4885 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8279) );
  AND2X2 AND2X2_4886 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8280) );
  AND2X2 AND2X2_4887 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8283) );
  AND2X2 AND2X2_4888 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8284) );
  AND2X2 AND2X2_4889 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8286) );
  AND2X2 AND2X2_489 ( .A(_abc_43815_n1522), .B(_abc_43815_n1527), .Y(_abc_43815_n1528) );
  AND2X2 AND2X2_4890 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8287) );
  AND2X2 AND2X2_4891 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8291) );
  AND2X2 AND2X2_4892 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8292) );
  AND2X2 AND2X2_4893 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8294) );
  AND2X2 AND2X2_4894 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8295) );
  AND2X2 AND2X2_4895 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8298) );
  AND2X2 AND2X2_4896 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8299) );
  AND2X2 AND2X2_4897 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8301) );
  AND2X2 AND2X2_4898 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8302) );
  AND2X2 AND2X2_4899 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8307) );
  AND2X2 AND2X2_49 ( .A(_abc_43815_n699), .B(_abc_43815_n686_1_bF_buf4), .Y(_abc_43815_n700) );
  AND2X2 AND2X2_490 ( .A(_abc_43815_n1507), .B(_abc_43815_n1529), .Y(_abc_43815_n1530) );
  AND2X2 AND2X2_4900 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8308) );
  AND2X2 AND2X2_4901 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8310) );
  AND2X2 AND2X2_4902 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8311) );
  AND2X2 AND2X2_4903 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8314) );
  AND2X2 AND2X2_4904 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8315) );
  AND2X2 AND2X2_4905 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8316) );
  AND2X2 AND2X2_4906 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8320) );
  AND2X2 AND2X2_4907 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8321) );
  AND2X2 AND2X2_4908 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8323) );
  AND2X2 AND2X2_4909 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8324) );
  AND2X2 AND2X2_491 ( .A(_abc_43815_n1531), .B(_abc_43815_n1532), .Y(_abc_43815_n1533) );
  AND2X2 AND2X2_4910 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8327) );
  AND2X2 AND2X2_4911 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8328) );
  AND2X2 AND2X2_4912 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8330) );
  AND2X2 AND2X2_4913 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8331) );
  AND2X2 AND2X2_4914 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8337) );
  AND2X2 AND2X2_4915 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8338) );
  AND2X2 AND2X2_4916 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8340) );
  AND2X2 AND2X2_4917 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8341) );
  AND2X2 AND2X2_4918 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8344) );
  AND2X2 AND2X2_4919 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8345) );
  AND2X2 AND2X2_492 ( .A(_abc_43815_n1535_1), .B(enable_i_bF_buf4), .Y(_abc_43815_n1536) );
  AND2X2 AND2X2_4920 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8347) );
  AND2X2 AND2X2_4921 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8348) );
  AND2X2 AND2X2_4922 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8352) );
  AND2X2 AND2X2_4923 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8353) );
  AND2X2 AND2X2_4924 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8355) );
  AND2X2 AND2X2_4925 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8356) );
  AND2X2 AND2X2_4926 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8359) );
  AND2X2 AND2X2_4927 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8360) );
  AND2X2 AND2X2_4928 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8362) );
  AND2X2 AND2X2_4929 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8363) );
  AND2X2 AND2X2_493 ( .A(_abc_43815_n1534_1), .B(_abc_43815_n1536), .Y(epc_q_3__FF_INPUT) );
  AND2X2 AND2X2_4930 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8368) );
  AND2X2 AND2X2_4931 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8369) );
  AND2X2 AND2X2_4932 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8371) );
  AND2X2 AND2X2_4933 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8372) );
  AND2X2 AND2X2_4934 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8375) );
  AND2X2 AND2X2_4935 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8376) );
  AND2X2 AND2X2_4936 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8377) );
  AND2X2 AND2X2_4937 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8381) );
  AND2X2 AND2X2_4938 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8382) );
  AND2X2 AND2X2_4939 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8384) );
  AND2X2 AND2X2_494 ( .A(_abc_43815_n1418_bF_buf2), .B(_abc_43815_n1539), .Y(_abc_43815_n1540) );
  AND2X2 AND2X2_4940 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8385) );
  AND2X2 AND2X2_4941 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8388) );
  AND2X2 AND2X2_4942 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8389) );
  AND2X2 AND2X2_4943 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8391) );
  AND2X2 AND2X2_4944 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8392) );
  AND2X2 AND2X2_4945 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8398) );
  AND2X2 AND2X2_4946 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8399) );
  AND2X2 AND2X2_4947 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8401) );
  AND2X2 AND2X2_4948 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8402) );
  AND2X2 AND2X2_4949 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8405) );
  AND2X2 AND2X2_495 ( .A(_abc_43815_n1541), .B(_abc_43815_n1538), .Y(_abc_43815_n1542) );
  AND2X2 AND2X2_4950 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8406) );
  AND2X2 AND2X2_4951 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8408) );
  AND2X2 AND2X2_4952 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8409) );
  AND2X2 AND2X2_4953 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8413) );
  AND2X2 AND2X2_4954 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8414) );
  AND2X2 AND2X2_4955 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8416) );
  AND2X2 AND2X2_4956 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8417) );
  AND2X2 AND2X2_4957 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8420) );
  AND2X2 AND2X2_4958 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8421) );
  AND2X2 AND2X2_4959 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8423) );
  AND2X2 AND2X2_496 ( .A(alu_op_r_2_), .B(pc_q_4_), .Y(_abc_43815_n1547_1) );
  AND2X2 AND2X2_4960 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8424) );
  AND2X2 AND2X2_4961 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8429) );
  AND2X2 AND2X2_4962 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8430) );
  AND2X2 AND2X2_4963 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8432) );
  AND2X2 AND2X2_4964 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8433) );
  AND2X2 AND2X2_4965 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8436) );
  AND2X2 AND2X2_4966 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8437) );
  AND2X2 AND2X2_4967 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8438) );
  AND2X2 AND2X2_4968 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8442) );
  AND2X2 AND2X2_4969 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8443) );
  AND2X2 AND2X2_497 ( .A(_abc_43815_n1548), .B(_abc_43815_n1546), .Y(_abc_43815_n1549) );
  AND2X2 AND2X2_4970 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8445) );
  AND2X2 AND2X2_4971 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8446) );
  AND2X2 AND2X2_4972 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8449) );
  AND2X2 AND2X2_4973 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8450) );
  AND2X2 AND2X2_4974 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8452) );
  AND2X2 AND2X2_4975 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8453) );
  AND2X2 AND2X2_4976 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8459) );
  AND2X2 AND2X2_4977 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8460) );
  AND2X2 AND2X2_4978 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8462) );
  AND2X2 AND2X2_4979 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8463) );
  AND2X2 AND2X2_498 ( .A(_abc_43815_n1545), .B(_abc_43815_n1549), .Y(_abc_43815_n1551) );
  AND2X2 AND2X2_4980 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8466) );
  AND2X2 AND2X2_4981 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8467) );
  AND2X2 AND2X2_4982 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8469) );
  AND2X2 AND2X2_4983 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8470) );
  AND2X2 AND2X2_4984 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8474) );
  AND2X2 AND2X2_4985 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8475) );
  AND2X2 AND2X2_4986 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8477) );
  AND2X2 AND2X2_4987 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8478) );
  AND2X2 AND2X2_4988 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8481) );
  AND2X2 AND2X2_4989 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8482) );
  AND2X2 AND2X2_499 ( .A(_abc_43815_n1552), .B(_abc_43815_n1550_1), .Y(_abc_43815_n1553) );
  AND2X2 AND2X2_4990 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8484) );
  AND2X2 AND2X2_4991 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8485) );
  AND2X2 AND2X2_4992 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8490) );
  AND2X2 AND2X2_4993 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8491) );
  AND2X2 AND2X2_4994 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8493) );
  AND2X2 AND2X2_4995 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8494) );
  AND2X2 AND2X2_4996 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8497) );
  AND2X2 AND2X2_4997 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8498) );
  AND2X2 AND2X2_4998 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8499) );
  AND2X2 AND2X2_4999 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8503) );
  AND2X2 AND2X2_5 ( .A(_abc_43815_n624_1), .B(_abc_43815_n626), .Y(_abc_43815_n627_1) );
  AND2X2 AND2X2_50 ( .A(_abc_43815_n689), .B(\mem_dat_i[24] ), .Y(_abc_43815_n701) );
  AND2X2 AND2X2_500 ( .A(_abc_43815_n1425_1_bF_buf0), .B(_abc_43815_n1553), .Y(_abc_43815_n1554) );
  AND2X2 AND2X2_5000 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8504) );
  AND2X2 AND2X2_5001 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8506) );
  AND2X2 AND2X2_5002 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8507) );
  AND2X2 AND2X2_5003 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8510) );
  AND2X2 AND2X2_5004 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8511) );
  AND2X2 AND2X2_5005 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8513) );
  AND2X2 AND2X2_5006 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8514) );
  AND2X2 AND2X2_5007 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8520) );
  AND2X2 AND2X2_5008 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8521) );
  AND2X2 AND2X2_5009 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8523) );
  AND2X2 AND2X2_501 ( .A(_abc_43815_n1065_1_bF_buf1), .B(epc_q_4_), .Y(_abc_43815_n1555) );
  AND2X2 AND2X2_5010 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8524) );
  AND2X2 AND2X2_5011 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8527) );
  AND2X2 AND2X2_5012 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8528) );
  AND2X2 AND2X2_5013 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8530) );
  AND2X2 AND2X2_5014 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8531) );
  AND2X2 AND2X2_5015 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8535) );
  AND2X2 AND2X2_5016 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8536) );
  AND2X2 AND2X2_5017 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8538) );
  AND2X2 AND2X2_5018 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8539) );
  AND2X2 AND2X2_5019 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8542) );
  AND2X2 AND2X2_502 ( .A(_abc_43815_n1557), .B(_abc_43815_n1544), .Y(_abc_43815_n1558) );
  AND2X2 AND2X2_5020 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8543) );
  AND2X2 AND2X2_5021 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8545) );
  AND2X2 AND2X2_5022 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8546) );
  AND2X2 AND2X2_5023 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8551) );
  AND2X2 AND2X2_5024 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8552) );
  AND2X2 AND2X2_5025 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8554) );
  AND2X2 AND2X2_5026 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8555) );
  AND2X2 AND2X2_5027 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8558) );
  AND2X2 AND2X2_5028 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8559) );
  AND2X2 AND2X2_5029 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8560) );
  AND2X2 AND2X2_503 ( .A(_abc_43815_n1524), .B(pc_q_4_), .Y(_abc_43815_n1561) );
  AND2X2 AND2X2_5030 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8564) );
  AND2X2 AND2X2_5031 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8565) );
  AND2X2 AND2X2_5032 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8567) );
  AND2X2 AND2X2_5033 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8568) );
  AND2X2 AND2X2_5034 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8571) );
  AND2X2 AND2X2_5035 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8572) );
  AND2X2 AND2X2_5036 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8574) );
  AND2X2 AND2X2_5037 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8575) );
  AND2X2 AND2X2_5038 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8581) );
  AND2X2 AND2X2_5039 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8582) );
  AND2X2 AND2X2_504 ( .A(_abc_43815_n1562), .B(_abc_43815_n1560), .Y(_abc_43815_n1563) );
  AND2X2 AND2X2_5040 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8584) );
  AND2X2 AND2X2_5041 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8585) );
  AND2X2 AND2X2_5042 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8588) );
  AND2X2 AND2X2_5043 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8589) );
  AND2X2 AND2X2_5044 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8591) );
  AND2X2 AND2X2_5045 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8592) );
  AND2X2 AND2X2_5046 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8596) );
  AND2X2 AND2X2_5047 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8597) );
  AND2X2 AND2X2_5048 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8599) );
  AND2X2 AND2X2_5049 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8600) );
  AND2X2 AND2X2_505 ( .A(_abc_43815_n1559), .B(_abc_43815_n1564), .Y(_abc_43815_n1565) );
  AND2X2 AND2X2_5050 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8603) );
  AND2X2 AND2X2_5051 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8604) );
  AND2X2 AND2X2_5052 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8606) );
  AND2X2 AND2X2_5053 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8607) );
  AND2X2 AND2X2_5054 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8612) );
  AND2X2 AND2X2_5055 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8613) );
  AND2X2 AND2X2_5056 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8615) );
  AND2X2 AND2X2_5057 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8616) );
  AND2X2 AND2X2_5058 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8619) );
  AND2X2 AND2X2_5059 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8620) );
  AND2X2 AND2X2_506 ( .A(_abc_43815_n1543), .B(_abc_43815_n1566_1), .Y(_abc_43815_n1567_1) );
  AND2X2 AND2X2_5060 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8621) );
  AND2X2 AND2X2_5061 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8625) );
  AND2X2 AND2X2_5062 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8626) );
  AND2X2 AND2X2_5063 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8628) );
  AND2X2 AND2X2_5064 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8629) );
  AND2X2 AND2X2_5065 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8632) );
  AND2X2 AND2X2_5066 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8633) );
  AND2X2 AND2X2_5067 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8635) );
  AND2X2 AND2X2_5068 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8636) );
  AND2X2 AND2X2_5069 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8642) );
  AND2X2 AND2X2_507 ( .A(_abc_43815_n1568), .B(_abc_43815_n1569), .Y(_abc_43815_n1570) );
  AND2X2 AND2X2_5070 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8643) );
  AND2X2 AND2X2_5071 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8645) );
  AND2X2 AND2X2_5072 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8646) );
  AND2X2 AND2X2_5073 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8649) );
  AND2X2 AND2X2_5074 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8650) );
  AND2X2 AND2X2_5075 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8652) );
  AND2X2 AND2X2_5076 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8653) );
  AND2X2 AND2X2_5077 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8657) );
  AND2X2 AND2X2_5078 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8658) );
  AND2X2 AND2X2_5079 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8660) );
  AND2X2 AND2X2_508 ( .A(_abc_43815_n1572), .B(enable_i_bF_buf3), .Y(_abc_43815_n1573) );
  AND2X2 AND2X2_5080 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8661) );
  AND2X2 AND2X2_5081 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8664) );
  AND2X2 AND2X2_5082 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8665) );
  AND2X2 AND2X2_5083 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8667) );
  AND2X2 AND2X2_5084 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8668) );
  AND2X2 AND2X2_5085 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8673) );
  AND2X2 AND2X2_5086 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8674) );
  AND2X2 AND2X2_5087 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8676) );
  AND2X2 AND2X2_5088 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8677) );
  AND2X2 AND2X2_5089 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8680) );
  AND2X2 AND2X2_509 ( .A(_abc_43815_n1571), .B(_abc_43815_n1573), .Y(epc_q_4__FF_INPUT) );
  AND2X2 AND2X2_5090 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8681) );
  AND2X2 AND2X2_5091 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8682) );
  AND2X2 AND2X2_5092 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8686) );
  AND2X2 AND2X2_5093 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8687) );
  AND2X2 AND2X2_5094 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8689) );
  AND2X2 AND2X2_5095 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8690) );
  AND2X2 AND2X2_5096 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8693) );
  AND2X2 AND2X2_5097 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8694) );
  AND2X2 AND2X2_5098 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8696) );
  AND2X2 AND2X2_5099 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8697) );
  AND2X2 AND2X2_51 ( .A(_abc_43815_n696), .B(\mem_dat_i[8] ), .Y(_abc_43815_n702) );
  AND2X2 AND2X2_510 ( .A(_abc_43815_n1418_bF_buf0), .B(_abc_43815_n1576), .Y(_abc_43815_n1577) );
  AND2X2 AND2X2_5100 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8703) );
  AND2X2 AND2X2_5101 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8704) );
  AND2X2 AND2X2_5102 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8706) );
  AND2X2 AND2X2_5103 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8707) );
  AND2X2 AND2X2_5104 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8710) );
  AND2X2 AND2X2_5105 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8711) );
  AND2X2 AND2X2_5106 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8713) );
  AND2X2 AND2X2_5107 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8714) );
  AND2X2 AND2X2_5108 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8718) );
  AND2X2 AND2X2_5109 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8719) );
  AND2X2 AND2X2_511 ( .A(_abc_43815_n1578), .B(_abc_43815_n1575), .Y(_abc_43815_n1579) );
  AND2X2 AND2X2_5110 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8721) );
  AND2X2 AND2X2_5111 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8722) );
  AND2X2 AND2X2_5112 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8725) );
  AND2X2 AND2X2_5113 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8726) );
  AND2X2 AND2X2_5114 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8728) );
  AND2X2 AND2X2_5115 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8729) );
  AND2X2 AND2X2_5116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8734) );
  AND2X2 AND2X2_5117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8735) );
  AND2X2 AND2X2_5118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8737) );
  AND2X2 AND2X2_5119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8738) );
  AND2X2 AND2X2_512 ( .A(alu_op_r_3_), .B(pc_q_5_), .Y(_abc_43815_n1582) );
  AND2X2 AND2X2_5120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8741) );
  AND2X2 AND2X2_5121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8742) );
  AND2X2 AND2X2_5122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8743) );
  AND2X2 AND2X2_5123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8747) );
  AND2X2 AND2X2_5124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8748) );
  AND2X2 AND2X2_5125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8750) );
  AND2X2 AND2X2_5126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8751) );
  AND2X2 AND2X2_5127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8754) );
  AND2X2 AND2X2_5128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8755) );
  AND2X2 AND2X2_5129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8757) );
  AND2X2 AND2X2_513 ( .A(_abc_43815_n1583_1), .B(_abc_43815_n1581), .Y(_abc_43815_n1584) );
  AND2X2 AND2X2_5130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8758) );
  AND2X2 AND2X2_5131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8764) );
  AND2X2 AND2X2_5132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8765) );
  AND2X2 AND2X2_5133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8767) );
  AND2X2 AND2X2_5134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8768) );
  AND2X2 AND2X2_5135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8771) );
  AND2X2 AND2X2_5136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8772) );
  AND2X2 AND2X2_5137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8774) );
  AND2X2 AND2X2_5138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8775) );
  AND2X2 AND2X2_5139 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8779) );
  AND2X2 AND2X2_514 ( .A(_abc_43815_n1584), .B(_abc_43815_n1547_1), .Y(_abc_43815_n1585) );
  AND2X2 AND2X2_5140 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8780) );
  AND2X2 AND2X2_5141 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8782) );
  AND2X2 AND2X2_5142 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8783) );
  AND2X2 AND2X2_5143 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8786) );
  AND2X2 AND2X2_5144 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8787) );
  AND2X2 AND2X2_5145 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8789) );
  AND2X2 AND2X2_5146 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8790) );
  AND2X2 AND2X2_5147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8795) );
  AND2X2 AND2X2_5148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8796) );
  AND2X2 AND2X2_5149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8798) );
  AND2X2 AND2X2_515 ( .A(_abc_43815_n1425_1_bF_buf4), .B(_abc_43815_n1586_1), .Y(_abc_43815_n1587) );
  AND2X2 AND2X2_5150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8799) );
  AND2X2 AND2X2_5151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8802) );
  AND2X2 AND2X2_5152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8803) );
  AND2X2 AND2X2_5153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8804) );
  AND2X2 AND2X2_5154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8808) );
  AND2X2 AND2X2_5155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8809) );
  AND2X2 AND2X2_5156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8811) );
  AND2X2 AND2X2_5157 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8812) );
  AND2X2 AND2X2_5158 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8815) );
  AND2X2 AND2X2_5159 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8816) );
  AND2X2 AND2X2_516 ( .A(_abc_43815_n1551), .B(_abc_43815_n1584), .Y(_abc_43815_n1590) );
  AND2X2 AND2X2_5160 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8818) );
  AND2X2 AND2X2_5161 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8819) );
  AND2X2 AND2X2_5162 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8825) );
  AND2X2 AND2X2_5163 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8826) );
  AND2X2 AND2X2_5164 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8828) );
  AND2X2 AND2X2_5165 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8829) );
  AND2X2 AND2X2_5166 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8832) );
  AND2X2 AND2X2_5167 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8833) );
  AND2X2 AND2X2_5168 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8835) );
  AND2X2 AND2X2_5169 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8836) );
  AND2X2 AND2X2_517 ( .A(_abc_43815_n1591), .B(_abc_43815_n1589), .Y(_abc_43815_n1592) );
  AND2X2 AND2X2_5170 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8840) );
  AND2X2 AND2X2_5171 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8841) );
  AND2X2 AND2X2_5172 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8843) );
  AND2X2 AND2X2_5173 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8844) );
  AND2X2 AND2X2_5174 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8847) );
  AND2X2 AND2X2_5175 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8848) );
  AND2X2 AND2X2_5176 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8850) );
  AND2X2 AND2X2_5177 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8851) );
  AND2X2 AND2X2_5178 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8856) );
  AND2X2 AND2X2_5179 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8857) );
  AND2X2 AND2X2_518 ( .A(_abc_43815_n1587), .B(_abc_43815_n1592), .Y(_abc_43815_n1593) );
  AND2X2 AND2X2_5180 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8859) );
  AND2X2 AND2X2_5181 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8860) );
  AND2X2 AND2X2_5182 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8863) );
  AND2X2 AND2X2_5183 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8864) );
  AND2X2 AND2X2_5184 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8865) );
  AND2X2 AND2X2_5185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8869) );
  AND2X2 AND2X2_5186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8870) );
  AND2X2 AND2X2_5187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8872) );
  AND2X2 AND2X2_5188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8873) );
  AND2X2 AND2X2_5189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8876) );
  AND2X2 AND2X2_519 ( .A(_abc_43815_n1065_1_bF_buf0), .B(epc_q_5_), .Y(_abc_43815_n1594) );
  AND2X2 AND2X2_5190 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8877) );
  AND2X2 AND2X2_5191 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8879) );
  AND2X2 AND2X2_5192 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8880) );
  AND2X2 AND2X2_5193 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8886) );
  AND2X2 AND2X2_5194 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8887) );
  AND2X2 AND2X2_5195 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8889) );
  AND2X2 AND2X2_5196 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8890) );
  AND2X2 AND2X2_5197 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8893) );
  AND2X2 AND2X2_5198 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8894) );
  AND2X2 AND2X2_5199 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8896) );
  AND2X2 AND2X2_52 ( .A(_abc_43815_n688), .B(mem_offset_q_0_), .Y(_abc_43815_n704) );
  AND2X2 AND2X2_520 ( .A(_abc_43815_n1596), .B(_abc_43815_n1597), .Y(_abc_43815_n1598) );
  AND2X2 AND2X2_5200 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8897) );
  AND2X2 AND2X2_5201 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8901) );
  AND2X2 AND2X2_5202 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8902) );
  AND2X2 AND2X2_5203 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8904) );
  AND2X2 AND2X2_5204 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8905) );
  AND2X2 AND2X2_5205 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8908) );
  AND2X2 AND2X2_5206 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8909) );
  AND2X2 AND2X2_5207 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8911) );
  AND2X2 AND2X2_5208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8912) );
  AND2X2 AND2X2_5209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8917) );
  AND2X2 AND2X2_521 ( .A(_abc_43815_n1561), .B(pc_q_5_), .Y(_abc_43815_n1601) );
  AND2X2 AND2X2_5210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8918) );
  AND2X2 AND2X2_5211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8920) );
  AND2X2 AND2X2_5212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8921) );
  AND2X2 AND2X2_5213 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8924) );
  AND2X2 AND2X2_5214 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8925) );
  AND2X2 AND2X2_5215 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8926) );
  AND2X2 AND2X2_5216 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8930) );
  AND2X2 AND2X2_5217 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8931) );
  AND2X2 AND2X2_5218 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8933) );
  AND2X2 AND2X2_5219 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8934) );
  AND2X2 AND2X2_522 ( .A(_abc_43815_n1602_1), .B(_abc_43815_n1600), .Y(_abc_43815_n1603_1) );
  AND2X2 AND2X2_5220 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8937) );
  AND2X2 AND2X2_5221 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8938) );
  AND2X2 AND2X2_5222 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8940) );
  AND2X2 AND2X2_5223 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8941) );
  AND2X2 AND2X2_5224 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8947) );
  AND2X2 AND2X2_5225 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8948) );
  AND2X2 AND2X2_5226 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8950) );
  AND2X2 AND2X2_5227 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8951) );
  AND2X2 AND2X2_5228 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8954) );
  AND2X2 AND2X2_5229 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8955) );
  AND2X2 AND2X2_523 ( .A(_abc_43815_n1599), .B(_abc_43815_n1604), .Y(_abc_43815_n1605) );
  AND2X2 AND2X2_5230 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8957) );
  AND2X2 AND2X2_5231 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8958) );
  AND2X2 AND2X2_5232 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8962) );
  AND2X2 AND2X2_5233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8963) );
  AND2X2 AND2X2_5234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8965) );
  AND2X2 AND2X2_5235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8966) );
  AND2X2 AND2X2_5236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8969) );
  AND2X2 AND2X2_5237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8970) );
  AND2X2 AND2X2_5238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8972) );
  AND2X2 AND2X2_5239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8973) );
  AND2X2 AND2X2_524 ( .A(_abc_43815_n1580), .B(_abc_43815_n1606), .Y(_abc_43815_n1607) );
  AND2X2 AND2X2_5240 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8978) );
  AND2X2 AND2X2_5241 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8979) );
  AND2X2 AND2X2_5242 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8981) );
  AND2X2 AND2X2_5243 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8982) );
  AND2X2 AND2X2_5244 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8985) );
  AND2X2 AND2X2_5245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8986) );
  AND2X2 AND2X2_5246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8987) );
  AND2X2 AND2X2_5247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8991) );
  AND2X2 AND2X2_5248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8992) );
  AND2X2 AND2X2_5249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8994) );
  AND2X2 AND2X2_525 ( .A(_abc_43815_n1608), .B(_abc_43815_n1609), .Y(_abc_43815_n1610) );
  AND2X2 AND2X2_5250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8995) );
  AND2X2 AND2X2_5251 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8998) );
  AND2X2 AND2X2_5252 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n8999) );
  AND2X2 AND2X2_5253 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9001) );
  AND2X2 AND2X2_5254 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9002) );
  AND2X2 AND2X2_5255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9008) );
  AND2X2 AND2X2_5256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9009) );
  AND2X2 AND2X2_5257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9011) );
  AND2X2 AND2X2_5258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9012) );
  AND2X2 AND2X2_5259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9015) );
  AND2X2 AND2X2_526 ( .A(_abc_43815_n1612), .B(enable_i_bF_buf2), .Y(_abc_43815_n1613) );
  AND2X2 AND2X2_5260 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9016) );
  AND2X2 AND2X2_5261 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9018) );
  AND2X2 AND2X2_5262 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9019) );
  AND2X2 AND2X2_5263 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9023) );
  AND2X2 AND2X2_5264 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9024) );
  AND2X2 AND2X2_5265 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9026) );
  AND2X2 AND2X2_5266 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9027) );
  AND2X2 AND2X2_5267 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9030) );
  AND2X2 AND2X2_5268 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9031) );
  AND2X2 AND2X2_5269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9033) );
  AND2X2 AND2X2_527 ( .A(_abc_43815_n1611), .B(_abc_43815_n1613), .Y(epc_q_5__FF_INPUT) );
  AND2X2 AND2X2_5270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9034) );
  AND2X2 AND2X2_5271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9039) );
  AND2X2 AND2X2_5272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9040) );
  AND2X2 AND2X2_5273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9042) );
  AND2X2 AND2X2_5274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9043) );
  AND2X2 AND2X2_5275 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9046) );
  AND2X2 AND2X2_5276 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9047) );
  AND2X2 AND2X2_5277 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9048) );
  AND2X2 AND2X2_5278 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9052) );
  AND2X2 AND2X2_5279 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9053) );
  AND2X2 AND2X2_528 ( .A(int32_r_4_), .B(pc_q_6_), .Y(_abc_43815_n1618_1) );
  AND2X2 AND2X2_5280 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9055) );
  AND2X2 AND2X2_5281 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9056) );
  AND2X2 AND2X2_5282 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9059) );
  AND2X2 AND2X2_5283 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9060) );
  AND2X2 AND2X2_5284 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9062) );
  AND2X2 AND2X2_5285 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9063) );
  AND2X2 AND2X2_5286 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9069) );
  AND2X2 AND2X2_5287 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9070) );
  AND2X2 AND2X2_5288 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9072) );
  AND2X2 AND2X2_5289 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9073) );
  AND2X2 AND2X2_529 ( .A(_abc_43815_n1619), .B(_abc_43815_n1617), .Y(_abc_43815_n1620) );
  AND2X2 AND2X2_5290 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9076) );
  AND2X2 AND2X2_5291 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9077) );
  AND2X2 AND2X2_5292 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9079) );
  AND2X2 AND2X2_5293 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9080) );
  AND2X2 AND2X2_5294 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9084) );
  AND2X2 AND2X2_5295 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9085) );
  AND2X2 AND2X2_5296 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9087) );
  AND2X2 AND2X2_5297 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9088) );
  AND2X2 AND2X2_5298 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9091) );
  AND2X2 AND2X2_5299 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9092) );
  AND2X2 AND2X2_53 ( .A(_abc_43815_n704), .B(\mem_dat_i[16] ), .Y(_abc_43815_n705) );
  AND2X2 AND2X2_530 ( .A(_abc_43815_n1616), .B(_abc_43815_n1620), .Y(_abc_43815_n1622) );
  AND2X2 AND2X2_5300 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9094) );
  AND2X2 AND2X2_5301 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9095) );
  AND2X2 AND2X2_5302 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9100) );
  AND2X2 AND2X2_5303 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9101) );
  AND2X2 AND2X2_5304 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9103) );
  AND2X2 AND2X2_5305 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9104) );
  AND2X2 AND2X2_5306 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9107) );
  AND2X2 AND2X2_5307 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9108) );
  AND2X2 AND2X2_5308 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9109) );
  AND2X2 AND2X2_5309 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9113) );
  AND2X2 AND2X2_531 ( .A(_abc_43815_n1623), .B(_abc_43815_n1425_1_bF_buf3), .Y(_abc_43815_n1624) );
  AND2X2 AND2X2_5310 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9114) );
  AND2X2 AND2X2_5311 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9116) );
  AND2X2 AND2X2_5312 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9117) );
  AND2X2 AND2X2_5313 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9120) );
  AND2X2 AND2X2_5314 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9121) );
  AND2X2 AND2X2_5315 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9123) );
  AND2X2 AND2X2_5316 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9124) );
  AND2X2 AND2X2_5317 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9130) );
  AND2X2 AND2X2_5318 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9131) );
  AND2X2 AND2X2_5319 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9133) );
  AND2X2 AND2X2_532 ( .A(_abc_43815_n1624), .B(_abc_43815_n1621), .Y(_abc_43815_n1625) );
  AND2X2 AND2X2_5320 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9134) );
  AND2X2 AND2X2_5321 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9137) );
  AND2X2 AND2X2_5322 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9138) );
  AND2X2 AND2X2_5323 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9140) );
  AND2X2 AND2X2_5324 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9141) );
  AND2X2 AND2X2_5325 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9145) );
  AND2X2 AND2X2_5326 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9146) );
  AND2X2 AND2X2_5327 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9148) );
  AND2X2 AND2X2_5328 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9149) );
  AND2X2 AND2X2_5329 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9152) );
  AND2X2 AND2X2_533 ( .A(_abc_43815_n1065_1_bF_buf4), .B(epc_q_6_), .Y(_abc_43815_n1626) );
  AND2X2 AND2X2_5330 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9153) );
  AND2X2 AND2X2_5331 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9155) );
  AND2X2 AND2X2_5332 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9156) );
  AND2X2 AND2X2_5333 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9161) );
  AND2X2 AND2X2_5334 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9162) );
  AND2X2 AND2X2_5335 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9164) );
  AND2X2 AND2X2_5336 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9165) );
  AND2X2 AND2X2_5337 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9168) );
  AND2X2 AND2X2_5338 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9169) );
  AND2X2 AND2X2_5339 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9170) );
  AND2X2 AND2X2_534 ( .A(_abc_43815_n1628), .B(_abc_43815_n1629), .Y(_abc_43815_n1630) );
  AND2X2 AND2X2_5340 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9174) );
  AND2X2 AND2X2_5341 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9175) );
  AND2X2 AND2X2_5342 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9177) );
  AND2X2 AND2X2_5343 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9178) );
  AND2X2 AND2X2_5344 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9181) );
  AND2X2 AND2X2_5345 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9182) );
  AND2X2 AND2X2_5346 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9184) );
  AND2X2 AND2X2_5347 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9185) );
  AND2X2 AND2X2_5348 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9191) );
  AND2X2 AND2X2_5349 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9192) );
  AND2X2 AND2X2_535 ( .A(_abc_43815_n1601), .B(pc_q_6_), .Y(_abc_43815_n1633) );
  AND2X2 AND2X2_5350 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9194) );
  AND2X2 AND2X2_5351 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9195) );
  AND2X2 AND2X2_5352 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9198) );
  AND2X2 AND2X2_5353 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9199) );
  AND2X2 AND2X2_5354 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9201) );
  AND2X2 AND2X2_5355 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9202) );
  AND2X2 AND2X2_5356 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9206) );
  AND2X2 AND2X2_5357 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9207) );
  AND2X2 AND2X2_5358 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9209) );
  AND2X2 AND2X2_5359 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9210) );
  AND2X2 AND2X2_536 ( .A(_abc_43815_n1634_1), .B(_abc_43815_n1632), .Y(_abc_43815_n1635_1) );
  AND2X2 AND2X2_5360 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9213) );
  AND2X2 AND2X2_5361 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9214) );
  AND2X2 AND2X2_5362 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9216) );
  AND2X2 AND2X2_5363 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9217) );
  AND2X2 AND2X2_5364 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9222) );
  AND2X2 AND2X2_5365 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9223) );
  AND2X2 AND2X2_5366 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9225) );
  AND2X2 AND2X2_5367 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9226) );
  AND2X2 AND2X2_5368 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9229) );
  AND2X2 AND2X2_5369 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9230) );
  AND2X2 AND2X2_537 ( .A(_abc_43815_n1631), .B(_abc_43815_n1636), .Y(_abc_43815_n1637) );
  AND2X2 AND2X2_5370 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9231) );
  AND2X2 AND2X2_5371 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9235) );
  AND2X2 AND2X2_5372 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9236) );
  AND2X2 AND2X2_5373 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9238) );
  AND2X2 AND2X2_5374 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9239) );
  AND2X2 AND2X2_5375 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9242) );
  AND2X2 AND2X2_5376 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9243) );
  AND2X2 AND2X2_5377 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9245) );
  AND2X2 AND2X2_5378 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9246) );
  AND2X2 AND2X2_5379 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9252) );
  AND2X2 AND2X2_538 ( .A(_abc_43815_n1418_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_43815_n1639) );
  AND2X2 AND2X2_5380 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9253) );
  AND2X2 AND2X2_5381 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9255) );
  AND2X2 AND2X2_5382 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9256) );
  AND2X2 AND2X2_5383 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9259) );
  AND2X2 AND2X2_5384 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9260) );
  AND2X2 AND2X2_5385 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9262) );
  AND2X2 AND2X2_5386 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9263) );
  AND2X2 AND2X2_5387 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9267) );
  AND2X2 AND2X2_5388 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9268) );
  AND2X2 AND2X2_5389 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9270) );
  AND2X2 AND2X2_539 ( .A(_abc_43815_n1489_bF_buf3), .B(epc_q_6_), .Y(_abc_43815_n1640) );
  AND2X2 AND2X2_5390 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9271) );
  AND2X2 AND2X2_5391 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9274) );
  AND2X2 AND2X2_5392 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9275) );
  AND2X2 AND2X2_5393 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9277) );
  AND2X2 AND2X2_5394 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9278) );
  AND2X2 AND2X2_5395 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9283) );
  AND2X2 AND2X2_5396 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9284) );
  AND2X2 AND2X2_5397 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9286) );
  AND2X2 AND2X2_5398 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9287) );
  AND2X2 AND2X2_5399 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9290) );
  AND2X2 AND2X2_54 ( .A(mem_offset_q_0_), .B(mem_offset_q_1_), .Y(_abc_43815_n706_1) );
  AND2X2 AND2X2_540 ( .A(_abc_43815_n1638), .B(_abc_43815_n1642), .Y(_abc_43815_n1643) );
  AND2X2 AND2X2_5400 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9291) );
  AND2X2 AND2X2_5401 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9292) );
  AND2X2 AND2X2_5402 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9296) );
  AND2X2 AND2X2_5403 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9297) );
  AND2X2 AND2X2_5404 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9299) );
  AND2X2 AND2X2_5405 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9300) );
  AND2X2 AND2X2_5406 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9303) );
  AND2X2 AND2X2_5407 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9304) );
  AND2X2 AND2X2_5408 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9306) );
  AND2X2 AND2X2_5409 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9307) );
  AND2X2 AND2X2_541 ( .A(_abc_43815_n1644), .B(_abc_43815_n1645), .Y(_abc_43815_n1646) );
  AND2X2 AND2X2_5410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9313) );
  AND2X2 AND2X2_5411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9314) );
  AND2X2 AND2X2_5412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9316) );
  AND2X2 AND2X2_5413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9317) );
  AND2X2 AND2X2_5414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9320) );
  AND2X2 AND2X2_5415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9321) );
  AND2X2 AND2X2_5416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9323) );
  AND2X2 AND2X2_5417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9324) );
  AND2X2 AND2X2_5418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9328) );
  AND2X2 AND2X2_5419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9329) );
  AND2X2 AND2X2_542 ( .A(_abc_43815_n1648), .B(enable_i_bF_buf1), .Y(_abc_43815_n1649) );
  AND2X2 AND2X2_5420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9331) );
  AND2X2 AND2X2_5421 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9332) );
  AND2X2 AND2X2_5422 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9335) );
  AND2X2 AND2X2_5423 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9336) );
  AND2X2 AND2X2_5424 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9338) );
  AND2X2 AND2X2_5425 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9339) );
  AND2X2 AND2X2_5426 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9344) );
  AND2X2 AND2X2_5427 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9345) );
  AND2X2 AND2X2_5428 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9347) );
  AND2X2 AND2X2_5429 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9348) );
  AND2X2 AND2X2_543 ( .A(_abc_43815_n1647), .B(_abc_43815_n1649), .Y(epc_q_6__FF_INPUT) );
  AND2X2 AND2X2_5430 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9351) );
  AND2X2 AND2X2_5431 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9352) );
  AND2X2 AND2X2_5432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9353) );
  AND2X2 AND2X2_5433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9357) );
  AND2X2 AND2X2_5434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9358) );
  AND2X2 AND2X2_5435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9360) );
  AND2X2 AND2X2_5436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9361) );
  AND2X2 AND2X2_5437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9364) );
  AND2X2 AND2X2_5438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9365) );
  AND2X2 AND2X2_5439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9367) );
  AND2X2 AND2X2_544 ( .A(_abc_43815_n1418_bF_buf3), .B(_abc_43815_n1652), .Y(_abc_43815_n1653) );
  AND2X2 AND2X2_5440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9368) );
  AND2X2 AND2X2_5441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9374) );
  AND2X2 AND2X2_5442 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9375) );
  AND2X2 AND2X2_5443 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9377) );
  AND2X2 AND2X2_5444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9378) );
  AND2X2 AND2X2_5445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9381) );
  AND2X2 AND2X2_5446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9382) );
  AND2X2 AND2X2_5447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9384) );
  AND2X2 AND2X2_5448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9385) );
  AND2X2 AND2X2_5449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9389) );
  AND2X2 AND2X2_545 ( .A(_abc_43815_n1654), .B(_abc_43815_n1651), .Y(_abc_43815_n1655_1) );
  AND2X2 AND2X2_5450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9390) );
  AND2X2 AND2X2_5451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9392) );
  AND2X2 AND2X2_5452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9393) );
  AND2X2 AND2X2_5453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9396) );
  AND2X2 AND2X2_5454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9397) );
  AND2X2 AND2X2_5455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9399) );
  AND2X2 AND2X2_5456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9400) );
  AND2X2 AND2X2_5457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9405) );
  AND2X2 AND2X2_5458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9406) );
  AND2X2 AND2X2_5459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9408) );
  AND2X2 AND2X2_546 ( .A(_abc_43815_n1350_bF_buf4), .B(_abc_43815_n1655_1), .Y(_abc_43815_n1656) );
  AND2X2 AND2X2_5460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9409) );
  AND2X2 AND2X2_5461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9412) );
  AND2X2 AND2X2_5462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9413) );
  AND2X2 AND2X2_5463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9414) );
  AND2X2 AND2X2_5464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9418) );
  AND2X2 AND2X2_5465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9419) );
  AND2X2 AND2X2_5466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9421) );
  AND2X2 AND2X2_5467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9422) );
  AND2X2 AND2X2_5468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9425) );
  AND2X2 AND2X2_5469 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9426) );
  AND2X2 AND2X2_547 ( .A(int32_r_5_), .B(pc_q_7_), .Y(_abc_43815_n1658_1) );
  AND2X2 AND2X2_5470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9428) );
  AND2X2 AND2X2_5471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9429) );
  AND2X2 AND2X2_5472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9435) );
  AND2X2 AND2X2_5473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9436) );
  AND2X2 AND2X2_5474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9438) );
  AND2X2 AND2X2_5475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9439) );
  AND2X2 AND2X2_5476 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9442) );
  AND2X2 AND2X2_5477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9443) );
  AND2X2 AND2X2_5478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9445) );
  AND2X2 AND2X2_5479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9446) );
  AND2X2 AND2X2_548 ( .A(_abc_43815_n1659), .B(_abc_43815_n1657), .Y(_abc_43815_n1660) );
  AND2X2 AND2X2_5480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9450) );
  AND2X2 AND2X2_5481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9451) );
  AND2X2 AND2X2_5482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9453) );
  AND2X2 AND2X2_5483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9454) );
  AND2X2 AND2X2_5484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9457) );
  AND2X2 AND2X2_5485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9458) );
  AND2X2 AND2X2_5486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9460) );
  AND2X2 AND2X2_5487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9461) );
  AND2X2 AND2X2_5488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9466) );
  AND2X2 AND2X2_5489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9467) );
  AND2X2 AND2X2_549 ( .A(_abc_43815_n1620), .B(_abc_43815_n1660), .Y(_abc_43815_n1663) );
  AND2X2 AND2X2_5490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9469) );
  AND2X2 AND2X2_5491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9470) );
  AND2X2 AND2X2_5492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9473) );
  AND2X2 AND2X2_5493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9474) );
  AND2X2 AND2X2_5494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9475) );
  AND2X2 AND2X2_5495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9479) );
  AND2X2 AND2X2_5496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9480) );
  AND2X2 AND2X2_5497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9482) );
  AND2X2 AND2X2_5498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9483) );
  AND2X2 AND2X2_5499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9486) );
  AND2X2 AND2X2_55 ( .A(_abc_43815_n706_1), .B(\mem_dat_i[0] ), .Y(_abc_43815_n707_1) );
  AND2X2 AND2X2_550 ( .A(_abc_43815_n1616), .B(_abc_43815_n1663), .Y(_abc_43815_n1664) );
  AND2X2 AND2X2_5500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9487) );
  AND2X2 AND2X2_5501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9489) );
  AND2X2 AND2X2_5502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9490) );
  AND2X2 AND2X2_5503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9496) );
  AND2X2 AND2X2_5504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9497) );
  AND2X2 AND2X2_5505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9499) );
  AND2X2 AND2X2_5506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9500) );
  AND2X2 AND2X2_5507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9503) );
  AND2X2 AND2X2_5508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9504) );
  AND2X2 AND2X2_5509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9506) );
  AND2X2 AND2X2_551 ( .A(_abc_43815_n1660), .B(_abc_43815_n1618_1), .Y(_abc_43815_n1666) );
  AND2X2 AND2X2_5510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9507) );
  AND2X2 AND2X2_5511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9511) );
  AND2X2 AND2X2_5512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9512) );
  AND2X2 AND2X2_5513 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9514) );
  AND2X2 AND2X2_5514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9515) );
  AND2X2 AND2X2_5515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9518) );
  AND2X2 AND2X2_5516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9519) );
  AND2X2 AND2X2_5517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9521) );
  AND2X2 AND2X2_5518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9522) );
  AND2X2 AND2X2_5519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9527) );
  AND2X2 AND2X2_552 ( .A(_abc_43815_n1425_1_bF_buf2), .B(_abc_43815_n1667), .Y(_abc_43815_n1668) );
  AND2X2 AND2X2_5520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9528) );
  AND2X2 AND2X2_5521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9530) );
  AND2X2 AND2X2_5522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9531) );
  AND2X2 AND2X2_5523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9534) );
  AND2X2 AND2X2_5524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9535) );
  AND2X2 AND2X2_5525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9536) );
  AND2X2 AND2X2_5526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9540) );
  AND2X2 AND2X2_5527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9541) );
  AND2X2 AND2X2_5528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9543) );
  AND2X2 AND2X2_5529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9544) );
  AND2X2 AND2X2_553 ( .A(_abc_43815_n1665), .B(_abc_43815_n1668), .Y(_abc_43815_n1669) );
  AND2X2 AND2X2_5530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9547) );
  AND2X2 AND2X2_5531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9548) );
  AND2X2 AND2X2_5532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9550) );
  AND2X2 AND2X2_5533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n9551) );
  AND2X2 AND2X2_5534 ( .A(alu_b_i_25_), .B(alu_a_i_25_), .Y(alu__abc_41358_n110) );
  AND2X2 AND2X2_5535 ( .A(alu__abc_41358_n112_1), .B(alu__abc_41358_n113_1), .Y(alu__abc_41358_n114) );
  AND2X2 AND2X2_5536 ( .A(alu__abc_41358_n115), .B(alu__abc_41358_n111), .Y(alu__abc_41358_n116) );
  AND2X2 AND2X2_5537 ( .A(alu_b_i_24_), .B(alu_a_i_24_), .Y(alu__abc_41358_n118) );
  AND2X2 AND2X2_5538 ( .A(alu__abc_41358_n120_1), .B(alu__abc_41358_n121), .Y(alu__abc_41358_n122) );
  AND2X2 AND2X2_5539 ( .A(alu__abc_41358_n123), .B(alu__abc_41358_n119_1), .Y(alu__abc_41358_n124_1) );
  AND2X2 AND2X2_554 ( .A(_abc_43815_n1669), .B(_abc_43815_n1662), .Y(_abc_43815_n1670) );
  AND2X2 AND2X2_5540 ( .A(alu__abc_41358_n117), .B(alu__abc_41358_n125_1), .Y(alu__abc_41358_n126) );
  AND2X2 AND2X2_5541 ( .A(alu_b_i_26_), .B(alu_a_i_26_), .Y(alu__abc_41358_n127) );
  AND2X2 AND2X2_5542 ( .A(alu__abc_41358_n129), .B(alu__abc_41358_n130_1), .Y(alu__abc_41358_n131_1) );
  AND2X2 AND2X2_5543 ( .A(alu__abc_41358_n132), .B(alu__abc_41358_n128), .Y(alu__abc_41358_n133) );
  AND2X2 AND2X2_5544 ( .A(alu_b_i_27_), .B(alu_a_i_27_), .Y(alu__abc_41358_n135_1) );
  AND2X2 AND2X2_5545 ( .A(alu__abc_41358_n137), .B(alu__abc_41358_n138), .Y(alu__abc_41358_n139) );
  AND2X2 AND2X2_5546 ( .A(alu__abc_41358_n140), .B(alu__abc_41358_n136_1), .Y(alu__abc_41358_n141) );
  AND2X2 AND2X2_5547 ( .A(alu__abc_41358_n134), .B(alu__abc_41358_n142), .Y(alu__abc_41358_n143_1) );
  AND2X2 AND2X2_5548 ( .A(alu__abc_41358_n126), .B(alu__abc_41358_n143_1), .Y(alu__abc_41358_n144_1) );
  AND2X2 AND2X2_5549 ( .A(alu_b_i_28_), .B(alu_a_i_28_), .Y(alu__abc_41358_n145) );
  AND2X2 AND2X2_555 ( .A(_abc_43815_n1065_1_bF_buf3), .B(epc_q_7_), .Y(_abc_43815_n1671) );
  AND2X2 AND2X2_5550 ( .A(alu__abc_41358_n147), .B(alu__abc_41358_n148_1), .Y(alu__abc_41358_n149_1) );
  AND2X2 AND2X2_5551 ( .A(alu__abc_41358_n150), .B(alu__abc_41358_n146), .Y(alu__abc_41358_n151) );
  AND2X2 AND2X2_5552 ( .A(alu_b_i_29_), .B(alu_a_i_29_), .Y(alu__abc_41358_n153) );
  AND2X2 AND2X2_5553 ( .A(alu__abc_41358_n155_1), .B(alu__abc_41358_n156), .Y(alu__abc_41358_n157) );
  AND2X2 AND2X2_5554 ( .A(alu__abc_41358_n158), .B(alu__abc_41358_n154_1), .Y(alu__abc_41358_n159_1) );
  AND2X2 AND2X2_5555 ( .A(alu__abc_41358_n152), .B(alu__abc_41358_n160_1), .Y(alu__abc_41358_n161) );
  AND2X2 AND2X2_5556 ( .A(alu_b_i_30_), .B(alu_a_i_30_), .Y(alu__abc_41358_n162) );
  AND2X2 AND2X2_5557 ( .A(alu__abc_41358_n164), .B(alu__abc_41358_n165), .Y(alu__abc_41358_n166_1) );
  AND2X2 AND2X2_5558 ( .A(alu__abc_41358_n167_1), .B(alu__abc_41358_n163), .Y(alu__abc_41358_n168) );
  AND2X2 AND2X2_5559 ( .A(alu_b_i_31_), .B(alu_a_i_31_), .Y(alu__abc_41358_n170) );
  AND2X2 AND2X2_556 ( .A(_abc_43815_n1673), .B(_abc_43815_n1674_1), .Y(_abc_43815_n1675_1) );
  AND2X2 AND2X2_5560 ( .A(alu__abc_41358_n171_1), .B(alu__abc_41358_n172_1), .Y(alu__abc_41358_n173) );
  AND2X2 AND2X2_5561 ( .A(alu__abc_41358_n169), .B(alu__abc_41358_n174), .Y(alu__abc_41358_n175) );
  AND2X2 AND2X2_5562 ( .A(alu__abc_41358_n161), .B(alu__abc_41358_n175), .Y(alu__abc_41358_n176) );
  AND2X2 AND2X2_5563 ( .A(alu__abc_41358_n144_1), .B(alu__abc_41358_n176), .Y(alu__abc_41358_n177_1) );
  AND2X2 AND2X2_5564 ( .A(alu_b_i_22_), .B(alu_a_i_22_), .Y(alu__abc_41358_n178_1) );
  AND2X2 AND2X2_5565 ( .A(alu__abc_41358_n180), .B(alu__abc_41358_n181), .Y(alu__abc_41358_n182_1) );
  AND2X2 AND2X2_5566 ( .A(alu__abc_41358_n183_1), .B(alu__abc_41358_n179), .Y(alu__abc_41358_n184) );
  AND2X2 AND2X2_5567 ( .A(alu_b_i_23_), .B(alu_a_i_23_), .Y(alu__abc_41358_n186) );
  AND2X2 AND2X2_5568 ( .A(alu__abc_41358_n188), .B(alu__abc_41358_n189), .Y(alu__abc_41358_n190) );
  AND2X2 AND2X2_5569 ( .A(alu__abc_41358_n191_1), .B(alu__abc_41358_n187), .Y(alu__abc_41358_n192_1) );
  AND2X2 AND2X2_557 ( .A(_abc_43815_n1633), .B(pc_q_7_), .Y(_abc_43815_n1678) );
  AND2X2 AND2X2_5570 ( .A(alu__abc_41358_n185), .B(alu__abc_41358_n193), .Y(alu__abc_41358_n194_1) );
  AND2X2 AND2X2_5571 ( .A(alu_b_i_20_), .B(alu_a_i_20_), .Y(alu__abc_41358_n195) );
  AND2X2 AND2X2_5572 ( .A(alu__abc_41358_n197), .B(alu__abc_41358_n198_1), .Y(alu__abc_41358_n199) );
  AND2X2 AND2X2_5573 ( .A(alu__abc_41358_n200), .B(alu__abc_41358_n196_1), .Y(alu__abc_41358_n201) );
  AND2X2 AND2X2_5574 ( .A(alu_b_i_21_), .B(alu_a_i_21_), .Y(alu__abc_41358_n203_1) );
  AND2X2 AND2X2_5575 ( .A(alu__abc_41358_n205), .B(alu__abc_41358_n206_1), .Y(alu__abc_41358_n207) );
  AND2X2 AND2X2_5576 ( .A(alu__abc_41358_n208), .B(alu__abc_41358_n204), .Y(alu__abc_41358_n209) );
  AND2X2 AND2X2_5577 ( .A(alu__abc_41358_n202), .B(alu__abc_41358_n210), .Y(alu__abc_41358_n211) );
  AND2X2 AND2X2_5578 ( .A(alu__abc_41358_n194_1), .B(alu__abc_41358_n211), .Y(alu__abc_41358_n212) );
  AND2X2 AND2X2_5579 ( .A(alu_b_i_18_), .B(alu_a_i_18_), .Y(alu__abc_41358_n213) );
  AND2X2 AND2X2_558 ( .A(_abc_43815_n1679), .B(_abc_43815_n1677), .Y(_abc_43815_n1680) );
  AND2X2 AND2X2_5580 ( .A(alu__abc_41358_n215), .B(alu__abc_41358_n216), .Y(alu__abc_41358_n217) );
  AND2X2 AND2X2_5581 ( .A(alu__abc_41358_n218), .B(alu__abc_41358_n214), .Y(alu__abc_41358_n219) );
  AND2X2 AND2X2_5582 ( .A(alu_b_i_19_), .B(alu_a_i_19_), .Y(alu__abc_41358_n221) );
  AND2X2 AND2X2_5583 ( .A(alu__abc_41358_n223), .B(alu__abc_41358_n224), .Y(alu__abc_41358_n225) );
  AND2X2 AND2X2_5584 ( .A(alu__abc_41358_n226), .B(alu__abc_41358_n222), .Y(alu__abc_41358_n227) );
  AND2X2 AND2X2_5585 ( .A(alu__abc_41358_n220), .B(alu__abc_41358_n228), .Y(alu__abc_41358_n229) );
  AND2X2 AND2X2_5586 ( .A(alu_b_i_16_), .B(alu_a_i_16_), .Y(alu__abc_41358_n230) );
  AND2X2 AND2X2_5587 ( .A(alu__abc_41358_n232), .B(alu__abc_41358_n233), .Y(alu__abc_41358_n234) );
  AND2X2 AND2X2_5588 ( .A(alu__abc_41358_n235), .B(alu__abc_41358_n231), .Y(alu__abc_41358_n236) );
  AND2X2 AND2X2_5589 ( .A(alu_b_i_17_), .B(alu_a_i_17_), .Y(alu__abc_41358_n238) );
  AND2X2 AND2X2_559 ( .A(_abc_43815_n1676), .B(_abc_43815_n1681), .Y(_abc_43815_n1682) );
  AND2X2 AND2X2_5590 ( .A(alu__abc_41358_n240), .B(alu__abc_41358_n241), .Y(alu__abc_41358_n242) );
  AND2X2 AND2X2_5591 ( .A(alu__abc_41358_n243), .B(alu__abc_41358_n239), .Y(alu__abc_41358_n244) );
  AND2X2 AND2X2_5592 ( .A(alu__abc_41358_n237), .B(alu__abc_41358_n245), .Y(alu__abc_41358_n246) );
  AND2X2 AND2X2_5593 ( .A(alu__abc_41358_n229), .B(alu__abc_41358_n246), .Y(alu__abc_41358_n247) );
  AND2X2 AND2X2_5594 ( .A(alu__abc_41358_n212), .B(alu__abc_41358_n247), .Y(alu__abc_41358_n248) );
  AND2X2 AND2X2_5595 ( .A(alu__abc_41358_n248), .B(alu__abc_41358_n177_1), .Y(alu__abc_41358_n249) );
  AND2X2 AND2X2_5596 ( .A(alu_a_i_1_), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n250) );
  AND2X2 AND2X2_5597 ( .A(alu__abc_41358_n251), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n253) );
  AND2X2 AND2X2_5598 ( .A(alu__abc_41358_n255), .B(alu_b_i_0_bF_buf4), .Y(alu__abc_41358_n256) );
  AND2X2 AND2X2_5599 ( .A(alu__abc_41358_n254), .B(alu__abc_41358_n257), .Y(alu__abc_41358_n258) );
  AND2X2 AND2X2_56 ( .A(_abc_43815_n709), .B(_abc_43815_n685), .Y(_abc_43815_n710) );
  AND2X2 AND2X2_560 ( .A(_abc_43815_n1682), .B(_abc_43815_n1413_bF_buf2), .Y(_abc_43815_n1683) );
  AND2X2 AND2X2_5600 ( .A(alu__abc_41358_n259_bF_buf4), .B(alu_a_i_0_), .Y(alu__abc_41358_n260) );
  AND2X2 AND2X2_5601 ( .A(alu__abc_41358_n258), .B(alu__abc_41358_n261), .Y(alu__abc_41358_n262) );
  AND2X2 AND2X2_5602 ( .A(alu_b_i_6_), .B(alu_a_i_6_), .Y(alu__abc_41358_n263) );
  AND2X2 AND2X2_5603 ( .A(alu__abc_41358_n265), .B(alu__abc_41358_n266), .Y(alu__abc_41358_n267) );
  AND2X2 AND2X2_5604 ( .A(alu__abc_41358_n268), .B(alu__abc_41358_n264), .Y(alu__abc_41358_n269) );
  AND2X2 AND2X2_5605 ( .A(alu_b_i_7_), .B(alu_a_i_7_), .Y(alu__abc_41358_n271) );
  AND2X2 AND2X2_5606 ( .A(alu__abc_41358_n272), .B(alu__abc_41358_n273), .Y(alu__abc_41358_n274) );
  AND2X2 AND2X2_5607 ( .A(alu__abc_41358_n270), .B(alu__abc_41358_n275), .Y(alu__abc_41358_n276) );
  AND2X2 AND2X2_5608 ( .A(alu_b_i_4_bF_buf4), .B(alu_a_i_4_), .Y(alu__abc_41358_n277) );
  AND2X2 AND2X2_5609 ( .A(alu__abc_41358_n279_bF_buf5), .B(alu__abc_41358_n280), .Y(alu__abc_41358_n281) );
  AND2X2 AND2X2_561 ( .A(_abc_43815_n1684), .B(_abc_43815_n1351_bF_buf4), .Y(_abc_43815_n1685) );
  AND2X2 AND2X2_5610 ( .A(alu__abc_41358_n282), .B(alu__abc_41358_n278), .Y(alu__abc_41358_n283) );
  AND2X2 AND2X2_5611 ( .A(alu_b_i_5_), .B(alu_a_i_5_), .Y(alu__abc_41358_n285) );
  AND2X2 AND2X2_5612 ( .A(alu__abc_41358_n286), .B(alu__abc_41358_n287), .Y(alu__abc_41358_n288) );
  AND2X2 AND2X2_5613 ( .A(alu__abc_41358_n284), .B(alu__abc_41358_n289), .Y(alu__abc_41358_n290) );
  AND2X2 AND2X2_5614 ( .A(alu__abc_41358_n276), .B(alu__abc_41358_n290), .Y(alu__abc_41358_n291) );
  AND2X2 AND2X2_5615 ( .A(alu_a_i_3_), .B(alu_b_i_3_bF_buf6), .Y(alu__abc_41358_n292) );
  AND2X2 AND2X2_5616 ( .A(alu__abc_41358_n293), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n295) );
  AND2X2 AND2X2_5617 ( .A(alu_a_i_2_), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n297) );
  AND2X2 AND2X2_5618 ( .A(alu__abc_41358_n298), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n300) );
  AND2X2 AND2X2_5619 ( .A(alu__abc_41358_n296), .B(alu__abc_41358_n301), .Y(alu__abc_41358_n302) );
  AND2X2 AND2X2_562 ( .A(_abc_43815_n1461_bF_buf2), .B(_abc_43815_n1680), .Y(_abc_43815_n1686_1) );
  AND2X2 AND2X2_5620 ( .A(alu__abc_41358_n291), .B(alu__abc_41358_n302), .Y(alu__abc_41358_n303) );
  AND2X2 AND2X2_5621 ( .A(alu__abc_41358_n303), .B(alu__abc_41358_n262), .Y(alu__abc_41358_n304) );
  AND2X2 AND2X2_5622 ( .A(alu_b_i_12_), .B(alu_a_i_12_), .Y(alu__abc_41358_n305) );
  AND2X2 AND2X2_5623 ( .A(alu__abc_41358_n307), .B(alu__abc_41358_n308), .Y(alu__abc_41358_n309) );
  AND2X2 AND2X2_5624 ( .A(alu__abc_41358_n310), .B(alu__abc_41358_n306), .Y(alu__abc_41358_n311) );
  AND2X2 AND2X2_5625 ( .A(alu_b_i_13_), .B(alu_a_i_13_), .Y(alu__abc_41358_n313) );
  AND2X2 AND2X2_5626 ( .A(alu__abc_41358_n315), .B(alu__abc_41358_n316), .Y(alu__abc_41358_n317) );
  AND2X2 AND2X2_5627 ( .A(alu__abc_41358_n318), .B(alu__abc_41358_n314), .Y(alu__abc_41358_n319) );
  AND2X2 AND2X2_5628 ( .A(alu__abc_41358_n312), .B(alu__abc_41358_n320), .Y(alu__abc_41358_n321) );
  AND2X2 AND2X2_5629 ( .A(alu_b_i_14_), .B(alu_a_i_14_), .Y(alu__abc_41358_n322) );
  AND2X2 AND2X2_563 ( .A(_abc_43815_n1689_1), .B(enable_i_bF_buf0), .Y(_abc_43815_n1690) );
  AND2X2 AND2X2_5630 ( .A(alu__abc_41358_n324), .B(alu__abc_41358_n325), .Y(alu__abc_41358_n326) );
  AND2X2 AND2X2_5631 ( .A(alu__abc_41358_n327), .B(alu__abc_41358_n323), .Y(alu__abc_41358_n328) );
  AND2X2 AND2X2_5632 ( .A(alu_b_i_15_), .B(alu_a_i_15_), .Y(alu__abc_41358_n330) );
  AND2X2 AND2X2_5633 ( .A(alu__abc_41358_n332), .B(alu__abc_41358_n333), .Y(alu__abc_41358_n334) );
  AND2X2 AND2X2_5634 ( .A(alu__abc_41358_n335), .B(alu__abc_41358_n331), .Y(alu__abc_41358_n336) );
  AND2X2 AND2X2_5635 ( .A(alu__abc_41358_n329_1), .B(alu__abc_41358_n337), .Y(alu__abc_41358_n338) );
  AND2X2 AND2X2_5636 ( .A(alu__abc_41358_n321), .B(alu__abc_41358_n338), .Y(alu__abc_41358_n339) );
  AND2X2 AND2X2_5637 ( .A(alu_b_i_10_), .B(alu_a_i_10_), .Y(alu__abc_41358_n340) );
  AND2X2 AND2X2_5638 ( .A(alu__abc_41358_n342), .B(alu__abc_41358_n343), .Y(alu__abc_41358_n344) );
  AND2X2 AND2X2_5639 ( .A(alu__abc_41358_n345), .B(alu__abc_41358_n341), .Y(alu__abc_41358_n346) );
  AND2X2 AND2X2_564 ( .A(_abc_43815_n1688), .B(_abc_43815_n1690), .Y(epc_q_7__FF_INPUT) );
  AND2X2 AND2X2_5640 ( .A(alu_b_i_11_), .B(alu_a_i_11_), .Y(alu__abc_41358_n348) );
  AND2X2 AND2X2_5641 ( .A(alu__abc_41358_n350), .B(alu__abc_41358_n351), .Y(alu__abc_41358_n352) );
  AND2X2 AND2X2_5642 ( .A(alu__abc_41358_n353), .B(alu__abc_41358_n349), .Y(alu__abc_41358_n354) );
  AND2X2 AND2X2_5643 ( .A(alu__abc_41358_n347), .B(alu__abc_41358_n355), .Y(alu__abc_41358_n356) );
  AND2X2 AND2X2_5644 ( .A(alu_b_i_8_), .B(alu_a_i_8_), .Y(alu__abc_41358_n357) );
  AND2X2 AND2X2_5645 ( .A(alu__abc_41358_n359), .B(alu__abc_41358_n360), .Y(alu__abc_41358_n361) );
  AND2X2 AND2X2_5646 ( .A(alu__abc_41358_n362), .B(alu__abc_41358_n358), .Y(alu__abc_41358_n363) );
  AND2X2 AND2X2_5647 ( .A(alu_b_i_9_), .B(alu_a_i_9_), .Y(alu__abc_41358_n365) );
  AND2X2 AND2X2_5648 ( .A(alu__abc_41358_n367), .B(alu__abc_41358_n368), .Y(alu__abc_41358_n369) );
  AND2X2 AND2X2_5649 ( .A(alu__abc_41358_n370), .B(alu__abc_41358_n366), .Y(alu__abc_41358_n371) );
  AND2X2 AND2X2_565 ( .A(_abc_43815_n1678), .B(pc_q_8_), .Y(_abc_43815_n1694) );
  AND2X2 AND2X2_5650 ( .A(alu__abc_41358_n364), .B(alu__abc_41358_n372), .Y(alu__abc_41358_n373) );
  AND2X2 AND2X2_5651 ( .A(alu__abc_41358_n356), .B(alu__abc_41358_n373), .Y(alu__abc_41358_n374) );
  AND2X2 AND2X2_5652 ( .A(alu__abc_41358_n339), .B(alu__abc_41358_n374), .Y(alu__abc_41358_n375) );
  AND2X2 AND2X2_5653 ( .A(alu__abc_41358_n304), .B(alu__abc_41358_n375), .Y(alu__abc_41358_n376) );
  AND2X2 AND2X2_5654 ( .A(alu__abc_41358_n376), .B(alu__abc_41358_n249), .Y(alu_equal_o) );
  AND2X2 AND2X2_5655 ( .A(alu__abc_41358_n379), .B(alu_op_i_2_), .Y(alu__abc_41358_n380) );
  AND2X2 AND2X2_5656 ( .A(alu__abc_41358_n380), .B(alu__abc_41358_n378), .Y(alu_c_update_o) );
  AND2X2 AND2X2_5657 ( .A(alu__abc_41358_n382), .B(alu_op_i_3_), .Y(alu__abc_41358_n383) );
  AND2X2 AND2X2_5658 ( .A(alu__abc_41358_n384), .B(alu_op_i_1_), .Y(alu__abc_41358_n385) );
  AND2X2 AND2X2_5659 ( .A(alu__abc_41358_n383), .B(alu__abc_41358_n385), .Y(alu_flag_update_o) );
  AND2X2 AND2X2_566 ( .A(_abc_43815_n1695), .B(_abc_43815_n1693), .Y(_abc_43815_n1696) );
  AND2X2 AND2X2_5660 ( .A(alu__abc_41358_n171_1), .B(alu_a_i_31_), .Y(alu__abc_41358_n387) );
  AND2X2 AND2X2_5661 ( .A(alu__abc_41358_n137), .B(alu_a_i_27_), .Y(alu__abc_41358_n388) );
  AND2X2 AND2X2_5662 ( .A(alu__abc_41358_n129), .B(alu_a_i_26_), .Y(alu__abc_41358_n389) );
  AND2X2 AND2X2_5663 ( .A(alu__abc_41358_n142), .B(alu__abc_41358_n389), .Y(alu__abc_41358_n390) );
  AND2X2 AND2X2_5664 ( .A(alu__abc_41358_n113_1), .B(alu_b_i_25_), .Y(alu__abc_41358_n394) );
  AND2X2 AND2X2_5665 ( .A(alu__abc_41358_n112_1), .B(alu_a_i_25_), .Y(alu__abc_41358_n395) );
  AND2X2 AND2X2_5666 ( .A(alu__abc_41358_n120_1), .B(alu_a_i_24_), .Y(alu__abc_41358_n397) );
  AND2X2 AND2X2_5667 ( .A(alu__abc_41358_n396), .B(alu__abc_41358_n398), .Y(alu__abc_41358_n399) );
  AND2X2 AND2X2_5668 ( .A(alu__abc_41358_n401), .B(alu__abc_41358_n392), .Y(alu__abc_41358_n402) );
  AND2X2 AND2X2_5669 ( .A(alu__abc_41358_n272), .B(alu_a_i_7_), .Y(alu__abc_41358_n404) );
  AND2X2 AND2X2_567 ( .A(_abc_43815_n1692), .B(_abc_43815_n1697), .Y(_abc_43815_n1698) );
  AND2X2 AND2X2_5670 ( .A(alu__abc_41358_n273), .B(alu_b_i_7_), .Y(alu__abc_41358_n405) );
  AND2X2 AND2X2_5671 ( .A(alu__abc_41358_n265), .B(alu_a_i_6_), .Y(alu__abc_41358_n407) );
  AND2X2 AND2X2_5672 ( .A(alu__abc_41358_n286), .B(alu_a_i_5_), .Y(alu__abc_41358_n408) );
  AND2X2 AND2X2_5673 ( .A(alu__abc_41358_n287), .B(alu_b_i_5_), .Y(alu__abc_41358_n409) );
  AND2X2 AND2X2_5674 ( .A(alu__abc_41358_n279_bF_buf4), .B(alu_a_i_4_), .Y(alu__abc_41358_n411) );
  AND2X2 AND2X2_5675 ( .A(alu__abc_41358_n294_bF_buf6), .B(alu_a_i_3_), .Y(alu__abc_41358_n412) );
  AND2X2 AND2X2_5676 ( .A(alu__abc_41358_n293), .B(alu_b_i_3_bF_buf4), .Y(alu__abc_41358_n413) );
  AND2X2 AND2X2_5677 ( .A(alu__abc_41358_n299_bF_buf6), .B(alu_a_i_2_), .Y(alu__abc_41358_n415) );
  AND2X2 AND2X2_5678 ( .A(alu__abc_41358_n252_bF_buf5), .B(alu_a_i_1_), .Y(alu__abc_41358_n416) );
  AND2X2 AND2X2_5679 ( .A(alu__abc_41358_n417), .B(alu__abc_41358_n301), .Y(alu__abc_41358_n418) );
  AND2X2 AND2X2_568 ( .A(_abc_43815_n1065_1_bF_buf2), .B(epc_q_8_), .Y(_abc_43815_n1700) );
  AND2X2 AND2X2_5680 ( .A(alu__abc_41358_n419), .B(alu__abc_41358_n414), .Y(alu__abc_41358_n420) );
  AND2X2 AND2X2_5681 ( .A(alu__abc_41358_n421), .B(alu__abc_41358_n284), .Y(alu__abc_41358_n422) );
  AND2X2 AND2X2_5682 ( .A(alu__abc_41358_n423), .B(alu__abc_41358_n410), .Y(alu__abc_41358_n424) );
  AND2X2 AND2X2_5683 ( .A(alu__abc_41358_n425), .B(alu__abc_41358_n270), .Y(alu__abc_41358_n426) );
  AND2X2 AND2X2_5684 ( .A(alu__abc_41358_n427), .B(alu__abc_41358_n406), .Y(alu__abc_41358_n428) );
  AND2X2 AND2X2_5685 ( .A(alu__abc_41358_n429), .B(alu__abc_41358_n375), .Y(alu__abc_41358_n430) );
  AND2X2 AND2X2_5686 ( .A(alu__abc_41358_n367), .B(alu_a_i_9_), .Y(alu__abc_41358_n431) );
  AND2X2 AND2X2_5687 ( .A(alu__abc_41358_n359), .B(alu_a_i_8_), .Y(alu__abc_41358_n433) );
  AND2X2 AND2X2_5688 ( .A(alu__abc_41358_n368), .B(alu_b_i_9_), .Y(alu__abc_41358_n435) );
  AND2X2 AND2X2_5689 ( .A(alu__abc_41358_n436), .B(alu__abc_41358_n432), .Y(alu__abc_41358_n437) );
  AND2X2 AND2X2_569 ( .A(_abc_43815_n1667), .B(_abc_43815_n1659), .Y(_abc_43815_n1701) );
  AND2X2 AND2X2_5690 ( .A(alu__abc_41358_n438), .B(alu__abc_41358_n356), .Y(alu__abc_41358_n439) );
  AND2X2 AND2X2_5691 ( .A(alu__abc_41358_n350), .B(alu_a_i_11_), .Y(alu__abc_41358_n440) );
  AND2X2 AND2X2_5692 ( .A(alu__abc_41358_n342), .B(alu_a_i_10_), .Y(alu__abc_41358_n441) );
  AND2X2 AND2X2_5693 ( .A(alu__abc_41358_n355), .B(alu__abc_41358_n441), .Y(alu__abc_41358_n442) );
  AND2X2 AND2X2_5694 ( .A(alu__abc_41358_n444), .B(alu__abc_41358_n339), .Y(alu__abc_41358_n445) );
  AND2X2 AND2X2_5695 ( .A(alu__abc_41358_n315), .B(alu_a_i_13_), .Y(alu__abc_41358_n446) );
  AND2X2 AND2X2_5696 ( .A(alu__abc_41358_n307), .B(alu_a_i_12_), .Y(alu__abc_41358_n448) );
  AND2X2 AND2X2_5697 ( .A(alu__abc_41358_n316), .B(alu_b_i_13_), .Y(alu__abc_41358_n450) );
  AND2X2 AND2X2_5698 ( .A(alu__abc_41358_n451), .B(alu__abc_41358_n447), .Y(alu__abc_41358_n452) );
  AND2X2 AND2X2_5699 ( .A(alu__abc_41358_n453), .B(alu__abc_41358_n338), .Y(alu__abc_41358_n454) );
  AND2X2 AND2X2_57 ( .A(_abc_43815_n711), .B(state_q_1_bF_buf1), .Y(_abc_43815_n712) );
  AND2X2 AND2X2_570 ( .A(alu_op_r_4_), .B(pc_q_8_), .Y(_abc_43815_n1705_1) );
  AND2X2 AND2X2_5700 ( .A(alu__abc_41358_n332), .B(alu_a_i_15_), .Y(alu__abc_41358_n455) );
  AND2X2 AND2X2_5701 ( .A(alu__abc_41358_n324), .B(alu_a_i_14_), .Y(alu__abc_41358_n456) );
  AND2X2 AND2X2_5702 ( .A(alu__abc_41358_n337), .B(alu__abc_41358_n456), .Y(alu__abc_41358_n457) );
  AND2X2 AND2X2_5703 ( .A(alu__abc_41358_n461), .B(alu__abc_41358_n248), .Y(alu__abc_41358_n462) );
  AND2X2 AND2X2_5704 ( .A(alu__abc_41358_n240), .B(alu_a_i_17_), .Y(alu__abc_41358_n463) );
  AND2X2 AND2X2_5705 ( .A(alu__abc_41358_n232), .B(alu_a_i_16_), .Y(alu__abc_41358_n465) );
  AND2X2 AND2X2_5706 ( .A(alu__abc_41358_n241), .B(alu_b_i_17_), .Y(alu__abc_41358_n467) );
  AND2X2 AND2X2_5707 ( .A(alu__abc_41358_n468), .B(alu__abc_41358_n464), .Y(alu__abc_41358_n469) );
  AND2X2 AND2X2_5708 ( .A(alu__abc_41358_n470), .B(alu__abc_41358_n229), .Y(alu__abc_41358_n471) );
  AND2X2 AND2X2_5709 ( .A(alu__abc_41358_n223), .B(alu_a_i_19_), .Y(alu__abc_41358_n472) );
  AND2X2 AND2X2_571 ( .A(_abc_43815_n1706_1), .B(_abc_43815_n1704), .Y(_abc_43815_n1707) );
  AND2X2 AND2X2_5710 ( .A(alu__abc_41358_n215), .B(alu_a_i_18_), .Y(alu__abc_41358_n473) );
  AND2X2 AND2X2_5711 ( .A(alu__abc_41358_n228), .B(alu__abc_41358_n473), .Y(alu__abc_41358_n474) );
  AND2X2 AND2X2_5712 ( .A(alu__abc_41358_n476), .B(alu__abc_41358_n212), .Y(alu__abc_41358_n477) );
  AND2X2 AND2X2_5713 ( .A(alu__abc_41358_n205), .B(alu_a_i_21_), .Y(alu__abc_41358_n478) );
  AND2X2 AND2X2_5714 ( .A(alu__abc_41358_n197), .B(alu_a_i_20_), .Y(alu__abc_41358_n480) );
  AND2X2 AND2X2_5715 ( .A(alu__abc_41358_n206_1), .B(alu_b_i_21_), .Y(alu__abc_41358_n482) );
  AND2X2 AND2X2_5716 ( .A(alu__abc_41358_n483), .B(alu__abc_41358_n479), .Y(alu__abc_41358_n484) );
  AND2X2 AND2X2_5717 ( .A(alu__abc_41358_n485), .B(alu__abc_41358_n194_1), .Y(alu__abc_41358_n486) );
  AND2X2 AND2X2_5718 ( .A(alu__abc_41358_n188), .B(alu_a_i_23_), .Y(alu__abc_41358_n487) );
  AND2X2 AND2X2_5719 ( .A(alu__abc_41358_n180), .B(alu_a_i_22_), .Y(alu__abc_41358_n488) );
  AND2X2 AND2X2_572 ( .A(_abc_43815_n1703), .B(_abc_43815_n1707), .Y(_abc_43815_n1709) );
  AND2X2 AND2X2_5720 ( .A(alu__abc_41358_n193), .B(alu__abc_41358_n488), .Y(alu__abc_41358_n489) );
  AND2X2 AND2X2_5721 ( .A(alu__abc_41358_n493), .B(alu__abc_41358_n144_1), .Y(alu__abc_41358_n494) );
  AND2X2 AND2X2_5722 ( .A(alu__abc_41358_n495), .B(alu__abc_41358_n161), .Y(alu__abc_41358_n496) );
  AND2X2 AND2X2_5723 ( .A(alu__abc_41358_n156), .B(alu_b_i_29_), .Y(alu__abc_41358_n497) );
  AND2X2 AND2X2_5724 ( .A(alu__abc_41358_n155_1), .B(alu_a_i_29_), .Y(alu__abc_41358_n498) );
  AND2X2 AND2X2_5725 ( .A(alu__abc_41358_n147), .B(alu_a_i_28_), .Y(alu__abc_41358_n500) );
  AND2X2 AND2X2_5726 ( .A(alu__abc_41358_n499), .B(alu__abc_41358_n501), .Y(alu__abc_41358_n502) );
  AND2X2 AND2X2_5727 ( .A(alu__abc_41358_n505), .B(alu__abc_41358_n169), .Y(alu__abc_41358_n506) );
  AND2X2 AND2X2_5728 ( .A(alu__abc_41358_n164), .B(alu_a_i_30_), .Y(alu__abc_41358_n508) );
  AND2X2 AND2X2_5729 ( .A(alu__abc_41358_n507), .B(alu__abc_41358_n509), .Y(alu__abc_41358_n510) );
  AND2X2 AND2X2_573 ( .A(_abc_43815_n1710), .B(_abc_43815_n1425_1_bF_buf1), .Y(_abc_43815_n1711) );
  AND2X2 AND2X2_5730 ( .A(alu__abc_41358_n510), .B(alu__abc_41358_n174), .Y(alu__abc_41358_n511) );
  AND2X2 AND2X2_5731 ( .A(alu__abc_41358_n133), .B(alu__abc_41358_n141), .Y(alu__abc_41358_n513) );
  AND2X2 AND2X2_5732 ( .A(alu__abc_41358_n111), .B(alu__abc_41358_n119_1), .Y(alu__abc_41358_n514) );
  AND2X2 AND2X2_5733 ( .A(alu__abc_41358_n516), .B(alu__abc_41358_n513), .Y(alu__abc_41358_n517) );
  AND2X2 AND2X2_5734 ( .A(alu__abc_41358_n140), .B(alu__abc_41358_n127), .Y(alu__abc_41358_n518) );
  AND2X2 AND2X2_5735 ( .A(alu__abc_41358_n151), .B(alu__abc_41358_n159_1), .Y(alu__abc_41358_n521) );
  AND2X2 AND2X2_5736 ( .A(alu__abc_41358_n522), .B(alu__abc_41358_n168), .Y(alu__abc_41358_n523) );
  AND2X2 AND2X2_5737 ( .A(alu__abc_41358_n523), .B(alu__abc_41358_n521), .Y(alu__abc_41358_n524) );
  AND2X2 AND2X2_5738 ( .A(alu__abc_41358_n520), .B(alu__abc_41358_n524), .Y(alu__abc_41358_n525) );
  AND2X2 AND2X2_5739 ( .A(alu__abc_41358_n146), .B(alu__abc_41358_n154_1), .Y(alu__abc_41358_n526) );
  AND2X2 AND2X2_574 ( .A(_abc_43815_n1711), .B(_abc_43815_n1708), .Y(_abc_43815_n1712) );
  AND2X2 AND2X2_5740 ( .A(alu__abc_41358_n528), .B(alu__abc_41358_n523), .Y(alu__abc_41358_n529) );
  AND2X2 AND2X2_5741 ( .A(alu__abc_41358_n530), .B(alu__abc_41358_n162), .Y(alu__abc_41358_n531) );
  AND2X2 AND2X2_5742 ( .A(alu__abc_41358_n184), .B(alu__abc_41358_n192_1), .Y(alu__abc_41358_n535) );
  AND2X2 AND2X2_5743 ( .A(alu__abc_41358_n201), .B(alu__abc_41358_n209), .Y(alu__abc_41358_n536) );
  AND2X2 AND2X2_5744 ( .A(alu__abc_41358_n535), .B(alu__abc_41358_n536), .Y(alu__abc_41358_n537) );
  AND2X2 AND2X2_5745 ( .A(alu__abc_41358_n219), .B(alu__abc_41358_n227), .Y(alu__abc_41358_n538) );
  AND2X2 AND2X2_5746 ( .A(alu__abc_41358_n231), .B(alu__abc_41358_n239), .Y(alu__abc_41358_n539) );
  AND2X2 AND2X2_5747 ( .A(alu__abc_41358_n541), .B(alu__abc_41358_n538), .Y(alu__abc_41358_n542) );
  AND2X2 AND2X2_5748 ( .A(alu__abc_41358_n214), .B(alu__abc_41358_n222), .Y(alu__abc_41358_n543) );
  AND2X2 AND2X2_5749 ( .A(alu__abc_41358_n546), .B(alu__abc_41358_n537), .Y(alu__abc_41358_n547) );
  AND2X2 AND2X2_575 ( .A(_abc_43815_n1713), .B(_abc_43815_n1431_1_bF_buf1), .Y(_abc_43815_n1714) );
  AND2X2 AND2X2_5750 ( .A(alu__abc_41358_n196_1), .B(alu__abc_41358_n204), .Y(alu__abc_41358_n548) );
  AND2X2 AND2X2_5751 ( .A(alu__abc_41358_n550), .B(alu__abc_41358_n535), .Y(alu__abc_41358_n551) );
  AND2X2 AND2X2_5752 ( .A(alu__abc_41358_n191_1), .B(alu__abc_41358_n178_1), .Y(alu__abc_41358_n552) );
  AND2X2 AND2X2_5753 ( .A(alu__abc_41358_n335), .B(alu__abc_41358_n322), .Y(alu__abc_41358_n556) );
  AND2X2 AND2X2_5754 ( .A(alu__abc_41358_n318), .B(alu__abc_41358_n305), .Y(alu__abc_41358_n558) );
  AND2X2 AND2X2_5755 ( .A(alu__abc_41358_n328), .B(alu__abc_41358_n336), .Y(alu__abc_41358_n560) );
  AND2X2 AND2X2_5756 ( .A(alu__abc_41358_n559), .B(alu__abc_41358_n560), .Y(alu__abc_41358_n561) );
  AND2X2 AND2X2_5757 ( .A(alu__abc_41358_n346), .B(alu__abc_41358_n354), .Y(alu__abc_41358_n563) );
  AND2X2 AND2X2_5758 ( .A(alu__abc_41358_n358), .B(alu__abc_41358_n366), .Y(alu__abc_41358_n564) );
  AND2X2 AND2X2_5759 ( .A(alu__abc_41358_n566), .B(alu__abc_41358_n563), .Y(alu__abc_41358_n567) );
  AND2X2 AND2X2_576 ( .A(_abc_43815_n1428_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_43815_n1715) );
  AND2X2 AND2X2_5760 ( .A(alu__abc_41358_n353), .B(alu__abc_41358_n340), .Y(alu__abc_41358_n568) );
  AND2X2 AND2X2_5761 ( .A(alu__abc_41358_n311), .B(alu__abc_41358_n319), .Y(alu__abc_41358_n571) );
  AND2X2 AND2X2_5762 ( .A(alu__abc_41358_n571), .B(alu__abc_41358_n560), .Y(alu__abc_41358_n572) );
  AND2X2 AND2X2_5763 ( .A(alu__abc_41358_n570), .B(alu__abc_41358_n572), .Y(alu__abc_41358_n573) );
  AND2X2 AND2X2_5764 ( .A(alu__abc_41358_n575), .B(alu__abc_41358_n576), .Y(alu__abc_41358_n577) );
  AND2X2 AND2X2_5765 ( .A(alu_b_i_0_bF_buf2), .B(alu_a_i_0_), .Y(alu__abc_41358_n578) );
  AND2X2 AND2X2_5766 ( .A(alu__abc_41358_n577), .B(alu__abc_41358_n578), .Y(alu__abc_41358_n579) );
  AND2X2 AND2X2_5767 ( .A(alu__abc_41358_n580), .B(alu__abc_41358_n582), .Y(alu__abc_41358_n583) );
  AND2X2 AND2X2_5768 ( .A(alu__abc_41358_n584), .B(alu__abc_41358_n297), .Y(alu__abc_41358_n585) );
  AND2X2 AND2X2_5769 ( .A(alu__abc_41358_n588), .B(alu__abc_41358_n269), .Y(alu__abc_41358_n589) );
  AND2X2 AND2X2_577 ( .A(_abc_43815_n1717), .B(_abc_43815_n1699), .Y(_abc_43815_n1718) );
  AND2X2 AND2X2_5770 ( .A(alu__abc_41358_n590), .B(alu__abc_41358_n283), .Y(alu__abc_41358_n591) );
  AND2X2 AND2X2_5771 ( .A(alu__abc_41358_n589), .B(alu__abc_41358_n591), .Y(alu__abc_41358_n592) );
  AND2X2 AND2X2_5772 ( .A(alu__abc_41358_n587), .B(alu__abc_41358_n592), .Y(alu__abc_41358_n593) );
  AND2X2 AND2X2_5773 ( .A(alu__abc_41358_n595), .B(alu__abc_41358_n594), .Y(alu__abc_41358_n596) );
  AND2X2 AND2X2_5774 ( .A(alu__abc_41358_n589), .B(alu__abc_41358_n596), .Y(alu__abc_41358_n597) );
  AND2X2 AND2X2_5775 ( .A(alu__abc_41358_n598), .B(alu__abc_41358_n263), .Y(alu__abc_41358_n599) );
  AND2X2 AND2X2_5776 ( .A(alu__abc_41358_n363), .B(alu__abc_41358_n371), .Y(alu__abc_41358_n603) );
  AND2X2 AND2X2_5777 ( .A(alu__abc_41358_n563), .B(alu__abc_41358_n603), .Y(alu__abc_41358_n604) );
  AND2X2 AND2X2_5778 ( .A(alu__abc_41358_n604), .B(alu__abc_41358_n572), .Y(alu__abc_41358_n605) );
  AND2X2 AND2X2_5779 ( .A(alu__abc_41358_n602), .B(alu__abc_41358_n605), .Y(alu__abc_41358_n606) );
  AND2X2 AND2X2_578 ( .A(_abc_43815_n1489_bF_buf2), .B(epc_q_8_), .Y(_abc_43815_n1720) );
  AND2X2 AND2X2_5780 ( .A(alu__abc_41358_n236), .B(alu__abc_41358_n244), .Y(alu__abc_41358_n608) );
  AND2X2 AND2X2_5781 ( .A(alu__abc_41358_n607), .B(alu__abc_41358_n608), .Y(alu__abc_41358_n609) );
  AND2X2 AND2X2_5782 ( .A(alu__abc_41358_n537), .B(alu__abc_41358_n538), .Y(alu__abc_41358_n610) );
  AND2X2 AND2X2_5783 ( .A(alu__abc_41358_n609), .B(alu__abc_41358_n610), .Y(alu__abc_41358_n611) );
  AND2X2 AND2X2_5784 ( .A(alu__abc_41358_n612), .B(alu__abc_41358_n124_1), .Y(alu__abc_41358_n613) );
  AND2X2 AND2X2_5785 ( .A(alu__abc_41358_n613), .B(alu__abc_41358_n116), .Y(alu__abc_41358_n614) );
  AND2X2 AND2X2_5786 ( .A(alu__abc_41358_n614), .B(alu__abc_41358_n513), .Y(alu__abc_41358_n615) );
  AND2X2 AND2X2_5787 ( .A(alu__abc_41358_n615), .B(alu__abc_41358_n524), .Y(alu__abc_41358_n616) );
  AND2X2 AND2X2_5788 ( .A(alu__abc_41358_n618), .B(alu__abc_41358_n521), .Y(alu__abc_41358_n619) );
  AND2X2 AND2X2_5789 ( .A(alu__abc_41358_n620_1), .B(alu__abc_41358_n168), .Y(alu__abc_41358_n621) );
  AND2X2 AND2X2_579 ( .A(_abc_43815_n1418_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_43815_n1721) );
  AND2X2 AND2X2_5790 ( .A(alu__abc_41358_n622), .B(alu__abc_41358_n163), .Y(alu__abc_41358_n623) );
  AND2X2 AND2X2_5791 ( .A(alu__abc_41358_n625), .B(alu__abc_41358_n626), .Y(alu__abc_41358_n627) );
  AND2X2 AND2X2_5792 ( .A(alu__abc_41358_n622), .B(alu__abc_41358_n628), .Y(alu__abc_41358_n629) );
  AND2X2 AND2X2_5793 ( .A(alu__abc_41358_n618), .B(alu__abc_41358_n151), .Y(alu__abc_41358_n630) );
  AND2X2 AND2X2_5794 ( .A(alu__abc_41358_n631), .B(alu__abc_41358_n146), .Y(alu__abc_41358_n632) );
  AND2X2 AND2X2_5795 ( .A(alu__abc_41358_n634), .B(alu__abc_41358_n635), .Y(alu__abc_41358_n636) );
  AND2X2 AND2X2_5796 ( .A(alu__abc_41358_n636), .B(alu__abc_41358_n629), .Y(alu__abc_41358_n637) );
  AND2X2 AND2X2_5797 ( .A(alu__abc_41358_n638), .B(alu__abc_41358_n538), .Y(alu__abc_41358_n639) );
  AND2X2 AND2X2_5798 ( .A(alu__abc_41358_n640), .B(alu__abc_41358_n536), .Y(alu__abc_41358_n641) );
  AND2X2 AND2X2_5799 ( .A(alu__abc_41358_n642), .B(alu__abc_41358_n184), .Y(alu__abc_41358_n643) );
  AND2X2 AND2X2_58 ( .A(_abc_43815_n682), .B(alu_p_o_1_), .Y(_abc_43815_n714) );
  AND2X2 AND2X2_580 ( .A(_abc_43815_n1723), .B(_abc_43815_n1351_bF_buf3), .Y(_abc_43815_n1724) );
  AND2X2 AND2X2_5800 ( .A(alu__abc_41358_n644), .B(alu__abc_41358_n179), .Y(alu__abc_41358_n645) );
  AND2X2 AND2X2_5801 ( .A(alu__abc_41358_n646), .B(alu__abc_41358_n193), .Y(alu__abc_41358_n647) );
  AND2X2 AND2X2_5802 ( .A(alu__abc_41358_n645), .B(alu__abc_41358_n192_1), .Y(alu__abc_41358_n648) );
  AND2X2 AND2X2_5803 ( .A(alu__abc_41358_n650), .B(alu__abc_41358_n133), .Y(alu__abc_41358_n651) );
  AND2X2 AND2X2_5804 ( .A(alu__abc_41358_n652), .B(alu__abc_41358_n128), .Y(alu__abc_41358_n653) );
  AND2X2 AND2X2_5805 ( .A(alu__abc_41358_n655), .B(alu__abc_41358_n656), .Y(alu__abc_41358_n657) );
  AND2X2 AND2X2_5806 ( .A(alu__abc_41358_n652), .B(alu__abc_41358_n658), .Y(alu__abc_41358_n659) );
  AND2X2 AND2X2_5807 ( .A(alu__abc_41358_n660), .B(alu__abc_41358_n119_1), .Y(alu__abc_41358_n661) );
  AND2X2 AND2X2_5808 ( .A(alu__abc_41358_n662), .B(alu__abc_41358_n117), .Y(alu__abc_41358_n663) );
  AND2X2 AND2X2_5809 ( .A(alu__abc_41358_n661), .B(alu__abc_41358_n116), .Y(alu__abc_41358_n664) );
  AND2X2 AND2X2_581 ( .A(_abc_43815_n1719_1), .B(_abc_43815_n1724), .Y(_abc_43815_n1725) );
  AND2X2 AND2X2_5810 ( .A(alu__abc_41358_n660), .B(alu__abc_41358_n666), .Y(alu__abc_41358_n667) );
  AND2X2 AND2X2_5811 ( .A(alu__abc_41358_n665), .B(alu__abc_41358_n667), .Y(alu__abc_41358_n668) );
  AND2X2 AND2X2_5812 ( .A(alu__abc_41358_n668), .B(alu__abc_41358_n659), .Y(alu__abc_41358_n669) );
  AND2X2 AND2X2_5813 ( .A(alu__abc_41358_n657), .B(alu__abc_41358_n669), .Y(alu__abc_41358_n670) );
  AND2X2 AND2X2_5814 ( .A(alu__abc_41358_n644), .B(alu__abc_41358_n671), .Y(alu__abc_41358_n672) );
  AND2X2 AND2X2_5815 ( .A(alu__abc_41358_n640), .B(alu__abc_41358_n201), .Y(alu__abc_41358_n673) );
  AND2X2 AND2X2_5816 ( .A(alu__abc_41358_n674), .B(alu__abc_41358_n675), .Y(alu__abc_41358_n676) );
  AND2X2 AND2X2_5817 ( .A(alu__abc_41358_n638), .B(alu__abc_41358_n219), .Y(alu__abc_41358_n677) );
  AND2X2 AND2X2_5818 ( .A(alu__abc_41358_n678), .B(alu__abc_41358_n214), .Y(alu__abc_41358_n679) );
  AND2X2 AND2X2_5819 ( .A(alu__abc_41358_n680), .B(alu__abc_41358_n228), .Y(alu__abc_41358_n681) );
  AND2X2 AND2X2_582 ( .A(_abc_43815_n1727), .B(enable_i_bF_buf7), .Y(_abc_43815_n1728) );
  AND2X2 AND2X2_5820 ( .A(alu__abc_41358_n679), .B(alu__abc_41358_n227), .Y(alu__abc_41358_n682) );
  AND2X2 AND2X2_5821 ( .A(alu__abc_41358_n678), .B(alu__abc_41358_n684), .Y(alu__abc_41358_n685) );
  AND2X2 AND2X2_5822 ( .A(alu__abc_41358_n607), .B(alu__abc_41358_n236), .Y(alu__abc_41358_n686) );
  AND2X2 AND2X2_5823 ( .A(alu__abc_41358_n687), .B(alu__abc_41358_n231), .Y(alu__abc_41358_n688) );
  AND2X2 AND2X2_5824 ( .A(alu__abc_41358_n688), .B(alu__abc_41358_n244), .Y(alu__abc_41358_n689) );
  AND2X2 AND2X2_5825 ( .A(alu__abc_41358_n690), .B(alu__abc_41358_n245), .Y(alu__abc_41358_n691) );
  AND2X2 AND2X2_5826 ( .A(alu__abc_41358_n687), .B(alu__abc_41358_n693), .Y(alu__abc_41358_n694) );
  AND2X2 AND2X2_5827 ( .A(alu__abc_41358_n602), .B(alu__abc_41358_n604), .Y(alu__abc_41358_n695) );
  AND2X2 AND2X2_5828 ( .A(alu__abc_41358_n696), .B(alu__abc_41358_n571), .Y(alu__abc_41358_n697) );
  AND2X2 AND2X2_5829 ( .A(alu__abc_41358_n698), .B(alu__abc_41358_n328), .Y(alu__abc_41358_n699) );
  AND2X2 AND2X2_583 ( .A(_abc_43815_n1726), .B(_abc_43815_n1728), .Y(epc_q_8__FF_INPUT) );
  AND2X2 AND2X2_5830 ( .A(alu__abc_41358_n701), .B(alu__abc_41358_n336), .Y(alu__abc_41358_n702) );
  AND2X2 AND2X2_5831 ( .A(alu__abc_41358_n700), .B(alu__abc_41358_n337), .Y(alu__abc_41358_n703) );
  AND2X2 AND2X2_5832 ( .A(alu__abc_41358_n602), .B(alu__abc_41358_n363), .Y(alu__abc_41358_n705) );
  AND2X2 AND2X2_5833 ( .A(alu__abc_41358_n707), .B(alu__abc_41358_n575), .Y(alu__abc_41358_n708) );
  AND2X2 AND2X2_5834 ( .A(alu__abc_41358_n709), .B(alu__abc_41358_n710), .Y(alu__abc_41358_n711) );
  AND2X2 AND2X2_5835 ( .A(alu__abc_41358_n713), .B(alu__abc_41358_n714), .Y(alu__abc_41358_n715) );
  AND2X2 AND2X2_5836 ( .A(alu__abc_41358_n715), .B(alu__abc_41358_n364), .Y(alu__abc_41358_n716) );
  AND2X2 AND2X2_5837 ( .A(alu__abc_41358_n587), .B(alu__abc_41358_n591), .Y(alu__abc_41358_n719) );
  AND2X2 AND2X2_5838 ( .A(alu__abc_41358_n720), .B(alu__abc_41358_n269), .Y(alu__abc_41358_n721) );
  AND2X2 AND2X2_5839 ( .A(alu__abc_41358_n722), .B(alu__abc_41358_n275), .Y(alu__abc_41358_n723) );
  AND2X2 AND2X2_584 ( .A(_abc_43815_n1694), .B(pc_q_9_), .Y(_abc_43815_n1731) );
  AND2X2 AND2X2_5840 ( .A(alu__abc_41358_n726), .B(alu__abc_41358_n724), .Y(alu__abc_41358_n727) );
  AND2X2 AND2X2_5841 ( .A(alu__abc_41358_n728), .B(alu__abc_41358_n264), .Y(alu__abc_41358_n729) );
  AND2X2 AND2X2_5842 ( .A(alu__abc_41358_n729), .B(alu__abc_41358_n588), .Y(alu__abc_41358_n730) );
  AND2X2 AND2X2_5843 ( .A(alu__abc_41358_n728), .B(alu__abc_41358_n732), .Y(alu__abc_41358_n733) );
  AND2X2 AND2X2_5844 ( .A(alu__abc_41358_n587), .B(alu__abc_41358_n283), .Y(alu__abc_41358_n734) );
  AND2X2 AND2X2_5845 ( .A(alu__abc_41358_n735), .B(alu__abc_41358_n289), .Y(alu__abc_41358_n736) );
  AND2X2 AND2X2_5846 ( .A(alu__abc_41358_n737), .B(alu__abc_41358_n278), .Y(alu__abc_41358_n738) );
  AND2X2 AND2X2_5847 ( .A(alu__abc_41358_n738), .B(alu__abc_41358_n590), .Y(alu__abc_41358_n739) );
  AND2X2 AND2X2_5848 ( .A(alu__abc_41358_n259_bF_buf3), .B(alu__abc_41358_n255), .Y(alu__abc_41358_n741) );
  AND2X2 AND2X2_5849 ( .A(alu__abc_41358_n742), .B(alu__abc_41358_n706), .Y(alu__abc_41358_n743) );
  AND2X2 AND2X2_585 ( .A(_abc_43815_n1732), .B(_abc_43815_n1730), .Y(_abc_43815_n1733) );
  AND2X2 AND2X2_5850 ( .A(alu__abc_41358_n743), .B(alu_c_i), .Y(alu__abc_41358_n744) );
  AND2X2 AND2X2_5851 ( .A(alu__abc_41358_n744), .B(alu__abc_41358_n577), .Y(alu__abc_41358_n745) );
  AND2X2 AND2X2_5852 ( .A(alu__abc_41358_n746), .B(alu__abc_41358_n748), .Y(alu__abc_41358_n749) );
  AND2X2 AND2X2_5853 ( .A(alu__abc_41358_n749), .B(alu__abc_41358_n745), .Y(alu__abc_41358_n750) );
  AND2X2 AND2X2_5854 ( .A(alu__abc_41358_n746), .B(alu__abc_41358_n752), .Y(alu__abc_41358_n753) );
  AND2X2 AND2X2_5855 ( .A(alu__abc_41358_n753), .B(alu__abc_41358_n751), .Y(alu__abc_41358_n754) );
  AND2X2 AND2X2_5856 ( .A(alu__abc_41358_n580), .B(alu__abc_41358_n747), .Y(alu__abc_41358_n755_1) );
  AND2X2 AND2X2_5857 ( .A(alu__abc_41358_n756), .B(alu__abc_41358_n296), .Y(alu__abc_41358_n757) );
  AND2X2 AND2X2_5858 ( .A(alu__abc_41358_n758), .B(alu__abc_41358_n750), .Y(alu__abc_41358_n759) );
  AND2X2 AND2X2_5859 ( .A(alu__abc_41358_n737), .B(alu__abc_41358_n760), .Y(alu__abc_41358_n761) );
  AND2X2 AND2X2_586 ( .A(_abc_43815_n1692), .B(_abc_43815_n1734), .Y(_abc_43815_n1735) );
  AND2X2 AND2X2_5860 ( .A(alu__abc_41358_n759), .B(alu__abc_41358_n761), .Y(alu__abc_41358_n762) );
  AND2X2 AND2X2_5861 ( .A(alu__abc_41358_n740), .B(alu__abc_41358_n762), .Y(alu__abc_41358_n763) );
  AND2X2 AND2X2_5862 ( .A(alu__abc_41358_n763), .B(alu__abc_41358_n733), .Y(alu__abc_41358_n764) );
  AND2X2 AND2X2_5863 ( .A(alu__abc_41358_n731), .B(alu__abc_41358_n764), .Y(alu__abc_41358_n765) );
  AND2X2 AND2X2_5864 ( .A(alu__abc_41358_n765), .B(alu__abc_41358_n718), .Y(alu__abc_41358_n766) );
  AND2X2 AND2X2_5865 ( .A(alu__abc_41358_n769), .B(alu__abc_41358_n767), .Y(alu__abc_41358_n770) );
  AND2X2 AND2X2_5866 ( .A(alu__abc_41358_n771), .B(alu__abc_41358_n772), .Y(alu__abc_41358_n773) );
  AND2X2 AND2X2_5867 ( .A(alu__abc_41358_n775), .B(alu__abc_41358_n565_1), .Y(alu__abc_41358_n776) );
  AND2X2 AND2X2_5868 ( .A(alu__abc_41358_n602), .B(alu__abc_41358_n603), .Y(alu__abc_41358_n778) );
  AND2X2 AND2X2_5869 ( .A(alu__abc_41358_n777), .B(alu__abc_41358_n780), .Y(alu__abc_41358_n781) );
  AND2X2 AND2X2_587 ( .A(_abc_43815_n1418_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n1736) );
  AND2X2 AND2X2_5870 ( .A(alu__abc_41358_n782), .B(alu__abc_41358_n372), .Y(alu__abc_41358_n783) );
  AND2X2 AND2X2_5871 ( .A(alu__abc_41358_n784), .B(alu__abc_41358_n358), .Y(alu__abc_41358_n785) );
  AND2X2 AND2X2_5872 ( .A(alu__abc_41358_n785), .B(alu__abc_41358_n371), .Y(alu__abc_41358_n786) );
  AND2X2 AND2X2_5873 ( .A(alu__abc_41358_n781), .B(alu__abc_41358_n787_1), .Y(alu__abc_41358_n788) );
  AND2X2 AND2X2_5874 ( .A(alu__abc_41358_n788), .B(alu__abc_41358_n773), .Y(alu__abc_41358_n789) );
  AND2X2 AND2X2_5875 ( .A(alu__abc_41358_n789), .B(alu__abc_41358_n766), .Y(alu__abc_41358_n790) );
  AND2X2 AND2X2_5876 ( .A(alu__abc_41358_n696), .B(alu__abc_41358_n311), .Y(alu__abc_41358_n791) );
  AND2X2 AND2X2_5877 ( .A(alu__abc_41358_n792), .B(alu__abc_41358_n320), .Y(alu__abc_41358_n793) );
  AND2X2 AND2X2_5878 ( .A(alu__abc_41358_n771), .B(alu__abc_41358_n306), .Y(alu__abc_41358_n794) );
  AND2X2 AND2X2_5879 ( .A(alu__abc_41358_n794), .B(alu__abc_41358_n319), .Y(alu__abc_41358_n795) );
  AND2X2 AND2X2_588 ( .A(_abc_43815_n1489_bF_buf1), .B(epc_q_9_), .Y(_abc_43815_n1737) );
  AND2X2 AND2X2_5880 ( .A(alu__abc_41358_n797), .B(alu__abc_41358_n798), .Y(alu__abc_41358_n799) );
  AND2X2 AND2X2_5881 ( .A(alu__abc_41358_n777), .B(alu__abc_41358_n341), .Y(alu__abc_41358_n800) );
  AND2X2 AND2X2_5882 ( .A(alu__abc_41358_n800), .B(alu__abc_41358_n354), .Y(alu__abc_41358_n801) );
  AND2X2 AND2X2_5883 ( .A(alu__abc_41358_n779), .B(alu__abc_41358_n346), .Y(alu__abc_41358_n802) );
  AND2X2 AND2X2_5884 ( .A(alu__abc_41358_n803), .B(alu__abc_41358_n355), .Y(alu__abc_41358_n804) );
  AND2X2 AND2X2_5885 ( .A(alu__abc_41358_n799), .B(alu__abc_41358_n805), .Y(alu__abc_41358_n806) );
  AND2X2 AND2X2_5886 ( .A(alu__abc_41358_n806), .B(alu__abc_41358_n796), .Y(alu__abc_41358_n807) );
  AND2X2 AND2X2_5887 ( .A(alu__abc_41358_n807), .B(alu__abc_41358_n790), .Y(alu__abc_41358_n808) );
  AND2X2 AND2X2_5888 ( .A(alu__abc_41358_n808), .B(alu__abc_41358_n704_1), .Y(alu__abc_41358_n809) );
  AND2X2 AND2X2_5889 ( .A(alu__abc_41358_n809), .B(alu__abc_41358_n694), .Y(alu__abc_41358_n810) );
  AND2X2 AND2X2_589 ( .A(_abc_43815_n1350_bF_buf2), .B(_abc_43815_n1738_1), .Y(_abc_43815_n1739_1) );
  AND2X2 AND2X2_5890 ( .A(alu__abc_41358_n810), .B(alu__abc_41358_n692), .Y(alu__abc_41358_n811) );
  AND2X2 AND2X2_5891 ( .A(alu__abc_41358_n811), .B(alu__abc_41358_n685), .Y(alu__abc_41358_n812) );
  AND2X2 AND2X2_5892 ( .A(alu__abc_41358_n812), .B(alu__abc_41358_n683), .Y(alu__abc_41358_n813) );
  AND2X2 AND2X2_5893 ( .A(alu__abc_41358_n813), .B(alu__abc_41358_n676), .Y(alu__abc_41358_n814) );
  AND2X2 AND2X2_5894 ( .A(alu__abc_41358_n814), .B(alu__abc_41358_n672), .Y(alu__abc_41358_n815) );
  AND2X2 AND2X2_5895 ( .A(alu__abc_41358_n674), .B(alu__abc_41358_n196_1), .Y(alu__abc_41358_n816) );
  AND2X2 AND2X2_5896 ( .A(alu__abc_41358_n816), .B(alu__abc_41358_n209), .Y(alu__abc_41358_n817) );
  AND2X2 AND2X2_5897 ( .A(alu__abc_41358_n818_1), .B(alu__abc_41358_n210), .Y(alu__abc_41358_n819) );
  AND2X2 AND2X2_5898 ( .A(alu__abc_41358_n631), .B(alu__abc_41358_n821), .Y(alu__abc_41358_n822) );
  AND2X2 AND2X2_5899 ( .A(alu__abc_41358_n822), .B(alu__abc_41358_n820), .Y(alu__abc_41358_n823) );
  AND2X2 AND2X2_59 ( .A(_abc_43815_n694), .B(\mem_dat_i[17] ), .Y(_abc_43815_n715) );
  AND2X2 AND2X2_590 ( .A(_abc_43815_n1740), .B(_abc_43815_n1066), .Y(_abc_43815_n1741) );
  AND2X2 AND2X2_5900 ( .A(alu__abc_41358_n815), .B(alu__abc_41358_n823), .Y(alu__abc_41358_n824) );
  AND2X2 AND2X2_5901 ( .A(alu__abc_41358_n824), .B(alu__abc_41358_n670), .Y(alu__abc_41358_n825) );
  AND2X2 AND2X2_5902 ( .A(alu__abc_41358_n825), .B(alu__abc_41358_n649), .Y(alu__abc_41358_n826) );
  AND2X2 AND2X2_5903 ( .A(alu__abc_41358_n826), .B(alu__abc_41358_n637), .Y(alu__abc_41358_n827) );
  AND2X2 AND2X2_5904 ( .A(alu__abc_41358_n827), .B(alu__abc_41358_n627), .Y(alu__abc_41358_n828) );
  AND2X2 AND2X2_5905 ( .A(alu__abc_41358_n828), .B(alu_op_i_0_bF_buf4), .Y(alu__abc_41358_n829) );
  AND2X2 AND2X2_5906 ( .A(alu__abc_41358_n830), .B(alu_c_update_o), .Y(alu_c_o) );
  AND2X2 AND2X2_5907 ( .A(alu__abc_41358_n382), .B(alu__abc_41358_n379), .Y(alu__abc_41358_n832) );
  AND2X2 AND2X2_5908 ( .A(alu__abc_41358_n832), .B(alu_op_i_1_), .Y(alu__abc_41358_n833) );
  AND2X2 AND2X2_5909 ( .A(alu__abc_41358_n742), .B(alu__abc_41358_n834), .Y(alu__abc_41358_n835) );
  AND2X2 AND2X2_591 ( .A(_abc_43815_n1710), .B(_abc_43815_n1706_1), .Y(_abc_43815_n1742) );
  AND2X2 AND2X2_5910 ( .A(alu__abc_41358_n835), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n836) );
  AND2X2 AND2X2_5911 ( .A(alu__abc_41358_n838), .B(alu__abc_41358_n837), .Y(alu__abc_41358_n839) );
  AND2X2 AND2X2_5912 ( .A(alu__abc_41358_n839), .B(alu_b_i_1_bF_buf4), .Y(alu__abc_41358_n840) );
  AND2X2 AND2X2_5913 ( .A(alu__abc_41358_n844), .B(alu__abc_41358_n843), .Y(alu__abc_41358_n845) );
  AND2X2 AND2X2_5914 ( .A(alu__abc_41358_n848), .B(alu__abc_41358_n847_1), .Y(alu__abc_41358_n849) );
  AND2X2 AND2X2_5915 ( .A(alu__abc_41358_n846), .B(alu__abc_41358_n850), .Y(alu__abc_41358_n851) );
  AND2X2 AND2X2_5916 ( .A(alu__abc_41358_n852), .B(alu__abc_41358_n842), .Y(alu__abc_41358_n853) );
  AND2X2 AND2X2_5917 ( .A(alu__abc_41358_n856), .B(alu__abc_41358_n855), .Y(alu__abc_41358_n857) );
  AND2X2 AND2X2_5918 ( .A(alu__abc_41358_n860), .B(alu__abc_41358_n859), .Y(alu__abc_41358_n861) );
  AND2X2 AND2X2_5919 ( .A(alu__abc_41358_n858), .B(alu__abc_41358_n862), .Y(alu__abc_41358_n863) );
  AND2X2 AND2X2_592 ( .A(alu_op_r_5_), .B(pc_q_9_), .Y(_abc_43815_n1745) );
  AND2X2 AND2X2_5920 ( .A(alu__abc_41358_n866), .B(alu__abc_41358_n865), .Y(alu__abc_41358_n867) );
  AND2X2 AND2X2_5921 ( .A(alu__abc_41358_n870), .B(alu__abc_41358_n869), .Y(alu__abc_41358_n871) );
  AND2X2 AND2X2_5922 ( .A(alu__abc_41358_n868), .B(alu__abc_41358_n872_1), .Y(alu__abc_41358_n873) );
  AND2X2 AND2X2_5923 ( .A(alu__abc_41358_n864), .B(alu__abc_41358_n874), .Y(alu__abc_41358_n875) );
  AND2X2 AND2X2_5924 ( .A(alu__abc_41358_n876), .B(alu__abc_41358_n854), .Y(alu__abc_41358_n877) );
  AND2X2 AND2X2_5925 ( .A(alu__abc_41358_n880), .B(alu__abc_41358_n879), .Y(alu__abc_41358_n881) );
  AND2X2 AND2X2_5926 ( .A(alu__abc_41358_n884), .B(alu__abc_41358_n883), .Y(alu__abc_41358_n885) );
  AND2X2 AND2X2_5927 ( .A(alu__abc_41358_n882), .B(alu__abc_41358_n886), .Y(alu__abc_41358_n887) );
  AND2X2 AND2X2_5928 ( .A(alu__abc_41358_n890), .B(alu__abc_41358_n889), .Y(alu__abc_41358_n891) );
  AND2X2 AND2X2_5929 ( .A(alu__abc_41358_n894), .B(alu__abc_41358_n893), .Y(alu__abc_41358_n895) );
  AND2X2 AND2X2_593 ( .A(_abc_43815_n1746), .B(_abc_43815_n1744), .Y(_abc_43815_n1747) );
  AND2X2 AND2X2_5930 ( .A(alu__abc_41358_n892), .B(alu__abc_41358_n896), .Y(alu__abc_41358_n897) );
  AND2X2 AND2X2_5931 ( .A(alu__abc_41358_n888), .B(alu__abc_41358_n898), .Y(alu__abc_41358_n899) );
  AND2X2 AND2X2_5932 ( .A(alu__abc_41358_n902), .B(alu__abc_41358_n901), .Y(alu__abc_41358_n903_1) );
  AND2X2 AND2X2_5933 ( .A(alu__abc_41358_n906), .B(alu__abc_41358_n905), .Y(alu__abc_41358_n907) );
  AND2X2 AND2X2_5934 ( .A(alu__abc_41358_n904), .B(alu__abc_41358_n908), .Y(alu__abc_41358_n909) );
  AND2X2 AND2X2_5935 ( .A(alu__abc_41358_n912), .B(alu__abc_41358_n911), .Y(alu__abc_41358_n913) );
  AND2X2 AND2X2_5936 ( .A(alu__abc_41358_n916), .B(alu__abc_41358_n915), .Y(alu__abc_41358_n917) );
  AND2X2 AND2X2_5937 ( .A(alu__abc_41358_n914), .B(alu__abc_41358_n918), .Y(alu__abc_41358_n919) );
  AND2X2 AND2X2_5938 ( .A(alu__abc_41358_n910), .B(alu__abc_41358_n920), .Y(alu__abc_41358_n921) );
  AND2X2 AND2X2_5939 ( .A(alu__abc_41358_n900), .B(alu__abc_41358_n922), .Y(alu__abc_41358_n923) );
  AND2X2 AND2X2_594 ( .A(_abc_43815_n1743), .B(_abc_43815_n1748), .Y(_abc_43815_n1749) );
  AND2X2 AND2X2_5940 ( .A(alu__abc_41358_n924), .B(alu__abc_41358_n878), .Y(alu__abc_41358_n925) );
  AND2X2 AND2X2_5941 ( .A(alu__abc_41358_n925), .B(alu__abc_41358_n833_bF_buf4), .Y(alu__abc_41358_n926) );
  AND2X2 AND2X2_5942 ( .A(alu__abc_41358_n383), .B(alu__abc_41358_n378), .Y(alu__abc_41358_n927) );
  AND2X2 AND2X2_5943 ( .A(alu__abc_41358_n378), .B(alu__abc_41358_n384), .Y(alu__abc_41358_n929) );
  AND2X2 AND2X2_5944 ( .A(alu__abc_41358_n929), .B(alu__abc_41358_n382), .Y(alu__abc_41358_n930) );
  AND2X2 AND2X2_5945 ( .A(alu__abc_41358_n931), .B(alu__abc_41358_n928), .Y(alu__abc_41358_n932) );
  AND2X2 AND2X2_5946 ( .A(alu__abc_41358_n932_bF_buf4), .B(alu_a_i_0_), .Y(alu__abc_41358_n933_1) );
  AND2X2 AND2X2_5947 ( .A(alu_op_i_1_), .B(alu_op_i_0_bF_buf3), .Y(alu__abc_41358_n934) );
  AND2X2 AND2X2_5948 ( .A(alu__abc_41358_n380), .B(alu__abc_41358_n934), .Y(alu__abc_41358_n935) );
  AND2X2 AND2X2_5949 ( .A(alu__abc_41358_n935_bF_buf4), .B(alu__abc_41358_n578), .Y(alu__abc_41358_n936) );
  AND2X2 AND2X2_595 ( .A(_abc_43815_n1742), .B(_abc_43815_n1747), .Y(_abc_43815_n1750_1) );
  AND2X2 AND2X2_5950 ( .A(alu__abc_41358_n380), .B(alu__abc_41358_n384), .Y(alu__abc_41358_n937) );
  AND2X2 AND2X2_5951 ( .A(alu__abc_41358_n743), .B(alu__abc_41358_n937), .Y(alu__abc_41358_n938) );
  AND2X2 AND2X2_5952 ( .A(alu__abc_41358_n378), .B(alu_op_i_0_bF_buf2), .Y(alu__abc_41358_n941) );
  AND2X2 AND2X2_5953 ( .A(alu__abc_41358_n380), .B(alu__abc_41358_n941), .Y(alu__abc_41358_n942) );
  AND2X2 AND2X2_5954 ( .A(alu__abc_41358_n943), .B(alu__abc_41358_n944), .Y(alu__abc_41358_n945) );
  AND2X2 AND2X2_5955 ( .A(alu__abc_41358_n945), .B(alu__abc_41358_n942_bF_buf4), .Y(alu__abc_41358_n946) );
  AND2X2 AND2X2_5956 ( .A(alu__abc_41358_n832), .B(alu__abc_41358_n941), .Y(alu__abc_41358_n947) );
  AND2X2 AND2X2_5957 ( .A(alu__abc_41358_n947), .B(alu__abc_41358_n279_bF_buf2), .Y(alu__abc_41358_n948) );
  AND2X2 AND2X2_5958 ( .A(alu__abc_41358_n260), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n949) );
  AND2X2 AND2X2_5959 ( .A(alu__abc_41358_n949), .B(alu__abc_41358_n299_bF_buf1), .Y(alu__abc_41358_n950) );
  AND2X2 AND2X2_596 ( .A(_abc_43815_n1752), .B(_abc_43815_n1741), .Y(_abc_43815_n1753_1) );
  AND2X2 AND2X2_5960 ( .A(alu__abc_41358_n950), .B(alu__abc_41358_n294_bF_buf3), .Y(alu__abc_41358_n951) );
  AND2X2 AND2X2_5961 ( .A(alu__abc_41358_n951), .B(alu__abc_41358_n948_bF_buf4), .Y(alu__abc_41358_n952) );
  AND2X2 AND2X2_5962 ( .A(alu__abc_41358_n742), .B(alu__abc_41358_n384), .Y(alu__abc_41358_n954) );
  AND2X2 AND2X2_5963 ( .A(alu__abc_41358_n743), .B(alu_op_i_0_bF_buf1), .Y(alu__abc_41358_n955) );
  AND2X2 AND2X2_5964 ( .A(alu__abc_41358_n956), .B(alu__abc_41358_n927_bF_buf3), .Y(alu__abc_41358_n957) );
  AND2X2 AND2X2_5965 ( .A(alu__abc_41358_n934), .B(alu_a_i_31_), .Y(alu__abc_41358_n961) );
  AND2X2 AND2X2_5966 ( .A(alu__abc_41358_n961), .B(alu__abc_41358_n832), .Y(alu__abc_41358_n962) );
  AND2X2 AND2X2_5967 ( .A(alu__abc_41358_n259_bF_buf1), .B(alu_a_i_31_), .Y(alu__abc_41358_n963) );
  AND2X2 AND2X2_5968 ( .A(alu__abc_41358_n964), .B(alu_b_i_1_bF_buf4), .Y(alu__abc_41358_n965) );
  AND2X2 AND2X2_5969 ( .A(alu_a_i_30_), .B(alu_b_i_0_bF_buf1), .Y(alu__abc_41358_n966) );
  AND2X2 AND2X2_597 ( .A(_abc_43815_n1065_1_bF_buf1), .B(epc_q_9_), .Y(_abc_43815_n1754) );
  AND2X2 AND2X2_5970 ( .A(alu__abc_41358_n259_bF_buf0), .B(alu_a_i_29_), .Y(alu__abc_41358_n967) );
  AND2X2 AND2X2_5971 ( .A(alu__abc_41358_n968), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n969) );
  AND2X2 AND2X2_5972 ( .A(alu__abc_41358_n970), .B(alu_b_i_2_bF_buf0), .Y(alu__abc_41358_n971) );
  AND2X2 AND2X2_5973 ( .A(alu__abc_41358_n973), .B(alu__abc_41358_n972), .Y(alu__abc_41358_n974) );
  AND2X2 AND2X2_5974 ( .A(alu__abc_41358_n977), .B(alu__abc_41358_n976), .Y(alu__abc_41358_n978) );
  AND2X2 AND2X2_5975 ( .A(alu__abc_41358_n975_1), .B(alu__abc_41358_n979), .Y(alu__abc_41358_n980) );
  AND2X2 AND2X2_5976 ( .A(alu__abc_41358_n980), .B(alu__abc_41358_n299_bF_buf0), .Y(alu__abc_41358_n981) );
  AND2X2 AND2X2_5977 ( .A(alu__abc_41358_n982), .B(alu_b_i_3_bF_buf1), .Y(alu__abc_41358_n983) );
  AND2X2 AND2X2_5978 ( .A(alu__abc_41358_n985), .B(alu__abc_41358_n984), .Y(alu__abc_41358_n986) );
  AND2X2 AND2X2_5979 ( .A(alu__abc_41358_n989), .B(alu__abc_41358_n988), .Y(alu__abc_41358_n990) );
  AND2X2 AND2X2_598 ( .A(_abc_43815_n1472_1_bF_buf1), .B(_abc_43815_n1757), .Y(_abc_43815_n1758) );
  AND2X2 AND2X2_5980 ( .A(alu__abc_41358_n987), .B(alu__abc_41358_n991), .Y(alu__abc_41358_n992) );
  AND2X2 AND2X2_5981 ( .A(alu__abc_41358_n995), .B(alu__abc_41358_n994), .Y(alu__abc_41358_n996) );
  AND2X2 AND2X2_5982 ( .A(alu__abc_41358_n999), .B(alu__abc_41358_n998), .Y(alu__abc_41358_n1000) );
  AND2X2 AND2X2_5983 ( .A(alu__abc_41358_n997), .B(alu__abc_41358_n1001_1), .Y(alu__abc_41358_n1002) );
  AND2X2 AND2X2_5984 ( .A(alu__abc_41358_n993), .B(alu__abc_41358_n1003), .Y(alu__abc_41358_n1004) );
  AND2X2 AND2X2_5985 ( .A(alu__abc_41358_n1004), .B(alu__abc_41358_n294_bF_buf2), .Y(alu__abc_41358_n1005) );
  AND2X2 AND2X2_5986 ( .A(alu__abc_41358_n1009), .B(alu__abc_41358_n252_bF_buf5), .Y(alu__abc_41358_n1010) );
  AND2X2 AND2X2_5987 ( .A(alu__abc_41358_n1010), .B(alu__abc_41358_n1008), .Y(alu__abc_41358_n1011) );
  AND2X2 AND2X2_5988 ( .A(alu__abc_41358_n1013), .B(alu__abc_41358_n1012), .Y(alu__abc_41358_n1014) );
  AND2X2 AND2X2_5989 ( .A(alu__abc_41358_n1014), .B(alu_b_i_1_bF_buf0), .Y(alu__abc_41358_n1015) );
  AND2X2 AND2X2_599 ( .A(_abc_43815_n1756), .B(_abc_43815_n1758), .Y(_abc_43815_n1759) );
  AND2X2 AND2X2_5990 ( .A(alu__abc_41358_n1019), .B(alu__abc_41358_n1018), .Y(alu__abc_41358_n1020) );
  AND2X2 AND2X2_5991 ( .A(alu__abc_41358_n1023), .B(alu__abc_41358_n1022), .Y(alu__abc_41358_n1024_1) );
  AND2X2 AND2X2_5992 ( .A(alu__abc_41358_n1021), .B(alu__abc_41358_n1025), .Y(alu__abc_41358_n1026) );
  AND2X2 AND2X2_5993 ( .A(alu__abc_41358_n1027), .B(alu__abc_41358_n1017), .Y(alu__abc_41358_n1028) );
  AND2X2 AND2X2_5994 ( .A(alu__abc_41358_n1031), .B(alu__abc_41358_n1030), .Y(alu__abc_41358_n1032) );
  AND2X2 AND2X2_5995 ( .A(alu__abc_41358_n1035), .B(alu__abc_41358_n1034), .Y(alu__abc_41358_n1036) );
  AND2X2 AND2X2_5996 ( .A(alu__abc_41358_n1033), .B(alu__abc_41358_n1037), .Y(alu__abc_41358_n1038) );
  AND2X2 AND2X2_5997 ( .A(alu__abc_41358_n1041), .B(alu__abc_41358_n1040), .Y(alu__abc_41358_n1042) );
  AND2X2 AND2X2_5998 ( .A(alu__abc_41358_n1045), .B(alu__abc_41358_n1044), .Y(alu__abc_41358_n1046) );
  AND2X2 AND2X2_5999 ( .A(alu__abc_41358_n1043), .B(alu__abc_41358_n1047), .Y(alu__abc_41358_n1048) );
  AND2X2 AND2X2_6 ( .A(_abc_43815_n627_1), .B(_abc_43815_n621), .Y(_abc_43815_n628) );
  AND2X2 AND2X2_60 ( .A(_abc_43815_n697), .B(\mem_dat_i[1] ), .Y(_abc_43815_n716) );
  AND2X2 AND2X2_600 ( .A(_abc_43815_n1473_bF_buf2), .B(_abc_43815_n1733), .Y(_abc_43815_n1760) );
  AND2X2 AND2X2_6000 ( .A(alu__abc_41358_n1039), .B(alu__abc_41358_n1049), .Y(alu__abc_41358_n1050_1) );
  AND2X2 AND2X2_6001 ( .A(alu__abc_41358_n1051), .B(alu__abc_41358_n1029), .Y(alu__abc_41358_n1052) );
  AND2X2 AND2X2_6002 ( .A(alu__abc_41358_n1053), .B(alu__abc_41358_n833_bF_buf3), .Y(alu__abc_41358_n1054) );
  AND2X2 AND2X2_6003 ( .A(alu__abc_41358_n1007), .B(alu__abc_41358_n1054), .Y(alu__abc_41358_n1055) );
  AND2X2 AND2X2_6004 ( .A(alu__abc_41358_n380), .B(alu__abc_41358_n385), .Y(alu__abc_41358_n1057) );
  AND2X2 AND2X2_6005 ( .A(alu__abc_41358_n1058), .B(alu__abc_41358_n1057_bF_buf4), .Y(alu__abc_41358_n1059) );
  AND2X2 AND2X2_6006 ( .A(alu__abc_41358_n1059), .B(alu__abc_41358_n1056), .Y(alu__abc_41358_n1060) );
  AND2X2 AND2X2_6007 ( .A(alu__abc_41358_n929), .B(alu__abc_41358_n380), .Y(alu__abc_41358_n1061) );
  AND2X2 AND2X2_6008 ( .A(alu__abc_41358_n707), .B(alu__abc_41358_n1062), .Y(alu__abc_41358_n1063) );
  AND2X2 AND2X2_6009 ( .A(alu__abc_41358_n1063), .B(alu__abc_41358_n1061_bF_buf4), .Y(alu__abc_41358_n1064) );
  AND2X2 AND2X2_601 ( .A(_abc_43815_n1761), .B(_abc_43815_n1413_bF_buf0), .Y(_abc_43815_n1762) );
  AND2X2 AND2X2_6010 ( .A(alu__abc_41358_n250), .B(alu_op_i_0_bF_buf0), .Y(alu__abc_41358_n1065) );
  AND2X2 AND2X2_6011 ( .A(alu__abc_41358_n927_bF_buf2), .B(alu__abc_41358_n576), .Y(alu__abc_41358_n1067) );
  AND2X2 AND2X2_6012 ( .A(alu__abc_41358_n1067), .B(alu__abc_41358_n1066), .Y(alu__abc_41358_n1068) );
  AND2X2 AND2X2_6013 ( .A(alu__abc_41358_n1072), .B(alu__abc_41358_n942_bF_buf3), .Y(alu__abc_41358_n1073) );
  AND2X2 AND2X2_6014 ( .A(alu__abc_41358_n1073), .B(alu__abc_41358_n1071), .Y(alu__abc_41358_n1074_1) );
  AND2X2 AND2X2_6015 ( .A(alu__abc_41358_n1010), .B(alu__abc_41358_n257), .Y(alu__abc_41358_n1075) );
  AND2X2 AND2X2_6016 ( .A(alu__abc_41358_n1075), .B(alu__abc_41358_n299_bF_buf4), .Y(alu__abc_41358_n1076) );
  AND2X2 AND2X2_6017 ( .A(alu__abc_41358_n1076), .B(alu__abc_41358_n294_bF_buf0), .Y(alu__abc_41358_n1077) );
  AND2X2 AND2X2_6018 ( .A(alu__abc_41358_n1077), .B(alu__abc_41358_n948_bF_buf3), .Y(alu__abc_41358_n1078) );
  AND2X2 AND2X2_6019 ( .A(alu__abc_41358_n932_bF_buf3), .B(alu_a_i_1_), .Y(alu__abc_41358_n1079) );
  AND2X2 AND2X2_602 ( .A(_abc_43815_n1763), .B(_abc_43815_n1351_bF_buf2), .Y(_abc_43815_n1764) );
  AND2X2 AND2X2_6020 ( .A(alu__abc_41358_n935_bF_buf3), .B(alu__abc_41358_n250), .Y(alu__abc_41358_n1080) );
  AND2X2 AND2X2_6021 ( .A(alu__abc_41358_n1087), .B(alu__abc_41358_n1086), .Y(alu__abc_41358_n1088) );
  AND2X2 AND2X2_6022 ( .A(alu__abc_41358_n1088), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n1089) );
  AND2X2 AND2X2_6023 ( .A(alu__abc_41358_n1090), .B(alu__abc_41358_n1091), .Y(alu__abc_41358_n1092) );
  AND2X2 AND2X2_6024 ( .A(alu__abc_41358_n1092), .B(alu__abc_41358_n299_bF_buf3), .Y(alu__abc_41358_n1093) );
  AND2X2 AND2X2_6025 ( .A(alu__abc_41358_n1094), .B(alu_b_i_3_bF_buf6), .Y(alu__abc_41358_n1095) );
  AND2X2 AND2X2_6026 ( .A(alu__abc_41358_n1096), .B(alu__abc_41358_n1097_1), .Y(alu__abc_41358_n1098) );
  AND2X2 AND2X2_6027 ( .A(alu__abc_41358_n1100), .B(alu__abc_41358_n1101), .Y(alu__abc_41358_n1102) );
  AND2X2 AND2X2_6028 ( .A(alu__abc_41358_n1099), .B(alu__abc_41358_n1103), .Y(alu__abc_41358_n1104) );
  AND2X2 AND2X2_6029 ( .A(alu__abc_41358_n1104), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n1105) );
  AND2X2 AND2X2_603 ( .A(_abc_43815_n1766), .B(enable_i_bF_buf6), .Y(_abc_43815_n1767) );
  AND2X2 AND2X2_6030 ( .A(alu__abc_41358_n839), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n1108) );
  AND2X2 AND2X2_6031 ( .A(alu__abc_41358_n845), .B(alu_b_i_1_bF_buf0), .Y(alu__abc_41358_n1109) );
  AND2X2 AND2X2_6032 ( .A(alu__abc_41358_n1112), .B(alu__abc_41358_n1113), .Y(alu__abc_41358_n1114) );
  AND2X2 AND2X2_6033 ( .A(alu__abc_41358_n1115), .B(alu__abc_41358_n1111), .Y(alu__abc_41358_n1116) );
  AND2X2 AND2X2_6034 ( .A(alu__abc_41358_n1116), .B(alu__abc_41358_n294_bF_buf6), .Y(alu__abc_41358_n1117_1) );
  AND2X2 AND2X2_6035 ( .A(alu__abc_41358_n1118), .B(alu__abc_41358_n1119), .Y(alu__abc_41358_n1120) );
  AND2X2 AND2X2_6036 ( .A(alu__abc_41358_n1122), .B(alu__abc_41358_n1123), .Y(alu__abc_41358_n1124) );
  AND2X2 AND2X2_6037 ( .A(alu__abc_41358_n1121), .B(alu__abc_41358_n1125), .Y(alu__abc_41358_n1126) );
  AND2X2 AND2X2_6038 ( .A(alu__abc_41358_n1126), .B(alu_b_i_3_bF_buf5), .Y(alu__abc_41358_n1127) );
  AND2X2 AND2X2_6039 ( .A(alu__abc_41358_n1129), .B(alu__abc_41358_n833_bF_buf2), .Y(alu__abc_41358_n1130) );
  AND2X2 AND2X2_604 ( .A(_abc_43815_n1765), .B(_abc_43815_n1767), .Y(epc_q_9__FF_INPUT) );
  AND2X2 AND2X2_6040 ( .A(alu__abc_41358_n1130), .B(alu__abc_41358_n1107), .Y(alu__abc_41358_n1131) );
  AND2X2 AND2X2_6041 ( .A(alu__abc_41358_n297), .B(alu_op_i_0_bF_buf5), .Y(alu__abc_41358_n1132) );
  AND2X2 AND2X2_6042 ( .A(alu__abc_41358_n927_bF_buf1), .B(alu__abc_41358_n1134), .Y(alu__abc_41358_n1135) );
  AND2X2 AND2X2_6043 ( .A(alu__abc_41358_n1135), .B(alu__abc_41358_n1133), .Y(alu__abc_41358_n1136) );
  AND2X2 AND2X2_6044 ( .A(alu__abc_41358_n1138), .B(alu__abc_41358_n1057_bF_buf3), .Y(alu__abc_41358_n1139) );
  AND2X2 AND2X2_6045 ( .A(alu__abc_41358_n1139), .B(alu__abc_41358_n1137_1), .Y(alu__abc_41358_n1140) );
  AND2X2 AND2X2_6046 ( .A(alu__abc_41358_n834), .B(alu__abc_41358_n837), .Y(alu__abc_41358_n1141) );
  AND2X2 AND2X2_6047 ( .A(alu__abc_41358_n261), .B(alu_b_i_1_bF_buf3), .Y(alu__abc_41358_n1143) );
  AND2X2 AND2X2_6048 ( .A(alu__abc_41358_n1142), .B(alu__abc_41358_n1144), .Y(alu__abc_41358_n1145) );
  AND2X2 AND2X2_6049 ( .A(alu__abc_41358_n1145), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n1146) );
  AND2X2 AND2X2_605 ( .A(_abc_43815_n1731), .B(pc_q_10_), .Y(_abc_43815_n1770) );
  AND2X2 AND2X2_6050 ( .A(alu__abc_41358_n1146), .B(alu__abc_41358_n294_bF_buf5), .Y(alu__abc_41358_n1147) );
  AND2X2 AND2X2_6051 ( .A(alu__abc_41358_n1147), .B(alu__abc_41358_n948_bF_buf2), .Y(alu__abc_41358_n1148) );
  AND2X2 AND2X2_6052 ( .A(alu__abc_41358_n1152), .B(alu__abc_41358_n942_bF_buf2), .Y(alu__abc_41358_n1153) );
  AND2X2 AND2X2_6053 ( .A(alu__abc_41358_n1153), .B(alu__abc_41358_n1151), .Y(alu__abc_41358_n1154) );
  AND2X2 AND2X2_6054 ( .A(alu__abc_41358_n749), .B(alu__abc_41358_n1061_bF_buf3), .Y(alu__abc_41358_n1155) );
  AND2X2 AND2X2_6055 ( .A(alu__abc_41358_n932_bF_buf2), .B(alu_a_i_2_), .Y(alu__abc_41358_n1156) );
  AND2X2 AND2X2_6056 ( .A(alu__abc_41358_n935_bF_buf2), .B(alu__abc_41358_n297), .Y(alu__abc_41358_n1157) );
  AND2X2 AND2X2_6057 ( .A(alu__abc_41358_n964), .B(alu__abc_41358_n1087), .Y(alu__abc_41358_n1163) );
  AND2X2 AND2X2_6058 ( .A(alu__abc_41358_n1163), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n1164) );
  AND2X2 AND2X2_6059 ( .A(alu__abc_41358_n1165), .B(alu__abc_41358_n1166), .Y(alu__abc_41358_n1167) );
  AND2X2 AND2X2_606 ( .A(_abc_43815_n1771), .B(_abc_43815_n1769_1), .Y(_abc_43815_n1772) );
  AND2X2 AND2X2_6060 ( .A(alu__abc_41358_n1167), .B(alu__abc_41358_n299_bF_buf6), .Y(alu__abc_41358_n1168) );
  AND2X2 AND2X2_6061 ( .A(alu__abc_41358_n1169), .B(alu_b_i_3_bF_buf4), .Y(alu__abc_41358_n1170) );
  AND2X2 AND2X2_6062 ( .A(alu__abc_41358_n1171), .B(alu__abc_41358_n1172), .Y(alu__abc_41358_n1173) );
  AND2X2 AND2X2_6063 ( .A(alu__abc_41358_n1175), .B(alu__abc_41358_n1176), .Y(alu__abc_41358_n1177) );
  AND2X2 AND2X2_6064 ( .A(alu__abc_41358_n1174), .B(alu__abc_41358_n1178), .Y(alu__abc_41358_n1179) );
  AND2X2 AND2X2_6065 ( .A(alu__abc_41358_n1179), .B(alu__abc_41358_n294_bF_buf4), .Y(alu__abc_41358_n1180) );
  AND2X2 AND2X2_6066 ( .A(alu__abc_41358_n1014), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n1183) );
  AND2X2 AND2X2_6067 ( .A(alu__abc_41358_n1020), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n1184) );
  AND2X2 AND2X2_6068 ( .A(alu__abc_41358_n1187), .B(alu__abc_41358_n1188), .Y(alu__abc_41358_n1189) );
  AND2X2 AND2X2_6069 ( .A(alu__abc_41358_n1190), .B(alu__abc_41358_n1186), .Y(alu__abc_41358_n1191) );
  AND2X2 AND2X2_607 ( .A(_abc_43815_n1692), .B(_abc_43815_n1773), .Y(_abc_43815_n1774) );
  AND2X2 AND2X2_6070 ( .A(alu__abc_41358_n1191), .B(alu__abc_41358_n294_bF_buf3), .Y(alu__abc_41358_n1192) );
  AND2X2 AND2X2_6071 ( .A(alu__abc_41358_n1193), .B(alu__abc_41358_n1194), .Y(alu__abc_41358_n1195) );
  AND2X2 AND2X2_6072 ( .A(alu__abc_41358_n1197), .B(alu__abc_41358_n1198), .Y(alu__abc_41358_n1199) );
  AND2X2 AND2X2_6073 ( .A(alu__abc_41358_n1196), .B(alu__abc_41358_n1200), .Y(alu__abc_41358_n1201) );
  AND2X2 AND2X2_6074 ( .A(alu__abc_41358_n1201), .B(alu_b_i_3_bF_buf3), .Y(alu__abc_41358_n1202_1) );
  AND2X2 AND2X2_6075 ( .A(alu__abc_41358_n1204), .B(alu__abc_41358_n833_bF_buf1), .Y(alu__abc_41358_n1205) );
  AND2X2 AND2X2_6076 ( .A(alu__abc_41358_n1205), .B(alu__abc_41358_n1182), .Y(alu__abc_41358_n1206) );
  AND2X2 AND2X2_6077 ( .A(alu__abc_41358_n1208), .B(alu__abc_41358_n942_bF_buf1), .Y(alu__abc_41358_n1209) );
  AND2X2 AND2X2_6078 ( .A(alu__abc_41358_n1209), .B(alu__abc_41358_n1207), .Y(alu__abc_41358_n1210) );
  AND2X2 AND2X2_6079 ( .A(alu__abc_41358_n1137_1), .B(alu__abc_41358_n1211), .Y(alu__abc_41358_n1212) );
  AND2X2 AND2X2_608 ( .A(_abc_43815_n1418_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_43815_n1775_1) );
  AND2X2 AND2X2_6080 ( .A(alu__abc_41358_n1214), .B(alu__abc_41358_n1057_bF_buf2), .Y(alu__abc_41358_n1215) );
  AND2X2 AND2X2_6081 ( .A(alu__abc_41358_n1215), .B(alu__abc_41358_n1213), .Y(alu__abc_41358_n1216) );
  AND2X2 AND2X2_6082 ( .A(alu__abc_41358_n758), .B(alu__abc_41358_n1061_bF_buf2), .Y(alu__abc_41358_n1217) );
  AND2X2 AND2X2_6083 ( .A(alu__abc_41358_n257), .B(alu__abc_41358_n1009), .Y(alu__abc_41358_n1218) );
  AND2X2 AND2X2_6084 ( .A(alu__abc_41358_n1008), .B(alu__abc_41358_n1012), .Y(alu__abc_41358_n1220) );
  AND2X2 AND2X2_6085 ( .A(alu__abc_41358_n1219), .B(alu__abc_41358_n1221), .Y(alu__abc_41358_n1222) );
  AND2X2 AND2X2_6086 ( .A(alu__abc_41358_n1222), .B(alu__abc_41358_n299_bF_buf2), .Y(alu__abc_41358_n1223_1) );
  AND2X2 AND2X2_6087 ( .A(alu__abc_41358_n1223_1), .B(alu__abc_41358_n294_bF_buf2), .Y(alu__abc_41358_n1224) );
  AND2X2 AND2X2_6088 ( .A(alu__abc_41358_n1224), .B(alu__abc_41358_n948_bF_buf1), .Y(alu__abc_41358_n1225) );
  AND2X2 AND2X2_6089 ( .A(alu__abc_41358_n292), .B(alu_op_i_0_bF_buf4), .Y(alu__abc_41358_n1226) );
  AND2X2 AND2X2_609 ( .A(_abc_43815_n1489_bF_buf0), .B(epc_q_10_), .Y(_abc_43815_n1776) );
  AND2X2 AND2X2_6090 ( .A(alu__abc_41358_n927_bF_buf0), .B(alu__abc_41358_n584), .Y(alu__abc_41358_n1228) );
  AND2X2 AND2X2_6091 ( .A(alu__abc_41358_n1228), .B(alu__abc_41358_n1227), .Y(alu__abc_41358_n1229) );
  AND2X2 AND2X2_6092 ( .A(alu__abc_41358_n932_bF_buf1), .B(alu_a_i_3_), .Y(alu__abc_41358_n1230) );
  AND2X2 AND2X2_6093 ( .A(alu__abc_41358_n935_bF_buf1), .B(alu__abc_41358_n292), .Y(alu__abc_41358_n1231) );
  AND2X2 AND2X2_6094 ( .A(alu__abc_41358_n1240), .B(alu__abc_41358_n942_bF_buf0), .Y(alu__abc_41358_n1241) );
  AND2X2 AND2X2_6095 ( .A(alu__abc_41358_n1241), .B(alu__abc_41358_n1239), .Y(alu__abc_41358_n1242) );
  AND2X2 AND2X2_6096 ( .A(alu__abc_41358_n1244), .B(alu__abc_41358_n294_bF_buf1), .Y(alu__abc_41358_n1245) );
  AND2X2 AND2X2_6097 ( .A(alu__abc_41358_n1245), .B(alu__abc_41358_n1243_1), .Y(alu__abc_41358_n1246) );
  AND2X2 AND2X2_6098 ( .A(alu__abc_41358_n1247), .B(alu__abc_41358_n1248), .Y(alu__abc_41358_n1249) );
  AND2X2 AND2X2_6099 ( .A(alu__abc_41358_n1249), .B(alu_b_i_3_bF_buf2), .Y(alu__abc_41358_n1250) );
  AND2X2 AND2X2_61 ( .A(_abc_43815_n706_1), .B(\mem_dat_i[1] ), .Y(_abc_43815_n719) );
  AND2X2 AND2X2_610 ( .A(_abc_43815_n1350_bF_buf1), .B(_abc_43815_n1777), .Y(_abc_43815_n1778_1) );
  AND2X2 AND2X2_6100 ( .A(alu__abc_41358_n1253), .B(alu__abc_41358_n1254), .Y(alu__abc_41358_n1255) );
  AND2X2 AND2X2_6101 ( .A(alu__abc_41358_n962), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n1257) );
  AND2X2 AND2X2_6102 ( .A(alu__abc_41358_n919), .B(alu__abc_41358_n299_bF_buf6), .Y(alu__abc_41358_n1258) );
  AND2X2 AND2X2_6103 ( .A(alu__abc_41358_n1256), .B(alu__abc_41358_n1260), .Y(alu__abc_41358_n1261) );
  AND2X2 AND2X2_6104 ( .A(alu__abc_41358_n1262), .B(alu__abc_41358_n833_bF_buf0), .Y(alu__abc_41358_n1263) );
  AND2X2 AND2X2_6105 ( .A(alu__abc_41358_n1263), .B(alu__abc_41358_n1252), .Y(alu__abc_41358_n1264_1) );
  AND2X2 AND2X2_6106 ( .A(alu__abc_41358_n1266), .B(alu__abc_41358_n1057_bF_buf1), .Y(alu__abc_41358_n1267) );
  AND2X2 AND2X2_6107 ( .A(alu__abc_41358_n1267), .B(alu__abc_41358_n1265), .Y(alu__abc_41358_n1268) );
  AND2X2 AND2X2_6108 ( .A(alu__abc_41358_n761), .B(alu__abc_41358_n1061_bF_buf1), .Y(alu__abc_41358_n1269) );
  AND2X2 AND2X2_6109 ( .A(alu__abc_41358_n838), .B(alu__abc_41358_n843), .Y(alu__abc_41358_n1271) );
  AND2X2 AND2X2_611 ( .A(alu_op_r_6_), .B(pc_q_10_), .Y(_abc_43815_n1781_1) );
  AND2X2 AND2X2_6110 ( .A(alu__abc_41358_n1272), .B(alu__abc_41358_n1273), .Y(alu__abc_41358_n1274) );
  AND2X2 AND2X2_6111 ( .A(alu__abc_41358_n1275), .B(alu__abc_41358_n1270), .Y(alu__abc_41358_n1276) );
  AND2X2 AND2X2_6112 ( .A(alu__abc_41358_n1276), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n1277) );
  AND2X2 AND2X2_6113 ( .A(alu__abc_41358_n1277), .B(alu__abc_41358_n948_bF_buf0), .Y(alu__abc_41358_n1278) );
  AND2X2 AND2X2_6114 ( .A(alu__abc_41358_n932_bF_buf0), .B(alu_a_i_4_), .Y(alu__abc_41358_n1279) );
  AND2X2 AND2X2_6115 ( .A(alu__abc_41358_n935_bF_buf0), .B(alu__abc_41358_n277), .Y(alu__abc_41358_n1280) );
  AND2X2 AND2X2_6116 ( .A(alu__abc_41358_n277), .B(alu_op_i_0_bF_buf3), .Y(alu__abc_41358_n1281) );
  AND2X2 AND2X2_6117 ( .A(alu__abc_41358_n927_bF_buf4), .B(alu__abc_41358_n282), .Y(alu__abc_41358_n1283) );
  AND2X2 AND2X2_6118 ( .A(alu__abc_41358_n1283), .B(alu__abc_41358_n1282), .Y(alu__abc_41358_n1284_1) );
  AND2X2 AND2X2_6119 ( .A(alu__abc_41358_n1293), .B(alu__abc_41358_n942_bF_buf4), .Y(alu__abc_41358_n1294) );
  AND2X2 AND2X2_612 ( .A(_abc_43815_n1782), .B(_abc_43815_n1780), .Y(_abc_43815_n1783) );
  AND2X2 AND2X2_6120 ( .A(alu__abc_41358_n1294), .B(alu__abc_41358_n1292), .Y(alu__abc_41358_n1295) );
  AND2X2 AND2X2_6121 ( .A(alu__abc_41358_n285), .B(alu_op_i_0_bF_buf2), .Y(alu__abc_41358_n1296) );
  AND2X2 AND2X2_6122 ( .A(alu__abc_41358_n927_bF_buf3), .B(alu__abc_41358_n594), .Y(alu__abc_41358_n1298) );
  AND2X2 AND2X2_6123 ( .A(alu__abc_41358_n1298), .B(alu__abc_41358_n1297), .Y(alu__abc_41358_n1299) );
  AND2X2 AND2X2_6124 ( .A(alu__abc_41358_n740), .B(alu__abc_41358_n1061_bF_buf0), .Y(alu__abc_41358_n1300) );
  AND2X2 AND2X2_6125 ( .A(alu__abc_41358_n1075), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n1301) );
  AND2X2 AND2X2_6126 ( .A(alu__abc_41358_n1013), .B(alu__abc_41358_n1018), .Y(alu__abc_41358_n1302) );
  AND2X2 AND2X2_6127 ( .A(alu__abc_41358_n1303), .B(alu__abc_41358_n1304_1), .Y(alu__abc_41358_n1305) );
  AND2X2 AND2X2_6128 ( .A(alu__abc_41358_n1305), .B(alu__abc_41358_n299_bF_buf4), .Y(alu__abc_41358_n1306) );
  AND2X2 AND2X2_6129 ( .A(alu__abc_41358_n1307), .B(alu__abc_41358_n294_bF_buf6), .Y(alu__abc_41358_n1308) );
  AND2X2 AND2X2_613 ( .A(_abc_43815_n1784), .B(_abc_43815_n1746), .Y(_abc_43815_n1785_1) );
  AND2X2 AND2X2_6130 ( .A(alu__abc_41358_n1308), .B(alu__abc_41358_n948_bF_buf4), .Y(alu__abc_41358_n1309) );
  AND2X2 AND2X2_6131 ( .A(alu__abc_41358_n932_bF_buf4), .B(alu_a_i_5_), .Y(alu__abc_41358_n1310) );
  AND2X2 AND2X2_6132 ( .A(alu__abc_41358_n935_bF_buf4), .B(alu__abc_41358_n285), .Y(alu__abc_41358_n1311) );
  AND2X2 AND2X2_6133 ( .A(alu__abc_41358_n1265), .B(alu__abc_41358_n1318), .Y(alu__abc_41358_n1319) );
  AND2X2 AND2X2_6134 ( .A(alu__abc_41358_n1320), .B(alu__abc_41358_n1057_bF_buf0), .Y(alu__abc_41358_n1321) );
  AND2X2 AND2X2_6135 ( .A(alu__abc_41358_n1321), .B(alu__abc_41358_n1317), .Y(alu__abc_41358_n1322) );
  AND2X2 AND2X2_6136 ( .A(alu__abc_41358_n970), .B(alu__abc_41358_n299_bF_buf3), .Y(alu__abc_41358_n1323_1) );
  AND2X2 AND2X2_6137 ( .A(alu__abc_41358_n1324), .B(alu_b_i_3_bF_buf0), .Y(alu__abc_41358_n1325) );
  AND2X2 AND2X2_6138 ( .A(alu__abc_41358_n1326), .B(alu__abc_41358_n1327), .Y(alu__abc_41358_n1328) );
  AND2X2 AND2X2_6139 ( .A(alu__abc_41358_n1328), .B(alu__abc_41358_n294_bF_buf5), .Y(alu__abc_41358_n1329) );
  AND2X2 AND2X2_614 ( .A(_abc_43815_n1707), .B(_abc_43815_n1747), .Y(_abc_43815_n1787) );
  AND2X2 AND2X2_6140 ( .A(alu__abc_41358_n1026), .B(alu__abc_41358_n299_bF_buf1), .Y(alu__abc_41358_n1332) );
  AND2X2 AND2X2_6141 ( .A(alu__abc_41358_n1038), .B(alu_b_i_2_bF_buf2), .Y(alu__abc_41358_n1333) );
  AND2X2 AND2X2_6142 ( .A(alu__abc_41358_n1336), .B(alu__abc_41358_n1337), .Y(alu__abc_41358_n1338) );
  AND2X2 AND2X2_6143 ( .A(alu__abc_41358_n1339), .B(alu__abc_41358_n1335), .Y(alu__abc_41358_n1340) );
  AND2X2 AND2X2_6144 ( .A(alu__abc_41358_n1341), .B(alu__abc_41358_n833_bF_buf4), .Y(alu__abc_41358_n1342) );
  AND2X2 AND2X2_6145 ( .A(alu__abc_41358_n1331), .B(alu__abc_41358_n1342), .Y(alu__abc_41358_n1343) );
  AND2X2 AND2X2_6146 ( .A(alu__abc_41358_n1347), .B(alu__abc_41358_n1057_bF_buf4), .Y(alu__abc_41358_n1348) );
  AND2X2 AND2X2_6147 ( .A(alu__abc_41358_n1348), .B(alu__abc_41358_n1346), .Y(alu__abc_41358_n1349) );
  AND2X2 AND2X2_6148 ( .A(alu__abc_41358_n1350), .B(alu__abc_41358_n1351), .Y(alu__abc_41358_n1352) );
  AND2X2 AND2X2_6149 ( .A(alu__abc_41358_n1352), .B(alu__abc_41358_n942_bF_buf3), .Y(alu__abc_41358_n1353) );
  AND2X2 AND2X2_615 ( .A(_abc_43815_n1703), .B(_abc_43815_n1787), .Y(_abc_43815_n1788_1) );
  AND2X2 AND2X2_6150 ( .A(alu__abc_41358_n1088), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n1354) );
  AND2X2 AND2X2_6151 ( .A(alu__abc_41358_n1357), .B(alu__abc_41358_n1358), .Y(alu__abc_41358_n1359) );
  AND2X2 AND2X2_6152 ( .A(alu__abc_41358_n1356), .B(alu__abc_41358_n1360), .Y(alu__abc_41358_n1361) );
  AND2X2 AND2X2_6153 ( .A(alu__abc_41358_n1363), .B(alu__abc_41358_n1364), .Y(alu__abc_41358_n1365) );
  AND2X2 AND2X2_6154 ( .A(alu__abc_41358_n1367), .B(alu__abc_41358_n1368), .Y(alu__abc_41358_n1369) );
  AND2X2 AND2X2_6155 ( .A(alu__abc_41358_n1366), .B(alu__abc_41358_n1370), .Y(alu__abc_41358_n1371) );
  AND2X2 AND2X2_6156 ( .A(alu__abc_41358_n1372), .B(alu__abc_41358_n833_bF_buf3), .Y(alu__abc_41358_n1373) );
  AND2X2 AND2X2_6157 ( .A(alu__abc_41358_n1373), .B(alu__abc_41358_n1362_1), .Y(alu__abc_41358_n1374) );
  AND2X2 AND2X2_6158 ( .A(alu__abc_41358_n733), .B(alu__abc_41358_n1061_bF_buf4), .Y(alu__abc_41358_n1375) );
  AND2X2 AND2X2_6159 ( .A(alu__abc_41358_n844), .B(alu__abc_41358_n847_1), .Y(alu__abc_41358_n1376) );
  AND2X2 AND2X2_616 ( .A(_abc_43815_n1789), .B(_abc_43815_n1783), .Y(_abc_43815_n1790) );
  AND2X2 AND2X2_6160 ( .A(alu__abc_41358_n1377), .B(alu__abc_41358_n1378), .Y(alu__abc_41358_n1379) );
  AND2X2 AND2X2_6161 ( .A(alu__abc_41358_n1380), .B(alu__abc_41358_n1381), .Y(alu__abc_41358_n1382_1) );
  AND2X2 AND2X2_6162 ( .A(alu__abc_41358_n1382_1), .B(alu__abc_41358_n294_bF_buf1), .Y(alu__abc_41358_n1383) );
  AND2X2 AND2X2_6163 ( .A(alu__abc_41358_n1383), .B(alu__abc_41358_n948_bF_buf3), .Y(alu__abc_41358_n1384) );
  AND2X2 AND2X2_6164 ( .A(alu__abc_41358_n932_bF_buf3), .B(alu_a_i_6_), .Y(alu__abc_41358_n1385) );
  AND2X2 AND2X2_6165 ( .A(alu__abc_41358_n935_bF_buf3), .B(alu__abc_41358_n263), .Y(alu__abc_41358_n1386) );
  AND2X2 AND2X2_6166 ( .A(alu__abc_41358_n263), .B(alu_op_i_0_bF_buf1), .Y(alu__abc_41358_n1387) );
  AND2X2 AND2X2_6167 ( .A(alu__abc_41358_n927_bF_buf2), .B(alu__abc_41358_n268), .Y(alu__abc_41358_n1389) );
  AND2X2 AND2X2_6168 ( .A(alu__abc_41358_n1389), .B(alu__abc_41358_n1388), .Y(alu__abc_41358_n1390) );
  AND2X2 AND2X2_6169 ( .A(alu__abc_41358_n1347), .B(alu__abc_41358_n1399), .Y(alu__abc_41358_n1400) );
  AND2X2 AND2X2_617 ( .A(_abc_43815_n1791_1), .B(_abc_43815_n1792), .Y(_abc_43815_n1793) );
  AND2X2 AND2X2_6170 ( .A(alu__abc_41358_n1401_1), .B(alu__abc_41358_n1057_bF_buf3), .Y(alu__abc_41358_n1402) );
  AND2X2 AND2X2_6171 ( .A(alu__abc_41358_n1402), .B(alu__abc_41358_n1398), .Y(alu__abc_41358_n1403) );
  AND2X2 AND2X2_6172 ( .A(alu__abc_41358_n1405), .B(alu__abc_41358_n942_bF_buf2), .Y(alu__abc_41358_n1406) );
  AND2X2 AND2X2_6173 ( .A(alu__abc_41358_n1406), .B(alu__abc_41358_n1404), .Y(alu__abc_41358_n1407) );
  AND2X2 AND2X2_6174 ( .A(alu__abc_41358_n731), .B(alu__abc_41358_n1061_bF_buf3), .Y(alu__abc_41358_n1408) );
  AND2X2 AND2X2_6175 ( .A(alu__abc_41358_n1163), .B(alu__abc_41358_n299_bF_buf2), .Y(alu__abc_41358_n1409) );
  AND2X2 AND2X2_6176 ( .A(alu__abc_41358_n1412), .B(alu__abc_41358_n1413), .Y(alu__abc_41358_n1414) );
  AND2X2 AND2X2_6177 ( .A(alu__abc_41358_n1411), .B(alu__abc_41358_n1415), .Y(alu__abc_41358_n1416) );
  AND2X2 AND2X2_6178 ( .A(alu__abc_41358_n1418), .B(alu__abc_41358_n1419_1), .Y(alu__abc_41358_n1420) );
  AND2X2 AND2X2_6179 ( .A(alu__abc_41358_n1420), .B(alu_b_i_3_bF_buf2), .Y(alu__abc_41358_n1421) );
  AND2X2 AND2X2_618 ( .A(_abc_43815_n1431_1_bF_buf4), .B(_abc_43815_n1795), .Y(_abc_43815_n1796) );
  AND2X2 AND2X2_6180 ( .A(alu__abc_41358_n1422), .B(alu__abc_41358_n1423), .Y(alu__abc_41358_n1424) );
  AND2X2 AND2X2_6181 ( .A(alu__abc_41358_n1424), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n1425) );
  AND2X2 AND2X2_6182 ( .A(alu__abc_41358_n1427), .B(alu__abc_41358_n833_bF_buf2), .Y(alu__abc_41358_n1428) );
  AND2X2 AND2X2_6183 ( .A(alu__abc_41358_n1428), .B(alu__abc_41358_n1417), .Y(alu__abc_41358_n1429) );
  AND2X2 AND2X2_6184 ( .A(alu__abc_41358_n1222), .B(alu_b_i_2_bF_buf0), .Y(alu__abc_41358_n1430) );
  AND2X2 AND2X2_6185 ( .A(alu__abc_41358_n1019), .B(alu__abc_41358_n1022), .Y(alu__abc_41358_n1431) );
  AND2X2 AND2X2_6186 ( .A(alu__abc_41358_n1432), .B(alu__abc_41358_n1433), .Y(alu__abc_41358_n1434) );
  AND2X2 AND2X2_6187 ( .A(alu__abc_41358_n1434), .B(alu__abc_41358_n299_bF_buf6), .Y(alu__abc_41358_n1435_1) );
  AND2X2 AND2X2_6188 ( .A(alu__abc_41358_n1436), .B(alu__abc_41358_n294_bF_buf6), .Y(alu__abc_41358_n1437) );
  AND2X2 AND2X2_6189 ( .A(alu__abc_41358_n1437), .B(alu__abc_41358_n948_bF_buf2), .Y(alu__abc_41358_n1438) );
  AND2X2 AND2X2_619 ( .A(_abc_43815_n1794_1), .B(_abc_43815_n1796), .Y(_abc_43815_n1797_1) );
  AND2X2 AND2X2_6190 ( .A(alu__abc_41358_n932_bF_buf2), .B(alu_a_i_7_), .Y(alu__abc_41358_n1439) );
  AND2X2 AND2X2_6191 ( .A(alu__abc_41358_n935_bF_buf2), .B(alu__abc_41358_n271), .Y(alu__abc_41358_n1440) );
  AND2X2 AND2X2_6192 ( .A(alu__abc_41358_n271), .B(alu_op_i_0_bF_buf0), .Y(alu__abc_41358_n1441) );
  AND2X2 AND2X2_6193 ( .A(alu__abc_41358_n927_bF_buf1), .B(alu__abc_41358_n598), .Y(alu__abc_41358_n1443) );
  AND2X2 AND2X2_6194 ( .A(alu__abc_41358_n1443), .B(alu__abc_41358_n1442), .Y(alu__abc_41358_n1444) );
  AND2X2 AND2X2_6195 ( .A(alu__abc_41358_n429), .B(alu__abc_41358_n364), .Y(alu__abc_41358_n1452) );
  AND2X2 AND2X2_6196 ( .A(alu__abc_41358_n1454), .B(alu__abc_41358_n1057_bF_buf2), .Y(alu__abc_41358_n1455) );
  AND2X2 AND2X2_6197 ( .A(alu__abc_41358_n1455), .B(alu__abc_41358_n1453), .Y(alu__abc_41358_n1456) );
  AND2X2 AND2X2_6198 ( .A(alu__abc_41358_n1457), .B(alu__abc_41358_n1458), .Y(alu__abc_41358_n1459) );
  AND2X2 AND2X2_6199 ( .A(alu__abc_41358_n1459), .B(alu__abc_41358_n942_bF_buf1), .Y(alu__abc_41358_n1460) );
  AND2X2 AND2X2_62 ( .A(_abc_43815_n696), .B(\mem_dat_i[9] ), .Y(_abc_43815_n720) );
  AND2X2 AND2X2_620 ( .A(_abc_43815_n1428_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_43815_n1798) );
  AND2X2 AND2X2_6200 ( .A(alu__abc_41358_n718), .B(alu__abc_41358_n1061_bF_buf2), .Y(alu__abc_41358_n1461) );
  AND2X2 AND2X2_6201 ( .A(alu__abc_41358_n1462), .B(alu__abc_41358_n1463), .Y(alu__abc_41358_n1464) );
  AND2X2 AND2X2_6202 ( .A(alu__abc_41358_n1467), .B(alu__abc_41358_n1466), .Y(alu__abc_41358_n1468) );
  AND2X2 AND2X2_6203 ( .A(alu__abc_41358_n1469), .B(alu__abc_41358_n833_bF_buf1), .Y(alu__abc_41358_n1470) );
  AND2X2 AND2X2_6204 ( .A(alu__abc_41358_n1470), .B(alu__abc_41358_n1465), .Y(alu__abc_41358_n1471) );
  AND2X2 AND2X2_6205 ( .A(alu__abc_41358_n848), .B(alu__abc_41358_n855), .Y(alu__abc_41358_n1473) );
  AND2X2 AND2X2_6206 ( .A(alu__abc_41358_n1474), .B(alu__abc_41358_n1475), .Y(alu__abc_41358_n1476) );
  AND2X2 AND2X2_6207 ( .A(alu__abc_41358_n1477), .B(alu__abc_41358_n1478), .Y(alu__abc_41358_n1479) );
  AND2X2 AND2X2_6208 ( .A(alu__abc_41358_n1480), .B(alu__abc_41358_n1472), .Y(alu__abc_41358_n1481) );
  AND2X2 AND2X2_6209 ( .A(alu__abc_41358_n1481), .B(alu__abc_41358_n948_bF_buf1), .Y(alu__abc_41358_n1482) );
  AND2X2 AND2X2_621 ( .A(_abc_43815_n1800), .B(_abc_43815_n1801), .Y(_abc_43815_n1802_1) );
  AND2X2 AND2X2_6210 ( .A(alu__abc_41358_n932_bF_buf1), .B(alu_a_i_8_), .Y(alu__abc_41358_n1483) );
  AND2X2 AND2X2_6211 ( .A(alu__abc_41358_n935_bF_buf1), .B(alu__abc_41358_n357), .Y(alu__abc_41358_n1484) );
  AND2X2 AND2X2_6212 ( .A(alu__abc_41358_n357), .B(alu_op_i_0_bF_buf5), .Y(alu__abc_41358_n1485) );
  AND2X2 AND2X2_6213 ( .A(alu__abc_41358_n927_bF_buf0), .B(alu__abc_41358_n362), .Y(alu__abc_41358_n1487) );
  AND2X2 AND2X2_6214 ( .A(alu__abc_41358_n1487), .B(alu__abc_41358_n1486), .Y(alu__abc_41358_n1488) );
  AND2X2 AND2X2_6215 ( .A(alu__abc_41358_n1453), .B(alu__abc_41358_n434), .Y(alu__abc_41358_n1496) );
  AND2X2 AND2X2_6216 ( .A(alu__abc_41358_n1499), .B(alu__abc_41358_n1057_bF_buf1), .Y(alu__abc_41358_n1500) );
  AND2X2 AND2X2_6217 ( .A(alu__abc_41358_n1500), .B(alu__abc_41358_n1498), .Y(alu__abc_41358_n1501) );
  AND2X2 AND2X2_6218 ( .A(alu__abc_41358_n766), .B(alu__abc_41358_n787_1), .Y(alu__abc_41358_n1502) );
  AND2X2 AND2X2_6219 ( .A(alu__abc_41358_n1504), .B(alu__abc_41358_n942_bF_buf0), .Y(alu__abc_41358_n1505) );
  AND2X2 AND2X2_622 ( .A(_abc_43815_n1802_1), .B(_abc_43815_n1413_bF_buf4), .Y(_abc_43815_n1803) );
  AND2X2 AND2X2_6220 ( .A(alu__abc_41358_n1505), .B(alu__abc_41358_n1503), .Y(alu__abc_41358_n1506) );
  AND2X2 AND2X2_6221 ( .A(alu__abc_41358_n787_1), .B(alu__abc_41358_n1061_bF_buf1), .Y(alu__abc_41358_n1507) );
  AND2X2 AND2X2_6222 ( .A(alu__abc_41358_n962), .B(alu_b_i_3_bF_buf5), .Y(alu__abc_41358_n1508) );
  AND2X2 AND2X2_6223 ( .A(alu__abc_41358_n982), .B(alu__abc_41358_n294_bF_buf2), .Y(alu__abc_41358_n1509) );
  AND2X2 AND2X2_6224 ( .A(alu__abc_41358_n1004), .B(alu_b_i_3_bF_buf4), .Y(alu__abc_41358_n1512) );
  AND2X2 AND2X2_6225 ( .A(alu__abc_41358_n1050_1), .B(alu__abc_41358_n294_bF_buf1), .Y(alu__abc_41358_n1513) );
  AND2X2 AND2X2_6226 ( .A(alu__abc_41358_n1515), .B(alu__abc_41358_n833_bF_buf0), .Y(alu__abc_41358_n1516) );
  AND2X2 AND2X2_6227 ( .A(alu__abc_41358_n1511), .B(alu__abc_41358_n1516), .Y(alu__abc_41358_n1517) );
  AND2X2 AND2X2_6228 ( .A(alu__abc_41358_n1076), .B(alu_b_i_3_bF_buf3), .Y(alu__abc_41358_n1518) );
  AND2X2 AND2X2_6229 ( .A(alu__abc_41358_n1023), .B(alu__abc_41358_n1030), .Y(alu__abc_41358_n1519) );
  AND2X2 AND2X2_623 ( .A(_abc_43815_n1804), .B(_abc_43815_n1351_bF_buf1), .Y(_abc_43815_n1805) );
  AND2X2 AND2X2_6230 ( .A(alu__abc_41358_n1520), .B(alu__abc_41358_n1521), .Y(alu__abc_41358_n1522) );
  AND2X2 AND2X2_6231 ( .A(alu__abc_41358_n1523), .B(alu__abc_41358_n1524), .Y(alu__abc_41358_n1525) );
  AND2X2 AND2X2_6232 ( .A(alu__abc_41358_n1525), .B(alu__abc_41358_n294_bF_buf0), .Y(alu__abc_41358_n1526) );
  AND2X2 AND2X2_6233 ( .A(alu__abc_41358_n1527), .B(alu__abc_41358_n948_bF_buf0), .Y(alu__abc_41358_n1528) );
  AND2X2 AND2X2_6234 ( .A(alu__abc_41358_n932_bF_buf0), .B(alu_a_i_9_), .Y(alu__abc_41358_n1529) );
  AND2X2 AND2X2_6235 ( .A(alu__abc_41358_n365), .B(alu_op_i_0_bF_buf4), .Y(alu__abc_41358_n1530) );
  AND2X2 AND2X2_6236 ( .A(alu__abc_41358_n927_bF_buf4), .B(alu__abc_41358_n370), .Y(alu__abc_41358_n1532) );
  AND2X2 AND2X2_6237 ( .A(alu__abc_41358_n1532), .B(alu__abc_41358_n1531), .Y(alu__abc_41358_n1533) );
  AND2X2 AND2X2_6238 ( .A(alu__abc_41358_n935_bF_buf0), .B(alu__abc_41358_n365), .Y(alu__abc_41358_n1534) );
  AND2X2 AND2X2_6239 ( .A(alu__abc_41358_n429), .B(alu__abc_41358_n373), .Y(alu__abc_41358_n1542) );
  AND2X2 AND2X2_624 ( .A(_abc_43815_n1807), .B(enable_i_bF_buf5), .Y(_abc_43815_n1808) );
  AND2X2 AND2X2_6240 ( .A(alu__abc_41358_n1543), .B(alu__abc_41358_n347), .Y(alu__abc_41358_n1545) );
  AND2X2 AND2X2_6241 ( .A(alu__abc_41358_n1546), .B(alu__abc_41358_n1057_bF_buf0), .Y(alu__abc_41358_n1547) );
  AND2X2 AND2X2_6242 ( .A(alu__abc_41358_n1547), .B(alu__abc_41358_n1544), .Y(alu__abc_41358_n1548) );
  AND2X2 AND2X2_6243 ( .A(alu__abc_41358_n1502), .B(alu__abc_41358_n781), .Y(alu__abc_41358_n1549) );
  AND2X2 AND2X2_6244 ( .A(alu__abc_41358_n1551), .B(alu__abc_41358_n942_bF_buf4), .Y(alu__abc_41358_n1552) );
  AND2X2 AND2X2_6245 ( .A(alu__abc_41358_n1552), .B(alu__abc_41358_n1550), .Y(alu__abc_41358_n1553) );
  AND2X2 AND2X2_6246 ( .A(alu__abc_41358_n781), .B(alu__abc_41358_n1061_bF_buf0), .Y(alu__abc_41358_n1554) );
  AND2X2 AND2X2_6247 ( .A(alu__abc_41358_n1094), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n1555) );
  AND2X2 AND2X2_6248 ( .A(alu__abc_41358_n1558), .B(alu__abc_41358_n1559), .Y(alu__abc_41358_n1560) );
  AND2X2 AND2X2_6249 ( .A(alu__abc_41358_n1561), .B(alu__abc_41358_n833_bF_buf4), .Y(alu__abc_41358_n1562) );
  AND2X2 AND2X2_625 ( .A(_abc_43815_n1806), .B(_abc_43815_n1808), .Y(epc_q_10__FF_INPUT) );
  AND2X2 AND2X2_6250 ( .A(alu__abc_41358_n1562), .B(alu__abc_41358_n1557), .Y(alu__abc_41358_n1563) );
  AND2X2 AND2X2_6251 ( .A(alu__abc_41358_n1146), .B(alu_b_i_3_bF_buf1), .Y(alu__abc_41358_n1564) );
  AND2X2 AND2X2_6252 ( .A(alu__abc_41358_n856), .B(alu__abc_41358_n859), .Y(alu__abc_41358_n1565) );
  AND2X2 AND2X2_6253 ( .A(alu__abc_41358_n1566), .B(alu__abc_41358_n1567), .Y(alu__abc_41358_n1568) );
  AND2X2 AND2X2_6254 ( .A(alu__abc_41358_n1569), .B(alu__abc_41358_n1570), .Y(alu__abc_41358_n1571) );
  AND2X2 AND2X2_6255 ( .A(alu__abc_41358_n1571), .B(alu__abc_41358_n294_bF_buf5), .Y(alu__abc_41358_n1572) );
  AND2X2 AND2X2_6256 ( .A(alu__abc_41358_n1573), .B(alu__abc_41358_n948_bF_buf4), .Y(alu__abc_41358_n1574) );
  AND2X2 AND2X2_6257 ( .A(alu__abc_41358_n932_bF_buf4), .B(alu_a_i_10_), .Y(alu__abc_41358_n1575) );
  AND2X2 AND2X2_6258 ( .A(alu__abc_41358_n340), .B(alu_op_i_0_bF_buf3), .Y(alu__abc_41358_n1576) );
  AND2X2 AND2X2_6259 ( .A(alu__abc_41358_n927_bF_buf3), .B(alu__abc_41358_n345), .Y(alu__abc_41358_n1578) );
  AND2X2 AND2X2_626 ( .A(_abc_43815_n1770), .B(pc_q_11_), .Y(_abc_43815_n1811) );
  AND2X2 AND2X2_6260 ( .A(alu__abc_41358_n1578), .B(alu__abc_41358_n1577), .Y(alu__abc_41358_n1579) );
  AND2X2 AND2X2_6261 ( .A(alu__abc_41358_n935_bF_buf4), .B(alu__abc_41358_n340), .Y(alu__abc_41358_n1580) );
  AND2X2 AND2X2_6262 ( .A(alu__abc_41358_n1591), .B(alu__abc_41358_n1057_bF_buf4), .Y(alu__abc_41358_n1592) );
  AND2X2 AND2X2_6263 ( .A(alu__abc_41358_n1592), .B(alu__abc_41358_n1590), .Y(alu__abc_41358_n1593) );
  AND2X2 AND2X2_6264 ( .A(alu__abc_41358_n1549), .B(alu__abc_41358_n805), .Y(alu__abc_41358_n1595) );
  AND2X2 AND2X2_6265 ( .A(alu__abc_41358_n1596), .B(alu__abc_41358_n942_bF_buf3), .Y(alu__abc_41358_n1597) );
  AND2X2 AND2X2_6266 ( .A(alu__abc_41358_n1597), .B(alu__abc_41358_n1594), .Y(alu__abc_41358_n1598) );
  AND2X2 AND2X2_6267 ( .A(alu__abc_41358_n348), .B(alu_op_i_0_bF_buf2), .Y(alu__abc_41358_n1599) );
  AND2X2 AND2X2_6268 ( .A(alu__abc_41358_n927_bF_buf2), .B(alu__abc_41358_n353), .Y(alu__abc_41358_n1601) );
  AND2X2 AND2X2_6269 ( .A(alu__abc_41358_n1601), .B(alu__abc_41358_n1600), .Y(alu__abc_41358_n1602) );
  AND2X2 AND2X2_627 ( .A(_abc_43815_n1812), .B(_abc_43815_n1810_1), .Y(_abc_43815_n1813) );
  AND2X2 AND2X2_6270 ( .A(alu__abc_41358_n805), .B(alu__abc_41358_n1061_bF_buf4), .Y(alu__abc_41358_n1603) );
  AND2X2 AND2X2_6271 ( .A(alu__abc_41358_n1169), .B(alu__abc_41358_n294_bF_buf4), .Y(alu__abc_41358_n1604) );
  AND2X2 AND2X2_6272 ( .A(alu__abc_41358_n1607), .B(alu__abc_41358_n1608), .Y(alu__abc_41358_n1609) );
  AND2X2 AND2X2_6273 ( .A(alu__abc_41358_n1610), .B(alu__abc_41358_n833_bF_buf3), .Y(alu__abc_41358_n1611) );
  AND2X2 AND2X2_6274 ( .A(alu__abc_41358_n1611), .B(alu__abc_41358_n1606), .Y(alu__abc_41358_n1612) );
  AND2X2 AND2X2_6275 ( .A(alu__abc_41358_n1223_1), .B(alu_b_i_3_bF_buf6), .Y(alu__abc_41358_n1613) );
  AND2X2 AND2X2_6276 ( .A(alu__abc_41358_n1031), .B(alu__abc_41358_n1034), .Y(alu__abc_41358_n1614) );
  AND2X2 AND2X2_6277 ( .A(alu__abc_41358_n1615), .B(alu__abc_41358_n1616), .Y(alu__abc_41358_n1617) );
  AND2X2 AND2X2_6278 ( .A(alu__abc_41358_n1618), .B(alu__abc_41358_n1619), .Y(alu__abc_41358_n1620) );
  AND2X2 AND2X2_6279 ( .A(alu__abc_41358_n1620), .B(alu__abc_41358_n294_bF_buf2), .Y(alu__abc_41358_n1621) );
  AND2X2 AND2X2_628 ( .A(_abc_43815_n1692), .B(_abc_43815_n1814), .Y(_abc_43815_n1815_1) );
  AND2X2 AND2X2_6280 ( .A(alu__abc_41358_n1622), .B(alu__abc_41358_n948_bF_buf3), .Y(alu__abc_41358_n1623) );
  AND2X2 AND2X2_6281 ( .A(alu__abc_41358_n932_bF_buf3), .B(alu_a_i_11_), .Y(alu__abc_41358_n1624) );
  AND2X2 AND2X2_6282 ( .A(alu__abc_41358_n935_bF_buf3), .B(alu__abc_41358_n348), .Y(alu__abc_41358_n1625) );
  AND2X2 AND2X2_6283 ( .A(alu__abc_41358_n429), .B(alu__abc_41358_n374), .Y(alu__abc_41358_n1633) );
  AND2X2 AND2X2_6284 ( .A(alu__abc_41358_n1634), .B(alu__abc_41358_n312), .Y(alu__abc_41358_n1636) );
  AND2X2 AND2X2_6285 ( .A(alu__abc_41358_n1637), .B(alu__abc_41358_n1057_bF_buf3), .Y(alu__abc_41358_n1638) );
  AND2X2 AND2X2_6286 ( .A(alu__abc_41358_n1638), .B(alu__abc_41358_n1635), .Y(alu__abc_41358_n1639) );
  AND2X2 AND2X2_6287 ( .A(alu__abc_41358_n1595), .B(alu__abc_41358_n773), .Y(alu__abc_41358_n1640) );
  AND2X2 AND2X2_6288 ( .A(alu__abc_41358_n1642), .B(alu__abc_41358_n942_bF_buf2), .Y(alu__abc_41358_n1643) );
  AND2X2 AND2X2_6289 ( .A(alu__abc_41358_n1643), .B(alu__abc_41358_n1641), .Y(alu__abc_41358_n1644) );
  AND2X2 AND2X2_629 ( .A(_abc_43815_n1065_1_bF_buf0), .B(epc_q_11_), .Y(_abc_43815_n1817) );
  AND2X2 AND2X2_6290 ( .A(alu__abc_41358_n773), .B(alu__abc_41358_n1061_bF_buf3), .Y(alu__abc_41358_n1645) );
  AND2X2 AND2X2_6291 ( .A(alu__abc_41358_n1647), .B(alu__abc_41358_n279_bF_buf2), .Y(alu__abc_41358_n1648) );
  AND2X2 AND2X2_6292 ( .A(alu__abc_41358_n1648), .B(alu__abc_41358_n1646), .Y(alu__abc_41358_n1649) );
  AND2X2 AND2X2_6293 ( .A(alu__abc_41358_n1650), .B(alu__abc_41358_n1466), .Y(alu__abc_41358_n1651) );
  AND2X2 AND2X2_6294 ( .A(alu__abc_41358_n1651), .B(alu_b_i_4_bF_buf0), .Y(alu__abc_41358_n1652) );
  AND2X2 AND2X2_6295 ( .A(alu__abc_41358_n1653), .B(alu__abc_41358_n833_bF_buf2), .Y(alu__abc_41358_n1654) );
  AND2X2 AND2X2_6296 ( .A(alu__abc_41358_n860), .B(alu__abc_41358_n865), .Y(alu__abc_41358_n1656) );
  AND2X2 AND2X2_6297 ( .A(alu__abc_41358_n1657), .B(alu__abc_41358_n1658), .Y(alu__abc_41358_n1659) );
  AND2X2 AND2X2_6298 ( .A(alu__abc_41358_n1660), .B(alu__abc_41358_n1661), .Y(alu__abc_41358_n1662) );
  AND2X2 AND2X2_6299 ( .A(alu__abc_41358_n1663), .B(alu__abc_41358_n1655), .Y(alu__abc_41358_n1664) );
  AND2X2 AND2X2_63 ( .A(_abc_43815_n689), .B(\mem_dat_i[25] ), .Y(_abc_43815_n722) );
  AND2X2 AND2X2_630 ( .A(_abc_43815_n1791_1), .B(_abc_43815_n1782), .Y(_abc_43815_n1818) );
  AND2X2 AND2X2_6300 ( .A(alu__abc_41358_n1664), .B(alu__abc_41358_n948_bF_buf2), .Y(alu__abc_41358_n1665) );
  AND2X2 AND2X2_6301 ( .A(alu__abc_41358_n932_bF_buf2), .B(alu_a_i_12_), .Y(alu__abc_41358_n1666) );
  AND2X2 AND2X2_6302 ( .A(alu__abc_41358_n935_bF_buf2), .B(alu__abc_41358_n305), .Y(alu__abc_41358_n1667) );
  AND2X2 AND2X2_6303 ( .A(alu__abc_41358_n305), .B(alu_op_i_0_bF_buf1), .Y(alu__abc_41358_n1668) );
  AND2X2 AND2X2_6304 ( .A(alu__abc_41358_n927_bF_buf1), .B(alu__abc_41358_n310), .Y(alu__abc_41358_n1670) );
  AND2X2 AND2X2_6305 ( .A(alu__abc_41358_n1670), .B(alu__abc_41358_n1669), .Y(alu__abc_41358_n1671) );
  AND2X2 AND2X2_6306 ( .A(alu__abc_41358_n1637), .B(alu__abc_41358_n449), .Y(alu__abc_41358_n1679) );
  AND2X2 AND2X2_6307 ( .A(alu__abc_41358_n1682), .B(alu__abc_41358_n1057_bF_buf2), .Y(alu__abc_41358_n1683) );
  AND2X2 AND2X2_6308 ( .A(alu__abc_41358_n1683), .B(alu__abc_41358_n1680), .Y(alu__abc_41358_n1684) );
  AND2X2 AND2X2_6309 ( .A(alu__abc_41358_n1640), .B(alu__abc_41358_n796), .Y(alu__abc_41358_n1685) );
  AND2X2 AND2X2_631 ( .A(alu_op_r_7_), .B(pc_q_11_), .Y(_abc_43815_n1821) );
  AND2X2 AND2X2_6310 ( .A(alu__abc_41358_n1687), .B(alu__abc_41358_n942_bF_buf1), .Y(alu__abc_41358_n1688) );
  AND2X2 AND2X2_6311 ( .A(alu__abc_41358_n1688), .B(alu__abc_41358_n1686), .Y(alu__abc_41358_n1689) );
  AND2X2 AND2X2_6312 ( .A(alu__abc_41358_n796), .B(alu__abc_41358_n1061_bF_buf2), .Y(alu__abc_41358_n1690) );
  AND2X2 AND2X2_6313 ( .A(alu__abc_41358_n1692), .B(alu__abc_41358_n279_bF_buf1), .Y(alu__abc_41358_n1693) );
  AND2X2 AND2X2_6314 ( .A(alu__abc_41358_n1693), .B(alu__abc_41358_n1691), .Y(alu__abc_41358_n1694) );
  AND2X2 AND2X2_6315 ( .A(alu__abc_41358_n1324), .B(alu__abc_41358_n294_bF_buf6), .Y(alu__abc_41358_n1695) );
  AND2X2 AND2X2_6316 ( .A(alu__abc_41358_n1696), .B(alu_b_i_4_bF_buf4), .Y(alu__abc_41358_n1697) );
  AND2X2 AND2X2_6317 ( .A(alu__abc_41358_n1698), .B(alu__abc_41358_n833_bF_buf1), .Y(alu__abc_41358_n1699) );
  AND2X2 AND2X2_6318 ( .A(alu__abc_41358_n1035), .B(alu__abc_41358_n1040), .Y(alu__abc_41358_n1700) );
  AND2X2 AND2X2_6319 ( .A(alu__abc_41358_n1701), .B(alu__abc_41358_n1702), .Y(alu__abc_41358_n1703) );
  AND2X2 AND2X2_632 ( .A(_abc_43815_n1822), .B(_abc_43815_n1820_1), .Y(_abc_43815_n1823_1) );
  AND2X2 AND2X2_6320 ( .A(alu__abc_41358_n1704), .B(alu__abc_41358_n1705), .Y(alu__abc_41358_n1706) );
  AND2X2 AND2X2_6321 ( .A(alu__abc_41358_n1707), .B(alu__abc_41358_n1708), .Y(alu__abc_41358_n1709) );
  AND2X2 AND2X2_6322 ( .A(alu__abc_41358_n1709), .B(alu__abc_41358_n948_bF_buf1), .Y(alu__abc_41358_n1710) );
  AND2X2 AND2X2_6323 ( .A(alu__abc_41358_n932_bF_buf1), .B(alu_a_i_13_), .Y(alu__abc_41358_n1711) );
  AND2X2 AND2X2_6324 ( .A(alu__abc_41358_n935_bF_buf1), .B(alu__abc_41358_n313), .Y(alu__abc_41358_n1712) );
  AND2X2 AND2X2_6325 ( .A(alu__abc_41358_n313), .B(alu_op_i_0_bF_buf0), .Y(alu__abc_41358_n1713) );
  AND2X2 AND2X2_6326 ( .A(alu__abc_41358_n927_bF_buf0), .B(alu__abc_41358_n318), .Y(alu__abc_41358_n1715) );
  AND2X2 AND2X2_6327 ( .A(alu__abc_41358_n1715), .B(alu__abc_41358_n1714), .Y(alu__abc_41358_n1716) );
  AND2X2 AND2X2_6328 ( .A(alu__abc_41358_n1634), .B(alu__abc_41358_n321), .Y(alu__abc_41358_n1724) );
  AND2X2 AND2X2_6329 ( .A(alu__abc_41358_n1725), .B(alu__abc_41358_n329_1), .Y(alu__abc_41358_n1727) );
  AND2X2 AND2X2_633 ( .A(_abc_43815_n1826_1), .B(_abc_43815_n1425_1_bF_buf4), .Y(_abc_43815_n1827) );
  AND2X2 AND2X2_6330 ( .A(alu__abc_41358_n1728), .B(alu__abc_41358_n1057_bF_buf1), .Y(alu__abc_41358_n1729) );
  AND2X2 AND2X2_6331 ( .A(alu__abc_41358_n1729), .B(alu__abc_41358_n1726), .Y(alu__abc_41358_n1730) );
  AND2X2 AND2X2_6332 ( .A(alu__abc_41358_n796), .B(alu__abc_41358_n805), .Y(alu__abc_41358_n1732) );
  AND2X2 AND2X2_6333 ( .A(alu__abc_41358_n1732), .B(alu__abc_41358_n790), .Y(alu__abc_41358_n1733) );
  AND2X2 AND2X2_6334 ( .A(alu__abc_41358_n1733), .B(alu__abc_41358_n799), .Y(alu__abc_41358_n1734) );
  AND2X2 AND2X2_6335 ( .A(alu__abc_41358_n1735), .B(alu__abc_41358_n942_bF_buf0), .Y(alu__abc_41358_n1736) );
  AND2X2 AND2X2_6336 ( .A(alu__abc_41358_n799), .B(alu__abc_41358_n1061_bF_buf1), .Y(alu__abc_41358_n1737) );
  AND2X2 AND2X2_6337 ( .A(alu__abc_41358_n1731), .B(alu__abc_41358_n1738), .Y(alu__abc_41358_n1739) );
  AND2X2 AND2X2_6338 ( .A(alu__abc_41358_n1741), .B(alu__abc_41358_n279_bF_buf0), .Y(alu__abc_41358_n1742) );
  AND2X2 AND2X2_6339 ( .A(alu__abc_41358_n1742), .B(alu__abc_41358_n1740), .Y(alu__abc_41358_n1743) );
  AND2X2 AND2X2_634 ( .A(_abc_43815_n1827), .B(_abc_43815_n1824), .Y(_abc_43815_n1828) );
  AND2X2 AND2X2_6340 ( .A(alu__abc_41358_n1355), .B(alu__abc_41358_n294_bF_buf3), .Y(alu__abc_41358_n1744) );
  AND2X2 AND2X2_6341 ( .A(alu__abc_41358_n1745), .B(alu_b_i_4_bF_buf3), .Y(alu__abc_41358_n1746) );
  AND2X2 AND2X2_6342 ( .A(alu__abc_41358_n1747), .B(alu__abc_41358_n833_bF_buf0), .Y(alu__abc_41358_n1748) );
  AND2X2 AND2X2_6343 ( .A(alu__abc_41358_n866), .B(alu__abc_41358_n869), .Y(alu__abc_41358_n1749) );
  AND2X2 AND2X2_6344 ( .A(alu__abc_41358_n1750), .B(alu__abc_41358_n1751), .Y(alu__abc_41358_n1752) );
  AND2X2 AND2X2_6345 ( .A(alu__abc_41358_n1753), .B(alu__abc_41358_n1754), .Y(alu__abc_41358_n1755) );
  AND2X2 AND2X2_6346 ( .A(alu__abc_41358_n1756), .B(alu__abc_41358_n1757), .Y(alu__abc_41358_n1758) );
  AND2X2 AND2X2_6347 ( .A(alu__abc_41358_n1758), .B(alu__abc_41358_n948_bF_buf0), .Y(alu__abc_41358_n1759) );
  AND2X2 AND2X2_6348 ( .A(alu__abc_41358_n932_bF_buf0), .B(alu_a_i_14_), .Y(alu__abc_41358_n1760) );
  AND2X2 AND2X2_6349 ( .A(alu__abc_41358_n935_bF_buf0), .B(alu__abc_41358_n322), .Y(alu__abc_41358_n1761) );
  AND2X2 AND2X2_635 ( .A(_abc_43815_n1829_1), .B(_abc_43815_n1431_1_bF_buf3), .Y(_abc_43815_n1830) );
  AND2X2 AND2X2_6350 ( .A(alu__abc_41358_n322), .B(alu_op_i_0_bF_buf5), .Y(alu__abc_41358_n1762) );
  AND2X2 AND2X2_6351 ( .A(alu__abc_41358_n927_bF_buf4), .B(alu__abc_41358_n327), .Y(alu__abc_41358_n1764) );
  AND2X2 AND2X2_6352 ( .A(alu__abc_41358_n1764), .B(alu__abc_41358_n1763), .Y(alu__abc_41358_n1765) );
  AND2X2 AND2X2_6353 ( .A(alu__abc_41358_n1775), .B(alu__abc_41358_n1057_bF_buf0), .Y(alu__abc_41358_n1776) );
  AND2X2 AND2X2_6354 ( .A(alu__abc_41358_n1776), .B(alu__abc_41358_n1774), .Y(alu__abc_41358_n1777) );
  AND2X2 AND2X2_6355 ( .A(alu__abc_41358_n1734), .B(alu__abc_41358_n704_1), .Y(alu__abc_41358_n1778) );
  AND2X2 AND2X2_6356 ( .A(alu__abc_41358_n1780), .B(alu__abc_41358_n942_bF_buf4), .Y(alu__abc_41358_n1781) );
  AND2X2 AND2X2_6357 ( .A(alu__abc_41358_n1781), .B(alu__abc_41358_n1779), .Y(alu__abc_41358_n1782) );
  AND2X2 AND2X2_6358 ( .A(alu__abc_41358_n330), .B(alu_op_i_0_bF_buf4), .Y(alu__abc_41358_n1783) );
  AND2X2 AND2X2_6359 ( .A(alu__abc_41358_n927_bF_buf3), .B(alu__abc_41358_n335), .Y(alu__abc_41358_n1785) );
  AND2X2 AND2X2_636 ( .A(_abc_43815_n1428_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_43815_n1831) );
  AND2X2 AND2X2_6360 ( .A(alu__abc_41358_n1785), .B(alu__abc_41358_n1784), .Y(alu__abc_41358_n1786) );
  AND2X2 AND2X2_6361 ( .A(alu__abc_41358_n704_1), .B(alu__abc_41358_n1061_bF_buf0), .Y(alu__abc_41358_n1787) );
  AND2X2 AND2X2_6362 ( .A(alu__abc_41358_n1789), .B(alu__abc_41358_n279_bF_buf5), .Y(alu__abc_41358_n1790) );
  AND2X2 AND2X2_6363 ( .A(alu__abc_41358_n1790), .B(alu__abc_41358_n1788), .Y(alu__abc_41358_n1791) );
  AND2X2 AND2X2_6364 ( .A(alu__abc_41358_n1410), .B(alu__abc_41358_n294_bF_buf0), .Y(alu__abc_41358_n1792) );
  AND2X2 AND2X2_6365 ( .A(alu__abc_41358_n1793), .B(alu_b_i_4_bF_buf2), .Y(alu__abc_41358_n1794) );
  AND2X2 AND2X2_6366 ( .A(alu__abc_41358_n1795), .B(alu__abc_41358_n833_bF_buf4), .Y(alu__abc_41358_n1796) );
  AND2X2 AND2X2_6367 ( .A(alu__abc_41358_n1436), .B(alu_b_i_3_bF_buf4), .Y(alu__abc_41358_n1797) );
  AND2X2 AND2X2_6368 ( .A(alu__abc_41358_n1041), .B(alu__abc_41358_n1044), .Y(alu__abc_41358_n1798) );
  AND2X2 AND2X2_6369 ( .A(alu__abc_41358_n1799), .B(alu__abc_41358_n1800), .Y(alu__abc_41358_n1801) );
  AND2X2 AND2X2_637 ( .A(_abc_43815_n1833), .B(_abc_43815_n1816), .Y(_abc_43815_n1834) );
  AND2X2 AND2X2_6370 ( .A(alu__abc_41358_n1802), .B(alu__abc_41358_n1803), .Y(alu__abc_41358_n1804) );
  AND2X2 AND2X2_6371 ( .A(alu__abc_41358_n1804), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n1805) );
  AND2X2 AND2X2_6372 ( .A(alu__abc_41358_n1806), .B(alu__abc_41358_n948_bF_buf4), .Y(alu__abc_41358_n1807) );
  AND2X2 AND2X2_6373 ( .A(alu__abc_41358_n932_bF_buf4), .B(alu_a_i_15_), .Y(alu__abc_41358_n1808) );
  AND2X2 AND2X2_6374 ( .A(alu__abc_41358_n935_bF_buf4), .B(alu__abc_41358_n330), .Y(alu__abc_41358_n1809) );
  AND2X2 AND2X2_6375 ( .A(alu__abc_41358_n1778), .B(alu__abc_41358_n694), .Y(alu__abc_41358_n1818) );
  AND2X2 AND2X2_6376 ( .A(alu__abc_41358_n1819), .B(alu__abc_41358_n1817), .Y(alu__abc_41358_n1820) );
  AND2X2 AND2X2_6377 ( .A(alu__abc_41358_n1820), .B(alu__abc_41358_n942_bF_buf3), .Y(alu__abc_41358_n1821) );
  AND2X2 AND2X2_6378 ( .A(alu__abc_41358_n461), .B(alu__abc_41358_n237), .Y(alu__abc_41358_n1823) );
  AND2X2 AND2X2_6379 ( .A(alu__abc_41358_n1824), .B(alu__abc_41358_n1057_bF_buf4), .Y(alu__abc_41358_n1825) );
  AND2X2 AND2X2_638 ( .A(_abc_43815_n1489_bF_buf4), .B(epc_q_11_), .Y(_abc_43815_n1836) );
  AND2X2 AND2X2_6380 ( .A(alu__abc_41358_n1825), .B(alu__abc_41358_n1822), .Y(alu__abc_41358_n1826) );
  AND2X2 AND2X2_6381 ( .A(alu__abc_41358_n694), .B(alu__abc_41358_n1061_bF_buf4), .Y(alu__abc_41358_n1827) );
  AND2X2 AND2X2_6382 ( .A(alu__abc_41358_n1829), .B(alu__abc_41358_n833_bF_buf3), .Y(alu__abc_41358_n1830) );
  AND2X2 AND2X2_6383 ( .A(alu__abc_41358_n1828), .B(alu__abc_41358_n1830), .Y(alu__abc_41358_n1831) );
  AND2X2 AND2X2_6384 ( .A(alu__abc_41358_n1479), .B(alu_b_i_3_bF_buf3), .Y(alu__abc_41358_n1832) );
  AND2X2 AND2X2_6385 ( .A(alu__abc_41358_n870), .B(alu__abc_41358_n879), .Y(alu__abc_41358_n1835) );
  AND2X2 AND2X2_6386 ( .A(alu__abc_41358_n1834), .B(alu__abc_41358_n1836), .Y(alu__abc_41358_n1837) );
  AND2X2 AND2X2_6387 ( .A(alu__abc_41358_n1833), .B(alu__abc_41358_n1838), .Y(alu__abc_41358_n1839) );
  AND2X2 AND2X2_6388 ( .A(alu__abc_41358_n1839), .B(alu__abc_41358_n294_bF_buf6), .Y(alu__abc_41358_n1840) );
  AND2X2 AND2X2_6389 ( .A(alu__abc_41358_n1841), .B(alu__abc_41358_n948_bF_buf3), .Y(alu__abc_41358_n1842) );
  AND2X2 AND2X2_639 ( .A(_abc_43815_n1418_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_43815_n1837) );
  AND2X2 AND2X2_6390 ( .A(alu__abc_41358_n932_bF_buf3), .B(alu_a_i_16_), .Y(alu__abc_41358_n1843) );
  AND2X2 AND2X2_6391 ( .A(alu__abc_41358_n935_bF_buf3), .B(alu__abc_41358_n230), .Y(alu__abc_41358_n1844) );
  AND2X2 AND2X2_6392 ( .A(alu__abc_41358_n230), .B(alu_op_i_0_bF_buf3), .Y(alu__abc_41358_n1845) );
  AND2X2 AND2X2_6393 ( .A(alu__abc_41358_n927_bF_buf2), .B(alu__abc_41358_n235), .Y(alu__abc_41358_n1847) );
  AND2X2 AND2X2_6394 ( .A(alu__abc_41358_n1847), .B(alu__abc_41358_n1846), .Y(alu__abc_41358_n1848) );
  AND2X2 AND2X2_6395 ( .A(alu__abc_41358_n947), .B(alu_b_i_4_bF_buf0), .Y(alu__abc_41358_n1850) );
  AND2X2 AND2X2_6396 ( .A(alu__abc_41358_n951), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n1851) );
  AND2X2 AND2X2_6397 ( .A(alu__abc_41358_n1824), .B(alu__abc_41358_n466), .Y(alu__abc_41358_n1859) );
  AND2X2 AND2X2_6398 ( .A(alu__abc_41358_n1862), .B(alu__abc_41358_n1057_bF_buf3), .Y(alu__abc_41358_n1863) );
  AND2X2 AND2X2_6399 ( .A(alu__abc_41358_n1863), .B(alu__abc_41358_n1861), .Y(alu__abc_41358_n1864) );
  AND2X2 AND2X2_64 ( .A(_abc_43815_n704), .B(\mem_dat_i[17] ), .Y(_abc_43815_n723) );
  AND2X2 AND2X2_640 ( .A(_abc_43815_n1839), .B(_abc_43815_n1351_bF_buf0), .Y(_abc_43815_n1840) );
  AND2X2 AND2X2_6400 ( .A(alu__abc_41358_n1866), .B(alu__abc_41358_n942_bF_buf2), .Y(alu__abc_41358_n1867) );
  AND2X2 AND2X2_6401 ( .A(alu__abc_41358_n1867), .B(alu__abc_41358_n1865), .Y(alu__abc_41358_n1868) );
  AND2X2 AND2X2_6402 ( .A(alu__abc_41358_n692), .B(alu__abc_41358_n1061_bF_buf3), .Y(alu__abc_41358_n1869) );
  AND2X2 AND2X2_6403 ( .A(alu__abc_41358_n1006), .B(alu__abc_41358_n279_bF_buf3), .Y(alu__abc_41358_n1870) );
  AND2X2 AND2X2_6404 ( .A(alu__abc_41358_n962), .B(alu_b_i_4_bF_buf4), .Y(alu__abc_41358_n1871) );
  AND2X2 AND2X2_6405 ( .A(alu__abc_41358_n1872), .B(alu__abc_41358_n833_bF_buf2), .Y(alu__abc_41358_n1873) );
  AND2X2 AND2X2_6406 ( .A(alu__abc_41358_n1045), .B(alu__abc_41358_n984), .Y(alu__abc_41358_n1874) );
  AND2X2 AND2X2_6407 ( .A(alu__abc_41358_n1875), .B(alu__abc_41358_n1876), .Y(alu__abc_41358_n1877) );
  AND2X2 AND2X2_6408 ( .A(alu__abc_41358_n1878), .B(alu__abc_41358_n1879), .Y(alu__abc_41358_n1880) );
  AND2X2 AND2X2_6409 ( .A(alu__abc_41358_n1880), .B(alu__abc_41358_n294_bF_buf5), .Y(alu__abc_41358_n1881) );
  AND2X2 AND2X2_641 ( .A(_abc_43815_n1835_1), .B(_abc_43815_n1840), .Y(_abc_43815_n1841_1) );
  AND2X2 AND2X2_6410 ( .A(alu__abc_41358_n1525), .B(alu_b_i_3_bF_buf2), .Y(alu__abc_41358_n1882) );
  AND2X2 AND2X2_6411 ( .A(alu__abc_41358_n1884), .B(alu__abc_41358_n1885), .Y(alu__abc_41358_n1886) );
  AND2X2 AND2X2_6412 ( .A(alu__abc_41358_n1886), .B(alu__abc_41358_n947), .Y(alu__abc_41358_n1887) );
  AND2X2 AND2X2_6413 ( .A(alu__abc_41358_n932_bF_buf2), .B(alu_a_i_17_), .Y(alu__abc_41358_n1888) );
  AND2X2 AND2X2_6414 ( .A(alu__abc_41358_n935_bF_buf2), .B(alu__abc_41358_n238), .Y(alu__abc_41358_n1889) );
  AND2X2 AND2X2_6415 ( .A(alu__abc_41358_n238), .B(alu_op_i_0_bF_buf2), .Y(alu__abc_41358_n1890) );
  AND2X2 AND2X2_6416 ( .A(alu__abc_41358_n927_bF_buf1), .B(alu__abc_41358_n243), .Y(alu__abc_41358_n1892) );
  AND2X2 AND2X2_6417 ( .A(alu__abc_41358_n1892), .B(alu__abc_41358_n1891), .Y(alu__abc_41358_n1893) );
  AND2X2 AND2X2_6418 ( .A(alu__abc_41358_n692), .B(alu__abc_41358_n685), .Y(alu__abc_41358_n1901) );
  AND2X2 AND2X2_6419 ( .A(alu__abc_41358_n1818), .B(alu__abc_41358_n1901), .Y(alu__abc_41358_n1902) );
  AND2X2 AND2X2_642 ( .A(_abc_43815_n1843), .B(enable_i_bF_buf4), .Y(_abc_43815_n1844_1) );
  AND2X2 AND2X2_6420 ( .A(alu__abc_41358_n1904), .B(alu__abc_41358_n942_bF_buf1), .Y(alu__abc_41358_n1905) );
  AND2X2 AND2X2_6421 ( .A(alu__abc_41358_n1905), .B(alu__abc_41358_n1903), .Y(alu__abc_41358_n1906) );
  AND2X2 AND2X2_6422 ( .A(alu__abc_41358_n461), .B(alu__abc_41358_n246), .Y(alu__abc_41358_n1907) );
  AND2X2 AND2X2_6423 ( .A(alu__abc_41358_n1908), .B(alu__abc_41358_n220), .Y(alu__abc_41358_n1910) );
  AND2X2 AND2X2_6424 ( .A(alu__abc_41358_n1911), .B(alu__abc_41358_n1057_bF_buf2), .Y(alu__abc_41358_n1912) );
  AND2X2 AND2X2_6425 ( .A(alu__abc_41358_n1912), .B(alu__abc_41358_n1909), .Y(alu__abc_41358_n1913) );
  AND2X2 AND2X2_6426 ( .A(alu__abc_41358_n685), .B(alu__abc_41358_n1061_bF_buf2), .Y(alu__abc_41358_n1914) );
  AND2X2 AND2X2_6427 ( .A(alu__abc_41358_n1106), .B(alu__abc_41358_n279_bF_buf1), .Y(alu__abc_41358_n1915) );
  AND2X2 AND2X2_6428 ( .A(alu__abc_41358_n1916), .B(alu__abc_41358_n833_bF_buf1), .Y(alu__abc_41358_n1917) );
  AND2X2 AND2X2_6429 ( .A(alu__abc_41358_n880), .B(alu__abc_41358_n883), .Y(alu__abc_41358_n1918) );
  AND2X2 AND2X2_643 ( .A(_abc_43815_n1842), .B(_abc_43815_n1844_1), .Y(epc_q_11__FF_INPUT) );
  AND2X2 AND2X2_6430 ( .A(alu__abc_41358_n1919), .B(alu__abc_41358_n1920), .Y(alu__abc_41358_n1921) );
  AND2X2 AND2X2_6431 ( .A(alu__abc_41358_n1922), .B(alu__abc_41358_n1923), .Y(alu__abc_41358_n1924) );
  AND2X2 AND2X2_6432 ( .A(alu__abc_41358_n1924), .B(alu__abc_41358_n294_bF_buf4), .Y(alu__abc_41358_n1925) );
  AND2X2 AND2X2_6433 ( .A(alu__abc_41358_n1571), .B(alu_b_i_3_bF_buf1), .Y(alu__abc_41358_n1926) );
  AND2X2 AND2X2_6434 ( .A(alu__abc_41358_n1929), .B(alu__abc_41358_n947), .Y(alu__abc_41358_n1930) );
  AND2X2 AND2X2_6435 ( .A(alu__abc_41358_n1928), .B(alu__abc_41358_n1930), .Y(alu__abc_41358_n1931) );
  AND2X2 AND2X2_6436 ( .A(alu__abc_41358_n932_bF_buf1), .B(alu_a_i_18_), .Y(alu__abc_41358_n1932) );
  AND2X2 AND2X2_6437 ( .A(alu__abc_41358_n935_bF_buf1), .B(alu__abc_41358_n213), .Y(alu__abc_41358_n1933) );
  AND2X2 AND2X2_6438 ( .A(alu__abc_41358_n213), .B(alu_op_i_0_bF_buf1), .Y(alu__abc_41358_n1934) );
  AND2X2 AND2X2_6439 ( .A(alu__abc_41358_n927_bF_buf0), .B(alu__abc_41358_n218), .Y(alu__abc_41358_n1936) );
  AND2X2 AND2X2_644 ( .A(_abc_43815_n1811), .B(pc_q_12_), .Y(_abc_43815_n1847_1) );
  AND2X2 AND2X2_6440 ( .A(alu__abc_41358_n1936), .B(alu__abc_41358_n1935), .Y(alu__abc_41358_n1937) );
  AND2X2 AND2X2_6441 ( .A(alu__abc_41358_n1948), .B(alu__abc_41358_n1057_bF_buf1), .Y(alu__abc_41358_n1949) );
  AND2X2 AND2X2_6442 ( .A(alu__abc_41358_n1949), .B(alu__abc_41358_n1946), .Y(alu__abc_41358_n1950) );
  AND2X2 AND2X2_6443 ( .A(alu__abc_41358_n1902), .B(alu__abc_41358_n683), .Y(alu__abc_41358_n1952) );
  AND2X2 AND2X2_6444 ( .A(alu__abc_41358_n1953), .B(alu__abc_41358_n1951), .Y(alu__abc_41358_n1954) );
  AND2X2 AND2X2_6445 ( .A(alu__abc_41358_n1954), .B(alu__abc_41358_n942_bF_buf0), .Y(alu__abc_41358_n1955) );
  AND2X2 AND2X2_6446 ( .A(alu__abc_41358_n683), .B(alu__abc_41358_n1061_bF_buf1), .Y(alu__abc_41358_n1956) );
  AND2X2 AND2X2_6447 ( .A(alu__abc_41358_n1181_1), .B(alu__abc_41358_n279_bF_buf5), .Y(alu__abc_41358_n1957) );
  AND2X2 AND2X2_6448 ( .A(alu__abc_41358_n1958), .B(alu__abc_41358_n833_bF_buf0), .Y(alu__abc_41358_n1959) );
  AND2X2 AND2X2_6449 ( .A(alu__abc_41358_n985), .B(alu__abc_41358_n988), .Y(alu__abc_41358_n1960) );
  AND2X2 AND2X2_645 ( .A(_abc_43815_n1848), .B(_abc_43815_n1846), .Y(_abc_43815_n1849) );
  AND2X2 AND2X2_6450 ( .A(alu__abc_41358_n1961), .B(alu__abc_41358_n1962), .Y(alu__abc_41358_n1963) );
  AND2X2 AND2X2_6451 ( .A(alu__abc_41358_n1964), .B(alu__abc_41358_n1965), .Y(alu__abc_41358_n1966) );
  AND2X2 AND2X2_6452 ( .A(alu__abc_41358_n1966), .B(alu__abc_41358_n294_bF_buf3), .Y(alu__abc_41358_n1967) );
  AND2X2 AND2X2_6453 ( .A(alu__abc_41358_n1620), .B(alu_b_i_3_bF_buf0), .Y(alu__abc_41358_n1968) );
  AND2X2 AND2X2_6454 ( .A(alu__abc_41358_n1971), .B(alu__abc_41358_n947), .Y(alu__abc_41358_n1972) );
  AND2X2 AND2X2_6455 ( .A(alu__abc_41358_n1970), .B(alu__abc_41358_n1972), .Y(alu__abc_41358_n1973) );
  AND2X2 AND2X2_6456 ( .A(alu__abc_41358_n932_bF_buf0), .B(alu_a_i_19_), .Y(alu__abc_41358_n1974) );
  AND2X2 AND2X2_6457 ( .A(alu__abc_41358_n935_bF_buf0), .B(alu__abc_41358_n221), .Y(alu__abc_41358_n1975) );
  AND2X2 AND2X2_6458 ( .A(alu__abc_41358_n221), .B(alu_op_i_0_bF_buf0), .Y(alu__abc_41358_n1976) );
  AND2X2 AND2X2_6459 ( .A(alu__abc_41358_n927_bF_buf4), .B(alu__abc_41358_n226), .Y(alu__abc_41358_n1978) );
  AND2X2 AND2X2_646 ( .A(_abc_43815_n1692), .B(_abc_43815_n1850_1), .Y(_abc_43815_n1851) );
  AND2X2 AND2X2_6460 ( .A(alu__abc_41358_n1978), .B(alu__abc_41358_n1977), .Y(alu__abc_41358_n1979) );
  AND2X2 AND2X2_6461 ( .A(alu__abc_41358_n1952), .B(alu__abc_41358_n676), .Y(alu__abc_41358_n1988) );
  AND2X2 AND2X2_6462 ( .A(alu__abc_41358_n1989), .B(alu__abc_41358_n1987), .Y(alu__abc_41358_n1990) );
  AND2X2 AND2X2_6463 ( .A(alu__abc_41358_n1990), .B(alu__abc_41358_n942_bF_buf4), .Y(alu__abc_41358_n1991) );
  AND2X2 AND2X2_6464 ( .A(alu__abc_41358_n461), .B(alu__abc_41358_n247), .Y(alu__abc_41358_n1992) );
  AND2X2 AND2X2_6465 ( .A(alu__abc_41358_n1993), .B(alu__abc_41358_n202), .Y(alu__abc_41358_n1994) );
  AND2X2 AND2X2_6466 ( .A(alu__abc_41358_n1996), .B(alu__abc_41358_n1057_bF_buf0), .Y(alu__abc_41358_n1997) );
  AND2X2 AND2X2_6467 ( .A(alu__abc_41358_n1997), .B(alu__abc_41358_n1995), .Y(alu__abc_41358_n1998) );
  AND2X2 AND2X2_6468 ( .A(alu__abc_41358_n676), .B(alu__abc_41358_n1061_bF_buf0), .Y(alu__abc_41358_n1999) );
  AND2X2 AND2X2_6469 ( .A(alu__abc_41358_n2000), .B(alu__abc_41358_n1830), .Y(alu__abc_41358_n2001) );
  AND2X2 AND2X2_647 ( .A(_abc_43815_n1418_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_43815_n1852) );
  AND2X2 AND2X2_6470 ( .A(alu__abc_41358_n1662), .B(alu_b_i_3_bF_buf6), .Y(alu__abc_41358_n2002) );
  AND2X2 AND2X2_6471 ( .A(alu__abc_41358_n884), .B(alu__abc_41358_n889), .Y(alu__abc_41358_n2005) );
  AND2X2 AND2X2_6472 ( .A(alu__abc_41358_n2004), .B(alu__abc_41358_n2006), .Y(alu__abc_41358_n2007) );
  AND2X2 AND2X2_6473 ( .A(alu__abc_41358_n2003), .B(alu__abc_41358_n2008), .Y(alu__abc_41358_n2009) );
  AND2X2 AND2X2_6474 ( .A(alu__abc_41358_n2009), .B(alu__abc_41358_n294_bF_buf2), .Y(alu__abc_41358_n2010) );
  AND2X2 AND2X2_6475 ( .A(alu__abc_41358_n2011), .B(alu__abc_41358_n948_bF_buf2), .Y(alu__abc_41358_n2012) );
  AND2X2 AND2X2_6476 ( .A(alu__abc_41358_n1277), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n2013) );
  AND2X2 AND2X2_6477 ( .A(alu__abc_41358_n932_bF_buf4), .B(alu_a_i_20_), .Y(alu__abc_41358_n2014) );
  AND2X2 AND2X2_6478 ( .A(alu__abc_41358_n195), .B(alu_op_i_0_bF_buf5), .Y(alu__abc_41358_n2015) );
  AND2X2 AND2X2_6479 ( .A(alu__abc_41358_n927_bF_buf3), .B(alu__abc_41358_n200), .Y(alu__abc_41358_n2017) );
  AND2X2 AND2X2_648 ( .A(_abc_43815_n1489_bF_buf3), .B(epc_q_12_), .Y(_abc_43815_n1853_1) );
  AND2X2 AND2X2_6480 ( .A(alu__abc_41358_n2017), .B(alu__abc_41358_n2016), .Y(alu__abc_41358_n2018) );
  AND2X2 AND2X2_6481 ( .A(alu__abc_41358_n935_bF_buf4), .B(alu__abc_41358_n195), .Y(alu__abc_41358_n2019) );
  AND2X2 AND2X2_6482 ( .A(alu__abc_41358_n1988), .B(alu__abc_41358_n820), .Y(alu__abc_41358_n2029) );
  AND2X2 AND2X2_6483 ( .A(alu__abc_41358_n2030), .B(alu__abc_41358_n2028), .Y(alu__abc_41358_n2031) );
  AND2X2 AND2X2_6484 ( .A(alu__abc_41358_n2031), .B(alu__abc_41358_n942_bF_buf3), .Y(alu__abc_41358_n2032) );
  AND2X2 AND2X2_6485 ( .A(alu__abc_41358_n1995), .B(alu__abc_41358_n481), .Y(alu__abc_41358_n2033) );
  AND2X2 AND2X2_6486 ( .A(alu__abc_41358_n2036), .B(alu__abc_41358_n1057_bF_buf4), .Y(alu__abc_41358_n2037) );
  AND2X2 AND2X2_6487 ( .A(alu__abc_41358_n2037), .B(alu__abc_41358_n2035), .Y(alu__abc_41358_n2038) );
  AND2X2 AND2X2_6488 ( .A(alu__abc_41358_n820), .B(alu__abc_41358_n1061_bF_buf4), .Y(alu__abc_41358_n2039) );
  AND2X2 AND2X2_6489 ( .A(alu__abc_41358_n1330), .B(alu__abc_41358_n279_bF_buf3), .Y(alu__abc_41358_n2040) );
  AND2X2 AND2X2_649 ( .A(_abc_43815_n1350_bF_buf4), .B(_abc_43815_n1854), .Y(_abc_43815_n1855) );
  AND2X2 AND2X2_6490 ( .A(alu__abc_41358_n2041), .B(alu__abc_41358_n833_bF_buf4), .Y(alu__abc_41358_n2042) );
  AND2X2 AND2X2_6491 ( .A(alu__abc_41358_n989), .B(alu__abc_41358_n994), .Y(alu__abc_41358_n2045) );
  AND2X2 AND2X2_6492 ( .A(alu__abc_41358_n2046), .B(alu__abc_41358_n2047), .Y(alu__abc_41358_n2048) );
  AND2X2 AND2X2_6493 ( .A(alu__abc_41358_n2049), .B(alu__abc_41358_n2050), .Y(alu__abc_41358_n2051) );
  AND2X2 AND2X2_6494 ( .A(alu__abc_41358_n2053), .B(alu__abc_41358_n947), .Y(alu__abc_41358_n2054) );
  AND2X2 AND2X2_6495 ( .A(alu__abc_41358_n2054), .B(alu__abc_41358_n2044), .Y(alu__abc_41358_n2055) );
  AND2X2 AND2X2_6496 ( .A(alu__abc_41358_n2055), .B(alu__abc_41358_n2043), .Y(alu__abc_41358_n2056) );
  AND2X2 AND2X2_6497 ( .A(alu__abc_41358_n932_bF_buf3), .B(alu_a_i_21_), .Y(alu__abc_41358_n2057) );
  AND2X2 AND2X2_6498 ( .A(alu__abc_41358_n203_1), .B(alu_op_i_0_bF_buf4), .Y(alu__abc_41358_n2058) );
  AND2X2 AND2X2_6499 ( .A(alu__abc_41358_n927_bF_buf2), .B(alu__abc_41358_n208), .Y(alu__abc_41358_n2060) );
  AND2X2 AND2X2_65 ( .A(_abc_43815_n726), .B(state_q_1_bF_buf0), .Y(_abc_43815_n727) );
  AND2X2 AND2X2_650 ( .A(_abc_43815_n1783), .B(_abc_43815_n1823_1), .Y(_abc_43815_n1857) );
  AND2X2 AND2X2_6500 ( .A(alu__abc_41358_n2060), .B(alu__abc_41358_n2059), .Y(alu__abc_41358_n2061) );
  AND2X2 AND2X2_6501 ( .A(alu__abc_41358_n935_bF_buf3), .B(alu__abc_41358_n203_1), .Y(alu__abc_41358_n2062) );
  AND2X2 AND2X2_6502 ( .A(alu__abc_41358_n2029), .B(alu__abc_41358_n672), .Y(alu__abc_41358_n2071) );
  AND2X2 AND2X2_6503 ( .A(alu__abc_41358_n2072), .B(alu__abc_41358_n2070), .Y(alu__abc_41358_n2073) );
  AND2X2 AND2X2_6504 ( .A(alu__abc_41358_n2073), .B(alu__abc_41358_n942_bF_buf2), .Y(alu__abc_41358_n2074) );
  AND2X2 AND2X2_6505 ( .A(alu__abc_41358_n1993), .B(alu__abc_41358_n211), .Y(alu__abc_41358_n2075) );
  AND2X2 AND2X2_6506 ( .A(alu__abc_41358_n2076), .B(alu__abc_41358_n185), .Y(alu__abc_41358_n2078) );
  AND2X2 AND2X2_6507 ( .A(alu__abc_41358_n2079), .B(alu__abc_41358_n1057_bF_buf3), .Y(alu__abc_41358_n2080) );
  AND2X2 AND2X2_6508 ( .A(alu__abc_41358_n2080), .B(alu__abc_41358_n2077), .Y(alu__abc_41358_n2081) );
  AND2X2 AND2X2_6509 ( .A(alu__abc_41358_n1361), .B(alu__abc_41358_n279_bF_buf1), .Y(alu__abc_41358_n2082) );
  AND2X2 AND2X2_651 ( .A(_abc_43815_n1787), .B(_abc_43815_n1857), .Y(_abc_43815_n1858) );
  AND2X2 AND2X2_6510 ( .A(alu__abc_41358_n2083), .B(alu__abc_41358_n833_bF_buf3), .Y(alu__abc_41358_n2084) );
  AND2X2 AND2X2_6511 ( .A(alu__abc_41358_n890), .B(alu__abc_41358_n893), .Y(alu__abc_41358_n2085) );
  AND2X2 AND2X2_6512 ( .A(alu__abc_41358_n2086), .B(alu__abc_41358_n2087), .Y(alu__abc_41358_n2088) );
  AND2X2 AND2X2_6513 ( .A(alu__abc_41358_n2089), .B(alu__abc_41358_n2090), .Y(alu__abc_41358_n2091) );
  AND2X2 AND2X2_6514 ( .A(alu__abc_41358_n2091), .B(alu__abc_41358_n294_bF_buf0), .Y(alu__abc_41358_n2092) );
  AND2X2 AND2X2_6515 ( .A(alu__abc_41358_n1755), .B(alu_b_i_3_bF_buf4), .Y(alu__abc_41358_n2093) );
  AND2X2 AND2X2_6516 ( .A(alu__abc_41358_n2096), .B(alu__abc_41358_n947), .Y(alu__abc_41358_n2097) );
  AND2X2 AND2X2_6517 ( .A(alu__abc_41358_n2095), .B(alu__abc_41358_n2097), .Y(alu__abc_41358_n2098) );
  AND2X2 AND2X2_6518 ( .A(alu__abc_41358_n932_bF_buf2), .B(alu_a_i_22_), .Y(alu__abc_41358_n2099) );
  AND2X2 AND2X2_6519 ( .A(alu__abc_41358_n935_bF_buf2), .B(alu__abc_41358_n178_1), .Y(alu__abc_41358_n2100) );
  AND2X2 AND2X2_652 ( .A(_abc_43815_n1703), .B(_abc_43815_n1858), .Y(_abc_43815_n1859_1) );
  AND2X2 AND2X2_6520 ( .A(alu__abc_41358_n178_1), .B(alu_op_i_0_bF_buf3), .Y(alu__abc_41358_n2101) );
  AND2X2 AND2X2_6521 ( .A(alu__abc_41358_n927_bF_buf1), .B(alu__abc_41358_n183_1), .Y(alu__abc_41358_n2103) );
  AND2X2 AND2X2_6522 ( .A(alu__abc_41358_n2103), .B(alu__abc_41358_n2102), .Y(alu__abc_41358_n2104) );
  AND2X2 AND2X2_6523 ( .A(alu__abc_41358_n672), .B(alu__abc_41358_n1061_bF_buf3), .Y(alu__abc_41358_n2109) );
  AND2X2 AND2X2_6524 ( .A(alu__abc_41358_n2071), .B(alu__abc_41358_n649), .Y(alu__abc_41358_n2114) );
  AND2X2 AND2X2_6525 ( .A(alu__abc_41358_n2115), .B(alu__abc_41358_n2113), .Y(alu__abc_41358_n2116) );
  AND2X2 AND2X2_6526 ( .A(alu__abc_41358_n2116), .B(alu__abc_41358_n942_bF_buf1), .Y(alu__abc_41358_n2117) );
  AND2X2 AND2X2_6527 ( .A(alu__abc_41358_n2121), .B(alu__abc_41358_n1057_bF_buf2), .Y(alu__abc_41358_n2122) );
  AND2X2 AND2X2_6528 ( .A(alu__abc_41358_n2122), .B(alu__abc_41358_n2120), .Y(alu__abc_41358_n2123) );
  AND2X2 AND2X2_6529 ( .A(alu__abc_41358_n1416), .B(alu__abc_41358_n279_bF_buf5), .Y(alu__abc_41358_n2124) );
  AND2X2 AND2X2_653 ( .A(_abc_43815_n1786), .B(_abc_43815_n1857), .Y(_abc_43815_n1860) );
  AND2X2 AND2X2_6530 ( .A(alu__abc_41358_n2125), .B(alu__abc_41358_n833_bF_buf2), .Y(alu__abc_41358_n2126) );
  AND2X2 AND2X2_6531 ( .A(alu__abc_41358_n995), .B(alu__abc_41358_n998), .Y(alu__abc_41358_n2127) );
  AND2X2 AND2X2_6532 ( .A(alu__abc_41358_n2128), .B(alu__abc_41358_n2129), .Y(alu__abc_41358_n2130) );
  AND2X2 AND2X2_6533 ( .A(alu__abc_41358_n2131), .B(alu__abc_41358_n2132), .Y(alu__abc_41358_n2133) );
  AND2X2 AND2X2_6534 ( .A(alu__abc_41358_n2133), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n2134) );
  AND2X2 AND2X2_6535 ( .A(alu__abc_41358_n1804), .B(alu_b_i_3_bF_buf3), .Y(alu__abc_41358_n2135) );
  AND2X2 AND2X2_6536 ( .A(alu__abc_41358_n2138), .B(alu__abc_41358_n947), .Y(alu__abc_41358_n2139) );
  AND2X2 AND2X2_6537 ( .A(alu__abc_41358_n2139), .B(alu__abc_41358_n2137), .Y(alu__abc_41358_n2140) );
  AND2X2 AND2X2_6538 ( .A(alu__abc_41358_n932_bF_buf1), .B(alu_a_i_23_), .Y(alu__abc_41358_n2141) );
  AND2X2 AND2X2_6539 ( .A(alu__abc_41358_n186), .B(alu_op_i_0_bF_buf2), .Y(alu__abc_41358_n2142) );
  AND2X2 AND2X2_654 ( .A(_abc_43815_n1862_1), .B(_abc_43815_n1822), .Y(_abc_43815_n1863) );
  AND2X2 AND2X2_6540 ( .A(alu__abc_41358_n927_bF_buf0), .B(alu__abc_41358_n191_1), .Y(alu__abc_41358_n2144) );
  AND2X2 AND2X2_6541 ( .A(alu__abc_41358_n2144), .B(alu__abc_41358_n2143), .Y(alu__abc_41358_n2145) );
  AND2X2 AND2X2_6542 ( .A(alu__abc_41358_n935_bF_buf1), .B(alu__abc_41358_n186), .Y(alu__abc_41358_n2146) );
  AND2X2 AND2X2_6543 ( .A(alu__abc_41358_n649), .B(alu__abc_41358_n1061_bF_buf2), .Y(alu__abc_41358_n2151) );
  AND2X2 AND2X2_6544 ( .A(alu__abc_41358_n2114), .B(alu__abc_41358_n667), .Y(alu__abc_41358_n2155) );
  AND2X2 AND2X2_6545 ( .A(alu__abc_41358_n2157), .B(alu__abc_41358_n942_bF_buf0), .Y(alu__abc_41358_n2158) );
  AND2X2 AND2X2_6546 ( .A(alu__abc_41358_n2158), .B(alu__abc_41358_n2156), .Y(alu__abc_41358_n2159) );
  AND2X2 AND2X2_6547 ( .A(alu__abc_41358_n493), .B(alu__abc_41358_n125_1), .Y(alu__abc_41358_n2161) );
  AND2X2 AND2X2_6548 ( .A(alu__abc_41358_n2162), .B(alu__abc_41358_n1057_bF_buf1), .Y(alu__abc_41358_n2163) );
  AND2X2 AND2X2_6549 ( .A(alu__abc_41358_n2163), .B(alu__abc_41358_n2160), .Y(alu__abc_41358_n2164) );
  AND2X2 AND2X2_655 ( .A(_abc_43815_n1861), .B(_abc_43815_n1863), .Y(_abc_43815_n1864) );
  AND2X2 AND2X2_6550 ( .A(alu__abc_41358_n667), .B(alu__abc_41358_n1061_bF_buf1), .Y(alu__abc_41358_n2165) );
  AND2X2 AND2X2_6551 ( .A(alu__abc_41358_n2166), .B(alu__abc_41358_n1830), .Y(alu__abc_41358_n2167) );
  AND2X2 AND2X2_6552 ( .A(alu__abc_41358_n1481), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n2168) );
  AND2X2 AND2X2_6553 ( .A(alu__abc_41358_n894), .B(alu__abc_41358_n901), .Y(alu__abc_41358_n2171) );
  AND2X2 AND2X2_6554 ( .A(alu__abc_41358_n2170), .B(alu__abc_41358_n2172), .Y(alu__abc_41358_n2173) );
  AND2X2 AND2X2_6555 ( .A(alu__abc_41358_n2174), .B(alu__abc_41358_n2175), .Y(alu__abc_41358_n2176) );
  AND2X2 AND2X2_6556 ( .A(alu__abc_41358_n2169), .B(alu__abc_41358_n2177), .Y(alu__abc_41358_n2178) );
  AND2X2 AND2X2_6557 ( .A(alu__abc_41358_n2178), .B(alu__abc_41358_n948_bF_buf1), .Y(alu__abc_41358_n2179) );
  AND2X2 AND2X2_6558 ( .A(alu__abc_41358_n118), .B(alu_op_i_0_bF_buf1), .Y(alu__abc_41358_n2180) );
  AND2X2 AND2X2_6559 ( .A(alu__abc_41358_n927_bF_buf4), .B(alu__abc_41358_n123), .Y(alu__abc_41358_n2182) );
  AND2X2 AND2X2_656 ( .A(int32_r_10_), .B(pc_q_12_), .Y(_abc_43815_n1868_1) );
  AND2X2 AND2X2_6560 ( .A(alu__abc_41358_n2182), .B(alu__abc_41358_n2181), .Y(alu__abc_41358_n2183) );
  AND2X2 AND2X2_6561 ( .A(alu__abc_41358_n932_bF_buf0), .B(alu_a_i_24_), .Y(alu__abc_41358_n2184) );
  AND2X2 AND2X2_6562 ( .A(alu__abc_41358_n935_bF_buf0), .B(alu__abc_41358_n118), .Y(alu__abc_41358_n2185) );
  AND2X2 AND2X2_6563 ( .A(alu__abc_41358_n2155), .B(alu__abc_41358_n665), .Y(alu__abc_41358_n2195) );
  AND2X2 AND2X2_6564 ( .A(alu__abc_41358_n2196), .B(alu__abc_41358_n2194), .Y(alu__abc_41358_n2197) );
  AND2X2 AND2X2_6565 ( .A(alu__abc_41358_n2197), .B(alu__abc_41358_n942_bF_buf4), .Y(alu__abc_41358_n2198) );
  AND2X2 AND2X2_6566 ( .A(alu__abc_41358_n2162), .B(alu__abc_41358_n398), .Y(alu__abc_41358_n2199) );
  AND2X2 AND2X2_6567 ( .A(alu__abc_41358_n2202), .B(alu__abc_41358_n1057_bF_buf0), .Y(alu__abc_41358_n2203) );
  AND2X2 AND2X2_6568 ( .A(alu__abc_41358_n2203), .B(alu__abc_41358_n2201), .Y(alu__abc_41358_n2204) );
  AND2X2 AND2X2_6569 ( .A(alu__abc_41358_n665), .B(alu__abc_41358_n1061_bF_buf0), .Y(alu__abc_41358_n2205) );
  AND2X2 AND2X2_657 ( .A(_abc_43815_n1869), .B(_abc_43815_n1867), .Y(_abc_43815_n1870) );
  AND2X2 AND2X2_6570 ( .A(alu__abc_41358_n1510), .B(alu__abc_41358_n279_bF_buf3), .Y(alu__abc_41358_n2206) );
  AND2X2 AND2X2_6571 ( .A(alu__abc_41358_n2207), .B(alu__abc_41358_n833_bF_buf1), .Y(alu__abc_41358_n2208) );
  AND2X2 AND2X2_6572 ( .A(alu__abc_41358_n1527), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n2209) );
  AND2X2 AND2X2_6573 ( .A(alu__abc_41358_n999), .B(alu__abc_41358_n972), .Y(alu__abc_41358_n2210) );
  AND2X2 AND2X2_6574 ( .A(alu__abc_41358_n2211), .B(alu__abc_41358_n2212), .Y(alu__abc_41358_n2213) );
  AND2X2 AND2X2_6575 ( .A(alu__abc_41358_n2213), .B(alu__abc_41358_n299_bF_buf4), .Y(alu__abc_41358_n2214) );
  AND2X2 AND2X2_6576 ( .A(alu__abc_41358_n2048), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n2215) );
  AND2X2 AND2X2_6577 ( .A(alu__abc_41358_n2218), .B(alu__abc_41358_n2217), .Y(alu__abc_41358_n2219) );
  AND2X2 AND2X2_6578 ( .A(alu__abc_41358_n2219), .B(alu__abc_41358_n948_bF_buf0), .Y(alu__abc_41358_n2220) );
  AND2X2 AND2X2_6579 ( .A(alu__abc_41358_n932_bF_buf4), .B(alu_a_i_25_), .Y(alu__abc_41358_n2221) );
  AND2X2 AND2X2_658 ( .A(_abc_43815_n1866), .B(_abc_43815_n1870), .Y(_abc_43815_n1871_1) );
  AND2X2 AND2X2_6580 ( .A(alu__abc_41358_n110), .B(alu_op_i_0_bF_buf0), .Y(alu__abc_41358_n2222) );
  AND2X2 AND2X2_6581 ( .A(alu__abc_41358_n927_bF_buf3), .B(alu__abc_41358_n115), .Y(alu__abc_41358_n2224) );
  AND2X2 AND2X2_6582 ( .A(alu__abc_41358_n2224), .B(alu__abc_41358_n2223), .Y(alu__abc_41358_n2225) );
  AND2X2 AND2X2_6583 ( .A(alu__abc_41358_n935_bF_buf4), .B(alu__abc_41358_n110), .Y(alu__abc_41358_n2226) );
  AND2X2 AND2X2_6584 ( .A(alu__abc_41358_n2195), .B(alu__abc_41358_n659), .Y(alu__abc_41358_n2236) );
  AND2X2 AND2X2_6585 ( .A(alu__abc_41358_n2237), .B(alu__abc_41358_n2235), .Y(alu__abc_41358_n2238) );
  AND2X2 AND2X2_6586 ( .A(alu__abc_41358_n2238), .B(alu__abc_41358_n942_bF_buf3), .Y(alu__abc_41358_n2239) );
  AND2X2 AND2X2_6587 ( .A(alu__abc_41358_n2162), .B(alu__abc_41358_n399), .Y(alu__abc_41358_n2240) );
  AND2X2 AND2X2_6588 ( .A(alu__abc_41358_n2242), .B(alu__abc_41358_n134), .Y(alu__abc_41358_n2244) );
  AND2X2 AND2X2_6589 ( .A(alu__abc_41358_n2245), .B(alu__abc_41358_n1057_bF_buf4), .Y(alu__abc_41358_n2246) );
  AND2X2 AND2X2_659 ( .A(_abc_43815_n1873), .B(_abc_43815_n1425_1_bF_buf3), .Y(_abc_43815_n1874_1) );
  AND2X2 AND2X2_6590 ( .A(alu__abc_41358_n2246), .B(alu__abc_41358_n2243), .Y(alu__abc_41358_n2247) );
  AND2X2 AND2X2_6591 ( .A(alu__abc_41358_n659), .B(alu__abc_41358_n1061_bF_buf4), .Y(alu__abc_41358_n2248) );
  AND2X2 AND2X2_6592 ( .A(alu__abc_41358_n1556), .B(alu__abc_41358_n279_bF_buf2), .Y(alu__abc_41358_n2249) );
  AND2X2 AND2X2_6593 ( .A(alu__abc_41358_n2250), .B(alu__abc_41358_n833_bF_buf0), .Y(alu__abc_41358_n2251) );
  AND2X2 AND2X2_6594 ( .A(alu__abc_41358_n1573), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n2252) );
  AND2X2 AND2X2_6595 ( .A(alu__abc_41358_n902), .B(alu__abc_41358_n905), .Y(alu__abc_41358_n2254) );
  AND2X2 AND2X2_6596 ( .A(alu__abc_41358_n2255), .B(alu__abc_41358_n2256), .Y(alu__abc_41358_n2257) );
  AND2X2 AND2X2_6597 ( .A(alu__abc_41358_n2253), .B(alu__abc_41358_n2258), .Y(alu__abc_41358_n2259) );
  AND2X2 AND2X2_6598 ( .A(alu__abc_41358_n2260), .B(alu__abc_41358_n2261), .Y(alu__abc_41358_n2262) );
  AND2X2 AND2X2_6599 ( .A(alu__abc_41358_n2262), .B(alu__abc_41358_n948_bF_buf4), .Y(alu__abc_41358_n2263) );
  AND2X2 AND2X2_66 ( .A(_abc_43815_n718), .B(_abc_43815_n727), .Y(_abc_43815_n728) );
  AND2X2 AND2X2_660 ( .A(_abc_43815_n1874_1), .B(_abc_43815_n1872), .Y(_abc_43815_n1875) );
  AND2X2 AND2X2_6600 ( .A(alu__abc_41358_n932_bF_buf3), .B(alu_a_i_26_), .Y(alu__abc_41358_n2264) );
  AND2X2 AND2X2_6601 ( .A(alu__abc_41358_n935_bF_buf3), .B(alu__abc_41358_n127), .Y(alu__abc_41358_n2265) );
  AND2X2 AND2X2_6602 ( .A(alu__abc_41358_n127), .B(alu_op_i_0_bF_buf5), .Y(alu__abc_41358_n2266) );
  AND2X2 AND2X2_6603 ( .A(alu__abc_41358_n927_bF_buf2), .B(alu__abc_41358_n132), .Y(alu__abc_41358_n2268) );
  AND2X2 AND2X2_6604 ( .A(alu__abc_41358_n2268), .B(alu__abc_41358_n2267), .Y(alu__abc_41358_n2269) );
  AND2X2 AND2X2_6605 ( .A(alu__abc_41358_n2236), .B(alu__abc_41358_n657), .Y(alu__abc_41358_n2279) );
  AND2X2 AND2X2_6606 ( .A(alu__abc_41358_n2280), .B(alu__abc_41358_n2278), .Y(alu__abc_41358_n2281) );
  AND2X2 AND2X2_6607 ( .A(alu__abc_41358_n2281), .B(alu__abc_41358_n942_bF_buf2), .Y(alu__abc_41358_n2282) );
  AND2X2 AND2X2_6608 ( .A(alu__abc_41358_n2286), .B(alu__abc_41358_n1057_bF_buf3), .Y(alu__abc_41358_n2287) );
  AND2X2 AND2X2_6609 ( .A(alu__abc_41358_n2287), .B(alu__abc_41358_n2285), .Y(alu__abc_41358_n2288) );
  AND2X2 AND2X2_661 ( .A(_abc_43815_n1065_1_bF_buf4), .B(epc_q_12_), .Y(_abc_43815_n1876) );
  AND2X2 AND2X2_6610 ( .A(alu__abc_41358_n657), .B(alu__abc_41358_n1061_bF_buf3), .Y(alu__abc_41358_n2289) );
  AND2X2 AND2X2_6611 ( .A(alu__abc_41358_n1605), .B(alu__abc_41358_n279_bF_buf1), .Y(alu__abc_41358_n2290) );
  AND2X2 AND2X2_6612 ( .A(alu__abc_41358_n2291), .B(alu__abc_41358_n833_bF_buf4), .Y(alu__abc_41358_n2292) );
  AND2X2 AND2X2_6613 ( .A(alu__abc_41358_n973), .B(alu__abc_41358_n976), .Y(alu__abc_41358_n2293) );
  AND2X2 AND2X2_6614 ( .A(alu__abc_41358_n2294), .B(alu__abc_41358_n2295), .Y(alu__abc_41358_n2296) );
  AND2X2 AND2X2_6615 ( .A(alu__abc_41358_n2297), .B(alu__abc_41358_n2298), .Y(alu__abc_41358_n2299) );
  AND2X2 AND2X2_6616 ( .A(alu__abc_41358_n2300), .B(alu__abc_41358_n2301), .Y(alu__abc_41358_n2302) );
  AND2X2 AND2X2_6617 ( .A(alu__abc_41358_n2302), .B(alu__abc_41358_n948_bF_buf3), .Y(alu__abc_41358_n2303) );
  AND2X2 AND2X2_6618 ( .A(alu__abc_41358_n1622), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n2304) );
  AND2X2 AND2X2_6619 ( .A(alu__abc_41358_n932_bF_buf2), .B(alu_a_i_27_), .Y(alu__abc_41358_n2305) );
  AND2X2 AND2X2_662 ( .A(_abc_43815_n1878), .B(_abc_43815_n1856_1), .Y(_abc_43815_n1879) );
  AND2X2 AND2X2_6620 ( .A(alu__abc_41358_n935_bF_buf2), .B(alu__abc_41358_n135_1), .Y(alu__abc_41358_n2306) );
  AND2X2 AND2X2_6621 ( .A(alu__abc_41358_n135_1), .B(alu_op_i_0_bF_buf4), .Y(alu__abc_41358_n2307) );
  AND2X2 AND2X2_6622 ( .A(alu__abc_41358_n927_bF_buf1), .B(alu__abc_41358_n140), .Y(alu__abc_41358_n2309) );
  AND2X2 AND2X2_6623 ( .A(alu__abc_41358_n2309), .B(alu__abc_41358_n2308), .Y(alu__abc_41358_n2310) );
  AND2X2 AND2X2_6624 ( .A(alu__abc_41358_n2319), .B(alu__abc_41358_n942_bF_buf1), .Y(alu__abc_41358_n2320) );
  AND2X2 AND2X2_6625 ( .A(alu__abc_41358_n2279), .B(alu__abc_41358_n822), .Y(alu__abc_41358_n2321) );
  AND2X2 AND2X2_6626 ( .A(alu__abc_41358_n2320), .B(alu__abc_41358_n2322), .Y(alu__abc_41358_n2323) );
  AND2X2 AND2X2_6627 ( .A(alu__abc_41358_n495), .B(alu__abc_41358_n152), .Y(alu__abc_41358_n2325) );
  AND2X2 AND2X2_6628 ( .A(alu__abc_41358_n2326), .B(alu__abc_41358_n1057_bF_buf2), .Y(alu__abc_41358_n2327) );
  AND2X2 AND2X2_6629 ( .A(alu__abc_41358_n2327), .B(alu__abc_41358_n2324), .Y(alu__abc_41358_n2328) );
  AND2X2 AND2X2_663 ( .A(_abc_43815_n1880_1), .B(_abc_43815_n1881), .Y(_abc_43815_n1882) );
  AND2X2 AND2X2_6630 ( .A(alu__abc_41358_n822), .B(alu__abc_41358_n1061_bF_buf2), .Y(alu__abc_41358_n2329) );
  AND2X2 AND2X2_6631 ( .A(alu__abc_41358_n2330), .B(alu__abc_41358_n1830), .Y(alu__abc_41358_n2331) );
  AND2X2 AND2X2_6632 ( .A(alu__abc_41358_n906), .B(alu__abc_41358_n911), .Y(alu__abc_41358_n2334) );
  AND2X2 AND2X2_6633 ( .A(alu__abc_41358_n2333), .B(alu__abc_41358_n2335), .Y(alu__abc_41358_n2336) );
  AND2X2 AND2X2_6634 ( .A(alu__abc_41358_n2337), .B(alu__abc_41358_n2338), .Y(alu__abc_41358_n2339) );
  AND2X2 AND2X2_6635 ( .A(alu__abc_41358_n2340), .B(alu__abc_41358_n948_bF_buf2), .Y(alu__abc_41358_n2341) );
  AND2X2 AND2X2_6636 ( .A(alu__abc_41358_n2341), .B(alu__abc_41358_n2332), .Y(alu__abc_41358_n2342) );
  AND2X2 AND2X2_6637 ( .A(alu__abc_41358_n1664), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n2343) );
  AND2X2 AND2X2_6638 ( .A(alu__abc_41358_n145), .B(alu_op_i_0_bF_buf3), .Y(alu__abc_41358_n2344) );
  AND2X2 AND2X2_6639 ( .A(alu__abc_41358_n927_bF_buf0), .B(alu__abc_41358_n150), .Y(alu__abc_41358_n2346) );
  AND2X2 AND2X2_664 ( .A(_abc_43815_n1882), .B(_abc_43815_n1413_bF_buf2), .Y(_abc_43815_n1883) );
  AND2X2 AND2X2_6640 ( .A(alu__abc_41358_n2346), .B(alu__abc_41358_n2345), .Y(alu__abc_41358_n2347) );
  AND2X2 AND2X2_6641 ( .A(alu__abc_41358_n932_bF_buf1), .B(alu_a_i_28_), .Y(alu__abc_41358_n2348) );
  AND2X2 AND2X2_6642 ( .A(alu__abc_41358_n935_bF_buf1), .B(alu__abc_41358_n145), .Y(alu__abc_41358_n2349) );
  AND2X2 AND2X2_6643 ( .A(alu__abc_41358_n2321), .B(alu__abc_41358_n636), .Y(alu__abc_41358_n2359) );
  AND2X2 AND2X2_6644 ( .A(alu__abc_41358_n2360), .B(alu__abc_41358_n2358), .Y(alu__abc_41358_n2361) );
  AND2X2 AND2X2_6645 ( .A(alu__abc_41358_n2361), .B(alu__abc_41358_n942_bF_buf0), .Y(alu__abc_41358_n2362) );
  AND2X2 AND2X2_6646 ( .A(alu__abc_41358_n2326), .B(alu__abc_41358_n501), .Y(alu__abc_41358_n2363) );
  AND2X2 AND2X2_6647 ( .A(alu__abc_41358_n2366), .B(alu__abc_41358_n1057_bF_buf1), .Y(alu__abc_41358_n2367) );
  AND2X2 AND2X2_6648 ( .A(alu__abc_41358_n2367), .B(alu__abc_41358_n2364), .Y(alu__abc_41358_n2368) );
  AND2X2 AND2X2_6649 ( .A(alu__abc_41358_n636), .B(alu__abc_41358_n1061_bF_buf1), .Y(alu__abc_41358_n2369) );
  AND2X2 AND2X2_665 ( .A(_abc_43815_n1884), .B(_abc_43815_n1351_bF_buf4), .Y(_abc_43815_n1885) );
  AND2X2 AND2X2_6650 ( .A(alu__abc_41358_n1696), .B(alu__abc_41358_n279_bF_buf0), .Y(alu__abc_41358_n2370) );
  AND2X2 AND2X2_6651 ( .A(alu__abc_41358_n2371), .B(alu__abc_41358_n833_bF_buf3), .Y(alu__abc_41358_n2372) );
  AND2X2 AND2X2_6652 ( .A(alu__abc_41358_n977), .B(alu__abc_41358_n2374), .Y(alu__abc_41358_n2375) );
  AND2X2 AND2X2_6653 ( .A(alu__abc_41358_n2376), .B(alu__abc_41358_n2377), .Y(alu__abc_41358_n2378) );
  AND2X2 AND2X2_6654 ( .A(alu__abc_41358_n2379), .B(alu__abc_41358_n2380), .Y(alu__abc_41358_n2381) );
  AND2X2 AND2X2_6655 ( .A(alu__abc_41358_n2381), .B(alu__abc_41358_n294_bF_buf1), .Y(alu__abc_41358_n2382) );
  AND2X2 AND2X2_6656 ( .A(alu__abc_41358_n2051), .B(alu_b_i_3_bF_buf4), .Y(alu__abc_41358_n2383) );
  AND2X2 AND2X2_6657 ( .A(alu__abc_41358_n2385), .B(alu__abc_41358_n947), .Y(alu__abc_41358_n2386) );
  AND2X2 AND2X2_6658 ( .A(alu__abc_41358_n2386), .B(alu__abc_41358_n2373), .Y(alu__abc_41358_n2387) );
  AND2X2 AND2X2_6659 ( .A(alu__abc_41358_n153), .B(alu_op_i_0_bF_buf2), .Y(alu__abc_41358_n2388) );
  AND2X2 AND2X2_666 ( .A(_abc_43815_n1887), .B(enable_i_bF_buf3), .Y(_abc_43815_n1888) );
  AND2X2 AND2X2_6660 ( .A(alu__abc_41358_n927_bF_buf4), .B(alu__abc_41358_n158), .Y(alu__abc_41358_n2390) );
  AND2X2 AND2X2_6661 ( .A(alu__abc_41358_n2390), .B(alu__abc_41358_n2389), .Y(alu__abc_41358_n2391) );
  AND2X2 AND2X2_6662 ( .A(alu__abc_41358_n932_bF_buf0), .B(alu_a_i_29_), .Y(alu__abc_41358_n2392) );
  AND2X2 AND2X2_6663 ( .A(alu__abc_41358_n935_bF_buf0), .B(alu__abc_41358_n153), .Y(alu__abc_41358_n2393) );
  AND2X2 AND2X2_6664 ( .A(alu__abc_41358_n2359), .B(alu__abc_41358_n629), .Y(alu__abc_41358_n2401) );
  AND2X2 AND2X2_6665 ( .A(alu__abc_41358_n2403), .B(alu__abc_41358_n942_bF_buf4), .Y(alu__abc_41358_n2404) );
  AND2X2 AND2X2_6666 ( .A(alu__abc_41358_n2404), .B(alu__abc_41358_n2402), .Y(alu__abc_41358_n2405) );
  AND2X2 AND2X2_6667 ( .A(alu__abc_41358_n507), .B(alu__abc_41358_n1057_bF_buf0), .Y(alu__abc_41358_n2407) );
  AND2X2 AND2X2_6668 ( .A(alu__abc_41358_n2407), .B(alu__abc_41358_n2406), .Y(alu__abc_41358_n2408) );
  AND2X2 AND2X2_6669 ( .A(alu__abc_41358_n629), .B(alu__abc_41358_n1061_bF_buf0), .Y(alu__abc_41358_n2409) );
  AND2X2 AND2X2_667 ( .A(_abc_43815_n1886), .B(_abc_43815_n1888), .Y(epc_q_12__FF_INPUT) );
  AND2X2 AND2X2_6670 ( .A(alu__abc_41358_n1745), .B(alu__abc_41358_n279_bF_buf4), .Y(alu__abc_41358_n2410) );
  AND2X2 AND2X2_6671 ( .A(alu__abc_41358_n2411), .B(alu__abc_41358_n833_bF_buf2), .Y(alu__abc_41358_n2412) );
  AND2X2 AND2X2_6672 ( .A(alu__abc_41358_n912), .B(alu__abc_41358_n915), .Y(alu__abc_41358_n2413) );
  AND2X2 AND2X2_6673 ( .A(alu__abc_41358_n2414), .B(alu__abc_41358_n2415), .Y(alu__abc_41358_n2416) );
  AND2X2 AND2X2_6674 ( .A(alu__abc_41358_n2417), .B(alu__abc_41358_n2418), .Y(alu__abc_41358_n2419) );
  AND2X2 AND2X2_6675 ( .A(alu__abc_41358_n2420), .B(alu__abc_41358_n2421), .Y(alu__abc_41358_n2422) );
  AND2X2 AND2X2_6676 ( .A(alu__abc_41358_n2422), .B(alu__abc_41358_n948_bF_buf1), .Y(alu__abc_41358_n2423) );
  AND2X2 AND2X2_6677 ( .A(alu__abc_41358_n1758), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n2424) );
  AND2X2 AND2X2_6678 ( .A(alu__abc_41358_n932_bF_buf4), .B(alu_a_i_30_), .Y(alu__abc_41358_n2425) );
  AND2X2 AND2X2_6679 ( .A(alu__abc_41358_n162), .B(alu_op_i_0_bF_buf1), .Y(alu__abc_41358_n2426) );
  AND2X2 AND2X2_668 ( .A(_abc_43815_n1847_1), .B(pc_q_13_), .Y(_abc_43815_n1891) );
  AND2X2 AND2X2_6680 ( .A(alu__abc_41358_n927_bF_buf3), .B(alu__abc_41358_n167_1), .Y(alu__abc_41358_n2428) );
  AND2X2 AND2X2_6681 ( .A(alu__abc_41358_n2428), .B(alu__abc_41358_n2427), .Y(alu__abc_41358_n2429) );
  AND2X2 AND2X2_6682 ( .A(alu__abc_41358_n935_bF_buf4), .B(alu__abc_41358_n162), .Y(alu__abc_41358_n2430) );
  AND2X2 AND2X2_6683 ( .A(alu__abc_41358_n2440), .B(alu__abc_41358_n942_bF_buf3), .Y(alu__abc_41358_n2441) );
  AND2X2 AND2X2_6684 ( .A(alu__abc_41358_n2439), .B(alu__abc_41358_n2441), .Y(alu__abc_41358_n2442) );
  AND2X2 AND2X2_6685 ( .A(alu__abc_41358_n2444), .B(alu__abc_41358_n2445), .Y(alu__abc_41358_n2446) );
  AND2X2 AND2X2_6686 ( .A(alu__abc_41358_n2446), .B(alu__abc_41358_n299_bF_buf6), .Y(alu__abc_41358_n2447) );
  AND2X2 AND2X2_6687 ( .A(alu__abc_41358_n2296), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n2448) );
  AND2X2 AND2X2_6688 ( .A(alu__abc_41358_n2451), .B(alu__abc_41358_n2450), .Y(alu__abc_41358_n2452) );
  AND2X2 AND2X2_6689 ( .A(alu__abc_41358_n2452), .B(alu__abc_41358_n948_bF_buf0), .Y(alu__abc_41358_n2453) );
  AND2X2 AND2X2_669 ( .A(_abc_43815_n1892), .B(_abc_43815_n1890), .Y(_abc_43815_n1893) );
  AND2X2 AND2X2_6690 ( .A(alu__abc_41358_n627), .B(alu__abc_41358_n1061_bF_buf4), .Y(alu__abc_41358_n2454) );
  AND2X2 AND2X2_6691 ( .A(alu__abc_41358_n2455), .B(alu__abc_41358_n522), .Y(alu__abc_41358_n2456) );
  AND2X2 AND2X2_6692 ( .A(alu__abc_41358_n2457), .B(alu__abc_41358_n1057_bF_buf4), .Y(alu__abc_41358_n2458) );
  AND2X2 AND2X2_6693 ( .A(alu__abc_41358_n1793), .B(alu__abc_41358_n279_bF_buf3), .Y(alu__abc_41358_n2459) );
  AND2X2 AND2X2_6694 ( .A(alu__abc_41358_n2460), .B(alu__abc_41358_n833_bF_buf1), .Y(alu__abc_41358_n2461) );
  AND2X2 AND2X2_6695 ( .A(alu__abc_41358_n1806), .B(alu__abc_41358_n1850), .Y(alu__abc_41358_n2462) );
  AND2X2 AND2X2_6696 ( .A(alu__abc_41358_n932_bF_buf3), .B(alu_a_i_31_), .Y(alu__abc_41358_n2463) );
  AND2X2 AND2X2_6697 ( .A(alu__abc_41358_n170), .B(alu_op_i_0_bF_buf0), .Y(alu__abc_41358_n2464) );
  AND2X2 AND2X2_6698 ( .A(alu__abc_41358_n927_bF_buf2), .B(alu__abc_41358_n530), .Y(alu__abc_41358_n2466) );
  AND2X2 AND2X2_6699 ( .A(alu__abc_41358_n2466), .B(alu__abc_41358_n2465), .Y(alu__abc_41358_n2467) );
  AND2X2 AND2X2_67 ( .A(_abc_43815_n682), .B(alu_p_o_2_), .Y(_abc_43815_n730_1) );
  AND2X2 AND2X2_670 ( .A(_abc_43815_n1692), .B(_abc_43815_n1894), .Y(_abc_43815_n1895) );
  AND2X2 AND2X2_6700 ( .A(alu__abc_41358_n935_bF_buf3), .B(alu__abc_41358_n170), .Y(alu__abc_41358_n2468) );
  AND2X2 AND2X2_6701 ( .A(alu__abc_41358_n1144), .B(alu__abc_41358_n2477), .Y(alu__abc_41358_n2478) );
  AND2X2 AND2X2_6702 ( .A(alu__abc_41358_n303), .B(alu__abc_41358_n2479), .Y(alu__abc_41358_n2480) );
  AND2X2 AND2X2_6703 ( .A(alu__abc_41358_n266), .B(alu_b_i_6_), .Y(alu__abc_41358_n2481) );
  AND2X2 AND2X2_6704 ( .A(alu__abc_41358_n275), .B(alu__abc_41358_n2481), .Y(alu__abc_41358_n2482) );
  AND2X2 AND2X2_6705 ( .A(alu__abc_41358_n280), .B(alu_b_i_4_bF_buf3), .Y(alu__abc_41358_n2484) );
  AND2X2 AND2X2_6706 ( .A(alu__abc_41358_n289), .B(alu__abc_41358_n2484), .Y(alu__abc_41358_n2485) );
  AND2X2 AND2X2_6707 ( .A(alu__abc_41358_n2486), .B(alu__abc_41358_n276), .Y(alu__abc_41358_n2487) );
  AND2X2 AND2X2_6708 ( .A(alu__abc_41358_n298), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n2489) );
  AND2X2 AND2X2_6709 ( .A(alu__abc_41358_n296), .B(alu__abc_41358_n2489), .Y(alu__abc_41358_n2490) );
  AND2X2 AND2X2_671 ( .A(_abc_43815_n1418_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_43815_n1896) );
  AND2X2 AND2X2_6710 ( .A(alu__abc_41358_n291), .B(alu__abc_41358_n2491), .Y(alu__abc_41358_n2492) );
  AND2X2 AND2X2_6711 ( .A(alu__abc_41358_n2494), .B(alu__abc_41358_n375), .Y(alu__abc_41358_n2495) );
  AND2X2 AND2X2_6712 ( .A(alu__abc_41358_n351), .B(alu_b_i_11_), .Y(alu__abc_41358_n2496) );
  AND2X2 AND2X2_6713 ( .A(alu__abc_41358_n343), .B(alu_b_i_10_), .Y(alu__abc_41358_n2497) );
  AND2X2 AND2X2_6714 ( .A(alu__abc_41358_n355), .B(alu__abc_41358_n2497), .Y(alu__abc_41358_n2498) );
  AND2X2 AND2X2_6715 ( .A(alu__abc_41358_n360), .B(alu_b_i_8_), .Y(alu__abc_41358_n2500) );
  AND2X2 AND2X2_6716 ( .A(alu__abc_41358_n2501), .B(alu__abc_41358_n432), .Y(alu__abc_41358_n2502) );
  AND2X2 AND2X2_6717 ( .A(alu__abc_41358_n356), .B(alu__abc_41358_n2502), .Y(alu__abc_41358_n2503) );
  AND2X2 AND2X2_6718 ( .A(alu__abc_41358_n2504), .B(alu__abc_41358_n339), .Y(alu__abc_41358_n2505) );
  AND2X2 AND2X2_6719 ( .A(alu__abc_41358_n333), .B(alu_b_i_15_), .Y(alu__abc_41358_n2506) );
  AND2X2 AND2X2_672 ( .A(_abc_43815_n1489_bF_buf2), .B(epc_q_13_), .Y(_abc_43815_n1897) );
  AND2X2 AND2X2_6720 ( .A(alu__abc_41358_n325), .B(alu_b_i_14_), .Y(alu__abc_41358_n2507) );
  AND2X2 AND2X2_6721 ( .A(alu__abc_41358_n337), .B(alu__abc_41358_n2507), .Y(alu__abc_41358_n2508) );
  AND2X2 AND2X2_6722 ( .A(alu__abc_41358_n308), .B(alu_b_i_12_), .Y(alu__abc_41358_n2510) );
  AND2X2 AND2X2_6723 ( .A(alu__abc_41358_n2511), .B(alu__abc_41358_n447), .Y(alu__abc_41358_n2512) );
  AND2X2 AND2X2_6724 ( .A(alu__abc_41358_n338), .B(alu__abc_41358_n2512), .Y(alu__abc_41358_n2513) );
  AND2X2 AND2X2_6725 ( .A(alu__abc_41358_n2516), .B(alu__abc_41358_n249), .Y(alu__abc_41358_n2517) );
  AND2X2 AND2X2_6726 ( .A(alu__abc_41358_n138), .B(alu_b_i_27_), .Y(alu__abc_41358_n2518) );
  AND2X2 AND2X2_6727 ( .A(alu__abc_41358_n130_1), .B(alu_b_i_26_), .Y(alu__abc_41358_n2519) );
  AND2X2 AND2X2_6728 ( .A(alu__abc_41358_n142), .B(alu__abc_41358_n2519), .Y(alu__abc_41358_n2520) );
  AND2X2 AND2X2_6729 ( .A(alu__abc_41358_n121), .B(alu_b_i_24_), .Y(alu__abc_41358_n2522) );
  AND2X2 AND2X2_673 ( .A(_abc_43815_n1350_bF_buf3), .B(_abc_43815_n1898), .Y(_abc_43815_n1899) );
  AND2X2 AND2X2_6730 ( .A(alu__abc_41358_n2523), .B(alu__abc_41358_n396), .Y(alu__abc_41358_n2524) );
  AND2X2 AND2X2_6731 ( .A(alu__abc_41358_n143_1), .B(alu__abc_41358_n2524), .Y(alu__abc_41358_n2525) );
  AND2X2 AND2X2_6732 ( .A(alu__abc_41358_n2526), .B(alu__abc_41358_n176), .Y(alu__abc_41358_n2527) );
  AND2X2 AND2X2_6733 ( .A(alu__abc_41358_n165), .B(alu_b_i_30_), .Y(alu__abc_41358_n2528) );
  AND2X2 AND2X2_6734 ( .A(alu__abc_41358_n174), .B(alu__abc_41358_n2528), .Y(alu__abc_41358_n2529) );
  AND2X2 AND2X2_6735 ( .A(alu__abc_41358_n172_1), .B(alu_b_i_31_), .Y(alu__abc_41358_n2530) );
  AND2X2 AND2X2_6736 ( .A(alu__abc_41358_n148_1), .B(alu_b_i_28_), .Y(alu__abc_41358_n2532) );
  AND2X2 AND2X2_6737 ( .A(alu__abc_41358_n2533), .B(alu__abc_41358_n499), .Y(alu__abc_41358_n2534) );
  AND2X2 AND2X2_6738 ( .A(alu__abc_41358_n175), .B(alu__abc_41358_n2534), .Y(alu__abc_41358_n2535) );
  AND2X2 AND2X2_6739 ( .A(alu__abc_41358_n224), .B(alu_b_i_19_), .Y(alu__abc_41358_n2538) );
  AND2X2 AND2X2_674 ( .A(pc_q_13_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_43815_n1902) );
  AND2X2 AND2X2_6740 ( .A(alu__abc_41358_n216), .B(alu_b_i_18_), .Y(alu__abc_41358_n2539) );
  AND2X2 AND2X2_6741 ( .A(alu__abc_41358_n228), .B(alu__abc_41358_n2539), .Y(alu__abc_41358_n2540) );
  AND2X2 AND2X2_6742 ( .A(alu__abc_41358_n233), .B(alu_b_i_16_), .Y(alu__abc_41358_n2542) );
  AND2X2 AND2X2_6743 ( .A(alu__abc_41358_n2543), .B(alu__abc_41358_n464), .Y(alu__abc_41358_n2544) );
  AND2X2 AND2X2_6744 ( .A(alu__abc_41358_n229), .B(alu__abc_41358_n2544), .Y(alu__abc_41358_n2545) );
  AND2X2 AND2X2_6745 ( .A(alu__abc_41358_n2546), .B(alu__abc_41358_n212), .Y(alu__abc_41358_n2547) );
  AND2X2 AND2X2_6746 ( .A(alu__abc_41358_n189), .B(alu_b_i_23_), .Y(alu__abc_41358_n2548) );
  AND2X2 AND2X2_6747 ( .A(alu__abc_41358_n181), .B(alu_b_i_22_), .Y(alu__abc_41358_n2549) );
  AND2X2 AND2X2_6748 ( .A(alu__abc_41358_n193), .B(alu__abc_41358_n2549), .Y(alu__abc_41358_n2550) );
  AND2X2 AND2X2_6749 ( .A(alu__abc_41358_n198_1), .B(alu_b_i_20_), .Y(alu__abc_41358_n2552) );
  AND2X2 AND2X2_675 ( .A(_abc_43815_n1903), .B(_abc_43815_n1901), .Y(_abc_43815_n1904) );
  AND2X2 AND2X2_6750 ( .A(alu__abc_41358_n2553), .B(alu__abc_41358_n479), .Y(alu__abc_41358_n2554) );
  AND2X2 AND2X2_6751 ( .A(alu__abc_41358_n194_1), .B(alu__abc_41358_n2554), .Y(alu__abc_41358_n2555) );
  AND2X2 AND2X2_6752 ( .A(alu__abc_41358_n2557), .B(alu__abc_41358_n177_1), .Y(alu__abc_41358_n2558) );
  AND2X2 AND2X2_6753 ( .A(alu__abc_41358_n2563), .B(alu__abc_41358_n2562), .Y(alu_greater_than_signed_o) );
  AND2X2 AND2X2_6754 ( .A(alu__abc_41358_n2560), .B(alu__abc_41358_n2562), .Y(alu_less_than_o) );
  AND2X2 AND2X2_676 ( .A(_abc_43815_n1870), .B(_abc_43815_n1904), .Y(_abc_43815_n1907) );
  AND2X2 AND2X2_677 ( .A(_abc_43815_n1866), .B(_abc_43815_n1907), .Y(_abc_43815_n1908) );
  AND2X2 AND2X2_678 ( .A(_abc_43815_n1904), .B(_abc_43815_n1868_1), .Y(_abc_43815_n1910) );
  AND2X2 AND2X2_679 ( .A(_abc_43815_n1425_1_bF_buf2), .B(_abc_43815_n1911), .Y(_abc_43815_n1912) );
  AND2X2 AND2X2_68 ( .A(_abc_43815_n694), .B(\mem_dat_i[18] ), .Y(_abc_43815_n731) );
  AND2X2 AND2X2_680 ( .A(_abc_43815_n1909), .B(_abc_43815_n1912), .Y(_abc_43815_n1913) );
  AND2X2 AND2X2_681 ( .A(_abc_43815_n1913), .B(_abc_43815_n1906), .Y(_abc_43815_n1914) );
  AND2X2 AND2X2_682 ( .A(_abc_43815_n1065_1_bF_buf3), .B(epc_q_13_), .Y(_abc_43815_n1915) );
  AND2X2 AND2X2_683 ( .A(_abc_43815_n1917), .B(_abc_43815_n1900), .Y(_abc_43815_n1918_1) );
  AND2X2 AND2X2_684 ( .A(_abc_43815_n1919), .B(_abc_43815_n1920_1), .Y(_abc_43815_n1921) );
  AND2X2 AND2X2_685 ( .A(_abc_43815_n1921), .B(_abc_43815_n1413_bF_buf1), .Y(_abc_43815_n1922_1) );
  AND2X2 AND2X2_686 ( .A(_abc_43815_n1923_1), .B(_abc_43815_n1351_bF_buf3), .Y(_abc_43815_n1924) );
  AND2X2 AND2X2_687 ( .A(_abc_43815_n1926), .B(enable_i_bF_buf2), .Y(_abc_43815_n1927) );
  AND2X2 AND2X2_688 ( .A(_abc_43815_n1925_1), .B(_abc_43815_n1927), .Y(epc_q_13__FF_INPUT) );
  AND2X2 AND2X2_689 ( .A(_abc_43815_n1891), .B(pc_q_14_), .Y(_abc_43815_n1930) );
  AND2X2 AND2X2_69 ( .A(_abc_43815_n697), .B(\mem_dat_i[2] ), .Y(_abc_43815_n732) );
  AND2X2 AND2X2_690 ( .A(_abc_43815_n1931), .B(_abc_43815_n1929), .Y(_abc_43815_n1932) );
  AND2X2 AND2X2_691 ( .A(_abc_43815_n1692), .B(_abc_43815_n1933), .Y(_abc_43815_n1934) );
  AND2X2 AND2X2_692 ( .A(_abc_43815_n1418_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_43815_n1935) );
  AND2X2 AND2X2_693 ( .A(_abc_43815_n1489_bF_buf1), .B(epc_q_14_), .Y(_abc_43815_n1936) );
  AND2X2 AND2X2_694 ( .A(_abc_43815_n1350_bF_buf2), .B(_abc_43815_n1937), .Y(_abc_43815_n1938) );
  AND2X2 AND2X2_695 ( .A(_abc_43815_n1911), .B(_abc_43815_n1903), .Y(_abc_43815_n1940) );
  AND2X2 AND2X2_696 ( .A(_abc_43815_n1909), .B(_abc_43815_n1940), .Y(_abc_43815_n1941) );
  AND2X2 AND2X2_697 ( .A(pc_q_14_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_43815_n1944) );
  AND2X2 AND2X2_698 ( .A(_abc_43815_n1945), .B(_abc_43815_n1943), .Y(_abc_43815_n1946) );
  AND2X2 AND2X2_699 ( .A(_abc_43815_n1942), .B(_abc_43815_n1946), .Y(_abc_43815_n1947) );
  AND2X2 AND2X2_7 ( .A(_abc_43815_n629), .B(_abc_43815_n630), .Y(_abc_43815_n631) );
  AND2X2 AND2X2_70 ( .A(_abc_43815_n733_1), .B(_abc_43815_n686_1_bF_buf2), .Y(_abc_43815_n734) );
  AND2X2 AND2X2_700 ( .A(_abc_43815_n1949), .B(_abc_43815_n1425_1_bF_buf1), .Y(_abc_43815_n1950) );
  AND2X2 AND2X2_701 ( .A(_abc_43815_n1950), .B(_abc_43815_n1948), .Y(_abc_43815_n1951) );
  AND2X2 AND2X2_702 ( .A(_abc_43815_n1065_1_bF_buf2), .B(epc_q_14_), .Y(_abc_43815_n1952) );
  AND2X2 AND2X2_703 ( .A(_abc_43815_n1954_1), .B(_abc_43815_n1939), .Y(_abc_43815_n1955) );
  AND2X2 AND2X2_704 ( .A(_abc_43815_n1956), .B(_abc_43815_n1957), .Y(_abc_43815_n1958) );
  AND2X2 AND2X2_705 ( .A(_abc_43815_n1958), .B(_abc_43815_n1413_bF_buf0), .Y(_abc_43815_n1959) );
  AND2X2 AND2X2_706 ( .A(_abc_43815_n1960), .B(_abc_43815_n1351_bF_buf2), .Y(_abc_43815_n1961) );
  AND2X2 AND2X2_707 ( .A(_abc_43815_n1963), .B(enable_i_bF_buf1), .Y(_abc_43815_n1964) );
  AND2X2 AND2X2_708 ( .A(_abc_43815_n1962), .B(_abc_43815_n1964), .Y(epc_q_14__FF_INPUT) );
  AND2X2 AND2X2_709 ( .A(_abc_43815_n1930), .B(pc_q_15_), .Y(_abc_43815_n1967) );
  AND2X2 AND2X2_71 ( .A(_abc_43815_n689), .B(\mem_dat_i[26] ), .Y(_abc_43815_n735) );
  AND2X2 AND2X2_710 ( .A(_abc_43815_n1968), .B(_abc_43815_n1966), .Y(_abc_43815_n1969) );
  AND2X2 AND2X2_711 ( .A(_abc_43815_n1692), .B(_abc_43815_n1970), .Y(_abc_43815_n1971) );
  AND2X2 AND2X2_712 ( .A(_abc_43815_n1948), .B(_abc_43815_n1945), .Y(_abc_43815_n1972) );
  AND2X2 AND2X2_713 ( .A(pc_q_15_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_43815_n1975) );
  AND2X2 AND2X2_714 ( .A(_abc_43815_n1976), .B(_abc_43815_n1974_1), .Y(_abc_43815_n1977) );
  AND2X2 AND2X2_715 ( .A(_abc_43815_n1980), .B(_abc_43815_n1425_1_bF_buf0), .Y(_abc_43815_n1981) );
  AND2X2 AND2X2_716 ( .A(_abc_43815_n1981), .B(_abc_43815_n1978), .Y(_abc_43815_n1982) );
  AND2X2 AND2X2_717 ( .A(_abc_43815_n1065_1_bF_buf1), .B(epc_q_15_), .Y(_abc_43815_n1983) );
  AND2X2 AND2X2_718 ( .A(_abc_43815_n1985), .B(_abc_43815_n1986), .Y(_abc_43815_n1987) );
  AND2X2 AND2X2_719 ( .A(_abc_43815_n1988), .B(_abc_43815_n1989), .Y(_abc_43815_n1990) );
  AND2X2 AND2X2_72 ( .A(_abc_43815_n696), .B(\mem_dat_i[10] ), .Y(_abc_43815_n736) );
  AND2X2 AND2X2_720 ( .A(_abc_43815_n1418_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_43815_n1992) );
  AND2X2 AND2X2_721 ( .A(_abc_43815_n1489_bF_buf0), .B(epc_q_15_), .Y(_abc_43815_n1993_1) );
  AND2X2 AND2X2_722 ( .A(_abc_43815_n1995), .B(_abc_43815_n1351_bF_buf1), .Y(_abc_43815_n1996) );
  AND2X2 AND2X2_723 ( .A(_abc_43815_n1991), .B(_abc_43815_n1996), .Y(_abc_43815_n1997) );
  AND2X2 AND2X2_724 ( .A(_abc_43815_n1999), .B(enable_i_bF_buf0), .Y(_abc_43815_n2000) );
  AND2X2 AND2X2_725 ( .A(_abc_43815_n1998), .B(_abc_43815_n2000), .Y(epc_q_15__FF_INPUT) );
  AND2X2 AND2X2_726 ( .A(_abc_43815_n1967), .B(pc_q_16_), .Y(_abc_43815_n2003) );
  AND2X2 AND2X2_727 ( .A(_abc_43815_n2004), .B(_abc_43815_n2002), .Y(_abc_43815_n2005) );
  AND2X2 AND2X2_728 ( .A(_abc_43815_n1692), .B(_abc_43815_n2006), .Y(_abc_43815_n2007) );
  AND2X2 AND2X2_729 ( .A(_abc_43815_n1418_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_43815_n2008) );
  AND2X2 AND2X2_73 ( .A(_abc_43815_n704), .B(\mem_dat_i[18] ), .Y(_abc_43815_n738) );
  AND2X2 AND2X2_730 ( .A(_abc_43815_n1489_bF_buf4), .B(epc_q_16_), .Y(_abc_43815_n2009) );
  AND2X2 AND2X2_731 ( .A(_abc_43815_n1350_bF_buf0), .B(_abc_43815_n2010), .Y(_abc_43815_n2011) );
  AND2X2 AND2X2_732 ( .A(_abc_43815_n1946), .B(_abc_43815_n1977), .Y(_abc_43815_n2012) );
  AND2X2 AND2X2_733 ( .A(_abc_43815_n1974_1), .B(_abc_43815_n1944), .Y(_abc_43815_n2015) );
  AND2X2 AND2X2_734 ( .A(_abc_43815_n2014), .B(_abc_43815_n2017), .Y(_abc_43815_n2018) );
  AND2X2 AND2X2_735 ( .A(_abc_43815_n1907), .B(_abc_43815_n2012), .Y(_abc_43815_n2020) );
  AND2X2 AND2X2_736 ( .A(_abc_43815_n1866), .B(_abc_43815_n2020), .Y(_abc_43815_n2021) );
  AND2X2 AND2X2_737 ( .A(pc_q_16_), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_43815_n2024) );
  AND2X2 AND2X2_738 ( .A(_abc_43815_n2025), .B(_abc_43815_n2023), .Y(_abc_43815_n2026) );
  AND2X2 AND2X2_739 ( .A(_abc_43815_n2022), .B(_abc_43815_n2026), .Y(_abc_43815_n2028) );
  AND2X2 AND2X2_74 ( .A(_abc_43815_n706_1), .B(\mem_dat_i[2] ), .Y(_abc_43815_n739) );
  AND2X2 AND2X2_740 ( .A(_abc_43815_n2029), .B(_abc_43815_n1425_1_bF_buf4), .Y(_abc_43815_n2030) );
  AND2X2 AND2X2_741 ( .A(_abc_43815_n2030), .B(_abc_43815_n2027), .Y(_abc_43815_n2031) );
  AND2X2 AND2X2_742 ( .A(_abc_43815_n1065_1_bF_buf0), .B(epc_q_16_), .Y(_abc_43815_n2032) );
  AND2X2 AND2X2_743 ( .A(_abc_43815_n2034_1), .B(_abc_43815_n2035), .Y(_abc_43815_n2036) );
  AND2X2 AND2X2_744 ( .A(_abc_43815_n2036), .B(_abc_43815_n1472_1_bF_buf4), .Y(_abc_43815_n2037) );
  AND2X2 AND2X2_745 ( .A(_abc_43815_n2005), .B(_abc_43815_n1473_bF_buf0), .Y(_abc_43815_n2038) );
  AND2X2 AND2X2_746 ( .A(_abc_43815_n2039), .B(_abc_43815_n1413_bF_buf3), .Y(_abc_43815_n2040) );
  AND2X2 AND2X2_747 ( .A(_abc_43815_n2041), .B(_abc_43815_n1351_bF_buf0), .Y(_abc_43815_n2042) );
  AND2X2 AND2X2_748 ( .A(_abc_43815_n2044), .B(enable_i_bF_buf7), .Y(_abc_43815_n2045) );
  AND2X2 AND2X2_749 ( .A(_abc_43815_n2043), .B(_abc_43815_n2045), .Y(epc_q_16__FF_INPUT) );
  AND2X2 AND2X2_75 ( .A(_abc_43815_n741), .B(_abc_43815_n685), .Y(_abc_43815_n742) );
  AND2X2 AND2X2_750 ( .A(_abc_43815_n2003), .B(pc_q_17_), .Y(_abc_43815_n2048) );
  AND2X2 AND2X2_751 ( .A(_abc_43815_n2049), .B(_abc_43815_n2047), .Y(_abc_43815_n2050) );
  AND2X2 AND2X2_752 ( .A(_abc_43815_n2050), .B(_abc_43815_n1461_bF_buf1), .Y(_abc_43815_n2051) );
  AND2X2 AND2X2_753 ( .A(_abc_43815_n1418_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_43815_n2053) );
  AND2X2 AND2X2_754 ( .A(_abc_43815_n1489_bF_buf3), .B(epc_q_17_), .Y(_abc_43815_n2054) );
  AND2X2 AND2X2_755 ( .A(_abc_43815_n1350_bF_buf4), .B(_abc_43815_n2055_1), .Y(_abc_43815_n2056) );
  AND2X2 AND2X2_756 ( .A(pc_q_17_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2), .Y(_abc_43815_n2059) );
  AND2X2 AND2X2_757 ( .A(_abc_43815_n2060), .B(_abc_43815_n2058), .Y(_abc_43815_n2061) );
  AND2X2 AND2X2_758 ( .A(_abc_43815_n2026), .B(_abc_43815_n2061), .Y(_abc_43815_n2064) );
  AND2X2 AND2X2_759 ( .A(_abc_43815_n2022), .B(_abc_43815_n2064), .Y(_abc_43815_n2065) );
  AND2X2 AND2X2_76 ( .A(_abc_43815_n743), .B(state_q_1_bF_buf4), .Y(_abc_43815_n744) );
  AND2X2 AND2X2_760 ( .A(_abc_43815_n2061), .B(_abc_43815_n2024), .Y(_abc_43815_n2067) );
  AND2X2 AND2X2_761 ( .A(_abc_43815_n1425_1_bF_buf3), .B(_abc_43815_n2068), .Y(_abc_43815_n2069) );
  AND2X2 AND2X2_762 ( .A(_abc_43815_n2066), .B(_abc_43815_n2069), .Y(_abc_43815_n2070) );
  AND2X2 AND2X2_763 ( .A(_abc_43815_n2070), .B(_abc_43815_n2063), .Y(_abc_43815_n2071) );
  AND2X2 AND2X2_764 ( .A(_abc_43815_n1065_1_bF_buf4), .B(epc_q_17_), .Y(_abc_43815_n2072) );
  AND2X2 AND2X2_765 ( .A(_abc_43815_n2074), .B(_abc_43815_n2057), .Y(_abc_43815_n2075) );
  AND2X2 AND2X2_766 ( .A(_abc_43815_n2076), .B(_abc_43815_n2077), .Y(_abc_43815_n2078) );
  AND2X2 AND2X2_767 ( .A(_abc_43815_n2078), .B(_abc_43815_n1413_bF_buf2), .Y(_abc_43815_n2079) );
  AND2X2 AND2X2_768 ( .A(_abc_43815_n2080), .B(_abc_43815_n1351_bF_buf4), .Y(_abc_43815_n2081) );
  AND2X2 AND2X2_769 ( .A(_abc_43815_n2083), .B(enable_i_bF_buf6), .Y(_abc_43815_n2084) );
  AND2X2 AND2X2_77 ( .A(_abc_43815_n682), .B(alu_p_o_3_), .Y(_abc_43815_n746) );
  AND2X2 AND2X2_770 ( .A(_abc_43815_n2082), .B(_abc_43815_n2084), .Y(epc_q_17__FF_INPUT) );
  AND2X2 AND2X2_771 ( .A(_abc_43815_n2048), .B(pc_q_18_), .Y(_abc_43815_n2087_1) );
  AND2X2 AND2X2_772 ( .A(_abc_43815_n2088), .B(_abc_43815_n2086), .Y(_abc_43815_n2089) );
  AND2X2 AND2X2_773 ( .A(_abc_43815_n2089), .B(_abc_43815_n1461_bF_buf0), .Y(_abc_43815_n2090) );
  AND2X2 AND2X2_774 ( .A(_abc_43815_n2068), .B(_abc_43815_n2060), .Y(_abc_43815_n2093) );
  AND2X2 AND2X2_775 ( .A(_abc_43815_n2066), .B(_abc_43815_n2093), .Y(_abc_43815_n2094) );
  AND2X2 AND2X2_776 ( .A(pc_q_18_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(_abc_43815_n2097) );
  AND2X2 AND2X2_777 ( .A(_abc_43815_n2098), .B(_abc_43815_n2096), .Y(_abc_43815_n2099) );
  AND2X2 AND2X2_778 ( .A(_abc_43815_n2095), .B(_abc_43815_n2099), .Y(_abc_43815_n2100) );
  AND2X2 AND2X2_779 ( .A(_abc_43815_n2102), .B(_abc_43815_n1425_1_bF_buf2), .Y(_abc_43815_n2103) );
  AND2X2 AND2X2_78 ( .A(_abc_43815_n694), .B(\mem_dat_i[19] ), .Y(_abc_43815_n747) );
  AND2X2 AND2X2_780 ( .A(_abc_43815_n2103), .B(_abc_43815_n2101_1), .Y(_abc_43815_n2104) );
  AND2X2 AND2X2_781 ( .A(_abc_43815_n1065_1_bF_buf3), .B(epc_q_18_), .Y(_abc_43815_n2105) );
  AND2X2 AND2X2_782 ( .A(_abc_43815_n2107), .B(_abc_43815_n2092), .Y(_abc_43815_n2108) );
  AND2X2 AND2X2_783 ( .A(_abc_43815_n2109), .B(_abc_43815_n2110), .Y(_abc_43815_n2111) );
  AND2X2 AND2X2_784 ( .A(_abc_43815_n1418_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_43815_n2113) );
  AND2X2 AND2X2_785 ( .A(_abc_43815_n1489_bF_buf2), .B(epc_q_18_), .Y(_abc_43815_n2114) );
  AND2X2 AND2X2_786 ( .A(_abc_43815_n2116), .B(_abc_43815_n1351_bF_buf3), .Y(_abc_43815_n2117) );
  AND2X2 AND2X2_787 ( .A(_abc_43815_n2112), .B(_abc_43815_n2117), .Y(_abc_43815_n2118) );
  AND2X2 AND2X2_788 ( .A(_abc_43815_n2120), .B(enable_i_bF_buf5), .Y(_abc_43815_n2121) );
  AND2X2 AND2X2_789 ( .A(_abc_43815_n2119), .B(_abc_43815_n2121), .Y(epc_q_18__FF_INPUT) );
  AND2X2 AND2X2_79 ( .A(_abc_43815_n697), .B(\mem_dat_i[3] ), .Y(_abc_43815_n748) );
  AND2X2 AND2X2_790 ( .A(_abc_43815_n2087_1), .B(pc_q_19_), .Y(_abc_43815_n2124) );
  AND2X2 AND2X2_791 ( .A(_abc_43815_n2125), .B(_abc_43815_n2123), .Y(_abc_43815_n2126) );
  AND2X2 AND2X2_792 ( .A(_abc_43815_n2126), .B(_abc_43815_n1461_bF_buf3), .Y(_abc_43815_n2127) );
  AND2X2 AND2X2_793 ( .A(_abc_43815_n2101_1), .B(_abc_43815_n2098), .Y(_abc_43815_n2129_1) );
  AND2X2 AND2X2_794 ( .A(pc_q_19_), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(_abc_43815_n2132) );
  AND2X2 AND2X2_795 ( .A(_abc_43815_n2133), .B(_abc_43815_n2131), .Y(_abc_43815_n2134) );
  AND2X2 AND2X2_796 ( .A(_abc_43815_n2137), .B(_abc_43815_n1425_1_bF_buf1), .Y(_abc_43815_n2138) );
  AND2X2 AND2X2_797 ( .A(_abc_43815_n2138), .B(_abc_43815_n2135), .Y(_abc_43815_n2139) );
  AND2X2 AND2X2_798 ( .A(_abc_43815_n1065_1_bF_buf2), .B(epc_q_19_), .Y(_abc_43815_n2140) );
  AND2X2 AND2X2_799 ( .A(_abc_43815_n1472_1_bF_buf1), .B(_abc_43815_n2143_1), .Y(_abc_43815_n2144) );
  AND2X2 AND2X2_8 ( .A(_abc_43815_n631), .B(opcode_q_24_), .Y(_abc_43815_n632) );
  AND2X2 AND2X2_80 ( .A(_abc_43815_n749), .B(_abc_43815_n686_1_bF_buf1), .Y(_abc_43815_n750) );
  AND2X2 AND2X2_800 ( .A(_abc_43815_n2142), .B(_abc_43815_n2144), .Y(_abc_43815_n2145) );
  AND2X2 AND2X2_801 ( .A(_abc_43815_n2126), .B(_abc_43815_n1473_bF_buf2), .Y(_abc_43815_n2146) );
  AND2X2 AND2X2_802 ( .A(_abc_43815_n1418_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_43815_n2149) );
  AND2X2 AND2X2_803 ( .A(_abc_43815_n1489_bF_buf1), .B(epc_q_19_), .Y(_abc_43815_n2150) );
  AND2X2 AND2X2_804 ( .A(_abc_43815_n2152), .B(_abc_43815_n1351_bF_buf2), .Y(_abc_43815_n2153) );
  AND2X2 AND2X2_805 ( .A(_abc_43815_n2148), .B(_abc_43815_n2153), .Y(_abc_43815_n2154) );
  AND2X2 AND2X2_806 ( .A(_abc_43815_n2156), .B(enable_i_bF_buf4), .Y(_abc_43815_n2157) );
  AND2X2 AND2X2_807 ( .A(_abc_43815_n2155), .B(_abc_43815_n2157), .Y(epc_q_19__FF_INPUT) );
  AND2X2 AND2X2_808 ( .A(_abc_43815_n2124), .B(pc_q_20_), .Y(_abc_43815_n2160) );
  AND2X2 AND2X2_809 ( .A(_abc_43815_n2161), .B(_abc_43815_n2159), .Y(_abc_43815_n2162) );
  AND2X2 AND2X2_81 ( .A(_abc_43815_n689), .B(\mem_dat_i[27] ), .Y(_abc_43815_n751) );
  AND2X2 AND2X2_810 ( .A(_abc_43815_n2162), .B(_abc_43815_n1461_bF_buf2), .Y(_abc_43815_n2163) );
  AND2X2 AND2X2_811 ( .A(_abc_43815_n2099), .B(_abc_43815_n2134), .Y(_abc_43815_n2165) );
  AND2X2 AND2X2_812 ( .A(_abc_43815_n2064), .B(_abc_43815_n2165), .Y(_abc_43815_n2166) );
  AND2X2 AND2X2_813 ( .A(_abc_43815_n2022), .B(_abc_43815_n2166), .Y(_abc_43815_n2167) );
  AND2X2 AND2X2_814 ( .A(_abc_43815_n2168), .B(_abc_43815_n2165), .Y(_abc_43815_n2169) );
  AND2X2 AND2X2_815 ( .A(_abc_43815_n2131), .B(_abc_43815_n2097), .Y(_abc_43815_n2170) );
  AND2X2 AND2X2_816 ( .A(pc_q_20_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(_abc_43815_n2175) );
  AND2X2 AND2X2_817 ( .A(_abc_43815_n2176), .B(_abc_43815_n2174), .Y(_abc_43815_n2177) );
  AND2X2 AND2X2_818 ( .A(_abc_43815_n2173_1), .B(_abc_43815_n2177), .Y(_abc_43815_n2179) );
  AND2X2 AND2X2_819 ( .A(_abc_43815_n2180), .B(_abc_43815_n1425_1_bF_buf0), .Y(_abc_43815_n2181) );
  AND2X2 AND2X2_82 ( .A(_abc_43815_n696), .B(\mem_dat_i[11] ), .Y(_abc_43815_n752) );
  AND2X2 AND2X2_820 ( .A(_abc_43815_n2181), .B(_abc_43815_n2178), .Y(_abc_43815_n2182) );
  AND2X2 AND2X2_821 ( .A(_abc_43815_n1065_1_bF_buf1), .B(epc_q_20_), .Y(_abc_43815_n2183) );
  AND2X2 AND2X2_822 ( .A(_abc_43815_n2185), .B(_abc_43815_n2186), .Y(_abc_43815_n2187) );
  AND2X2 AND2X2_823 ( .A(_abc_43815_n2187), .B(_abc_43815_n1472_1_bF_buf0), .Y(_abc_43815_n2188_1) );
  AND2X2 AND2X2_824 ( .A(_abc_43815_n2162), .B(_abc_43815_n1473_bF_buf1), .Y(_abc_43815_n2189) );
  AND2X2 AND2X2_825 ( .A(_abc_43815_n1418_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_43815_n2192) );
  AND2X2 AND2X2_826 ( .A(_abc_43815_n1489_bF_buf0), .B(epc_q_20_), .Y(_abc_43815_n2193) );
  AND2X2 AND2X2_827 ( .A(_abc_43815_n2195), .B(_abc_43815_n1351_bF_buf1), .Y(_abc_43815_n2196) );
  AND2X2 AND2X2_828 ( .A(_abc_43815_n2191), .B(_abc_43815_n2196), .Y(_abc_43815_n2197) );
  AND2X2 AND2X2_829 ( .A(_abc_43815_n2199), .B(enable_i_bF_buf3), .Y(_abc_43815_n2200) );
  AND2X2 AND2X2_83 ( .A(_abc_43815_n704), .B(\mem_dat_i[19] ), .Y(_abc_43815_n754_1) );
  AND2X2 AND2X2_830 ( .A(_abc_43815_n2198), .B(_abc_43815_n2200), .Y(epc_q_20__FF_INPUT) );
  AND2X2 AND2X2_831 ( .A(_abc_43815_n2160), .B(pc_q_21_), .Y(_abc_43815_n2203_1) );
  AND2X2 AND2X2_832 ( .A(_abc_43815_n2204), .B(_abc_43815_n2202), .Y(_abc_43815_n2205) );
  AND2X2 AND2X2_833 ( .A(_abc_43815_n2205), .B(_abc_43815_n1461_bF_buf1), .Y(_abc_43815_n2206) );
  AND2X2 AND2X2_834 ( .A(pc_q_21_), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(_abc_43815_n2210) );
  AND2X2 AND2X2_835 ( .A(_abc_43815_n2211), .B(_abc_43815_n2209), .Y(_abc_43815_n2212) );
  AND2X2 AND2X2_836 ( .A(_abc_43815_n2177), .B(_abc_43815_n2212), .Y(_abc_43815_n2215) );
  AND2X2 AND2X2_837 ( .A(_abc_43815_n2173_1), .B(_abc_43815_n2215), .Y(_abc_43815_n2216) );
  AND2X2 AND2X2_838 ( .A(_abc_43815_n2212), .B(_abc_43815_n2175), .Y(_abc_43815_n2217) );
  AND2X2 AND2X2_839 ( .A(_abc_43815_n2219), .B(_abc_43815_n1425_1_bF_buf4), .Y(_abc_43815_n2220) );
  AND2X2 AND2X2_84 ( .A(_abc_43815_n706_1), .B(\mem_dat_i[3] ), .Y(_abc_43815_n755) );
  AND2X2 AND2X2_840 ( .A(_abc_43815_n2220), .B(_abc_43815_n2214), .Y(_abc_43815_n2221) );
  AND2X2 AND2X2_841 ( .A(_abc_43815_n1065_1_bF_buf0), .B(epc_q_21_), .Y(_abc_43815_n2222_1) );
  AND2X2 AND2X2_842 ( .A(_abc_43815_n2224), .B(_abc_43815_n2208), .Y(_abc_43815_n2225) );
  AND2X2 AND2X2_843 ( .A(_abc_43815_n2226), .B(_abc_43815_n2227), .Y(_abc_43815_n2228) );
  AND2X2 AND2X2_844 ( .A(_abc_43815_n1418_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_43815_n2230) );
  AND2X2 AND2X2_845 ( .A(_abc_43815_n1489_bF_buf4), .B(epc_q_21_), .Y(_abc_43815_n2231) );
  AND2X2 AND2X2_846 ( .A(_abc_43815_n2233), .B(_abc_43815_n1351_bF_buf0), .Y(_abc_43815_n2234) );
  AND2X2 AND2X2_847 ( .A(_abc_43815_n2229), .B(_abc_43815_n2234), .Y(_abc_43815_n2235) );
  AND2X2 AND2X2_848 ( .A(_abc_43815_n2237), .B(enable_i_bF_buf2), .Y(_abc_43815_n2238) );
  AND2X2 AND2X2_849 ( .A(_abc_43815_n2236), .B(_abc_43815_n2238), .Y(epc_q_21__FF_INPUT) );
  AND2X2 AND2X2_85 ( .A(_abc_43815_n757), .B(_abc_43815_n685), .Y(_abc_43815_n758) );
  AND2X2 AND2X2_850 ( .A(_abc_43815_n2203_1), .B(pc_q_22_), .Y(_abc_43815_n2241) );
  AND2X2 AND2X2_851 ( .A(_abc_43815_n2242_1), .B(_abc_43815_n2240), .Y(_abc_43815_n2243) );
  AND2X2 AND2X2_852 ( .A(_abc_43815_n2243), .B(_abc_43815_n1461_bF_buf0), .Y(_abc_43815_n2244) );
  AND2X2 AND2X2_853 ( .A(_abc_43815_n2219), .B(_abc_43815_n2211), .Y(_abc_43815_n2247) );
  AND2X2 AND2X2_854 ( .A(pc_q_22_), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(_abc_43815_n2250) );
  AND2X2 AND2X2_855 ( .A(_abc_43815_n2251), .B(_abc_43815_n2249), .Y(_abc_43815_n2252_1) );
  AND2X2 AND2X2_856 ( .A(_abc_43815_n2248), .B(_abc_43815_n2252_1), .Y(_abc_43815_n2253) );
  AND2X2 AND2X2_857 ( .A(_abc_43815_n2255), .B(_abc_43815_n1425_1_bF_buf3), .Y(_abc_43815_n2256) );
  AND2X2 AND2X2_858 ( .A(_abc_43815_n2256), .B(_abc_43815_n2254), .Y(_abc_43815_n2257) );
  AND2X2 AND2X2_859 ( .A(_abc_43815_n1065_1_bF_buf4), .B(epc_q_22_), .Y(_abc_43815_n2258) );
  AND2X2 AND2X2_86 ( .A(_abc_43815_n759), .B(state_q_1_bF_buf3), .Y(_abc_43815_n760_1) );
  AND2X2 AND2X2_860 ( .A(_abc_43815_n2260), .B(_abc_43815_n2261), .Y(_abc_43815_n2262_1) );
  AND2X2 AND2X2_861 ( .A(_abc_43815_n2263), .B(_abc_43815_n2246), .Y(_abc_43815_n2264) );
  AND2X2 AND2X2_862 ( .A(_abc_43815_n1418_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_43815_n2266) );
  AND2X2 AND2X2_863 ( .A(_abc_43815_n1489_bF_buf3), .B(epc_q_22_), .Y(_abc_43815_n2267) );
  AND2X2 AND2X2_864 ( .A(_abc_43815_n2269), .B(_abc_43815_n1351_bF_buf4), .Y(_abc_43815_n2270) );
  AND2X2 AND2X2_865 ( .A(_abc_43815_n2265), .B(_abc_43815_n2270), .Y(_abc_43815_n2271) );
  AND2X2 AND2X2_866 ( .A(_abc_43815_n2273), .B(enable_i_bF_buf1), .Y(_abc_43815_n2274) );
  AND2X2 AND2X2_867 ( .A(_abc_43815_n2272_1), .B(_abc_43815_n2274), .Y(epc_q_22__FF_INPUT) );
  AND2X2 AND2X2_868 ( .A(_abc_43815_n2241), .B(pc_q_23_), .Y(_abc_43815_n2277) );
  AND2X2 AND2X2_869 ( .A(_abc_43815_n2278), .B(_abc_43815_n2276), .Y(_abc_43815_n2279) );
  AND2X2 AND2X2_87 ( .A(_abc_43815_n682), .B(alu_p_o_4_), .Y(_abc_43815_n762) );
  AND2X2 AND2X2_870 ( .A(_abc_43815_n2279), .B(_abc_43815_n1461_bF_buf3), .Y(_abc_43815_n2280) );
  AND2X2 AND2X2_871 ( .A(opcode_q_21_), .B(pc_q_23_), .Y(_abc_43815_n2285) );
  AND2X2 AND2X2_872 ( .A(_abc_43815_n2286), .B(_abc_43815_n2284), .Y(_abc_43815_n2287) );
  AND2X2 AND2X2_873 ( .A(_abc_43815_n2290), .B(_abc_43815_n1425_1_bF_buf2), .Y(_abc_43815_n2291) );
  AND2X2 AND2X2_874 ( .A(_abc_43815_n2291), .B(_abc_43815_n2289), .Y(_abc_43815_n2292_1) );
  AND2X2 AND2X2_875 ( .A(_abc_43815_n1065_1_bF_buf3), .B(epc_q_23_), .Y(_abc_43815_n2293) );
  AND2X2 AND2X2_876 ( .A(_abc_43815_n2295), .B(_abc_43815_n2296), .Y(_abc_43815_n2297) );
  AND2X2 AND2X2_877 ( .A(_abc_43815_n2298), .B(_abc_43815_n2299), .Y(_abc_43815_n2300) );
  AND2X2 AND2X2_878 ( .A(_abc_43815_n1418_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_43815_n2302_1) );
  AND2X2 AND2X2_879 ( .A(_abc_43815_n1489_bF_buf2), .B(epc_q_23_), .Y(_abc_43815_n2303) );
  AND2X2 AND2X2_88 ( .A(_abc_43815_n694), .B(\mem_dat_i[20] ), .Y(_abc_43815_n763) );
  AND2X2 AND2X2_880 ( .A(_abc_43815_n2305), .B(_abc_43815_n1351_bF_buf3), .Y(_abc_43815_n2306) );
  AND2X2 AND2X2_881 ( .A(_abc_43815_n2301), .B(_abc_43815_n2306), .Y(_abc_43815_n2307) );
  AND2X2 AND2X2_882 ( .A(_abc_43815_n2309), .B(enable_i_bF_buf0), .Y(_abc_43815_n2310) );
  AND2X2 AND2X2_883 ( .A(_abc_43815_n2308), .B(_abc_43815_n2310), .Y(epc_q_23__FF_INPUT) );
  AND2X2 AND2X2_884 ( .A(_abc_43815_n2277), .B(pc_q_24_), .Y(_abc_43815_n2313) );
  AND2X2 AND2X2_885 ( .A(_abc_43815_n2314), .B(_abc_43815_n2312_1), .Y(_abc_43815_n2315) );
  AND2X2 AND2X2_886 ( .A(_abc_43815_n2315), .B(_abc_43815_n1461_bF_buf2), .Y(_abc_43815_n2316) );
  AND2X2 AND2X2_887 ( .A(_abc_43815_n2252_1), .B(_abc_43815_n2287), .Y(_abc_43815_n2319) );
  AND2X2 AND2X2_888 ( .A(_abc_43815_n2318), .B(_abc_43815_n2319), .Y(_abc_43815_n2320) );
  AND2X2 AND2X2_889 ( .A(_abc_43815_n2284), .B(_abc_43815_n2250), .Y(_abc_43815_n2321) );
  AND2X2 AND2X2_89 ( .A(_abc_43815_n697), .B(\mem_dat_i[4] ), .Y(_abc_43815_n764) );
  AND2X2 AND2X2_890 ( .A(_abc_43815_n2215), .B(_abc_43815_n2319), .Y(_abc_43815_n2324) );
  AND2X2 AND2X2_891 ( .A(_abc_43815_n2173_1), .B(_abc_43815_n2324), .Y(_abc_43815_n2325) );
  AND2X2 AND2X2_892 ( .A(opcode_q_22_), .B(pc_q_24_), .Y(_abc_43815_n2328) );
  AND2X2 AND2X2_893 ( .A(_abc_43815_n2329), .B(_abc_43815_n2327), .Y(_abc_43815_n2330) );
  AND2X2 AND2X2_894 ( .A(_abc_43815_n2326), .B(_abc_43815_n2330), .Y(_abc_43815_n2331) );
  AND2X2 AND2X2_895 ( .A(_abc_43815_n2333), .B(_abc_43815_n1425_1_bF_buf1), .Y(_abc_43815_n2334) );
  AND2X2 AND2X2_896 ( .A(_abc_43815_n2334), .B(_abc_43815_n2332_1), .Y(_abc_43815_n2335) );
  AND2X2 AND2X2_897 ( .A(_abc_43815_n1065_1_bF_buf2), .B(epc_q_24_), .Y(_abc_43815_n2336) );
  AND2X2 AND2X2_898 ( .A(_abc_43815_n2338), .B(_abc_43815_n2339), .Y(_abc_43815_n2340) );
  AND2X2 AND2X2_899 ( .A(_abc_43815_n2341), .B(_abc_43815_n2342_1), .Y(_abc_43815_n2343) );
  AND2X2 AND2X2_9 ( .A(_abc_43815_n628), .B(_abc_43815_n632), .Y(inst_trap_w) );
  AND2X2 AND2X2_90 ( .A(_abc_43815_n765_1), .B(_abc_43815_n686_1_bF_buf0), .Y(_abc_43815_n766) );
  AND2X2 AND2X2_900 ( .A(_abc_43815_n1418_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_43815_n2345) );
  AND2X2 AND2X2_901 ( .A(_abc_43815_n1489_bF_buf1), .B(epc_q_24_), .Y(_abc_43815_n2346) );
  AND2X2 AND2X2_902 ( .A(_abc_43815_n2348), .B(_abc_43815_n1351_bF_buf2), .Y(_abc_43815_n2349) );
  AND2X2 AND2X2_903 ( .A(_abc_43815_n2344), .B(_abc_43815_n2349), .Y(_abc_43815_n2350) );
  AND2X2 AND2X2_904 ( .A(_abc_43815_n2352_1), .B(enable_i_bF_buf7), .Y(_abc_43815_n2353) );
  AND2X2 AND2X2_905 ( .A(_abc_43815_n2351), .B(_abc_43815_n2353), .Y(epc_q_24__FF_INPUT) );
  AND2X2 AND2X2_906 ( .A(_abc_43815_n2313), .B(pc_q_25_), .Y(_abc_43815_n2356) );
  AND2X2 AND2X2_907 ( .A(_abc_43815_n2357), .B(_abc_43815_n2355), .Y(_abc_43815_n2358) );
  AND2X2 AND2X2_908 ( .A(_abc_43815_n2358), .B(_abc_43815_n1461_bF_buf1), .Y(_abc_43815_n2359) );
  AND2X2 AND2X2_909 ( .A(opcode_q_23_), .B(pc_q_25_), .Y(_abc_43815_n2362_1) );
  AND2X2 AND2X2_91 ( .A(_abc_43815_n689), .B(\mem_dat_i[28] ), .Y(_abc_43815_n767) );
  AND2X2 AND2X2_910 ( .A(_abc_43815_n2363), .B(_abc_43815_n2361), .Y(_abc_43815_n2364) );
  AND2X2 AND2X2_911 ( .A(_abc_43815_n2330), .B(_abc_43815_n2364), .Y(_abc_43815_n2367) );
  AND2X2 AND2X2_912 ( .A(_abc_43815_n2326), .B(_abc_43815_n2367), .Y(_abc_43815_n2368) );
  AND2X2 AND2X2_913 ( .A(_abc_43815_n2364), .B(_abc_43815_n2328), .Y(_abc_43815_n2370) );
  AND2X2 AND2X2_914 ( .A(_abc_43815_n1425_1_bF_buf0), .B(_abc_43815_n2371), .Y(_abc_43815_n2372_1) );
  AND2X2 AND2X2_915 ( .A(_abc_43815_n2369), .B(_abc_43815_n2372_1), .Y(_abc_43815_n2373) );
  AND2X2 AND2X2_916 ( .A(_abc_43815_n2373), .B(_abc_43815_n2366), .Y(_abc_43815_n2374) );
  AND2X2 AND2X2_917 ( .A(_abc_43815_n1065_1_bF_buf1), .B(epc_q_25_), .Y(_abc_43815_n2375) );
  AND2X2 AND2X2_918 ( .A(_abc_43815_n2377), .B(_abc_43815_n2378), .Y(_abc_43815_n2379) );
  AND2X2 AND2X2_919 ( .A(_abc_43815_n2381), .B(_abc_43815_n2380), .Y(_abc_43815_n2382) );
  AND2X2 AND2X2_92 ( .A(_abc_43815_n696), .B(\mem_dat_i[12] ), .Y(_abc_43815_n768) );
  AND2X2 AND2X2_920 ( .A(_abc_43815_n1418_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_43815_n2384) );
  AND2X2 AND2X2_921 ( .A(_abc_43815_n1489_bF_buf0), .B(epc_q_25_), .Y(_abc_43815_n2385) );
  AND2X2 AND2X2_922 ( .A(_abc_43815_n2387), .B(_abc_43815_n1351_bF_buf1), .Y(_abc_43815_n2388) );
  AND2X2 AND2X2_923 ( .A(_abc_43815_n2383), .B(_abc_43815_n2388), .Y(_abc_43815_n2389) );
  AND2X2 AND2X2_924 ( .A(_abc_43815_n2391), .B(enable_i_bF_buf6), .Y(_abc_43815_n2392) );
  AND2X2 AND2X2_925 ( .A(_abc_43815_n2390), .B(_abc_43815_n2392), .Y(epc_q_25__FF_INPUT) );
  AND2X2 AND2X2_926 ( .A(_abc_43815_n2356), .B(pc_q_26_), .Y(_abc_43815_n2395) );
  AND2X2 AND2X2_927 ( .A(_abc_43815_n2396_1), .B(_abc_43815_n2394), .Y(_abc_43815_n2397) );
  AND2X2 AND2X2_928 ( .A(_abc_43815_n2397), .B(_abc_43815_n1461_bF_buf0), .Y(_abc_43815_n2398) );
  AND2X2 AND2X2_929 ( .A(_abc_43815_n2371), .B(_abc_43815_n2363), .Y(_abc_43815_n2400) );
  AND2X2 AND2X2_93 ( .A(_abc_43815_n704), .B(\mem_dat_i[20] ), .Y(_abc_43815_n770) );
  AND2X2 AND2X2_930 ( .A(_abc_43815_n2369), .B(_abc_43815_n2400), .Y(_abc_43815_n2401) );
  AND2X2 AND2X2_931 ( .A(opcode_q_24_), .B(pc_q_26_), .Y(_abc_43815_n2404) );
  AND2X2 AND2X2_932 ( .A(_abc_43815_n2405), .B(_abc_43815_n2403), .Y(_abc_43815_n2406) );
  AND2X2 AND2X2_933 ( .A(_abc_43815_n2402), .B(_abc_43815_n2406), .Y(_abc_43815_n2407) );
  AND2X2 AND2X2_934 ( .A(_abc_43815_n2409), .B(_abc_43815_n1425_1_bF_buf4), .Y(_abc_43815_n2410) );
  AND2X2 AND2X2_935 ( .A(_abc_43815_n2410), .B(_abc_43815_n2408), .Y(_abc_43815_n2411) );
  AND2X2 AND2X2_936 ( .A(_abc_43815_n1065_1_bF_buf0), .B(epc_q_26_), .Y(_abc_43815_n2412) );
  AND2X2 AND2X2_937 ( .A(_abc_43815_n2414), .B(_abc_43815_n2415), .Y(_abc_43815_n2416) );
  AND2X2 AND2X2_938 ( .A(_abc_43815_n2417), .B(_abc_43815_n2418), .Y(_abc_43815_n2419) );
  AND2X2 AND2X2_939 ( .A(_abc_43815_n1418_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_43815_n2421) );
  AND2X2 AND2X2_94 ( .A(_abc_43815_n706_1), .B(\mem_dat_i[4] ), .Y(_abc_43815_n771) );
  AND2X2 AND2X2_940 ( .A(_abc_43815_n1489_bF_buf4), .B(epc_q_26_), .Y(_abc_43815_n2422) );
  AND2X2 AND2X2_941 ( .A(_abc_43815_n2424), .B(_abc_43815_n1351_bF_buf0), .Y(_abc_43815_n2425) );
  AND2X2 AND2X2_942 ( .A(_abc_43815_n2420_1), .B(_abc_43815_n2425), .Y(_abc_43815_n2426) );
  AND2X2 AND2X2_943 ( .A(_abc_43815_n2428), .B(enable_i_bF_buf5), .Y(_abc_43815_n2429) );
  AND2X2 AND2X2_944 ( .A(_abc_43815_n2427), .B(_abc_43815_n2429), .Y(epc_q_26__FF_INPUT) );
  AND2X2 AND2X2_945 ( .A(_abc_43815_n2395), .B(pc_q_27_), .Y(_abc_43815_n2432) );
  AND2X2 AND2X2_946 ( .A(_abc_43815_n2433), .B(_abc_43815_n2431), .Y(_abc_43815_n2434) );
  AND2X2 AND2X2_947 ( .A(_abc_43815_n2434), .B(_abc_43815_n1461_bF_buf3), .Y(_abc_43815_n2435) );
  AND2X2 AND2X2_948 ( .A(opcode_q_25_), .B(pc_q_27_), .Y(_abc_43815_n2438) );
  AND2X2 AND2X2_949 ( .A(_abc_43815_n2439), .B(_abc_43815_n2437), .Y(_abc_43815_n2440) );
  AND2X2 AND2X2_95 ( .A(_abc_43815_n773), .B(_abc_43815_n685), .Y(_abc_43815_n774) );
  AND2X2 AND2X2_950 ( .A(_abc_43815_n2406), .B(_abc_43815_n2440), .Y(_abc_43815_n2443) );
  AND2X2 AND2X2_951 ( .A(_abc_43815_n2440), .B(_abc_43815_n2404), .Y(_abc_43815_n2446) );
  AND2X2 AND2X2_952 ( .A(_abc_43815_n1425_1_bF_buf3), .B(_abc_43815_n2447), .Y(_abc_43815_n2448) );
  AND2X2 AND2X2_953 ( .A(_abc_43815_n2445_1), .B(_abc_43815_n2448), .Y(_abc_43815_n2449) );
  AND2X2 AND2X2_954 ( .A(_abc_43815_n2442), .B(_abc_43815_n2449), .Y(_abc_43815_n2450) );
  AND2X2 AND2X2_955 ( .A(_abc_43815_n1065_1_bF_buf4), .B(epc_q_27_), .Y(_abc_43815_n2451) );
  AND2X2 AND2X2_956 ( .A(_abc_43815_n2453), .B(_abc_43815_n2454), .Y(_abc_43815_n2455) );
  AND2X2 AND2X2_957 ( .A(_abc_43815_n2456), .B(_abc_43815_n2457), .Y(_abc_43815_n2458) );
  AND2X2 AND2X2_958 ( .A(_abc_43815_n1418_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_43815_n2460) );
  AND2X2 AND2X2_959 ( .A(_abc_43815_n1489_bF_buf3), .B(epc_q_27_), .Y(_abc_43815_n2461) );
  AND2X2 AND2X2_96 ( .A(_abc_43815_n775), .B(state_q_1_bF_buf2), .Y(_abc_43815_n776) );
  AND2X2 AND2X2_960 ( .A(_abc_43815_n2463), .B(_abc_43815_n1351_bF_buf4), .Y(_abc_43815_n2464) );
  AND2X2 AND2X2_961 ( .A(_abc_43815_n2459), .B(_abc_43815_n2464), .Y(_abc_43815_n2465) );
  AND2X2 AND2X2_962 ( .A(_abc_43815_n2467), .B(enable_i_bF_buf4), .Y(_abc_43815_n2468) );
  AND2X2 AND2X2_963 ( .A(_abc_43815_n2466), .B(_abc_43815_n2468), .Y(epc_q_27__FF_INPUT) );
  AND2X2 AND2X2_964 ( .A(_abc_43815_n2432), .B(pc_q_28_), .Y(_abc_43815_n2471) );
  AND2X2 AND2X2_965 ( .A(_abc_43815_n2472), .B(_abc_43815_n2470), .Y(_abc_43815_n2473) );
  AND2X2 AND2X2_966 ( .A(_abc_43815_n2473), .B(_abc_43815_n1461_bF_buf2), .Y(_abc_43815_n2474) );
  AND2X2 AND2X2_967 ( .A(_abc_43815_n2447), .B(_abc_43815_n2439), .Y(_abc_43815_n2476) );
  AND2X2 AND2X2_968 ( .A(_abc_43815_n2477), .B(_abc_43815_n2476), .Y(_abc_43815_n2478) );
  AND2X2 AND2X2_969 ( .A(_abc_43815_n2367), .B(_abc_43815_n2443), .Y(_abc_43815_n2480) );
  AND2X2 AND2X2_97 ( .A(_abc_43815_n682), .B(alu_p_o_5_), .Y(_abc_43815_n778) );
  AND2X2 AND2X2_970 ( .A(_abc_43815_n2326), .B(_abc_43815_n2480), .Y(_abc_43815_n2481) );
  AND2X2 AND2X2_971 ( .A(opcode_q_25_), .B(pc_q_28_), .Y(_abc_43815_n2484) );
  AND2X2 AND2X2_972 ( .A(_abc_43815_n2485), .B(_abc_43815_n2483), .Y(_abc_43815_n2486) );
  AND2X2 AND2X2_973 ( .A(_abc_43815_n2482), .B(_abc_43815_n2486), .Y(_abc_43815_n2487) );
  AND2X2 AND2X2_974 ( .A(_abc_43815_n2489), .B(_abc_43815_n1425_1_bF_buf2), .Y(_abc_43815_n2490) );
  AND2X2 AND2X2_975 ( .A(_abc_43815_n2490), .B(_abc_43815_n2488), .Y(_abc_43815_n2491) );
  AND2X2 AND2X2_976 ( .A(_abc_43815_n1065_1_bF_buf3), .B(epc_q_28_), .Y(_abc_43815_n2492) );
  AND2X2 AND2X2_977 ( .A(_abc_43815_n2494), .B(_abc_43815_n2495), .Y(_abc_43815_n2496) );
  AND2X2 AND2X2_978 ( .A(_abc_43815_n2498), .B(_abc_43815_n2497), .Y(_abc_43815_n2499) );
  AND2X2 AND2X2_979 ( .A(_abc_43815_n1418_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_43815_n2501) );
  AND2X2 AND2X2_98 ( .A(_abc_43815_n694), .B(\mem_dat_i[21] ), .Y(_abc_43815_n779) );
  AND2X2 AND2X2_980 ( .A(_abc_43815_n1489_bF_buf2), .B(epc_q_28_), .Y(_abc_43815_n2502) );
  AND2X2 AND2X2_981 ( .A(_abc_43815_n2504), .B(_abc_43815_n1351_bF_buf3), .Y(_abc_43815_n2505) );
  AND2X2 AND2X2_982 ( .A(_abc_43815_n2500), .B(_abc_43815_n2505), .Y(_abc_43815_n2506) );
  AND2X2 AND2X2_983 ( .A(_abc_43815_n2508), .B(enable_i_bF_buf3), .Y(_abc_43815_n2509) );
  AND2X2 AND2X2_984 ( .A(_abc_43815_n2507), .B(_abc_43815_n2509), .Y(epc_q_28__FF_INPUT) );
  AND2X2 AND2X2_985 ( .A(_abc_43815_n2471), .B(pc_q_29_), .Y(_abc_43815_n2512) );
  AND2X2 AND2X2_986 ( .A(_abc_43815_n2513), .B(_abc_43815_n2511), .Y(_abc_43815_n2514) );
  AND2X2 AND2X2_987 ( .A(_abc_43815_n2514), .B(_abc_43815_n1461_bF_buf1), .Y(_abc_43815_n2515) );
  AND2X2 AND2X2_988 ( .A(opcode_q_25_), .B(pc_q_29_), .Y(_abc_43815_n2520) );
  AND2X2 AND2X2_989 ( .A(_abc_43815_n2521), .B(_abc_43815_n2519), .Y(_abc_43815_n2522) );
  AND2X2 AND2X2_99 ( .A(_abc_43815_n697), .B(\mem_dat_i[5] ), .Y(_abc_43815_n780) );
  AND2X2 AND2X2_990 ( .A(_abc_43815_n2525), .B(_abc_43815_n1425_1_bF_buf1), .Y(_abc_43815_n2526) );
  AND2X2 AND2X2_991 ( .A(_abc_43815_n2526), .B(_abc_43815_n2524), .Y(_abc_43815_n2527) );
  AND2X2 AND2X2_992 ( .A(_abc_43815_n1065_1_bF_buf2), .B(epc_q_29_), .Y(_abc_43815_n2528) );
  AND2X2 AND2X2_993 ( .A(_abc_43815_n2530), .B(_abc_43815_n2531), .Y(_abc_43815_n2532) );
  AND2X2 AND2X2_994 ( .A(_abc_43815_n2534), .B(_abc_43815_n2533), .Y(_abc_43815_n2535) );
  AND2X2 AND2X2_995 ( .A(_abc_43815_n1418_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_43815_n2537) );
  AND2X2 AND2X2_996 ( .A(_abc_43815_n1489_bF_buf1), .B(epc_q_29_), .Y(_abc_43815_n2538) );
  AND2X2 AND2X2_997 ( .A(_abc_43815_n2540), .B(_abc_43815_n1351_bF_buf2), .Y(_abc_43815_n2541_1) );
  AND2X2 AND2X2_998 ( .A(_abc_43815_n2536), .B(_abc_43815_n2541_1), .Y(_abc_43815_n2542) );
  AND2X2 AND2X2_999 ( .A(_abc_43815_n2544), .B(enable_i_bF_buf2), .Y(_abc_43815_n2545) );
  BUFX2 BUFX2_1 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8) );
  BUFX2 BUFX2_10 ( .A(_abc_43815_n4167_bF_buf15), .Y(_abc_43815_n4167_bF_buf15_bF_buf3) );
  BUFX2 BUFX2_100 ( .A(_abc_43815_n1431_1), .Y(_abc_43815_n1431_1_bF_buf1) );
  BUFX2 BUFX2_1000 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606), .Y(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf3) );
  BUFX2 BUFX2_1001 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606), .Y(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf2) );
  BUFX2 BUFX2_1002 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606), .Y(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf1) );
  BUFX2 BUFX2_1003 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606), .Y(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf0) );
  BUFX2 BUFX2_1004 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609), .Y(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf4) );
  BUFX2 BUFX2_1005 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609), .Y(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf3) );
  BUFX2 BUFX2_1006 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609), .Y(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf2) );
  BUFX2 BUFX2_1007 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609), .Y(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf1) );
  BUFX2 BUFX2_1008 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7609), .Y(REGFILE_SIM_reg_bank__abc_33898_n7609_bF_buf0) );
  BUFX2 BUFX2_1009 ( .A(alu__abc_41358_n927), .Y(alu__abc_41358_n927_bF_buf4) );
  BUFX2 BUFX2_101 ( .A(_abc_43815_n1431_1), .Y(_abc_43815_n1431_1_bF_buf0) );
  BUFX2 BUFX2_1010 ( .A(alu__abc_41358_n927), .Y(alu__abc_41358_n927_bF_buf3) );
  BUFX2 BUFX2_1011 ( .A(alu__abc_41358_n927), .Y(alu__abc_41358_n927_bF_buf2) );
  BUFX2 BUFX2_1012 ( .A(alu__abc_41358_n927), .Y(alu__abc_41358_n927_bF_buf1) );
  BUFX2 BUFX2_1013 ( .A(alu__abc_41358_n927), .Y(alu__abc_41358_n927_bF_buf0) );
  BUFX2 BUFX2_1014 ( .A(_abc_43815_n650), .Y(_abc_43815_n650_bF_buf4) );
  BUFX2 BUFX2_1015 ( .A(_abc_43815_n650), .Y(_abc_43815_n650_bF_buf3) );
  BUFX2 BUFX2_1016 ( .A(_abc_43815_n650), .Y(_abc_43815_n650_bF_buf2) );
  BUFX2 BUFX2_1017 ( .A(_abc_43815_n650), .Y(_abc_43815_n650_bF_buf1) );
  BUFX2 BUFX2_1018 ( .A(_abc_43815_n650), .Y(_abc_43815_n650_bF_buf0) );
  BUFX2 BUFX2_1019 ( .A(_abc_27555_n4367), .Y(_abc_27555_n4367_bF_buf7) );
  BUFX2 BUFX2_102 ( .A(_abc_43815_n1065_1), .Y(_abc_43815_n1065_1_bF_buf4) );
  BUFX2 BUFX2_1020 ( .A(_abc_27555_n4367), .Y(_abc_27555_n4367_bF_buf6) );
  BUFX2 BUFX2_1021 ( .A(_abc_27555_n4367), .Y(_abc_27555_n4367_bF_buf5) );
  BUFX2 BUFX2_1022 ( .A(_abc_27555_n4367), .Y(_abc_27555_n4367_bF_buf4) );
  BUFX2 BUFX2_1023 ( .A(_abc_27555_n4367), .Y(_abc_27555_n4367_bF_buf3) );
  BUFX2 BUFX2_1024 ( .A(_abc_27555_n4367), .Y(_abc_27555_n4367_bF_buf2) );
  BUFX2 BUFX2_1025 ( .A(_abc_27555_n4367), .Y(_abc_27555_n4367_bF_buf1) );
  BUFX2 BUFX2_1026 ( .A(_abc_27555_n4367), .Y(_abc_27555_n4367_bF_buf0) );
  BUFX2 BUFX2_1027 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574), .Y(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf4) );
  BUFX2 BUFX2_1028 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574), .Y(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf3) );
  BUFX2 BUFX2_1029 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574), .Y(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf2) );
  BUFX2 BUFX2_103 ( .A(_abc_43815_n1065_1), .Y(_abc_43815_n1065_1_bF_buf3) );
  BUFX2 BUFX2_1030 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574), .Y(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf1) );
  BUFX2 BUFX2_1031 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7574), .Y(REGFILE_SIM_reg_bank__abc_33898_n7574_bF_buf0) );
  BUFX2 BUFX2_1032 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577), .Y(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf4) );
  BUFX2 BUFX2_1033 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577), .Y(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf3) );
  BUFX2 BUFX2_1034 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577), .Y(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf2) );
  BUFX2 BUFX2_1035 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577), .Y(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf1) );
  BUFX2 BUFX2_1036 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7577), .Y(REGFILE_SIM_reg_bank__abc_33898_n7577_bF_buf0) );
  BUFX2 BUFX2_1037 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693), .Y(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4) );
  BUFX2 BUFX2_1038 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693), .Y(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3) );
  BUFX2 BUFX2_1039 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693), .Y(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2) );
  BUFX2 BUFX2_104 ( .A(_abc_43815_n1065_1), .Y(_abc_43815_n1065_1_bF_buf2) );
  BUFX2 BUFX2_1040 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693), .Y(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf1) );
  BUFX2 BUFX2_1041 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693), .Y(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf0) );
  BUFX2 BUFX2_1042 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695), .Y(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4) );
  BUFX2 BUFX2_1043 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695), .Y(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3) );
  BUFX2 BUFX2_1044 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695), .Y(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf2) );
  BUFX2 BUFX2_1045 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695), .Y(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf1) );
  BUFX2 BUFX2_1046 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695), .Y(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf0) );
  BUFX2 BUFX2_1047 ( .A(_abc_43815_n1171), .Y(_abc_43815_n1171_bF_buf5) );
  BUFX2 BUFX2_1048 ( .A(_abc_43815_n1171), .Y(_abc_43815_n1171_bF_buf4) );
  BUFX2 BUFX2_1049 ( .A(_abc_43815_n1171), .Y(_abc_43815_n1171_bF_buf3) );
  BUFX2 BUFX2_105 ( .A(_abc_43815_n1065_1), .Y(_abc_43815_n1065_1_bF_buf1) );
  BUFX2 BUFX2_1050 ( .A(_abc_43815_n1171), .Y(_abc_43815_n1171_bF_buf2) );
  BUFX2 BUFX2_1051 ( .A(_abc_43815_n1171), .Y(_abc_43815_n1171_bF_buf1) );
  BUFX2 BUFX2_1052 ( .A(_abc_43815_n1171), .Y(_abc_43815_n1171_bF_buf0) );
  BUFX2 BUFX2_1053 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3) );
  BUFX2 BUFX2_1054 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2) );
  BUFX2 BUFX2_1055 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1) );
  BUFX2 BUFX2_1056 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0) );
  BUFX2 BUFX2_1057 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632), .Y(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf4) );
  BUFX2 BUFX2_1058 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632), .Y(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf3) );
  BUFX2 BUFX2_1059 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632), .Y(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf2) );
  BUFX2 BUFX2_106 ( .A(_abc_43815_n1065_1), .Y(_abc_43815_n1065_1_bF_buf0) );
  BUFX2 BUFX2_1060 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632), .Y(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf1) );
  BUFX2 BUFX2_1061 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5632), .Y(REGFILE_SIM_reg_bank__abc_33898_n5632_bF_buf0) );
  BUFX2 BUFX2_1062 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634), .Y(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf4) );
  BUFX2 BUFX2_1063 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634), .Y(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf3) );
  BUFX2 BUFX2_1064 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634), .Y(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf2) );
  BUFX2 BUFX2_1065 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634), .Y(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf1) );
  BUFX2 BUFX2_1066 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5634), .Y(REGFILE_SIM_reg_bank__abc_33898_n5634_bF_buf0) );
  BUFX2 BUFX2_1067 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637), .Y(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf4) );
  BUFX2 BUFX2_1068 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637), .Y(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf3) );
  BUFX2 BUFX2_1069 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637), .Y(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf2) );
  BUFX2 BUFX2_107 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3) );
  BUFX2 BUFX2_1070 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637), .Y(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf1) );
  BUFX2 BUFX2_1071 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5637), .Y(REGFILE_SIM_reg_bank__abc_33898_n5637_bF_buf0) );
  BUFX2 BUFX2_1072 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639), .Y(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf4) );
  BUFX2 BUFX2_1073 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639), .Y(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf3) );
  BUFX2 BUFX2_1074 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639), .Y(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf2) );
  BUFX2 BUFX2_1075 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639), .Y(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf1) );
  BUFX2 BUFX2_1076 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5639), .Y(REGFILE_SIM_reg_bank__abc_33898_n5639_bF_buf0) );
  BUFX2 BUFX2_1077 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370), .Y(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4) );
  BUFX2 BUFX2_1078 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370), .Y(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3) );
  BUFX2 BUFX2_1079 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370), .Y(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf2) );
  BUFX2 BUFX2_108 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2) );
  BUFX2 BUFX2_1080 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370), .Y(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf1) );
  BUFX2 BUFX2_1081 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370), .Y(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf0) );
  BUFX2 BUFX2_1082 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4) );
  BUFX2 BUFX2_1083 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3) );
  BUFX2 BUFX2_1084 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf2) );
  BUFX2 BUFX2_1085 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf1) );
  BUFX2 BUFX2_1086 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf0) );
  BUFX2 BUFX2_1087 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4) );
  BUFX2 BUFX2_1088 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3) );
  BUFX2 BUFX2_1089 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf2) );
  BUFX2 BUFX2_109 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1) );
  BUFX2 BUFX2_1090 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf1) );
  BUFX2 BUFX2_1091 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf0) );
  BUFX2 BUFX2_1092 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3) );
  BUFX2 BUFX2_1093 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2) );
  BUFX2 BUFX2_1094 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1) );
  BUFX2 BUFX2_1095 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0) );
  BUFX2 BUFX2_1096 ( .A(_abc_43815_n2840), .Y(_abc_43815_n2840_bF_buf4) );
  BUFX2 BUFX2_1097 ( .A(_abc_43815_n2840), .Y(_abc_43815_n2840_bF_buf3) );
  BUFX2 BUFX2_1098 ( .A(_abc_43815_n2840), .Y(_abc_43815_n2840_bF_buf2) );
  BUFX2 BUFX2_1099 ( .A(_abc_43815_n2840), .Y(_abc_43815_n2840_bF_buf1) );
  BUFX2 BUFX2_11 ( .A(_abc_43815_n4167_bF_buf15), .Y(_abc_43815_n4167_bF_buf15_bF_buf2) );
  BUFX2 BUFX2_110 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0) );
  BUFX2 BUFX2_1100 ( .A(_abc_43815_n2840), .Y(_abc_43815_n2840_bF_buf0) );
  BUFX2 BUFX2_1101 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600), .Y(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf4) );
  BUFX2 BUFX2_1102 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600), .Y(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf3) );
  BUFX2 BUFX2_1103 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600), .Y(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf2) );
  BUFX2 BUFX2_1104 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600), .Y(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf1) );
  BUFX2 BUFX2_1105 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5600), .Y(REGFILE_SIM_reg_bank__abc_33898_n5600_bF_buf0) );
  BUFX2 BUFX2_1106 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603), .Y(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf4) );
  BUFX2 BUFX2_1107 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603), .Y(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf3) );
  BUFX2 BUFX2_1108 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603), .Y(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf2) );
  BUFX2 BUFX2_1109 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603), .Y(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf1) );
  BUFX2 BUFX2_111 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98) );
  BUFX2 BUFX2_1110 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5603), .Y(REGFILE_SIM_reg_bank__abc_33898_n5603_bF_buf0) );
  BUFX2 BUFX2_1111 ( .A(alu__abc_41358_n833), .Y(alu__abc_41358_n833_bF_buf4) );
  BUFX2 BUFX2_1112 ( .A(alu__abc_41358_n833), .Y(alu__abc_41358_n833_bF_buf3) );
  BUFX2 BUFX2_1113 ( .A(alu__abc_41358_n833), .Y(alu__abc_41358_n833_bF_buf2) );
  BUFX2 BUFX2_1114 ( .A(alu__abc_41358_n833), .Y(alu__abc_41358_n833_bF_buf1) );
  BUFX2 BUFX2_1115 ( .A(alu__abc_41358_n833), .Y(alu__abc_41358_n833_bF_buf0) );
  BUFX2 BUFX2_1116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7) );
  BUFX2 BUFX2_1117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf6) );
  BUFX2 BUFX2_1118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5) );
  BUFX2 BUFX2_1119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf4) );
  BUFX2 BUFX2_112 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97) );
  BUFX2 BUFX2_1120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3) );
  BUFX2 BUFX2_1121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf2) );
  BUFX2 BUFX2_1122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1) );
  BUFX2 BUFX2_1123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288), .Y(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf0) );
  BUFX2 BUFX2_1124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4) );
  BUFX2 BUFX2_1125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3) );
  BUFX2 BUFX2_1126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf2) );
  BUFX2 BUFX2_1127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf1) );
  BUFX2 BUFX2_1128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf0) );
  BUFX2 BUFX2_1129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573), .Y(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf4) );
  BUFX2 BUFX2_113 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96) );
  BUFX2 BUFX2_1130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573), .Y(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf3) );
  BUFX2 BUFX2_1131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573), .Y(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf2) );
  BUFX2 BUFX2_1132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573), .Y(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf1) );
  BUFX2 BUFX2_1133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5573), .Y(REGFILE_SIM_reg_bank__abc_33898_n5573_bF_buf0) );
  BUFX2 BUFX2_1134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576), .Y(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf4) );
  BUFX2 BUFX2_1135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576), .Y(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf3) );
  BUFX2 BUFX2_1136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576), .Y(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf2) );
  BUFX2 BUFX2_1137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576), .Y(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf1) );
  BUFX2 BUFX2_1138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5576), .Y(REGFILE_SIM_reg_bank__abc_33898_n5576_bF_buf0) );
  BUFX2 BUFX2_1139 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3) );
  BUFX2 BUFX2_114 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95) );
  BUFX2 BUFX2_1140 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2) );
  BUFX2 BUFX2_1141 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1) );
  BUFX2 BUFX2_1142 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0) );
  BUFX2 BUFX2_1143 ( .A(_abc_43815_n1461), .Y(_abc_43815_n1461_bF_buf3) );
  BUFX2 BUFX2_1144 ( .A(_abc_43815_n1461), .Y(_abc_43815_n1461_bF_buf2) );
  BUFX2 BUFX2_1145 ( .A(_abc_43815_n1461), .Y(_abc_43815_n1461_bF_buf1) );
  BUFX2 BUFX2_1146 ( .A(_abc_43815_n1461), .Y(_abc_43815_n1461_bF_buf0) );
  BUFX2 BUFX2_1147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545), .Y(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf4) );
  BUFX2 BUFX2_1148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545), .Y(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf3) );
  BUFX2 BUFX2_1149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545), .Y(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf2) );
  BUFX2 BUFX2_115 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94) );
  BUFX2 BUFX2_1150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545), .Y(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf1) );
  BUFX2 BUFX2_1151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5545), .Y(REGFILE_SIM_reg_bank__abc_33898_n5545_bF_buf0) );
  BUFX2 BUFX2_1152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548), .Y(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf4) );
  BUFX2 BUFX2_1153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548), .Y(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf3) );
  BUFX2 BUFX2_1154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548), .Y(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf2) );
  BUFX2 BUFX2_1155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548), .Y(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf1) );
  BUFX2 BUFX2_1156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5548), .Y(REGFILE_SIM_reg_bank__abc_33898_n5548_bF_buf0) );
  BUFX2 BUFX2_1157 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3) );
  BUFX2 BUFX2_1158 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2) );
  BUFX2 BUFX2_1159 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1) );
  BUFX2 BUFX2_116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93) );
  BUFX2 BUFX2_1160 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0) );
  BUFX2 BUFX2_1161 ( .A(_abc_43815_n3317), .Y(_abc_43815_n3317_bF_buf3) );
  BUFX2 BUFX2_1162 ( .A(_abc_43815_n3317), .Y(_abc_43815_n3317_bF_buf2) );
  BUFX2 BUFX2_1163 ( .A(_abc_43815_n3317), .Y(_abc_43815_n3317_bF_buf1) );
  BUFX2 BUFX2_1164 ( .A(_abc_43815_n3317), .Y(_abc_43815_n3317_bF_buf0) );
  BUFX2 BUFX2_1165 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3) );
  BUFX2 BUFX2_1166 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2) );
  BUFX2 BUFX2_1167 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1) );
  BUFX2 BUFX2_1168 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0) );
  BUFX2 BUFX2_1169 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf5) );
  BUFX2 BUFX2_117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92) );
  BUFX2 BUFX2_1170 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf4) );
  BUFX2 BUFX2_1171 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf3) );
  BUFX2 BUFX2_1172 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf2) );
  BUFX2 BUFX2_1173 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf1) );
  BUFX2 BUFX2_1174 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf0) );
  BUFX2 BUFX2_1175 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3) );
  BUFX2 BUFX2_1176 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2) );
  BUFX2 BUFX2_1177 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1) );
  BUFX2 BUFX2_1178 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0) );
  BUFX2 BUFX2_1179 ( .A(alu_op_i_0_), .Y(alu_op_i_0_bF_buf5) );
  BUFX2 BUFX2_118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91) );
  BUFX2 BUFX2_1180 ( .A(alu_op_i_0_), .Y(alu_op_i_0_bF_buf4) );
  BUFX2 BUFX2_1181 ( .A(alu_op_i_0_), .Y(alu_op_i_0_bF_buf3) );
  BUFX2 BUFX2_1182 ( .A(alu_op_i_0_), .Y(alu_op_i_0_bF_buf2) );
  BUFX2 BUFX2_1183 ( .A(alu_op_i_0_), .Y(alu_op_i_0_bF_buf1) );
  BUFX2 BUFX2_1184 ( .A(alu_op_i_0_), .Y(alu_op_i_0_bF_buf0) );
  BUFX2 BUFX2_1185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958), .Y(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4) );
  BUFX2 BUFX2_1186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958), .Y(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3) );
  BUFX2 BUFX2_1187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958), .Y(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2) );
  BUFX2 BUFX2_1188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958), .Y(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf1) );
  BUFX2 BUFX2_1189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958), .Y(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf0) );
  BUFX2 BUFX2_119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90) );
  BUFX2 BUFX2_1190 ( .A(_abc_43815_n3521_1), .Y(_abc_43815_n3521_1_bF_buf3) );
  BUFX2 BUFX2_1191 ( .A(_abc_43815_n3521_1), .Y(_abc_43815_n3521_1_bF_buf2) );
  BUFX2 BUFX2_1192 ( .A(_abc_43815_n3521_1), .Y(_abc_43815_n3521_1_bF_buf1) );
  BUFX2 BUFX2_1193 ( .A(_abc_43815_n3521_1), .Y(_abc_43815_n3521_1_bF_buf0) );
  BUFX2 BUFX2_1194 ( .A(alu__abc_41358_n279), .Y(alu__abc_41358_n279_bF_buf5) );
  BUFX2 BUFX2_1195 ( .A(alu__abc_41358_n279), .Y(alu__abc_41358_n279_bF_buf4) );
  BUFX2 BUFX2_1196 ( .A(alu__abc_41358_n279), .Y(alu__abc_41358_n279_bF_buf3) );
  BUFX2 BUFX2_1197 ( .A(alu__abc_41358_n279), .Y(alu__abc_41358_n279_bF_buf2) );
  BUFX2 BUFX2_1198 ( .A(alu__abc_41358_n279), .Y(alu__abc_41358_n279_bF_buf1) );
  BUFX2 BUFX2_1199 ( .A(alu__abc_41358_n279), .Y(alu__abc_41358_n279_bF_buf0) );
  BUFX2 BUFX2_12 ( .A(_abc_43815_n4167_bF_buf15), .Y(_abc_43815_n4167_bF_buf15_bF_buf1) );
  BUFX2 BUFX2_120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89) );
  BUFX2 BUFX2_1200 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3) );
  BUFX2 BUFX2_1201 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2) );
  BUFX2 BUFX2_1202 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1) );
  BUFX2 BUFX2_1203 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0) );
  BUFX2 BUFX2_1204 ( .A(_abc_43815_n832_1), .Y(_abc_43815_n832_1_bF_buf3) );
  BUFX2 BUFX2_1205 ( .A(_abc_43815_n832_1), .Y(_abc_43815_n832_1_bF_buf2) );
  BUFX2 BUFX2_1206 ( .A(_abc_43815_n832_1), .Y(_abc_43815_n832_1_bF_buf1) );
  BUFX2 BUFX2_1207 ( .A(_abc_43815_n832_1), .Y(_abc_43815_n832_1_bF_buf0) );
  BUFX2 BUFX2_1208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519), .Y(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4) );
  BUFX2 BUFX2_1209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519), .Y(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3) );
  BUFX2 BUFX2_121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88) );
  BUFX2 BUFX2_1210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519), .Y(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf2) );
  BUFX2 BUFX2_1211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519), .Y(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf1) );
  BUFX2 BUFX2_1212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519), .Y(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf0) );
  BUFX2 BUFX2_1213 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3) );
  BUFX2 BUFX2_1214 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2) );
  BUFX2 BUFX2_1215 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1) );
  BUFX2 BUFX2_1216 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0) );
  BUFX2 BUFX2_1217 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf15) );
  BUFX2 BUFX2_1218 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf14) );
  BUFX2 BUFX2_1219 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf13) );
  BUFX2 BUFX2_122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87) );
  BUFX2 BUFX2_1220 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf12) );
  BUFX2 BUFX2_1221 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf11) );
  BUFX2 BUFX2_1222 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf10) );
  BUFX2 BUFX2_1223 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf9) );
  BUFX2 BUFX2_1224 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf8) );
  BUFX2 BUFX2_1225 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf7) );
  BUFX2 BUFX2_1226 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf6) );
  BUFX2 BUFX2_1227 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf5) );
  BUFX2 BUFX2_1228 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf4) );
  BUFX2 BUFX2_1229 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf3) );
  BUFX2 BUFX2_123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86) );
  BUFX2 BUFX2_1230 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf2) );
  BUFX2 BUFX2_1231 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf1) );
  BUFX2 BUFX2_1232 ( .A(_abc_43815_n4167), .Y(_abc_43815_n4167_bF_buf0) );
  BUFX2 BUFX2_1233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7) );
  BUFX2 BUFX2_1234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf6) );
  BUFX2 BUFX2_1235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5) );
  BUFX2 BUFX2_1236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf4) );
  BUFX2 BUFX2_1237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3) );
  BUFX2 BUFX2_1238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf2) );
  BUFX2 BUFX2_1239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1) );
  BUFX2 BUFX2_124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85) );
  BUFX2 BUFX2_1240 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018), .Y(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf0) );
  BUFX2 BUFX2_1241 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042), .Y(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4) );
  BUFX2 BUFX2_1242 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042), .Y(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3) );
  BUFX2 BUFX2_1243 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042), .Y(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2) );
  BUFX2 BUFX2_1244 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042), .Y(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf1) );
  BUFX2 BUFX2_1245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042), .Y(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf0) );
  BUFX2 BUFX2_1246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044), .Y(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4) );
  BUFX2 BUFX2_1247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044), .Y(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3) );
  BUFX2 BUFX2_1248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044), .Y(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf2) );
  BUFX2 BUFX2_1249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044), .Y(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf1) );
  BUFX2 BUFX2_125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84) );
  BUFX2 BUFX2_1250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044), .Y(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf0) );
  BUFX2 BUFX2_1251 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3) );
  BUFX2 BUFX2_1252 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2) );
  BUFX2 BUFX2_1253 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1) );
  BUFX2 BUFX2_1254 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0) );
  BUFX2 BUFX2_1255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652), .Y(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf4) );
  BUFX2 BUFX2_1256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652), .Y(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf3) );
  BUFX2 BUFX2_1257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652), .Y(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf2) );
  BUFX2 BUFX2_1258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652), .Y(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf1) );
  BUFX2 BUFX2_1259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7652), .Y(REGFILE_SIM_reg_bank__abc_33898_n7652_bF_buf0) );
  BUFX2 BUFX2_126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83) );
  BUFX2 BUFX2_1260 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654), .Y(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf4) );
  BUFX2 BUFX2_1261 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654), .Y(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf3) );
  BUFX2 BUFX2_1262 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654), .Y(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf2) );
  BUFX2 BUFX2_1263 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654), .Y(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf1) );
  BUFX2 BUFX2_1264 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7654), .Y(REGFILE_SIM_reg_bank__abc_33898_n7654_bF_buf0) );
  BUFX2 BUFX2_1265 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657), .Y(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf4) );
  BUFX2 BUFX2_1266 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657), .Y(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf3) );
  BUFX2 BUFX2_1267 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657), .Y(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf2) );
  BUFX2 BUFX2_1268 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657), .Y(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf1) );
  BUFX2 BUFX2_1269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7657), .Y(REGFILE_SIM_reg_bank__abc_33898_n7657_bF_buf0) );
  BUFX2 BUFX2_127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82) );
  BUFX2 BUFX2_1270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659), .Y(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf4) );
  BUFX2 BUFX2_1271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659), .Y(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf3) );
  BUFX2 BUFX2_1272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659), .Y(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf2) );
  BUFX2 BUFX2_1273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659), .Y(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf1) );
  BUFX2 BUFX2_1274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7659), .Y(REGFILE_SIM_reg_bank__abc_33898_n7659_bF_buf0) );
  BUFX2 BUFX2_1275 ( .A(_abc_43815_n680_1), .Y(_abc_43815_n680_1_bF_buf4) );
  BUFX2 BUFX2_1276 ( .A(_abc_43815_n680_1), .Y(_abc_43815_n680_1_bF_buf3) );
  BUFX2 BUFX2_1277 ( .A(_abc_43815_n680_1), .Y(_abc_43815_n680_1_bF_buf2) );
  BUFX2 BUFX2_1278 ( .A(_abc_43815_n680_1), .Y(_abc_43815_n680_1_bF_buf1) );
  BUFX2 BUFX2_1279 ( .A(_abc_43815_n680_1), .Y(_abc_43815_n680_1_bF_buf0) );
  BUFX2 BUFX2_128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81) );
  BUFX2 BUFX2_1280 ( .A(_abc_43815_n3549), .Y(_abc_43815_n3549_bF_buf4) );
  BUFX2 BUFX2_1281 ( .A(_abc_43815_n3549), .Y(_abc_43815_n3549_bF_buf3) );
  BUFX2 BUFX2_1282 ( .A(_abc_43815_n3549), .Y(_abc_43815_n3549_bF_buf2) );
  BUFX2 BUFX2_1283 ( .A(_abc_43815_n3549), .Y(_abc_43815_n3549_bF_buf1) );
  BUFX2 BUFX2_1284 ( .A(_abc_43815_n3549), .Y(_abc_43815_n3549_bF_buf0) );
  BUFX2 BUFX2_1285 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf6) );
  BUFX2 BUFX2_1286 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf5) );
  BUFX2 BUFX2_1287 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf4) );
  BUFX2 BUFX2_1288 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf3) );
  BUFX2 BUFX2_1289 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf2) );
  BUFX2 BUFX2_129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80) );
  BUFX2 BUFX2_1290 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf1) );
  BUFX2 BUFX2_1291 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf0) );
  BUFX2 BUFX2_1292 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3) );
  BUFX2 BUFX2_1293 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2) );
  BUFX2 BUFX2_1294 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1) );
  BUFX2 BUFX2_1295 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0) );
  BUFX2 BUFX2_1296 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622), .Y(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf4) );
  BUFX2 BUFX2_1297 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622), .Y(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf3) );
  BUFX2 BUFX2_1298 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622), .Y(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf2) );
  BUFX2 BUFX2_1299 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622), .Y(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf1) );
  BUFX2 BUFX2_13 ( .A(_abc_43815_n4167_bF_buf15), .Y(_abc_43815_n4167_bF_buf15_bF_buf0) );
  BUFX2 BUFX2_130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79) );
  BUFX2 BUFX2_1300 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7622), .Y(REGFILE_SIM_reg_bank__abc_33898_n7622_bF_buf0) );
  BUFX2 BUFX2_1301 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625), .Y(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf4) );
  BUFX2 BUFX2_1302 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625), .Y(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf3) );
  BUFX2 BUFX2_1303 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625), .Y(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf2) );
  BUFX2 BUFX2_1304 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625), .Y(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf1) );
  BUFX2 BUFX2_1305 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7625), .Y(REGFILE_SIM_reg_bank__abc_33898_n7625_bF_buf0) );
  BUFX2 BUFX2_1306 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627), .Y(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf4) );
  BUFX2 BUFX2_1307 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627), .Y(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf3) );
  BUFX2 BUFX2_1308 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627), .Y(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf2) );
  BUFX2 BUFX2_1309 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627), .Y(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf1) );
  BUFX2 BUFX2_131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78) );
  BUFX2 BUFX2_1310 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7627), .Y(REGFILE_SIM_reg_bank__abc_33898_n7627_bF_buf0) );
  BUFX2 BUFX2_1311 ( .A(alu__abc_41358_n942), .Y(alu__abc_41358_n942_bF_buf4) );
  BUFX2 BUFX2_1312 ( .A(alu__abc_41358_n942), .Y(alu__abc_41358_n942_bF_buf3) );
  BUFX2 BUFX2_1313 ( .A(alu__abc_41358_n942), .Y(alu__abc_41358_n942_bF_buf2) );
  BUFX2 BUFX2_1314 ( .A(alu__abc_41358_n942), .Y(alu__abc_41358_n942_bF_buf1) );
  BUFX2 BUFX2_1315 ( .A(alu__abc_41358_n942), .Y(alu__abc_41358_n942_bF_buf0) );
  BUFX2 BUFX2_1316 ( .A(alu__abc_41358_n948), .Y(alu__abc_41358_n948_bF_buf4) );
  BUFX2 BUFX2_1317 ( .A(alu__abc_41358_n948), .Y(alu__abc_41358_n948_bF_buf3) );
  BUFX2 BUFX2_1318 ( .A(alu__abc_41358_n948), .Y(alu__abc_41358_n948_bF_buf2) );
  BUFX2 BUFX2_1319 ( .A(alu__abc_41358_n948), .Y(alu__abc_41358_n948_bF_buf1) );
  BUFX2 BUFX2_132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77) );
  BUFX2 BUFX2_1320 ( .A(alu__abc_41358_n948), .Y(alu__abc_41358_n948_bF_buf0) );
  BUFX2 BUFX2_1321 ( .A(_auto_iopadmap_cc_313_execute_47726), .Y(break_o) );
  BUFX2 BUFX2_1322 ( .A(_auto_iopadmap_cc_313_execute_47728), .Y(fault_o) );
  BUFX2 BUFX2_1323 ( .A(_auto_iopadmap_cc_313_execute_47730_0_), .Y(\mem_addr_o[0] ) );
  BUFX2 BUFX2_1324 ( .A(_auto_iopadmap_cc_313_execute_47730_1_), .Y(\mem_addr_o[1] ) );
  BUFX2 BUFX2_1325 ( .A(_auto_iopadmap_cc_313_execute_47730_2_), .Y(\mem_addr_o[2] ) );
  BUFX2 BUFX2_1326 ( .A(_auto_iopadmap_cc_313_execute_47730_3_), .Y(\mem_addr_o[3] ) );
  BUFX2 BUFX2_1327 ( .A(_auto_iopadmap_cc_313_execute_47730_4_), .Y(\mem_addr_o[4] ) );
  BUFX2 BUFX2_1328 ( .A(_auto_iopadmap_cc_313_execute_47730_5_), .Y(\mem_addr_o[5] ) );
  BUFX2 BUFX2_1329 ( .A(_auto_iopadmap_cc_313_execute_47730_6_), .Y(\mem_addr_o[6] ) );
  BUFX2 BUFX2_133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76) );
  BUFX2 BUFX2_1330 ( .A(_auto_iopadmap_cc_313_execute_47730_7_), .Y(\mem_addr_o[7] ) );
  BUFX2 BUFX2_1331 ( .A(_auto_iopadmap_cc_313_execute_47730_8_), .Y(\mem_addr_o[8] ) );
  BUFX2 BUFX2_1332 ( .A(_auto_iopadmap_cc_313_execute_47730_9_), .Y(\mem_addr_o[9] ) );
  BUFX2 BUFX2_1333 ( .A(_auto_iopadmap_cc_313_execute_47730_10_), .Y(\mem_addr_o[10] ) );
  BUFX2 BUFX2_1334 ( .A(_auto_iopadmap_cc_313_execute_47730_11_), .Y(\mem_addr_o[11] ) );
  BUFX2 BUFX2_1335 ( .A(_auto_iopadmap_cc_313_execute_47730_12_), .Y(\mem_addr_o[12] ) );
  BUFX2 BUFX2_1336 ( .A(_auto_iopadmap_cc_313_execute_47730_13_), .Y(\mem_addr_o[13] ) );
  BUFX2 BUFX2_1337 ( .A(_auto_iopadmap_cc_313_execute_47730_14_), .Y(\mem_addr_o[14] ) );
  BUFX2 BUFX2_1338 ( .A(_auto_iopadmap_cc_313_execute_47730_15_), .Y(\mem_addr_o[15] ) );
  BUFX2 BUFX2_1339 ( .A(_auto_iopadmap_cc_313_execute_47730_16_), .Y(\mem_addr_o[16] ) );
  BUFX2 BUFX2_134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75) );
  BUFX2 BUFX2_1340 ( .A(_auto_iopadmap_cc_313_execute_47730_17_), .Y(\mem_addr_o[17] ) );
  BUFX2 BUFX2_1341 ( .A(_auto_iopadmap_cc_313_execute_47730_18_), .Y(\mem_addr_o[18] ) );
  BUFX2 BUFX2_1342 ( .A(_auto_iopadmap_cc_313_execute_47730_19_), .Y(\mem_addr_o[19] ) );
  BUFX2 BUFX2_1343 ( .A(_auto_iopadmap_cc_313_execute_47730_20_), .Y(\mem_addr_o[20] ) );
  BUFX2 BUFX2_1344 ( .A(_auto_iopadmap_cc_313_execute_47730_21_), .Y(\mem_addr_o[21] ) );
  BUFX2 BUFX2_1345 ( .A(_auto_iopadmap_cc_313_execute_47730_22_), .Y(\mem_addr_o[22] ) );
  BUFX2 BUFX2_1346 ( .A(_auto_iopadmap_cc_313_execute_47730_23_), .Y(\mem_addr_o[23] ) );
  BUFX2 BUFX2_1347 ( .A(_auto_iopadmap_cc_313_execute_47730_24_), .Y(\mem_addr_o[24] ) );
  BUFX2 BUFX2_1348 ( .A(_auto_iopadmap_cc_313_execute_47730_25_), .Y(\mem_addr_o[25] ) );
  BUFX2 BUFX2_1349 ( .A(_auto_iopadmap_cc_313_execute_47730_26_), .Y(\mem_addr_o[26] ) );
  BUFX2 BUFX2_135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74) );
  BUFX2 BUFX2_1350 ( .A(_auto_iopadmap_cc_313_execute_47730_27_), .Y(\mem_addr_o[27] ) );
  BUFX2 BUFX2_1351 ( .A(_auto_iopadmap_cc_313_execute_47730_28_), .Y(\mem_addr_o[28] ) );
  BUFX2 BUFX2_1352 ( .A(_auto_iopadmap_cc_313_execute_47730_29_), .Y(\mem_addr_o[29] ) );
  BUFX2 BUFX2_1353 ( .A(_auto_iopadmap_cc_313_execute_47730_30_), .Y(\mem_addr_o[30] ) );
  BUFX2 BUFX2_1354 ( .A(_auto_iopadmap_cc_313_execute_47730_31_), .Y(\mem_addr_o[31] ) );
  BUFX2 BUFX2_1355 ( .A(1'b1), .Y(\mem_cti_o[0] ) );
  BUFX2 BUFX2_1356 ( .A(1'b1), .Y(\mem_cti_o[1] ) );
  BUFX2 BUFX2_1357 ( .A(1'b1), .Y(\mem_cti_o[2] ) );
  BUFX2 BUFX2_1358 ( .A(_auto_iopadmap_cc_313_execute_47767), .Y(mem_cyc_o) );
  BUFX2 BUFX2_1359 ( .A(_auto_iopadmap_cc_313_execute_47769_0_), .Y(\mem_dat_o[0] ) );
  BUFX2 BUFX2_136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73) );
  BUFX2 BUFX2_1360 ( .A(_auto_iopadmap_cc_313_execute_47769_1_), .Y(\mem_dat_o[1] ) );
  BUFX2 BUFX2_1361 ( .A(_auto_iopadmap_cc_313_execute_47769_2_), .Y(\mem_dat_o[2] ) );
  BUFX2 BUFX2_1362 ( .A(_auto_iopadmap_cc_313_execute_47769_3_), .Y(\mem_dat_o[3] ) );
  BUFX2 BUFX2_1363 ( .A(_auto_iopadmap_cc_313_execute_47769_4_), .Y(\mem_dat_o[4] ) );
  BUFX2 BUFX2_1364 ( .A(_auto_iopadmap_cc_313_execute_47769_5_), .Y(\mem_dat_o[5] ) );
  BUFX2 BUFX2_1365 ( .A(_auto_iopadmap_cc_313_execute_47769_6_), .Y(\mem_dat_o[6] ) );
  BUFX2 BUFX2_1366 ( .A(_auto_iopadmap_cc_313_execute_47769_7_), .Y(\mem_dat_o[7] ) );
  BUFX2 BUFX2_1367 ( .A(_auto_iopadmap_cc_313_execute_47769_8_), .Y(\mem_dat_o[8] ) );
  BUFX2 BUFX2_1368 ( .A(_auto_iopadmap_cc_313_execute_47769_9_), .Y(\mem_dat_o[9] ) );
  BUFX2 BUFX2_1369 ( .A(_auto_iopadmap_cc_313_execute_47769_10_), .Y(\mem_dat_o[10] ) );
  BUFX2 BUFX2_137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72) );
  BUFX2 BUFX2_1370 ( .A(_auto_iopadmap_cc_313_execute_47769_11_), .Y(\mem_dat_o[11] ) );
  BUFX2 BUFX2_1371 ( .A(_auto_iopadmap_cc_313_execute_47769_12_), .Y(\mem_dat_o[12] ) );
  BUFX2 BUFX2_1372 ( .A(_auto_iopadmap_cc_313_execute_47769_13_), .Y(\mem_dat_o[13] ) );
  BUFX2 BUFX2_1373 ( .A(_auto_iopadmap_cc_313_execute_47769_14_), .Y(\mem_dat_o[14] ) );
  BUFX2 BUFX2_1374 ( .A(_auto_iopadmap_cc_313_execute_47769_15_), .Y(\mem_dat_o[15] ) );
  BUFX2 BUFX2_1375 ( .A(_auto_iopadmap_cc_313_execute_47769_16_), .Y(\mem_dat_o[16] ) );
  BUFX2 BUFX2_1376 ( .A(_auto_iopadmap_cc_313_execute_47769_17_), .Y(\mem_dat_o[17] ) );
  BUFX2 BUFX2_1377 ( .A(_auto_iopadmap_cc_313_execute_47769_18_), .Y(\mem_dat_o[18] ) );
  BUFX2 BUFX2_1378 ( .A(_auto_iopadmap_cc_313_execute_47769_19_), .Y(\mem_dat_o[19] ) );
  BUFX2 BUFX2_1379 ( .A(_auto_iopadmap_cc_313_execute_47769_20_), .Y(\mem_dat_o[20] ) );
  BUFX2 BUFX2_138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71) );
  BUFX2 BUFX2_1380 ( .A(_auto_iopadmap_cc_313_execute_47769_21_), .Y(\mem_dat_o[21] ) );
  BUFX2 BUFX2_1381 ( .A(_auto_iopadmap_cc_313_execute_47769_22_), .Y(\mem_dat_o[22] ) );
  BUFX2 BUFX2_1382 ( .A(_auto_iopadmap_cc_313_execute_47769_23_), .Y(\mem_dat_o[23] ) );
  BUFX2 BUFX2_1383 ( .A(_auto_iopadmap_cc_313_execute_47769_24_), .Y(\mem_dat_o[24] ) );
  BUFX2 BUFX2_1384 ( .A(_auto_iopadmap_cc_313_execute_47769_25_), .Y(\mem_dat_o[25] ) );
  BUFX2 BUFX2_1385 ( .A(_auto_iopadmap_cc_313_execute_47769_26_), .Y(\mem_dat_o[26] ) );
  BUFX2 BUFX2_1386 ( .A(_auto_iopadmap_cc_313_execute_47769_27_), .Y(\mem_dat_o[27] ) );
  BUFX2 BUFX2_1387 ( .A(_auto_iopadmap_cc_313_execute_47769_28_), .Y(\mem_dat_o[28] ) );
  BUFX2 BUFX2_1388 ( .A(_auto_iopadmap_cc_313_execute_47769_29_), .Y(\mem_dat_o[29] ) );
  BUFX2 BUFX2_1389 ( .A(_auto_iopadmap_cc_313_execute_47769_30_), .Y(\mem_dat_o[30] ) );
  BUFX2 BUFX2_139 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70) );
  BUFX2 BUFX2_1390 ( .A(_auto_iopadmap_cc_313_execute_47769_31_), .Y(\mem_dat_o[31] ) );
  BUFX2 BUFX2_1391 ( .A(_auto_iopadmap_cc_313_execute_47802_0_), .Y(\mem_sel_o[0] ) );
  BUFX2 BUFX2_1392 ( .A(_auto_iopadmap_cc_313_execute_47802_1_), .Y(\mem_sel_o[1] ) );
  BUFX2 BUFX2_1393 ( .A(_auto_iopadmap_cc_313_execute_47802_2_), .Y(\mem_sel_o[2] ) );
  BUFX2 BUFX2_1394 ( .A(_auto_iopadmap_cc_313_execute_47802_3_), .Y(\mem_sel_o[3] ) );
  BUFX2 BUFX2_1395 ( .A(_auto_iopadmap_cc_313_execute_47807), .Y(mem_stb_o) );
  BUFX2 BUFX2_1396 ( .A(_auto_iopadmap_cc_313_execute_47809), .Y(mem_we_o) );
  BUFX2 BUFX2_14 ( .A(clk_i), .Y(clk_i_hier0_bF_buf9) );
  BUFX2 BUFX2_140 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69) );
  BUFX2 BUFX2_141 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68) );
  BUFX2 BUFX2_142 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67) );
  BUFX2 BUFX2_143 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66) );
  BUFX2 BUFX2_144 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65) );
  BUFX2 BUFX2_145 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64) );
  BUFX2 BUFX2_146 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63) );
  BUFX2 BUFX2_147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62) );
  BUFX2 BUFX2_148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61) );
  BUFX2 BUFX2_149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60) );
  BUFX2 BUFX2_15 ( .A(clk_i), .Y(clk_i_hier0_bF_buf8) );
  BUFX2 BUFX2_150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59) );
  BUFX2 BUFX2_151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58) );
  BUFX2 BUFX2_152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57) );
  BUFX2 BUFX2_153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56) );
  BUFX2 BUFX2_154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55) );
  BUFX2 BUFX2_155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54) );
  BUFX2 BUFX2_156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53) );
  BUFX2 BUFX2_157 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52) );
  BUFX2 BUFX2_158 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51) );
  BUFX2 BUFX2_159 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50) );
  BUFX2 BUFX2_16 ( .A(clk_i), .Y(clk_i_hier0_bF_buf7) );
  BUFX2 BUFX2_160 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49) );
  BUFX2 BUFX2_161 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48) );
  BUFX2 BUFX2_162 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47) );
  BUFX2 BUFX2_163 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46) );
  BUFX2 BUFX2_164 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45) );
  BUFX2 BUFX2_165 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44) );
  BUFX2 BUFX2_166 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43) );
  BUFX2 BUFX2_167 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42) );
  BUFX2 BUFX2_168 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41) );
  BUFX2 BUFX2_169 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40) );
  BUFX2 BUFX2_17 ( .A(clk_i), .Y(clk_i_hier0_bF_buf6) );
  BUFX2 BUFX2_170 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39) );
  BUFX2 BUFX2_171 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38) );
  BUFX2 BUFX2_172 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37) );
  BUFX2 BUFX2_173 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36) );
  BUFX2 BUFX2_174 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35) );
  BUFX2 BUFX2_175 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34) );
  BUFX2 BUFX2_176 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33) );
  BUFX2 BUFX2_177 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32) );
  BUFX2 BUFX2_178 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31) );
  BUFX2 BUFX2_179 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30) );
  BUFX2 BUFX2_18 ( .A(clk_i), .Y(clk_i_hier0_bF_buf5) );
  BUFX2 BUFX2_180 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29) );
  BUFX2 BUFX2_181 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28) );
  BUFX2 BUFX2_182 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27) );
  BUFX2 BUFX2_183 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26) );
  BUFX2 BUFX2_184 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25) );
  BUFX2 BUFX2_185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24) );
  BUFX2 BUFX2_186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23) );
  BUFX2 BUFX2_187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22) );
  BUFX2 BUFX2_188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21) );
  BUFX2 BUFX2_189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20) );
  BUFX2 BUFX2_19 ( .A(clk_i), .Y(clk_i_hier0_bF_buf4) );
  BUFX2 BUFX2_190 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19) );
  BUFX2 BUFX2_191 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18) );
  BUFX2 BUFX2_192 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17) );
  BUFX2 BUFX2_193 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16) );
  BUFX2 BUFX2_194 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15) );
  BUFX2 BUFX2_195 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14) );
  BUFX2 BUFX2_196 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13) );
  BUFX2 BUFX2_197 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12) );
  BUFX2 BUFX2_198 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11) );
  BUFX2 BUFX2_199 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10) );
  BUFX2 BUFX2_2 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7) );
  BUFX2 BUFX2_20 ( .A(clk_i), .Y(clk_i_hier0_bF_buf3) );
  BUFX2 BUFX2_200 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9) );
  BUFX2 BUFX2_201 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8) );
  BUFX2 BUFX2_202 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7) );
  BUFX2 BUFX2_203 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6) );
  BUFX2 BUFX2_204 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5) );
  BUFX2 BUFX2_205 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4) );
  BUFX2 BUFX2_206 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3) );
  BUFX2 BUFX2_207 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2) );
  BUFX2 BUFX2_208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1) );
  BUFX2 BUFX2_209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0) );
  BUFX2 BUFX2_21 ( .A(clk_i), .Y(clk_i_hier0_bF_buf2) );
  BUFX2 BUFX2_210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247), .Y(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4) );
  BUFX2 BUFX2_211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247), .Y(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3) );
  BUFX2 BUFX2_212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247), .Y(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf2) );
  BUFX2 BUFX2_213 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247), .Y(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf1) );
  BUFX2 BUFX2_214 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247), .Y(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf0) );
  BUFX2 BUFX2_215 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623), .Y(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf4) );
  BUFX2 BUFX2_216 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623), .Y(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf3) );
  BUFX2 BUFX2_217 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623), .Y(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf2) );
  BUFX2 BUFX2_218 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623), .Y(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf1) );
  BUFX2 BUFX2_219 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5623), .Y(REGFILE_SIM_reg_bank__abc_33898_n5623_bF_buf0) );
  BUFX2 BUFX2_22 ( .A(clk_i), .Y(clk_i_hier0_bF_buf1) );
  BUFX2 BUFX2_220 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625), .Y(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf4) );
  BUFX2 BUFX2_221 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625), .Y(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf3) );
  BUFX2 BUFX2_222 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625), .Y(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf2) );
  BUFX2 BUFX2_223 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625), .Y(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf1) );
  BUFX2 BUFX2_224 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5625), .Y(REGFILE_SIM_reg_bank__abc_33898_n5625_bF_buf0) );
  BUFX2 BUFX2_225 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627), .Y(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf4) );
  BUFX2 BUFX2_226 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627), .Y(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf3) );
  BUFX2 BUFX2_227 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627), .Y(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf2) );
  BUFX2 BUFX2_228 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627), .Y(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf1) );
  BUFX2 BUFX2_229 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5627), .Y(REGFILE_SIM_reg_bank__abc_33898_n5627_bF_buf0) );
  BUFX2 BUFX2_23 ( .A(clk_i), .Y(clk_i_hier0_bF_buf0) );
  BUFX2 BUFX2_230 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715), .Y(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4) );
  BUFX2 BUFX2_231 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715), .Y(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3) );
  BUFX2 BUFX2_232 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715), .Y(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2) );
  BUFX2 BUFX2_233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715), .Y(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf1) );
  BUFX2 BUFX2_234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715), .Y(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf0) );
  BUFX2 BUFX2_235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717), .Y(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4) );
  BUFX2 BUFX2_236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717), .Y(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3) );
  BUFX2 BUFX2_237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717), .Y(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf2) );
  BUFX2 BUFX2_238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717), .Y(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf1) );
  BUFX2 BUFX2_239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717), .Y(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf0) );
  BUFX2 BUFX2_24 ( .A(_abc_43815_n671), .Y(_abc_43815_n671_bF_buf4) );
  BUFX2 BUFX2_240 ( .A(_abc_43815_n1172_1), .Y(_abc_43815_n1172_1_bF_buf4) );
  BUFX2 BUFX2_241 ( .A(_abc_43815_n1172_1), .Y(_abc_43815_n1172_1_bF_buf3) );
  BUFX2 BUFX2_242 ( .A(_abc_43815_n1172_1), .Y(_abc_43815_n1172_1_bF_buf2) );
  BUFX2 BUFX2_243 ( .A(_abc_43815_n1172_1), .Y(_abc_43815_n1172_1_bF_buf1) );
  BUFX2 BUFX2_244 ( .A(_abc_43815_n1172_1), .Y(_abc_43815_n1172_1_bF_buf0) );
  BUFX2 BUFX2_245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590), .Y(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf4) );
  BUFX2 BUFX2_246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590), .Y(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf3) );
  BUFX2 BUFX2_247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590), .Y(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf2) );
  BUFX2 BUFX2_248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590), .Y(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf1) );
  BUFX2 BUFX2_249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5590), .Y(REGFILE_SIM_reg_bank__abc_33898_n5590_bF_buf0) );
  BUFX2 BUFX2_25 ( .A(_abc_43815_n671), .Y(_abc_43815_n671_bF_buf3) );
  BUFX2 BUFX2_250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594), .Y(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf4) );
  BUFX2 BUFX2_251 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594), .Y(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf3) );
  BUFX2 BUFX2_252 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594), .Y(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf2) );
  BUFX2 BUFX2_253 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594), .Y(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf1) );
  BUFX2 BUFX2_254 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5594), .Y(REGFILE_SIM_reg_bank__abc_33898_n5594_bF_buf0) );
  BUFX2 BUFX2_255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597), .Y(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf4) );
  BUFX2 BUFX2_256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597), .Y(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf3) );
  BUFX2 BUFX2_257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597), .Y(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf2) );
  BUFX2 BUFX2_258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597), .Y(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf1) );
  BUFX2 BUFX2_259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5597), .Y(REGFILE_SIM_reg_bank__abc_33898_n5597_bF_buf0) );
  BUFX2 BUFX2_26 ( .A(_abc_43815_n671), .Y(_abc_43815_n671_bF_buf2) );
  BUFX2 BUFX2_260 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3) );
  BUFX2 BUFX2_261 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2) );
  BUFX2 BUFX2_262 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1) );
  BUFX2 BUFX2_263 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0) );
  BUFX2 BUFX2_264 ( .A(_abc_43815_n1489), .Y(_abc_43815_n1489_bF_buf4) );
  BUFX2 BUFX2_265 ( .A(_abc_43815_n1489), .Y(_abc_43815_n1489_bF_buf3) );
  BUFX2 BUFX2_266 ( .A(_abc_43815_n1489), .Y(_abc_43815_n1489_bF_buf2) );
  BUFX2 BUFX2_267 ( .A(_abc_43815_n1489), .Y(_abc_43815_n1489_bF_buf1) );
  BUFX2 BUFX2_268 ( .A(_abc_43815_n1489), .Y(_abc_43815_n1489_bF_buf0) );
  BUFX2 BUFX2_269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241), .Y(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4) );
  BUFX2 BUFX2_27 ( .A(_abc_43815_n671), .Y(_abc_43815_n671_bF_buf1) );
  BUFX2 BUFX2_270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241), .Y(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3) );
  BUFX2 BUFX2_271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241), .Y(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf2) );
  BUFX2 BUFX2_272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241), .Y(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf1) );
  BUFX2 BUFX2_273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241), .Y(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf0) );
  BUFX2 BUFX2_274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565), .Y(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf4) );
  BUFX2 BUFX2_275 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565), .Y(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf3) );
  BUFX2 BUFX2_276 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565), .Y(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf2) );
  BUFX2 BUFX2_277 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565), .Y(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf1) );
  BUFX2 BUFX2_278 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5565), .Y(REGFILE_SIM_reg_bank__abc_33898_n5565_bF_buf0) );
  BUFX2 BUFX2_279 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568), .Y(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf4) );
  BUFX2 BUFX2_28 ( .A(_abc_43815_n671), .Y(_abc_43815_n671_bF_buf0) );
  BUFX2 BUFX2_280 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568), .Y(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf3) );
  BUFX2 BUFX2_281 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568), .Y(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf2) );
  BUFX2 BUFX2_282 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568), .Y(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf1) );
  BUFX2 BUFX2_283 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5568), .Y(REGFILE_SIM_reg_bank__abc_33898_n5568_bF_buf0) );
  BUFX2 BUFX2_284 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3) );
  BUFX2 BUFX2_285 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2) );
  BUFX2 BUFX2_286 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1) );
  BUFX2 BUFX2_287 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0) );
  BUFX2 BUFX2_288 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf114) );
  BUFX2 BUFX2_289 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf113) );
  BUFX2 BUFX2_29 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590), .Y(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf4) );
  BUFX2 BUFX2_290 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf112) );
  BUFX2 BUFX2_291 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf111) );
  BUFX2 BUFX2_292 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf110) );
  BUFX2 BUFX2_293 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf109) );
  BUFX2 BUFX2_294 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf108) );
  BUFX2 BUFX2_295 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf107) );
  BUFX2 BUFX2_296 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf106) );
  BUFX2 BUFX2_297 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf105) );
  BUFX2 BUFX2_298 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf104) );
  BUFX2 BUFX2_299 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf103) );
  BUFX2 BUFX2_3 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf6) );
  BUFX2 BUFX2_30 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590), .Y(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf3) );
  BUFX2 BUFX2_300 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf102) );
  BUFX2 BUFX2_301 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf101) );
  BUFX2 BUFX2_302 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf100) );
  BUFX2 BUFX2_303 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf99) );
  BUFX2 BUFX2_304 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf98) );
  BUFX2 BUFX2_305 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf97) );
  BUFX2 BUFX2_306 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf96) );
  BUFX2 BUFX2_307 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf95) );
  BUFX2 BUFX2_308 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf94) );
  BUFX2 BUFX2_309 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf93) );
  BUFX2 BUFX2_31 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590), .Y(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf2) );
  BUFX2 BUFX2_310 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf92) );
  BUFX2 BUFX2_311 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf91) );
  BUFX2 BUFX2_312 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf90) );
  BUFX2 BUFX2_313 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf89) );
  BUFX2 BUFX2_314 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf88) );
  BUFX2 BUFX2_315 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf87) );
  BUFX2 BUFX2_316 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf86) );
  BUFX2 BUFX2_317 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf85) );
  BUFX2 BUFX2_318 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf84) );
  BUFX2 BUFX2_319 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf83) );
  BUFX2 BUFX2_32 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590), .Y(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf1) );
  BUFX2 BUFX2_320 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf82) );
  BUFX2 BUFX2_321 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf81) );
  BUFX2 BUFX2_322 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf80) );
  BUFX2 BUFX2_323 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf79) );
  BUFX2 BUFX2_324 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf78) );
  BUFX2 BUFX2_325 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf77) );
  BUFX2 BUFX2_326 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf76) );
  BUFX2 BUFX2_327 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf75) );
  BUFX2 BUFX2_328 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf74) );
  BUFX2 BUFX2_329 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf73) );
  BUFX2 BUFX2_33 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7590), .Y(REGFILE_SIM_reg_bank__abc_33898_n7590_bF_buf0) );
  BUFX2 BUFX2_330 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf72) );
  BUFX2 BUFX2_331 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf71) );
  BUFX2 BUFX2_332 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf70) );
  BUFX2 BUFX2_333 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf69) );
  BUFX2 BUFX2_334 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf68) );
  BUFX2 BUFX2_335 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf67) );
  BUFX2 BUFX2_336 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf66) );
  BUFX2 BUFX2_337 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf65) );
  BUFX2 BUFX2_338 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf64) );
  BUFX2 BUFX2_339 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf63) );
  BUFX2 BUFX2_34 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592), .Y(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf4) );
  BUFX2 BUFX2_340 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf62) );
  BUFX2 BUFX2_341 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf61) );
  BUFX2 BUFX2_342 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf60) );
  BUFX2 BUFX2_343 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf59) );
  BUFX2 BUFX2_344 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf58) );
  BUFX2 BUFX2_345 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf57) );
  BUFX2 BUFX2_346 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf56) );
  BUFX2 BUFX2_347 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf55) );
  BUFX2 BUFX2_348 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf54) );
  BUFX2 BUFX2_349 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf53) );
  BUFX2 BUFX2_35 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592), .Y(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf3) );
  BUFX2 BUFX2_350 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf52) );
  BUFX2 BUFX2_351 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf51) );
  BUFX2 BUFX2_352 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf50) );
  BUFX2 BUFX2_353 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf49) );
  BUFX2 BUFX2_354 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf48) );
  BUFX2 BUFX2_355 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf47) );
  BUFX2 BUFX2_356 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf46) );
  BUFX2 BUFX2_357 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf45) );
  BUFX2 BUFX2_358 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf44) );
  BUFX2 BUFX2_359 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf43) );
  BUFX2 BUFX2_36 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592), .Y(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf2) );
  BUFX2 BUFX2_360 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf42) );
  BUFX2 BUFX2_361 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf41) );
  BUFX2 BUFX2_362 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf40) );
  BUFX2 BUFX2_363 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf39) );
  BUFX2 BUFX2_364 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf38) );
  BUFX2 BUFX2_365 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf37) );
  BUFX2 BUFX2_366 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf36) );
  BUFX2 BUFX2_367 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf35) );
  BUFX2 BUFX2_368 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf34) );
  BUFX2 BUFX2_369 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf33) );
  BUFX2 BUFX2_37 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592), .Y(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf1) );
  BUFX2 BUFX2_370 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf32) );
  BUFX2 BUFX2_371 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf31) );
  BUFX2 BUFX2_372 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf30) );
  BUFX2 BUFX2_373 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf29) );
  BUFX2 BUFX2_374 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf28) );
  BUFX2 BUFX2_375 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf27) );
  BUFX2 BUFX2_376 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf26) );
  BUFX2 BUFX2_377 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf25) );
  BUFX2 BUFX2_378 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf24) );
  BUFX2 BUFX2_379 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf23) );
  BUFX2 BUFX2_38 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7592), .Y(REGFILE_SIM_reg_bank__abc_33898_n7592_bF_buf0) );
  BUFX2 BUFX2_380 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf22) );
  BUFX2 BUFX2_381 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf21) );
  BUFX2 BUFX2_382 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf20) );
  BUFX2 BUFX2_383 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf19) );
  BUFX2 BUFX2_384 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf18) );
  BUFX2 BUFX2_385 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf17) );
  BUFX2 BUFX2_386 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf16) );
  BUFX2 BUFX2_387 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf15) );
  BUFX2 BUFX2_388 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf14) );
  BUFX2 BUFX2_389 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf13) );
  BUFX2 BUFX2_39 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596), .Y(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf4) );
  BUFX2 BUFX2_390 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf12) );
  BUFX2 BUFX2_391 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf11) );
  BUFX2 BUFX2_392 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf10) );
  BUFX2 BUFX2_393 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf9) );
  BUFX2 BUFX2_394 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf8) );
  BUFX2 BUFX2_395 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf7) );
  BUFX2 BUFX2_396 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf6) );
  BUFX2 BUFX2_397 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf5) );
  BUFX2 BUFX2_398 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf4) );
  BUFX2 BUFX2_399 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf3) );
  BUFX2 BUFX2_4 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf5) );
  BUFX2 BUFX2_40 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596), .Y(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf3) );
  BUFX2 BUFX2_400 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf2) );
  BUFX2 BUFX2_401 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf1) );
  BUFX2 BUFX2_402 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf0) );
  BUFX2 BUFX2_403 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4) );
  BUFX2 BUFX2_404 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3) );
  BUFX2 BUFX2_405 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2) );
  BUFX2 BUFX2_406 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf1) );
  BUFX2 BUFX2_407 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf0) );
  BUFX2 BUFX2_408 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4) );
  BUFX2 BUFX2_409 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3) );
  BUFX2 BUFX2_41 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596), .Y(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf2) );
  BUFX2 BUFX2_410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2) );
  BUFX2 BUFX2_411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf1) );
  BUFX2 BUFX2_412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf0) );
  BUFX2 BUFX2_413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7) );
  BUFX2 BUFX2_414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf6) );
  BUFX2 BUFX2_415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5) );
  BUFX2 BUFX2_416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf4) );
  BUFX2 BUFX2_417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3) );
  BUFX2 BUFX2_418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf2) );
  BUFX2 BUFX2_419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1) );
  BUFX2 BUFX2_42 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596), .Y(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf1) );
  BUFX2 BUFX2_420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564), .Y(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf0) );
  BUFX2 BUFX2_421 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3) );
  BUFX2 BUFX2_422 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2) );
  BUFX2 BUFX2_423 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1) );
  BUFX2 BUFX2_424 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0) );
  BUFX2 BUFX2_425 ( .A(_abc_43815_n1428), .Y(_abc_43815_n1428_bF_buf4) );
  BUFX2 BUFX2_426 ( .A(_abc_43815_n1428), .Y(_abc_43815_n1428_bF_buf3) );
  BUFX2 BUFX2_427 ( .A(_abc_43815_n1428), .Y(_abc_43815_n1428_bF_buf2) );
  BUFX2 BUFX2_428 ( .A(_abc_43815_n1428), .Y(_abc_43815_n1428_bF_buf1) );
  BUFX2 BUFX2_429 ( .A(_abc_43815_n1428), .Y(_abc_43815_n1428_bF_buf0) );
  BUFX2 BUFX2_43 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7596), .Y(REGFILE_SIM_reg_bank__abc_33898_n7596_bF_buf0) );
  BUFX2 BUFX2_430 ( .A(alu__abc_41358_n1061), .Y(alu__abc_41358_n1061_bF_buf4) );
  BUFX2 BUFX2_431 ( .A(alu__abc_41358_n1061), .Y(alu__abc_41358_n1061_bF_buf3) );
  BUFX2 BUFX2_432 ( .A(alu__abc_41358_n1061), .Y(alu__abc_41358_n1061_bF_buf2) );
  BUFX2 BUFX2_433 ( .A(alu__abc_41358_n1061), .Y(alu__abc_41358_n1061_bF_buf1) );
  BUFX2 BUFX2_434 ( .A(alu__abc_41358_n1061), .Y(alu__abc_41358_n1061_bF_buf0) );
  BUFX2 BUFX2_435 ( .A(_abc_43815_n1399), .Y(_abc_43815_n1399_bF_buf4) );
  BUFX2 BUFX2_436 ( .A(_abc_43815_n1399), .Y(_abc_43815_n1399_bF_buf3) );
  BUFX2 BUFX2_437 ( .A(_abc_43815_n1399), .Y(_abc_43815_n1399_bF_buf2) );
  BUFX2 BUFX2_438 ( .A(_abc_43815_n1399), .Y(_abc_43815_n1399_bF_buf1) );
  BUFX2 BUFX2_439 ( .A(_abc_43815_n1399), .Y(_abc_43815_n1399_bF_buf0) );
  BUFX2 BUFX2_44 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599), .Y(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf4) );
  BUFX2 BUFX2_440 ( .A(_abc_43815_n3985_1), .Y(_abc_43815_n3985_1_bF_buf4) );
  BUFX2 BUFX2_441 ( .A(_abc_43815_n3985_1), .Y(_abc_43815_n3985_1_bF_buf3) );
  BUFX2 BUFX2_442 ( .A(_abc_43815_n3985_1), .Y(_abc_43815_n3985_1_bF_buf2) );
  BUFX2 BUFX2_443 ( .A(_abc_43815_n3985_1), .Y(_abc_43815_n3985_1_bF_buf1) );
  BUFX2 BUFX2_444 ( .A(_abc_43815_n3985_1), .Y(_abc_43815_n3985_1_bF_buf0) );
  BUFX2 BUFX2_445 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3) );
  BUFX2 BUFX2_446 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2) );
  BUFX2 BUFX2_447 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1) );
  BUFX2 BUFX2_448 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0) );
  BUFX2 BUFX2_449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7) );
  BUFX2 BUFX2_45 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599), .Y(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf3) );
  BUFX2 BUFX2_450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf6) );
  BUFX2 BUFX2_451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5) );
  BUFX2 BUFX2_452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf4) );
  BUFX2 BUFX2_453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3) );
  BUFX2 BUFX2_454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf2) );
  BUFX2 BUFX2_455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1) );
  BUFX2 BUFX2_456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889), .Y(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf0) );
  BUFX2 BUFX2_457 ( .A(state_q_1_), .Y(state_q_1_bF_buf4) );
  BUFX2 BUFX2_458 ( .A(state_q_1_), .Y(state_q_1_bF_buf3) );
  BUFX2 BUFX2_459 ( .A(state_q_1_), .Y(state_q_1_bF_buf2) );
  BUFX2 BUFX2_46 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599), .Y(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf2) );
  BUFX2 BUFX2_460 ( .A(state_q_1_), .Y(state_q_1_bF_buf1) );
  BUFX2 BUFX2_461 ( .A(state_q_1_), .Y(state_q_1_bF_buf0) );
  BUFX2 BUFX2_462 ( .A(alu__abc_41358_n294), .Y(alu__abc_41358_n294_bF_buf7) );
  BUFX2 BUFX2_463 ( .A(alu__abc_41358_n294), .Y(alu__abc_41358_n294_bF_buf6) );
  BUFX2 BUFX2_464 ( .A(alu__abc_41358_n294), .Y(alu__abc_41358_n294_bF_buf5) );
  BUFX2 BUFX2_465 ( .A(alu__abc_41358_n294), .Y(alu__abc_41358_n294_bF_buf4) );
  BUFX2 BUFX2_466 ( .A(alu__abc_41358_n294), .Y(alu__abc_41358_n294_bF_buf3) );
  BUFX2 BUFX2_467 ( .A(alu__abc_41358_n294), .Y(alu__abc_41358_n294_bF_buf2) );
  BUFX2 BUFX2_468 ( .A(alu__abc_41358_n294), .Y(alu__abc_41358_n294_bF_buf1) );
  BUFX2 BUFX2_469 ( .A(alu__abc_41358_n294), .Y(alu__abc_41358_n294_bF_buf0) );
  BUFX2 BUFX2_47 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599), .Y(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf1) );
  BUFX2 BUFX2_470 ( .A(alu__abc_41358_n299), .Y(alu__abc_41358_n299_bF_buf7) );
  BUFX2 BUFX2_471 ( .A(alu__abc_41358_n299), .Y(alu__abc_41358_n299_bF_buf6) );
  BUFX2 BUFX2_472 ( .A(alu__abc_41358_n299), .Y(alu__abc_41358_n299_bF_buf5) );
  BUFX2 BUFX2_473 ( .A(alu__abc_41358_n299), .Y(alu__abc_41358_n299_bF_buf4) );
  BUFX2 BUFX2_474 ( .A(alu__abc_41358_n299), .Y(alu__abc_41358_n299_bF_buf3) );
  BUFX2 BUFX2_475 ( .A(alu__abc_41358_n299), .Y(alu__abc_41358_n299_bF_buf2) );
  BUFX2 BUFX2_476 ( .A(alu__abc_41358_n299), .Y(alu__abc_41358_n299_bF_buf1) );
  BUFX2 BUFX2_477 ( .A(alu__abc_41358_n299), .Y(alu__abc_41358_n299_bF_buf0) );
  BUFX2 BUFX2_478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7) );
  BUFX2 BUFX2_479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf6) );
  BUFX2 BUFX2_48 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7599), .Y(REGFILE_SIM_reg_bank__abc_33898_n7599_bF_buf0) );
  BUFX2 BUFX2_480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5) );
  BUFX2 BUFX2_481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf4) );
  BUFX2 BUFX2_482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3) );
  BUFX2 BUFX2_483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf2) );
  BUFX2 BUFX2_484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1) );
  BUFX2 BUFX2_485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158), .Y(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf0) );
  BUFX2 BUFX2_486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441), .Y(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4) );
  BUFX2 BUFX2_487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441), .Y(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3) );
  BUFX2 BUFX2_488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441), .Y(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2) );
  BUFX2 BUFX2_489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441), .Y(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf1) );
  BUFX2 BUFX2_49 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf4) );
  BUFX2 BUFX2_490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441), .Y(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf0) );
  BUFX2 BUFX2_491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443), .Y(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4) );
  BUFX2 BUFX2_492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443), .Y(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3) );
  BUFX2 BUFX2_493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443), .Y(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf2) );
  BUFX2 BUFX2_494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443), .Y(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf1) );
  BUFX2 BUFX2_495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443), .Y(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf0) );
  BUFX2 BUFX2_496 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3) );
  BUFX2 BUFX2_497 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2) );
  BUFX2 BUFX2_498 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1) );
  BUFX2 BUFX2_499 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0) );
  BUFX2 BUFX2_5 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf4) );
  BUFX2 BUFX2_50 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf3) );
  BUFX2 BUFX2_500 ( .A(_abc_43815_n4217), .Y(_abc_43815_n4217_bF_buf4) );
  BUFX2 BUFX2_501 ( .A(_abc_43815_n4217), .Y(_abc_43815_n4217_bF_buf3) );
  BUFX2 BUFX2_502 ( .A(_abc_43815_n4217), .Y(_abc_43815_n4217_bF_buf2) );
  BUFX2 BUFX2_503 ( .A(_abc_43815_n4217), .Y(_abc_43815_n4217_bF_buf1) );
  BUFX2 BUFX2_504 ( .A(_abc_43815_n4217), .Y(_abc_43815_n4217_bF_buf0) );
  BUFX2 BUFX2_505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7) );
  BUFX2 BUFX2_506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf6) );
  BUFX2 BUFX2_507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5) );
  BUFX2 BUFX2_508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf4) );
  BUFX2 BUFX2_509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3) );
  BUFX2 BUFX2_51 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf2) );
  BUFX2 BUFX2_510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf2) );
  BUFX2 BUFX2_511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1) );
  BUFX2 BUFX2_512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913), .Y(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf0) );
  BUFX2 BUFX2_513 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3) );
  BUFX2 BUFX2_514 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2) );
  BUFX2 BUFX2_515 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1) );
  BUFX2 BUFX2_516 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0) );
  BUFX2 BUFX2_517 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3) );
  BUFX2 BUFX2_518 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2) );
  BUFX2 BUFX2_519 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1) );
  BUFX2 BUFX2_52 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf1) );
  BUFX2 BUFX2_520 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0) );
  BUFX2 BUFX2_521 ( .A(_abc_43815_n642_1), .Y(_abc_43815_n642_1_bF_buf5) );
  BUFX2 BUFX2_522 ( .A(_abc_43815_n642_1), .Y(_abc_43815_n642_1_bF_buf4) );
  BUFX2 BUFX2_523 ( .A(_abc_43815_n642_1), .Y(_abc_43815_n642_1_bF_buf3) );
  BUFX2 BUFX2_524 ( .A(_abc_43815_n642_1), .Y(_abc_43815_n642_1_bF_buf2) );
  BUFX2 BUFX2_525 ( .A(_abc_43815_n642_1), .Y(_abc_43815_n642_1_bF_buf1) );
  BUFX2 BUFX2_526 ( .A(_abc_43815_n642_1), .Y(_abc_43815_n642_1_bF_buf0) );
  BUFX2 BUFX2_527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791), .Y(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4) );
  BUFX2 BUFX2_528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791), .Y(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3) );
  BUFX2 BUFX2_529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791), .Y(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2) );
  BUFX2 BUFX2_53 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf0) );
  BUFX2 BUFX2_530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791), .Y(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf1) );
  BUFX2 BUFX2_531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791), .Y(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf0) );
  BUFX2 BUFX2_532 ( .A(_abc_43815_n1278), .Y(_abc_43815_n1278_bF_buf7) );
  BUFX2 BUFX2_533 ( .A(_abc_43815_n1278), .Y(_abc_43815_n1278_bF_buf6) );
  BUFX2 BUFX2_534 ( .A(_abc_43815_n1278), .Y(_abc_43815_n1278_bF_buf5) );
  BUFX2 BUFX2_535 ( .A(_abc_43815_n1278), .Y(_abc_43815_n1278_bF_buf4) );
  BUFX2 BUFX2_536 ( .A(_abc_43815_n1278), .Y(_abc_43815_n1278_bF_buf3) );
  BUFX2 BUFX2_537 ( .A(_abc_43815_n1278), .Y(_abc_43815_n1278_bF_buf2) );
  BUFX2 BUFX2_538 ( .A(_abc_43815_n1278), .Y(_abc_43815_n1278_bF_buf1) );
  BUFX2 BUFX2_539 ( .A(_abc_43815_n1278), .Y(_abc_43815_n1278_bF_buf0) );
  BUFX2 BUFX2_54 ( .A(_abc_43815_n645_1), .Y(_abc_43815_n645_1_bF_buf4) );
  BUFX2 BUFX2_540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061), .Y(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4) );
  BUFX2 BUFX2_541 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061), .Y(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3) );
  BUFX2 BUFX2_542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061), .Y(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf2) );
  BUFX2 BUFX2_543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061), .Y(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf1) );
  BUFX2 BUFX2_544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061), .Y(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf0) );
  BUFX2 BUFX2_545 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3) );
  BUFX2 BUFX2_546 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2) );
  BUFX2 BUFX2_547 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1) );
  BUFX2 BUFX2_548 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0) );
  BUFX2 BUFX2_549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641), .Y(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf4) );
  BUFX2 BUFX2_55 ( .A(_abc_43815_n645_1), .Y(_abc_43815_n645_1_bF_buf3) );
  BUFX2 BUFX2_550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641), .Y(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf3) );
  BUFX2 BUFX2_551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641), .Y(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf2) );
  BUFX2 BUFX2_552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641), .Y(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf1) );
  BUFX2 BUFX2_553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7641), .Y(REGFILE_SIM_reg_bank__abc_33898_n7641_bF_buf0) );
  BUFX2 BUFX2_554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643), .Y(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf4) );
  BUFX2 BUFX2_555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643), .Y(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf3) );
  BUFX2 BUFX2_556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643), .Y(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf2) );
  BUFX2 BUFX2_557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643), .Y(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf1) );
  BUFX2 BUFX2_558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7643), .Y(REGFILE_SIM_reg_bank__abc_33898_n7643_bF_buf0) );
  BUFX2 BUFX2_559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646), .Y(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf4) );
  BUFX2 BUFX2_56 ( .A(_abc_43815_n645_1), .Y(_abc_43815_n645_1_bF_buf2) );
  BUFX2 BUFX2_560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646), .Y(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf3) );
  BUFX2 BUFX2_561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646), .Y(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf2) );
  BUFX2 BUFX2_562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646), .Y(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf1) );
  BUFX2 BUFX2_563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7646), .Y(REGFILE_SIM_reg_bank__abc_33898_n7646_bF_buf0) );
  BUFX2 BUFX2_564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648), .Y(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf4) );
  BUFX2 BUFX2_565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648), .Y(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf3) );
  BUFX2 BUFX2_566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648), .Y(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf2) );
  BUFX2 BUFX2_567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648), .Y(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf1) );
  BUFX2 BUFX2_568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7648), .Y(REGFILE_SIM_reg_bank__abc_33898_n7648_bF_buf0) );
  BUFX2 BUFX2_569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7) );
  BUFX2 BUFX2_57 ( .A(_abc_43815_n645_1), .Y(_abc_43815_n645_1_bF_buf1) );
  BUFX2 BUFX2_570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf6) );
  BUFX2 BUFX2_571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5) );
  BUFX2 BUFX2_572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf4) );
  BUFX2 BUFX2_573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3) );
  BUFX2 BUFX2_574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf2) );
  BUFX2 BUFX2_575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1) );
  BUFX2 BUFX2_576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf0) );
  BUFX2 BUFX2_577 ( .A(_abc_43815_n692), .Y(_abc_43815_n692_bF_buf3) );
  BUFX2 BUFX2_578 ( .A(_abc_43815_n692), .Y(_abc_43815_n692_bF_buf2) );
  BUFX2 BUFX2_579 ( .A(_abc_43815_n692), .Y(_abc_43815_n692_bF_buf1) );
  BUFX2 BUFX2_58 ( .A(_abc_43815_n645_1), .Y(_abc_43815_n645_1_bF_buf0) );
  BUFX2 BUFX2_580 ( .A(_abc_43815_n692), .Y(_abc_43815_n692_bF_buf0) );
  BUFX2 BUFX2_581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7) );
  BUFX2 BUFX2_582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf6) );
  BUFX2 BUFX2_583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5) );
  BUFX2 BUFX2_584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf4) );
  BUFX2 BUFX2_585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3) );
  BUFX2 BUFX2_586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf2) );
  BUFX2 BUFX2_587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1) );
  BUFX2 BUFX2_588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf0) );
  BUFX2 BUFX2_589 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf6) );
  BUFX2 BUFX2_59 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3) );
  BUFX2 BUFX2_590 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf5) );
  BUFX2 BUFX2_591 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf4) );
  BUFX2 BUFX2_592 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf3) );
  BUFX2 BUFX2_593 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf2) );
  BUFX2 BUFX2_594 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf1) );
  BUFX2 BUFX2_595 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf0) );
  BUFX2 BUFX2_596 ( .A(_abc_43815_n2993_1), .Y(_abc_43815_n2993_1_bF_buf4) );
  BUFX2 BUFX2_597 ( .A(_abc_43815_n2993_1), .Y(_abc_43815_n2993_1_bF_buf3) );
  BUFX2 BUFX2_598 ( .A(_abc_43815_n2993_1), .Y(_abc_43815_n2993_1_bF_buf2) );
  BUFX2 BUFX2_599 ( .A(_abc_43815_n2993_1), .Y(_abc_43815_n2993_1_bF_buf1) );
  BUFX2 BUFX2_6 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf3) );
  BUFX2 BUFX2_60 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2) );
  BUFX2 BUFX2_600 ( .A(_abc_43815_n2993_1), .Y(_abc_43815_n2993_1_bF_buf0) );
  BUFX2 BUFX2_601 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3) );
  BUFX2 BUFX2_602 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2) );
  BUFX2 BUFX2_603 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1) );
  BUFX2 BUFX2_604 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0) );
  BUFX2 BUFX2_605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612), .Y(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf4) );
  BUFX2 BUFX2_606 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612), .Y(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf3) );
  BUFX2 BUFX2_607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612), .Y(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf2) );
  BUFX2 BUFX2_608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612), .Y(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf1) );
  BUFX2 BUFX2_609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7612), .Y(REGFILE_SIM_reg_bank__abc_33898_n7612_bF_buf0) );
  BUFX2 BUFX2_61 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1) );
  BUFX2 BUFX2_610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417), .Y(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4) );
  BUFX2 BUFX2_611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417), .Y(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3) );
  BUFX2 BUFX2_612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417), .Y(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2) );
  BUFX2 BUFX2_613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417), .Y(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf1) );
  BUFX2 BUFX2_614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417), .Y(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf0) );
  BUFX2 BUFX2_615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619), .Y(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf4) );
  BUFX2 BUFX2_616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619), .Y(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf3) );
  BUFX2 BUFX2_617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619), .Y(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf2) );
  BUFX2 BUFX2_618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619), .Y(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf1) );
  BUFX2 BUFX2_619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7619), .Y(REGFILE_SIM_reg_bank__abc_33898_n7619_bF_buf0) );
  BUFX2 BUFX2_62 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0) );
  BUFX2 BUFX2_620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419), .Y(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4) );
  BUFX2 BUFX2_621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419), .Y(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3) );
  BUFX2 BUFX2_622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419), .Y(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf2) );
  BUFX2 BUFX2_623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419), .Y(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf1) );
  BUFX2 BUFX2_624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419), .Y(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf0) );
  BUFX2 BUFX2_625 ( .A(alu__abc_41358_n932), .Y(alu__abc_41358_n932_bF_buf4) );
  BUFX2 BUFX2_626 ( .A(alu__abc_41358_n932), .Y(alu__abc_41358_n932_bF_buf3) );
  BUFX2 BUFX2_627 ( .A(alu__abc_41358_n932), .Y(alu__abc_41358_n932_bF_buf2) );
  BUFX2 BUFX2_628 ( .A(alu__abc_41358_n932), .Y(alu__abc_41358_n932_bF_buf1) );
  BUFX2 BUFX2_629 ( .A(alu__abc_41358_n932), .Y(alu__abc_41358_n932_bF_buf0) );
  BUFX2 BUFX2_63 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337), .Y(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4) );
  BUFX2 BUFX2_630 ( .A(alu__abc_41358_n935), .Y(alu__abc_41358_n935_bF_buf4) );
  BUFX2 BUFX2_631 ( .A(alu__abc_41358_n935), .Y(alu__abc_41358_n935_bF_buf3) );
  BUFX2 BUFX2_632 ( .A(alu__abc_41358_n935), .Y(alu__abc_41358_n935_bF_buf2) );
  BUFX2 BUFX2_633 ( .A(alu__abc_41358_n935), .Y(alu__abc_41358_n935_bF_buf1) );
  BUFX2 BUFX2_634 ( .A(alu__abc_41358_n935), .Y(alu__abc_41358_n935_bF_buf0) );
  BUFX2 BUFX2_635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582), .Y(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf4) );
  BUFX2 BUFX2_636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582), .Y(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf3) );
  BUFX2 BUFX2_637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582), .Y(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf2) );
  BUFX2 BUFX2_638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582), .Y(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf1) );
  BUFX2 BUFX2_639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7582), .Y(REGFILE_SIM_reg_bank__abc_33898_n7582_bF_buf0) );
  BUFX2 BUFX2_64 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337), .Y(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3) );
  BUFX2 BUFX2_640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585), .Y(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf4) );
  BUFX2 BUFX2_641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585), .Y(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf3) );
  BUFX2 BUFX2_642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585), .Y(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf2) );
  BUFX2 BUFX2_643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585), .Y(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf1) );
  BUFX2 BUFX2_644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7585), .Y(REGFILE_SIM_reg_bank__abc_33898_n7585_bF_buf0) );
  BUFX2 BUFX2_645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4) );
  BUFX2 BUFX2_646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3) );
  BUFX2 BUFX2_647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf2) );
  BUFX2 BUFX2_648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf1) );
  BUFX2 BUFX2_649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf0) );
  BUFX2 BUFX2_65 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337), .Y(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2) );
  BUFX2 BUFX2_650 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3) );
  BUFX2 BUFX2_651 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2) );
  BUFX2 BUFX2_652 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1) );
  BUFX2 BUFX2_653 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0) );
  BUFX2 BUFX2_654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7) );
  BUFX2 BUFX2_655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf6) );
  BUFX2 BUFX2_656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5) );
  BUFX2 BUFX2_657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf4) );
  BUFX2 BUFX2_658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3) );
  BUFX2 BUFX2_659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf2) );
  BUFX2 BUFX2_66 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337), .Y(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf1) );
  BUFX2 BUFX2_660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1) );
  BUFX2 BUFX2_661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf0) );
  BUFX2 BUFX2_662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554), .Y(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf4) );
  BUFX2 BUFX2_663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554), .Y(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf3) );
  BUFX2 BUFX2_664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554), .Y(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf2) );
  BUFX2 BUFX2_665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554), .Y(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf1) );
  BUFX2 BUFX2_666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7554), .Y(REGFILE_SIM_reg_bank__abc_33898_n7554_bF_buf0) );
  BUFX2 BUFX2_667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557), .Y(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf4) );
  BUFX2 BUFX2_668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557), .Y(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf3) );
  BUFX2 BUFX2_669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557), .Y(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf2) );
  BUFX2 BUFX2_67 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337), .Y(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf0) );
  BUFX2 BUFX2_670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557), .Y(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf1) );
  BUFX2 BUFX2_671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7557), .Y(REGFILE_SIM_reg_bank__abc_33898_n7557_bF_buf0) );
  BUFX2 BUFX2_672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643), .Y(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf4) );
  BUFX2 BUFX2_673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643), .Y(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf3) );
  BUFX2 BUFX2_674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643), .Y(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf2) );
  BUFX2 BUFX2_675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643), .Y(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf1) );
  BUFX2 BUFX2_676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5643), .Y(REGFILE_SIM_reg_bank__abc_33898_n5643_bF_buf0) );
  BUFX2 BUFX2_677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645), .Y(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf4) );
  BUFX2 BUFX2_678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645), .Y(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf3) );
  BUFX2 BUFX2_679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645), .Y(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf2) );
  BUFX2 BUFX2_68 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339), .Y(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4) );
  BUFX2 BUFX2_680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645), .Y(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf1) );
  BUFX2 BUFX2_681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5645), .Y(REGFILE_SIM_reg_bank__abc_33898_n5645_bF_buf0) );
  BUFX2 BUFX2_682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648), .Y(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf4) );
  BUFX2 BUFX2_683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648), .Y(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf3) );
  BUFX2 BUFX2_684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648), .Y(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf2) );
  BUFX2 BUFX2_685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648), .Y(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf1) );
  BUFX2 BUFX2_686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5648), .Y(REGFILE_SIM_reg_bank__abc_33898_n5648_bF_buf0) );
  BUFX2 BUFX2_687 ( .A(_abc_43815_n986), .Y(_abc_43815_n986_bF_buf4) );
  BUFX2 BUFX2_688 ( .A(_abc_43815_n986), .Y(_abc_43815_n986_bF_buf3) );
  BUFX2 BUFX2_689 ( .A(_abc_43815_n986), .Y(_abc_43815_n986_bF_buf2) );
  BUFX2 BUFX2_69 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339), .Y(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3) );
  BUFX2 BUFX2_690 ( .A(_abc_43815_n986), .Y(_abc_43815_n986_bF_buf1) );
  BUFX2 BUFX2_691 ( .A(_abc_43815_n986), .Y(_abc_43815_n986_bF_buf0) );
  BUFX2 BUFX2_692 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3) );
  BUFX2 BUFX2_693 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2) );
  BUFX2 BUFX2_694 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1) );
  BUFX2 BUFX2_695 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0) );
  BUFX2 BUFX2_696 ( .A(_abc_43815_n1425_1), .Y(_abc_43815_n1425_1_bF_buf4) );
  BUFX2 BUFX2_697 ( .A(_abc_43815_n1425_1), .Y(_abc_43815_n1425_1_bF_buf3) );
  BUFX2 BUFX2_698 ( .A(_abc_43815_n1425_1), .Y(_abc_43815_n1425_1_bF_buf2) );
  BUFX2 BUFX2_699 ( .A(_abc_43815_n1425_1), .Y(_abc_43815_n1425_1_bF_buf1) );
  BUFX2 BUFX2_7 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf2) );
  BUFX2 BUFX2_70 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339), .Y(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf2) );
  BUFX2 BUFX2_700 ( .A(_abc_43815_n1425_1), .Y(_abc_43815_n1425_1_bF_buf0) );
  BUFX2 BUFX2_701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610), .Y(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf4) );
  BUFX2 BUFX2_702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610), .Y(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf3) );
  BUFX2 BUFX2_703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610), .Y(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf2) );
  BUFX2 BUFX2_704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610), .Y(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf1) );
  BUFX2 BUFX2_705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5610), .Y(REGFILE_SIM_reg_bank__abc_33898_n5610_bF_buf0) );
  BUFX2 BUFX2_706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613), .Y(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf4) );
  BUFX2 BUFX2_707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613), .Y(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf3) );
  BUFX2 BUFX2_708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613), .Y(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf2) );
  BUFX2 BUFX2_709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613), .Y(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf1) );
  BUFX2 BUFX2_71 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339), .Y(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf1) );
  BUFX2 BUFX2_710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5613), .Y(REGFILE_SIM_reg_bank__abc_33898_n5613_bF_buf0) );
  BUFX2 BUFX2_711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616), .Y(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf4) );
  BUFX2 BUFX2_712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616), .Y(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf3) );
  BUFX2 BUFX2_713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616), .Y(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf2) );
  BUFX2 BUFX2_714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616), .Y(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf1) );
  BUFX2 BUFX2_715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5616), .Y(REGFILE_SIM_reg_bank__abc_33898_n5616_bF_buf0) );
  BUFX2 BUFX2_716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618), .Y(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf4) );
  BUFX2 BUFX2_717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618), .Y(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf3) );
  BUFX2 BUFX2_718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618), .Y(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf2) );
  BUFX2 BUFX2_719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618), .Y(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf1) );
  BUFX2 BUFX2_72 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339), .Y(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf0) );
  BUFX2 BUFX2_720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5618), .Y(REGFILE_SIM_reg_bank__abc_33898_n5618_bF_buf0) );
  BUFX2 BUFX2_721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581), .Y(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf4) );
  BUFX2 BUFX2_722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581), .Y(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf3) );
  BUFX2 BUFX2_723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581), .Y(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf2) );
  BUFX2 BUFX2_724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581), .Y(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf1) );
  BUFX2 BUFX2_725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5581), .Y(REGFILE_SIM_reg_bank__abc_33898_n5581_bF_buf0) );
  BUFX2 BUFX2_726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583), .Y(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf4) );
  BUFX2 BUFX2_727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583), .Y(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf3) );
  BUFX2 BUFX2_728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583), .Y(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf2) );
  BUFX2 BUFX2_729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583), .Y(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf1) );
  BUFX2 BUFX2_73 ( .A(_abc_43815_n641), .Y(_abc_43815_n641_bF_buf3) );
  BUFX2 BUFX2_730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5583), .Y(REGFILE_SIM_reg_bank__abc_33898_n5583_bF_buf0) );
  BUFX2 BUFX2_731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587), .Y(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf4) );
  BUFX2 BUFX2_732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587), .Y(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf3) );
  BUFX2 BUFX2_733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587), .Y(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf2) );
  BUFX2 BUFX2_734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587), .Y(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf1) );
  BUFX2 BUFX2_735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5587), .Y(REGFILE_SIM_reg_bank__abc_33898_n5587_bF_buf0) );
  BUFX2 BUFX2_736 ( .A(_abc_43815_n686_1), .Y(_abc_43815_n686_1_bF_buf4) );
  BUFX2 BUFX2_737 ( .A(_abc_43815_n686_1), .Y(_abc_43815_n686_1_bF_buf3) );
  BUFX2 BUFX2_738 ( .A(_abc_43815_n686_1), .Y(_abc_43815_n686_1_bF_buf2) );
  BUFX2 BUFX2_739 ( .A(_abc_43815_n686_1), .Y(_abc_43815_n686_1_bF_buf1) );
  BUFX2 BUFX2_74 ( .A(_abc_43815_n641), .Y(_abc_43815_n641_bF_buf2) );
  BUFX2 BUFX2_740 ( .A(_abc_43815_n686_1), .Y(_abc_43815_n686_1_bF_buf0) );
  BUFX2 BUFX2_741 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3) );
  BUFX2 BUFX2_742 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2) );
  BUFX2 BUFX2_743 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1) );
  BUFX2 BUFX2_744 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0) );
  BUFX2 BUFX2_745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7) );
  BUFX2 BUFX2_746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf6) );
  BUFX2 BUFX2_747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5) );
  BUFX2 BUFX2_748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf4) );
  BUFX2 BUFX2_749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3) );
  BUFX2 BUFX2_75 ( .A(_abc_43815_n641), .Y(_abc_43815_n641_bF_buf1) );
  BUFX2 BUFX2_750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf2) );
  BUFX2 BUFX2_751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1) );
  BUFX2 BUFX2_752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf0) );
  BUFX2 BUFX2_753 ( .A(_abc_43815_n1473), .Y(_abc_43815_n1473_bF_buf4) );
  BUFX2 BUFX2_754 ( .A(_abc_43815_n1473), .Y(_abc_43815_n1473_bF_buf3) );
  BUFX2 BUFX2_755 ( .A(_abc_43815_n1473), .Y(_abc_43815_n1473_bF_buf2) );
  BUFX2 BUFX2_756 ( .A(_abc_43815_n1473), .Y(_abc_43815_n1473_bF_buf1) );
  BUFX2 BUFX2_757 ( .A(_abc_43815_n1473), .Y(_abc_43815_n1473_bF_buf0) );
  BUFX2 BUFX2_758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239), .Y(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4) );
  BUFX2 BUFX2_759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239), .Y(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3) );
  BUFX2 BUFX2_76 ( .A(_abc_43815_n641), .Y(_abc_43815_n641_bF_buf0) );
  BUFX2 BUFX2_760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239), .Y(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2) );
  BUFX2 BUFX2_761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239), .Y(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf1) );
  BUFX2 BUFX2_762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239), .Y(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf0) );
  BUFX2 BUFX2_763 ( .A(_abc_43815_n3002), .Y(_abc_43815_n3002_bF_buf4) );
  BUFX2 BUFX2_764 ( .A(_abc_43815_n3002), .Y(_abc_43815_n3002_bF_buf3) );
  BUFX2 BUFX2_765 ( .A(_abc_43815_n3002), .Y(_abc_43815_n3002_bF_buf2) );
  BUFX2 BUFX2_766 ( .A(_abc_43815_n3002), .Y(_abc_43815_n3002_bF_buf1) );
  BUFX2 BUFX2_767 ( .A(_abc_43815_n3002), .Y(_abc_43815_n3002_bF_buf0) );
  BUFX2 BUFX2_768 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554), .Y(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf4) );
  BUFX2 BUFX2_769 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554), .Y(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf3) );
  BUFX2 BUFX2_77 ( .A(_abc_43815_n649), .Y(_abc_43815_n649_bF_buf4) );
  BUFX2 BUFX2_770 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554), .Y(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf2) );
  BUFX2 BUFX2_771 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554), .Y(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf1) );
  BUFX2 BUFX2_772 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5554), .Y(REGFILE_SIM_reg_bank__abc_33898_n5554_bF_buf0) );
  BUFX2 BUFX2_773 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557), .Y(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf4) );
  BUFX2 BUFX2_774 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557), .Y(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf3) );
  BUFX2 BUFX2_775 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557), .Y(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf2) );
  BUFX2 BUFX2_776 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557), .Y(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf1) );
  BUFX2 BUFX2_777 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5557), .Y(REGFILE_SIM_reg_bank__abc_33898_n5557_bF_buf0) );
  BUFX2 BUFX2_778 ( .A(_abc_43815_n1060), .Y(_abc_43815_n1060_bF_buf3) );
  BUFX2 BUFX2_779 ( .A(_abc_43815_n1060), .Y(_abc_43815_n1060_bF_buf2) );
  BUFX2 BUFX2_78 ( .A(_abc_43815_n649), .Y(_abc_43815_n649_bF_buf3) );
  BUFX2 BUFX2_780 ( .A(_abc_43815_n1060), .Y(_abc_43815_n1060_bF_buf1) );
  BUFX2 BUFX2_781 ( .A(_abc_43815_n1060), .Y(_abc_43815_n1060_bF_buf0) );
  BUFX2 BUFX2_782 ( .A(_abc_43815_n1472_1), .Y(_abc_43815_n1472_1_bF_buf4) );
  BUFX2 BUFX2_783 ( .A(_abc_43815_n1472_1), .Y(_abc_43815_n1472_1_bF_buf3) );
  BUFX2 BUFX2_784 ( .A(_abc_43815_n1472_1), .Y(_abc_43815_n1472_1_bF_buf2) );
  BUFX2 BUFX2_785 ( .A(_abc_43815_n1472_1), .Y(_abc_43815_n1472_1_bF_buf1) );
  BUFX2 BUFX2_786 ( .A(_abc_43815_n1472_1), .Y(_abc_43815_n1472_1_bF_buf0) );
  BUFX2 BUFX2_787 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4) );
  BUFX2 BUFX2_788 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3) );
  BUFX2 BUFX2_789 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2) );
  BUFX2 BUFX2_79 ( .A(_abc_43815_n649), .Y(_abc_43815_n649_bF_buf2) );
  BUFX2 BUFX2_790 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf1) );
  BUFX2 BUFX2_791 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf0) );
  BUFX2 BUFX2_792 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147), .Y(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4) );
  BUFX2 BUFX2_793 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147), .Y(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3) );
  BUFX2 BUFX2_794 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147), .Y(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2) );
  BUFX2 BUFX2_795 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147), .Y(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf1) );
  BUFX2 BUFX2_796 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147), .Y(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf0) );
  BUFX2 BUFX2_797 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149), .Y(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4) );
  BUFX2 BUFX2_798 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149), .Y(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3) );
  BUFX2 BUFX2_799 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149), .Y(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf2) );
  BUFX2 BUFX2_8 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf1) );
  BUFX2 BUFX2_80 ( .A(_abc_43815_n649), .Y(_abc_43815_n649_bF_buf1) );
  BUFX2 BUFX2_800 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149), .Y(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf1) );
  BUFX2 BUFX2_801 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149), .Y(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf0) );
  BUFX2 BUFX2_802 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3) );
  BUFX2 BUFX2_803 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2) );
  BUFX2 BUFX2_804 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1) );
  BUFX2 BUFX2_805 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0) );
  BUFX2 BUFX2_806 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616), .Y(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4) );
  BUFX2 BUFX2_807 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616), .Y(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3) );
  BUFX2 BUFX2_808 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616), .Y(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2) );
  BUFX2 BUFX2_809 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616), .Y(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf1) );
  BUFX2 BUFX2_81 ( .A(_abc_43815_n649), .Y(_abc_43815_n649_bF_buf0) );
  BUFX2 BUFX2_810 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616), .Y(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf0) );
  BUFX2 BUFX2_811 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618), .Y(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4) );
  BUFX2 BUFX2_812 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618), .Y(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3) );
  BUFX2 BUFX2_813 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618), .Y(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf2) );
  BUFX2 BUFX2_814 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618), .Y(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf1) );
  BUFX2 BUFX2_815 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618), .Y(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf0) );
  BUFX2 BUFX2_816 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267), .Y(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4) );
  BUFX2 BUFX2_817 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267), .Y(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3) );
  BUFX2 BUFX2_818 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267), .Y(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2) );
  BUFX2 BUFX2_819 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267), .Y(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf1) );
  BUFX2 BUFX2_82 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563), .Y(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf4) );
  BUFX2 BUFX2_820 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267), .Y(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf0) );
  BUFX2 BUFX2_821 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3) );
  BUFX2 BUFX2_822 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2) );
  BUFX2 BUFX2_823 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1) );
  BUFX2 BUFX2_824 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0) );
  BUFX2 BUFX2_825 ( .A(_abc_43815_n1413), .Y(_abc_43815_n1413_bF_buf4) );
  BUFX2 BUFX2_826 ( .A(_abc_43815_n1413), .Y(_abc_43815_n1413_bF_buf3) );
  BUFX2 BUFX2_827 ( .A(_abc_43815_n1413), .Y(_abc_43815_n1413_bF_buf2) );
  BUFX2 BUFX2_828 ( .A(_abc_43815_n1413), .Y(_abc_43815_n1413_bF_buf1) );
  BUFX2 BUFX2_829 ( .A(_abc_43815_n1413), .Y(_abc_43815_n1413_bF_buf0) );
  BUFX2 BUFX2_83 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563), .Y(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf3) );
  BUFX2 BUFX2_830 ( .A(_abc_43815_n1418), .Y(_abc_43815_n1418_bF_buf5) );
  BUFX2 BUFX2_831 ( .A(_abc_43815_n1418), .Y(_abc_43815_n1418_bF_buf4) );
  BUFX2 BUFX2_832 ( .A(_abc_43815_n1418), .Y(_abc_43815_n1418_bF_buf3) );
  BUFX2 BUFX2_833 ( .A(_abc_43815_n1418), .Y(_abc_43815_n1418_bF_buf2) );
  BUFX2 BUFX2_834 ( .A(_abc_43815_n1418), .Y(_abc_43815_n1418_bF_buf1) );
  BUFX2 BUFX2_835 ( .A(_abc_43815_n1418), .Y(_abc_43815_n1418_bF_buf0) );
  BUFX2 BUFX2_836 ( .A(alu__abc_41358_n1057), .Y(alu__abc_41358_n1057_bF_buf4) );
  BUFX2 BUFX2_837 ( .A(alu__abc_41358_n1057), .Y(alu__abc_41358_n1057_bF_buf3) );
  BUFX2 BUFX2_838 ( .A(alu__abc_41358_n1057), .Y(alu__abc_41358_n1057_bF_buf2) );
  BUFX2 BUFX2_839 ( .A(alu__abc_41358_n1057), .Y(alu__abc_41358_n1057_bF_buf1) );
  BUFX2 BUFX2_84 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563), .Y(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf2) );
  BUFX2 BUFX2_840 ( .A(alu__abc_41358_n1057), .Y(alu__abc_41358_n1057_bF_buf0) );
  BUFX2 BUFX2_841 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140), .Y(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4) );
  BUFX2 BUFX2_842 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140), .Y(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3) );
  BUFX2 BUFX2_843 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140), .Y(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2) );
  BUFX2 BUFX2_844 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140), .Y(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf1) );
  BUFX2 BUFX2_845 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140), .Y(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf0) );
  BUFX2 BUFX2_846 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142), .Y(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4) );
  BUFX2 BUFX2_847 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142), .Y(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3) );
  BUFX2 BUFX2_848 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142), .Y(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf2) );
  BUFX2 BUFX2_849 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142), .Y(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf1) );
  BUFX2 BUFX2_85 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563), .Y(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf1) );
  BUFX2 BUFX2_850 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142), .Y(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf0) );
  BUFX2 BUFX2_851 ( .A(state_q_3_), .Y(state_q_3_bF_buf5) );
  BUFX2 BUFX2_852 ( .A(state_q_3_), .Y(state_q_3_bF_buf4) );
  BUFX2 BUFX2_853 ( .A(state_q_3_), .Y(state_q_3_bF_buf3) );
  BUFX2 BUFX2_854 ( .A(state_q_3_), .Y(state_q_3_bF_buf2) );
  BUFX2 BUFX2_855 ( .A(state_q_3_), .Y(state_q_3_bF_buf1) );
  BUFX2 BUFX2_856 ( .A(state_q_3_), .Y(state_q_3_bF_buf0) );
  BUFX2 BUFX2_857 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3) );
  BUFX2 BUFX2_858 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2) );
  BUFX2 BUFX2_859 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1) );
  BUFX2 BUFX2_86 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7563), .Y(REGFILE_SIM_reg_bank__abc_33898_n7563_bF_buf0) );
  BUFX2 BUFX2_860 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0) );
  BUFX2 BUFX2_861 ( .A(_abc_43815_n1350), .Y(_abc_43815_n1350_bF_buf4) );
  BUFX2 BUFX2_862 ( .A(_abc_43815_n1350), .Y(_abc_43815_n1350_bF_buf3) );
  BUFX2 BUFX2_863 ( .A(_abc_43815_n1350), .Y(_abc_43815_n1350_bF_buf2) );
  BUFX2 BUFX2_864 ( .A(_abc_43815_n1350), .Y(_abc_43815_n1350_bF_buf1) );
  BUFX2 BUFX2_865 ( .A(_abc_43815_n1350), .Y(_abc_43815_n1350_bF_buf0) );
  BUFX2 BUFX2_866 ( .A(_abc_43815_n1351), .Y(_abc_43815_n1351_bF_buf4) );
  BUFX2 BUFX2_867 ( .A(_abc_43815_n1351), .Y(_abc_43815_n1351_bF_buf3) );
  BUFX2 BUFX2_868 ( .A(_abc_43815_n1351), .Y(_abc_43815_n1351_bF_buf2) );
  BUFX2 BUFX2_869 ( .A(_abc_43815_n1351), .Y(_abc_43815_n1351_bF_buf1) );
  BUFX2 BUFX2_87 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566), .Y(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf4) );
  BUFX2 BUFX2_870 ( .A(_abc_43815_n1351), .Y(_abc_43815_n1351_bF_buf0) );
  BUFX2 BUFX2_871 ( .A(enable_i), .Y(enable_i_bF_buf7) );
  BUFX2 BUFX2_872 ( .A(enable_i), .Y(enable_i_bF_buf6) );
  BUFX2 BUFX2_873 ( .A(enable_i), .Y(enable_i_bF_buf5) );
  BUFX2 BUFX2_874 ( .A(enable_i), .Y(enable_i_bF_buf4) );
  BUFX2 BUFX2_875 ( .A(enable_i), .Y(enable_i_bF_buf3) );
  BUFX2 BUFX2_876 ( .A(enable_i), .Y(enable_i_bF_buf2) );
  BUFX2 BUFX2_877 ( .A(enable_i), .Y(enable_i_bF_buf1) );
  BUFX2 BUFX2_878 ( .A(enable_i), .Y(enable_i_bF_buf0) );
  BUFX2 BUFX2_879 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3) );
  BUFX2 BUFX2_88 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566), .Y(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf3) );
  BUFX2 BUFX2_880 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2) );
  BUFX2 BUFX2_881 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1) );
  BUFX2 BUFX2_882 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0) );
  BUFX2 BUFX2_883 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4) );
  BUFX2 BUFX2_884 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3) );
  BUFX2 BUFX2_885 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2) );
  BUFX2 BUFX2_886 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf1) );
  BUFX2 BUFX2_887 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf0) );
  BUFX2 BUFX2_888 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4) );
  BUFX2 BUFX2_889 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3) );
  BUFX2 BUFX2_89 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566), .Y(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf2) );
  BUFX2 BUFX2_890 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2) );
  BUFX2 BUFX2_891 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf1) );
  BUFX2 BUFX2_892 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf0) );
  BUFX2 BUFX2_893 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3) );
  BUFX2 BUFX2_894 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2) );
  BUFX2 BUFX2_895 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1) );
  BUFX2 BUFX2_896 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0) );
  BUFX2 BUFX2_897 ( .A(_abc_43815_n646_1), .Y(_abc_43815_n646_1_bF_buf3) );
  BUFX2 BUFX2_898 ( .A(_abc_43815_n646_1), .Y(_abc_43815_n646_1_bF_buf2) );
  BUFX2 BUFX2_899 ( .A(_abc_43815_n646_1), .Y(_abc_43815_n646_1_bF_buf1) );
  BUFX2 BUFX2_9 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245_hier0_bF_buf0) );
  BUFX2 BUFX2_90 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566), .Y(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf1) );
  BUFX2 BUFX2_900 ( .A(_abc_43815_n646_1), .Y(_abc_43815_n646_1_bF_buf0) );
  BUFX2 BUFX2_901 ( .A(alu__abc_41358_n252), .Y(alu__abc_41358_n252_bF_buf6) );
  BUFX2 BUFX2_902 ( .A(alu__abc_41358_n252), .Y(alu__abc_41358_n252_bF_buf5) );
  BUFX2 BUFX2_903 ( .A(alu__abc_41358_n252), .Y(alu__abc_41358_n252_bF_buf4) );
  BUFX2 BUFX2_904 ( .A(alu__abc_41358_n252), .Y(alu__abc_41358_n252_bF_buf3) );
  BUFX2 BUFX2_905 ( .A(alu__abc_41358_n252), .Y(alu__abc_41358_n252_bF_buf2) );
  BUFX2 BUFX2_906 ( .A(alu__abc_41358_n252), .Y(alu__abc_41358_n252_bF_buf1) );
  BUFX2 BUFX2_907 ( .A(alu__abc_41358_n252), .Y(alu__abc_41358_n252_bF_buf0) );
  BUFX2 BUFX2_908 ( .A(alu__abc_41358_n259), .Y(alu__abc_41358_n259_bF_buf4) );
  BUFX2 BUFX2_909 ( .A(alu__abc_41358_n259), .Y(alu__abc_41358_n259_bF_buf3) );
  BUFX2 BUFX2_91 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7566), .Y(REGFILE_SIM_reg_bank__abc_33898_n7566_bF_buf0) );
  BUFX2 BUFX2_910 ( .A(alu__abc_41358_n259), .Y(alu__abc_41358_n259_bF_buf2) );
  BUFX2 BUFX2_911 ( .A(alu__abc_41358_n259), .Y(alu__abc_41358_n259_bF_buf1) );
  BUFX2 BUFX2_912 ( .A(alu__abc_41358_n259), .Y(alu__abc_41358_n259_bF_buf0) );
  BUFX2 BUFX2_913 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7) );
  BUFX2 BUFX2_914 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf6) );
  BUFX2 BUFX2_915 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5) );
  BUFX2 BUFX2_916 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf4) );
  BUFX2 BUFX2_917 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3) );
  BUFX2 BUFX2_918 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf2) );
  BUFX2 BUFX2_919 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1) );
  BUFX2 BUFX2_92 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650), .Y(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf4) );
  BUFX2 BUFX2_920 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435), .Y(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf0) );
  BUFX2 BUFX2_921 ( .A(_abc_43815_n2991), .Y(_abc_43815_n2991_bF_buf4) );
  BUFX2 BUFX2_922 ( .A(_abc_43815_n2991), .Y(_abc_43815_n2991_bF_buf3) );
  BUFX2 BUFX2_923 ( .A(_abc_43815_n2991), .Y(_abc_43815_n2991_bF_buf2) );
  BUFX2 BUFX2_924 ( .A(_abc_43815_n2991), .Y(_abc_43815_n2991_bF_buf1) );
  BUFX2 BUFX2_925 ( .A(_abc_43815_n2991), .Y(_abc_43815_n2991_bF_buf0) );
  BUFX2 BUFX2_926 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3) );
  BUFX2 BUFX2_927 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2) );
  BUFX2 BUFX2_928 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1) );
  BUFX2 BUFX2_929 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0) );
  BUFX2 BUFX2_93 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650), .Y(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf3) );
  BUFX2 BUFX2_930 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3) );
  BUFX2 BUFX2_931 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2) );
  BUFX2 BUFX2_932 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1) );
  BUFX2 BUFX2_933 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0) );
  BUFX2 BUFX2_934 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf4) );
  BUFX2 BUFX2_935 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf3) );
  BUFX2 BUFX2_936 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf2) );
  BUFX2 BUFX2_937 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf1) );
  BUFX2 BUFX2_938 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf0) );
  BUFX2 BUFX2_939 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343), .Y(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4) );
  BUFX2 BUFX2_94 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650), .Y(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf2) );
  BUFX2 BUFX2_940 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343), .Y(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3) );
  BUFX2 BUFX2_941 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343), .Y(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2) );
  BUFX2 BUFX2_942 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343), .Y(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf1) );
  BUFX2 BUFX2_943 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343), .Y(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf0) );
  BUFX2 BUFX2_944 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345), .Y(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4) );
  BUFX2 BUFX2_945 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345), .Y(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3) );
  BUFX2 BUFX2_946 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345), .Y(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf2) );
  BUFX2 BUFX2_947 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345), .Y(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf1) );
  BUFX2 BUFX2_948 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345), .Y(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf0) );
  BUFX2 BUFX2_949 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3) );
  BUFX2 BUFX2_95 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650), .Y(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf1) );
  BUFX2 BUFX2_950 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2) );
  BUFX2 BUFX2_951 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1) );
  BUFX2 BUFX2_952 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0) );
  BUFX2 BUFX2_953 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632), .Y(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf4) );
  BUFX2 BUFX2_954 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632), .Y(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf3) );
  BUFX2 BUFX2_955 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632), .Y(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf2) );
  BUFX2 BUFX2_956 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632), .Y(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf1) );
  BUFX2 BUFX2_957 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7632), .Y(REGFILE_SIM_reg_bank__abc_33898_n7632_bF_buf0) );
  BUFX2 BUFX2_958 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634), .Y(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf4) );
  BUFX2 BUFX2_959 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634), .Y(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf3) );
  BUFX2 BUFX2_96 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5650), .Y(REGFILE_SIM_reg_bank__abc_33898_n5650_bF_buf0) );
  BUFX2 BUFX2_960 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634), .Y(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf2) );
  BUFX2 BUFX2_961 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634), .Y(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf1) );
  BUFX2 BUFX2_962 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7634), .Y(REGFILE_SIM_reg_bank__abc_33898_n7634_bF_buf0) );
  BUFX2 BUFX2_963 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636), .Y(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf4) );
  BUFX2 BUFX2_964 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636), .Y(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf3) );
  BUFX2 BUFX2_965 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636), .Y(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf2) );
  BUFX2 BUFX2_966 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636), .Y(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf1) );
  BUFX2 BUFX2_967 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7636), .Y(REGFILE_SIM_reg_bank__abc_33898_n7636_bF_buf0) );
  BUFX2 BUFX2_968 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813), .Y(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4) );
  BUFX2 BUFX2_969 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813), .Y(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3) );
  BUFX2 BUFX2_97 ( .A(_abc_43815_n1431_1), .Y(_abc_43815_n1431_1_bF_buf4) );
  BUFX2 BUFX2_970 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813), .Y(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2) );
  BUFX2 BUFX2_971 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813), .Y(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf1) );
  BUFX2 BUFX2_972 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813), .Y(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf0) );
  BUFX2 BUFX2_973 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815), .Y(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4) );
  BUFX2 BUFX2_974 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815), .Y(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3) );
  BUFX2 BUFX2_975 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815), .Y(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf2) );
  BUFX2 BUFX2_976 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815), .Y(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf1) );
  BUFX2 BUFX2_977 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815), .Y(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf0) );
  BUFX2 BUFX2_978 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf7) );
  BUFX2 BUFX2_979 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf6) );
  BUFX2 BUFX2_98 ( .A(_abc_43815_n1431_1), .Y(_abc_43815_n1431_1_bF_buf3) );
  BUFX2 BUFX2_980 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf5) );
  BUFX2 BUFX2_981 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf4) );
  BUFX2 BUFX2_982 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf3) );
  BUFX2 BUFX2_983 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf2) );
  BUFX2 BUFX2_984 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf1) );
  BUFX2 BUFX2_985 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf0) );
  BUFX2 BUFX2_986 ( .A(_abc_43815_n3496), .Y(_abc_43815_n3496_bF_buf3) );
  BUFX2 BUFX2_987 ( .A(_abc_43815_n3496), .Y(_abc_43815_n3496_bF_buf2) );
  BUFX2 BUFX2_988 ( .A(_abc_43815_n3496), .Y(_abc_43815_n3496_bF_buf1) );
  BUFX2 BUFX2_989 ( .A(_abc_43815_n3496), .Y(_abc_43815_n3496_bF_buf0) );
  BUFX2 BUFX2_99 ( .A(_abc_43815_n1431_1), .Y(_abc_43815_n1431_1_bF_buf2) );
  BUFX2 BUFX2_990 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3) );
  BUFX2 BUFX2_991 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2) );
  BUFX2 BUFX2_992 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1) );
  BUFX2 BUFX2_993 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0) );
  BUFX2 BUFX2_994 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603), .Y(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf4) );
  BUFX2 BUFX2_995 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603), .Y(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf3) );
  BUFX2 BUFX2_996 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603), .Y(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf2) );
  BUFX2 BUFX2_997 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603), .Y(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf1) );
  BUFX2 BUFX2_998 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7603), .Y(REGFILE_SIM_reg_bank__abc_33898_n7603_bF_buf0) );
  BUFX2 BUFX2_999 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7606), .Y(REGFILE_SIM_reg_bank__abc_33898_n7606_bF_buf4) );
  DFFSR DFFSR_1 ( .CLK(clk_i_bF_buf114), .D(_abc_27555_n4360), .Q(state_q_0_), .R(1'b1), .S(_abc_43815_n4167_bF_buf15_bF_buf3) );
  DFFSR DFFSR_10 ( .CLK(clk_i_bF_buf105), .D(pc_q_1__FF_INPUT), .Q(next_pc_r_1_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_100 ( .CLK(clk_i_bF_buf15), .D(alu_input_a_r_15_), .Q(alu_a_i_15_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_1000 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r24_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_1001 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r24_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_1002 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r24_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_1003 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r24_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_1004 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r24_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_1005 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r24_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_1006 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r24_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_1007 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r24_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_1008 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r24_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_1009 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r24_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_101 ( .CLK(clk_i_bF_buf14), .D(alu_input_a_r_16_), .Q(alu_a_i_16_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_1010 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r24_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_1011 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r24_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_1012 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r24_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_1013 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r24_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_1014 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r24_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_1015 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r24_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_1016 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r24_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_1017 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r24_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_1018 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r24_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_1019 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r24_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_102 ( .CLK(clk_i_bF_buf13), .D(alu_input_a_r_17_), .Q(alu_a_i_17_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_1020 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank_reg_r24_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_1021 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank_reg_r24_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_1022 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank_reg_r24_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_1023 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank_reg_r24_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_1024 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank_reg_r24_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_1025 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank_reg_r24_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_1026 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank_reg_r25_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_1027 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank_reg_r25_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_1028 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank_reg_r25_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_1029 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank_reg_r25_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_103 ( .CLK(clk_i_bF_buf12), .D(alu_input_a_r_18_), .Q(alu_a_i_18_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_1030 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank_reg_r25_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_1031 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank_reg_r25_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_1032 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank_reg_r25_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_1033 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank_reg_r25_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_1034 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank_reg_r25_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_1035 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank_reg_r25_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_1036 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank_reg_r25_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_1037 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank_reg_r25_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_1038 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank_reg_r25_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_1039 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank_reg_r25_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_104 ( .CLK(clk_i_bF_buf11), .D(alu_input_a_r_19_), .Q(alu_a_i_19_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_1040 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank_reg_r25_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_1041 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank_reg_r25_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_1042 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank_reg_r25_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_1043 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank_reg_r25_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_1044 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank_reg_r25_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_1045 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank_reg_r25_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_1046 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank_reg_r25_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_1047 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank_reg_r25_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_1048 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank_reg_r25_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_1049 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank_reg_r25_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_105 ( .CLK(clk_i_bF_buf10), .D(alu_input_a_r_20_), .Q(alu_a_i_20_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_1050 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank_reg_r25_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_1051 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank_reg_r25_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_1052 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank_reg_r25_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_1053 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank_reg_r25_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_1054 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank_reg_r25_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_1055 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank_reg_r25_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_1056 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank_reg_r25_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_1057 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank_reg_r25_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r25_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_1058 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank_reg_r26_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_1059 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank_reg_r26_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_106 ( .CLK(clk_i_bF_buf9), .D(alu_input_a_r_21_), .Q(alu_a_i_21_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_1060 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank_reg_r26_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_1061 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank_reg_r26_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_1062 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank_reg_r26_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_1063 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r26_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_1064 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r26_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_1065 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r26_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_1066 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r26_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_1067 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r26_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_1068 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r26_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_1069 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r26_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_107 ( .CLK(clk_i_bF_buf8), .D(alu_input_a_r_22_), .Q(alu_a_i_22_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_1070 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r26_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_1071 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r26_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_1072 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r26_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_1073 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r26_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_1074 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r26_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_1075 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r26_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_1076 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r26_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_1077 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r26_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_1078 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r26_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_1079 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r26_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_108 ( .CLK(clk_i_bF_buf7), .D(alu_input_a_r_23_), .Q(alu_a_i_23_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_1080 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r26_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_1081 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r26_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_1082 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r26_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_1083 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r26_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_1084 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r26_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_1085 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r26_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_1086 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r26_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_1087 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r26_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_1088 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r26_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_1089 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r26_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r26_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_109 ( .CLK(clk_i_bF_buf6), .D(alu_input_a_r_24_), .Q(alu_a_i_24_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_1090 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r27_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_1091 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r27_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_1092 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r27_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_1093 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r27_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_1094 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r27_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_1095 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r27_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_1096 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r27_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_1097 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r27_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_1098 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r27_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_1099 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r27_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_11 ( .CLK(clk_i_bF_buf104), .D(pc_q_2__FF_INPUT), .Q(pc_q_2_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_110 ( .CLK(clk_i_bF_buf5), .D(alu_input_a_r_25_), .Q(alu_a_i_25_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_1100 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r27_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_1101 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r27_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_1102 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r27_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_1103 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r27_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_1104 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r27_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_1105 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r27_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_1106 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r27_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_1107 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r27_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_1108 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r27_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_1109 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r27_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_111 ( .CLK(clk_i_bF_buf4), .D(alu_input_a_r_26_), .Q(alu_a_i_26_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_1110 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r27_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_1111 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r27_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_1112 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r27_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_1113 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r27_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_1114 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r27_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_1115 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r27_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_1116 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r27_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_1117 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r27_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_1118 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r27_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_1119 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r27_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_112 ( .CLK(clk_i_bF_buf3), .D(alu_input_a_r_27_), .Q(alu_a_i_27_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_1120 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r27_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_1121 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r27_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r27_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_1122 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r28_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_1123 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r28_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_1124 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r28_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_1125 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r28_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_1126 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r28_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_1127 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r28_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_1128 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r28_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_1129 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r28_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_113 ( .CLK(clk_i_bF_buf2), .D(alu_input_a_r_28_), .Q(alu_a_i_28_), .R(_abc_43815_n4167_bF_buf15_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_1130 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r28_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_1131 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r28_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_1132 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r28_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_1133 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r28_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_1134 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r28_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_1135 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank_reg_r28_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_1136 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank_reg_r28_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_1137 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank_reg_r28_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_1138 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank_reg_r28_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_1139 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank_reg_r28_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_114 ( .CLK(clk_i_bF_buf1), .D(alu_input_a_r_29_), .Q(alu_a_i_29_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_1140 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank_reg_r28_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_1141 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank_reg_r28_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_1142 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank_reg_r28_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_1143 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank_reg_r28_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_1144 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank_reg_r28_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_1145 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank_reg_r28_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_1146 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank_reg_r28_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_1147 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank_reg_r28_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_1148 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank_reg_r28_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_1149 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank_reg_r28_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_115 ( .CLK(clk_i_bF_buf0), .D(alu_input_a_r_30_), .Q(alu_a_i_30_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_1150 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank_reg_r28_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_1151 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank_reg_r28_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_1152 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank_reg_r28_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_1153 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank_reg_r28_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r28_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_1154 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank_reg_r29_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_1155 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank_reg_r29_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_1156 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank_reg_r29_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_1157 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank_reg_r29_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_1158 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank_reg_r29_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_1159 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank_reg_r29_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_116 ( .CLK(clk_i_bF_buf114), .D(alu_input_a_r_31_), .Q(alu_a_i_31_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_1160 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank_reg_r29_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_1161 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank_reg_r29_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_1162 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank_reg_r29_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_1163 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank_reg_r29_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_1164 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank_reg_r29_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_1165 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank_reg_r29_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_1166 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank_reg_r29_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_1167 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank_reg_r29_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_1168 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank_reg_r29_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_1169 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank_reg_r29_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_117 ( .CLK(clk_i_bF_buf113), .D(alu_input_b_r_0_), .Q(alu_b_i_0_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_1170 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank_reg_r29_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_1171 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank_reg_r29_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_1172 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank_reg_r29_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_1173 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank_reg_r29_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_1174 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank_reg_r29_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_1175 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank_reg_r29_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_1176 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank_reg_r29_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_1177 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank_reg_r29_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_1178 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r29_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_1179 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r29_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_118 ( .CLK(clk_i_bF_buf112), .D(alu_input_b_r_1_), .Q(alu_b_i_1_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_1180 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r29_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_1181 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r29_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_1182 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r29_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_1183 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r29_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_1184 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r29_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_1185 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r29_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r29_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_1186 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r30_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_1187 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r30_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_1188 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r30_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_1189 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r30_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_119 ( .CLK(clk_i_bF_buf111), .D(alu_input_b_r_2_), .Q(alu_b_i_2_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_1190 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r30_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_1191 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r30_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_1192 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r30_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_1193 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r30_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_1194 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r30_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_1195 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r30_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_1196 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r30_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_1197 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r30_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_1198 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r30_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_1199 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r30_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_12 ( .CLK(clk_i_bF_buf103), .D(pc_q_3__FF_INPUT), .Q(pc_q_3_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_120 ( .CLK(clk_i_bF_buf110), .D(alu_input_b_r_3_), .Q(alu_b_i_3_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_1200 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r30_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_1201 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r30_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_1202 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r30_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_1203 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r30_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_1204 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r30_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_1205 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r30_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_1206 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r30_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_1207 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r30_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_1208 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r30_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_1209 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r30_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_121 ( .CLK(clk_i_bF_buf109), .D(alu_input_b_r_4_), .Q(alu_b_i_4_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_1210 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r30_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_1211 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r30_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_1212 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r30_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_1213 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r30_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_1214 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r30_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_1215 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r30_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_1216 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r30_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_1217 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r30_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r30_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_1218 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r31_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_1219 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r31_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_122 ( .CLK(clk_i_bF_buf108), .D(alu_input_b_r_5_), .Q(alu_b_i_5_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_1220 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r31_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_1221 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r31_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_1222 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r31_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_1223 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r31_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_1224 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r31_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_1225 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r31_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_1226 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r31_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_1227 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r31_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_1228 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r31_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_1229 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r31_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_123 ( .CLK(clk_i_bF_buf107), .D(alu_input_b_r_6_), .Q(alu_b_i_6_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_1230 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r31_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_1231 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r31_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_1232 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r31_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_1233 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r31_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_1234 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r31_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_1235 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r31_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_1236 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r31_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_1237 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r31_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_1238 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r31_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_1239 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r31_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_124 ( .CLK(clk_i_bF_buf106), .D(alu_input_b_r_7_), .Q(alu_b_i_7_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_1240 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r31_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_1241 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r31_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_1242 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r31_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_1243 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r31_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_1244 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r31_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_1245 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r31_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_1246 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r31_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_1247 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r31_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_1248 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r31_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_1249 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r31_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r31_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_125 ( .CLK(clk_i_bF_buf105), .D(alu_input_b_r_8_), .Q(alu_b_i_8_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_126 ( .CLK(clk_i_bF_buf104), .D(alu_input_b_r_9_), .Q(alu_b_i_9_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_127 ( .CLK(clk_i_bF_buf103), .D(alu_input_b_r_10_), .Q(alu_b_i_10_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_128 ( .CLK(clk_i_bF_buf102), .D(alu_input_b_r_11_), .Q(alu_b_i_11_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_129 ( .CLK(clk_i_bF_buf101), .D(alu_input_b_r_12_), .Q(alu_b_i_12_), .R(_abc_43815_n4167_bF_buf15_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_13 ( .CLK(clk_i_bF_buf102), .D(pc_q_4__FF_INPUT), .Q(pc_q_4_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_130 ( .CLK(clk_i_bF_buf100), .D(alu_input_b_r_13_), .Q(alu_b_i_13_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_131 ( .CLK(clk_i_bF_buf99), .D(alu_input_b_r_14_), .Q(alu_b_i_14_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_132 ( .CLK(clk_i_bF_buf98), .D(alu_input_b_r_15_), .Q(alu_b_i_15_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_133 ( .CLK(clk_i_bF_buf97), .D(alu_input_b_r_16_), .Q(alu_b_i_16_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_134 ( .CLK(clk_i_bF_buf96), .D(alu_input_b_r_17_), .Q(alu_b_i_17_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_135 ( .CLK(clk_i_bF_buf95), .D(alu_input_b_r_18_), .Q(alu_b_i_18_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_136 ( .CLK(clk_i_bF_buf94), .D(alu_input_b_r_19_), .Q(alu_b_i_19_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_137 ( .CLK(clk_i_bF_buf93), .D(alu_input_b_r_20_), .Q(alu_b_i_20_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_138 ( .CLK(clk_i_bF_buf92), .D(alu_input_b_r_21_), .Q(alu_b_i_21_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_139 ( .CLK(clk_i_bF_buf91), .D(alu_input_b_r_22_), .Q(alu_b_i_22_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_14 ( .CLK(clk_i_bF_buf101), .D(pc_q_5__FF_INPUT), .Q(pc_q_5_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_140 ( .CLK(clk_i_bF_buf90), .D(alu_input_b_r_23_), .Q(alu_b_i_23_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_141 ( .CLK(clk_i_bF_buf89), .D(alu_input_b_r_24_), .Q(alu_b_i_24_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_142 ( .CLK(clk_i_bF_buf88), .D(alu_input_b_r_25_), .Q(alu_b_i_25_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_143 ( .CLK(clk_i_bF_buf87), .D(alu_input_b_r_26_), .Q(alu_b_i_26_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_144 ( .CLK(clk_i_bF_buf86), .D(alu_input_b_r_27_), .Q(alu_b_i_27_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_145 ( .CLK(clk_i_bF_buf85), .D(alu_input_b_r_28_), .Q(alu_b_i_28_), .R(_abc_43815_n4167_bF_buf15_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_146 ( .CLK(clk_i_bF_buf84), .D(alu_input_b_r_29_), .Q(alu_b_i_29_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_147 ( .CLK(clk_i_bF_buf83), .D(alu_input_b_r_30_), .Q(alu_b_i_30_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_148 ( .CLK(clk_i_bF_buf82), .D(alu_input_b_r_31_), .Q(alu_b_i_31_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_149 ( .CLK(clk_i_bF_buf81), .D(alu_func_r_0_), .Q(alu_op_i_0_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_15 ( .CLK(clk_i_bF_buf100), .D(pc_q_6__FF_INPUT), .Q(pc_q_6_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_150 ( .CLK(clk_i_bF_buf80), .D(alu_func_r_1_), .Q(alu_op_i_1_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_151 ( .CLK(clk_i_bF_buf79), .D(alu_func_r_2_), .Q(alu_op_i_2_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_152 ( .CLK(clk_i_bF_buf78), .D(alu_func_r_3_), .Q(alu_op_i_3_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_153 ( .CLK(clk_i_bF_buf77), .D(mem_addr_o_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_0_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_154 ( .CLK(clk_i_bF_buf76), .D(mem_addr_o_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_1_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_155 ( .CLK(clk_i_bF_buf75), .D(mem_addr_o_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_2_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_156 ( .CLK(clk_i_bF_buf74), .D(mem_addr_o_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_3_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_157 ( .CLK(clk_i_bF_buf73), .D(mem_addr_o_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_4_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_158 ( .CLK(clk_i_bF_buf72), .D(mem_addr_o_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_5_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_159 ( .CLK(clk_i_bF_buf71), .D(mem_addr_o_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_6_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_16 ( .CLK(clk_i_bF_buf99), .D(pc_q_7__FF_INPUT), .Q(pc_q_7_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_160 ( .CLK(clk_i_bF_buf70), .D(mem_addr_o_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_7_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_161 ( .CLK(clk_i_bF_buf69), .D(mem_addr_o_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_8_), .R(_abc_43815_n4167_bF_buf15_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_162 ( .CLK(clk_i_bF_buf68), .D(mem_addr_o_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_9_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_163 ( .CLK(clk_i_bF_buf67), .D(mem_addr_o_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_10_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_164 ( .CLK(clk_i_bF_buf66), .D(mem_addr_o_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_11_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_165 ( .CLK(clk_i_bF_buf65), .D(mem_addr_o_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_12_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_166 ( .CLK(clk_i_bF_buf64), .D(mem_addr_o_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_13_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_167 ( .CLK(clk_i_bF_buf63), .D(mem_addr_o_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_14_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_168 ( .CLK(clk_i_bF_buf62), .D(mem_addr_o_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_15_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_169 ( .CLK(clk_i_bF_buf61), .D(mem_addr_o_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_16_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_17 ( .CLK(clk_i_bF_buf98), .D(pc_q_8__FF_INPUT), .Q(pc_q_8_), .R(1'b1), .S(_abc_43815_n4167_bF_buf15_bF_buf2) );
  DFFSR DFFSR_170 ( .CLK(clk_i_bF_buf60), .D(mem_addr_o_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_17_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_171 ( .CLK(clk_i_bF_buf59), .D(mem_addr_o_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_18_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_172 ( .CLK(clk_i_bF_buf58), .D(mem_addr_o_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_19_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_173 ( .CLK(clk_i_bF_buf57), .D(mem_addr_o_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_20_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_174 ( .CLK(clk_i_bF_buf56), .D(mem_addr_o_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_21_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_175 ( .CLK(clk_i_bF_buf55), .D(mem_addr_o_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_22_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_176 ( .CLK(clk_i_bF_buf54), .D(mem_addr_o_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_23_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_177 ( .CLK(clk_i_bF_buf53), .D(mem_addr_o_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_24_), .R(_abc_43815_n4167_bF_buf15_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_178 ( .CLK(clk_i_bF_buf52), .D(mem_addr_o_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_25_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_179 ( .CLK(clk_i_bF_buf51), .D(mem_addr_o_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_26_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_18 ( .CLK(clk_i_bF_buf97), .D(pc_q_9__FF_INPUT), .Q(pc_q_9_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_180 ( .CLK(clk_i_bF_buf50), .D(mem_addr_o_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_27_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_181 ( .CLK(clk_i_bF_buf49), .D(mem_addr_o_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_28_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_182 ( .CLK(clk_i_bF_buf48), .D(mem_addr_o_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_29_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_183 ( .CLK(clk_i_bF_buf47), .D(mem_addr_o_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_30_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_184 ( .CLK(clk_i_bF_buf46), .D(mem_addr_o_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47730_31_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_185 ( .CLK(clk_i_bF_buf45), .D(mem_dat_o_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_0_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_186 ( .CLK(clk_i_bF_buf44), .D(mem_dat_o_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_1_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_187 ( .CLK(clk_i_bF_buf43), .D(mem_dat_o_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_2_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_188 ( .CLK(clk_i_bF_buf42), .D(mem_dat_o_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_3_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_189 ( .CLK(clk_i_bF_buf41), .D(mem_dat_o_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_4_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_19 ( .CLK(clk_i_bF_buf96), .D(pc_q_10__FF_INPUT), .Q(pc_q_10_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_190 ( .CLK(clk_i_bF_buf40), .D(mem_dat_o_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_5_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_191 ( .CLK(clk_i_bF_buf39), .D(mem_dat_o_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_6_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_192 ( .CLK(clk_i_bF_buf38), .D(mem_dat_o_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_7_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_193 ( .CLK(clk_i_bF_buf37), .D(mem_dat_o_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_8_), .R(_abc_43815_n4167_bF_buf15_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_194 ( .CLK(clk_i_bF_buf36), .D(mem_dat_o_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_9_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_195 ( .CLK(clk_i_bF_buf35), .D(mem_dat_o_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_10_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_196 ( .CLK(clk_i_bF_buf34), .D(mem_dat_o_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_11_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_197 ( .CLK(clk_i_bF_buf33), .D(mem_dat_o_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_12_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_198 ( .CLK(clk_i_bF_buf32), .D(mem_dat_o_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_13_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_199 ( .CLK(clk_i_bF_buf31), .D(mem_dat_o_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_14_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_2 ( .CLK(clk_i_bF_buf113), .D(_abc_27555_n353), .Q(state_q_1_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_20 ( .CLK(clk_i_bF_buf95), .D(pc_q_11__FF_INPUT), .Q(pc_q_11_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_200 ( .CLK(clk_i_bF_buf30), .D(mem_dat_o_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_15_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_201 ( .CLK(clk_i_bF_buf29), .D(mem_dat_o_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_16_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_202 ( .CLK(clk_i_bF_buf28), .D(mem_dat_o_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_17_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_203 ( .CLK(clk_i_bF_buf27), .D(mem_dat_o_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_18_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_204 ( .CLK(clk_i_bF_buf26), .D(mem_dat_o_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_19_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_205 ( .CLK(clk_i_bF_buf25), .D(mem_dat_o_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_20_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_206 ( .CLK(clk_i_bF_buf24), .D(mem_dat_o_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_21_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_207 ( .CLK(clk_i_bF_buf23), .D(mem_dat_o_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_22_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_208 ( .CLK(clk_i_bF_buf22), .D(mem_dat_o_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_23_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_209 ( .CLK(clk_i_bF_buf21), .D(mem_dat_o_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_24_), .R(_abc_43815_n4167_bF_buf15_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_21 ( .CLK(clk_i_bF_buf94), .D(pc_q_12__FF_INPUT), .Q(pc_q_12_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_210 ( .CLK(clk_i_bF_buf20), .D(mem_dat_o_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_25_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_211 ( .CLK(clk_i_bF_buf19), .D(mem_dat_o_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_26_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_212 ( .CLK(clk_i_bF_buf18), .D(mem_dat_o_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_27_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_213 ( .CLK(clk_i_bF_buf17), .D(mem_dat_o_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_28_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_214 ( .CLK(clk_i_bF_buf16), .D(mem_dat_o_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_29_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_215 ( .CLK(clk_i_bF_buf15), .D(mem_dat_o_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_30_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_216 ( .CLK(clk_i_bF_buf14), .D(mem_dat_o_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47769_31_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_217 ( .CLK(clk_i_bF_buf13), .D(mem_cyc_o_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47767), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_218 ( .CLK(clk_i_bF_buf12), .D(mem_stb_o_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47807), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_219 ( .CLK(clk_i_bF_buf11), .D(mem_we_o_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47809), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_22 ( .CLK(clk_i_bF_buf93), .D(pc_q_13__FF_INPUT), .Q(pc_q_13_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_220 ( .CLK(clk_i_bF_buf10), .D(mem_sel_o_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47802_0_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_221 ( .CLK(clk_i_bF_buf9), .D(mem_sel_o_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47802_1_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_222 ( .CLK(clk_i_bF_buf8), .D(mem_sel_o_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47802_2_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_223 ( .CLK(clk_i_bF_buf7), .D(mem_sel_o_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47802_3_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_224 ( .CLK(clk_i_bF_buf6), .D(opcode_q_0__FF_INPUT), .Q(alu_op_r_0_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_225 ( .CLK(clk_i_bF_buf5), .D(opcode_q_1__FF_INPUT), .Q(alu_op_r_1_), .R(_abc_43815_n4167_bF_buf15_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_226 ( .CLK(clk_i_bF_buf4), .D(opcode_q_2__FF_INPUT), .Q(alu_op_r_2_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_227 ( .CLK(clk_i_bF_buf3), .D(opcode_q_3__FF_INPUT), .Q(alu_op_r_3_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_228 ( .CLK(clk_i_bF_buf2), .D(opcode_q_4__FF_INPUT), .Q(int32_r_4_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_229 ( .CLK(clk_i_bF_buf1), .D(opcode_q_5__FF_INPUT), .Q(int32_r_5_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_23 ( .CLK(clk_i_bF_buf92), .D(pc_q_14__FF_INPUT), .Q(pc_q_14_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_230 ( .CLK(clk_i_bF_buf0), .D(opcode_q_6__FF_INPUT), .Q(alu_op_r_4_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_231 ( .CLK(clk_i_bF_buf114), .D(opcode_q_7__FF_INPUT), .Q(alu_op_r_5_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_232 ( .CLK(clk_i_bF_buf113), .D(opcode_q_8__FF_INPUT), .Q(alu_op_r_6_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_233 ( .CLK(clk_i_bF_buf112), .D(opcode_q_9__FF_INPUT), .Q(alu_op_r_7_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_234 ( .CLK(clk_i_bF_buf111), .D(opcode_q_10__FF_INPUT), .Q(int32_r_10_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_235 ( .CLK(clk_i_bF_buf110), .D(opcode_q_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rb_i_0_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_236 ( .CLK(clk_i_bF_buf109), .D(opcode_q_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rb_i_1_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_237 ( .CLK(clk_i_bF_buf108), .D(opcode_q_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rb_i_2_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_238 ( .CLK(clk_i_bF_buf107), .D(opcode_q_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rb_i_3_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_239 ( .CLK(clk_i_bF_buf106), .D(opcode_q_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rb_i_4_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_24 ( .CLK(clk_i_bF_buf91), .D(pc_q_15__FF_INPUT), .Q(pc_q_15_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_240 ( .CLK(clk_i_bF_buf105), .D(opcode_q_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_ra_i_0_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_241 ( .CLK(clk_i_bF_buf104), .D(opcode_q_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_ra_i_1_), .R(_abc_43815_n4167_bF_buf15_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_242 ( .CLK(clk_i_bF_buf103), .D(opcode_q_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_ra_i_2_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_243 ( .CLK(clk_i_bF_buf102), .D(opcode_q_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_ra_i_3_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_244 ( .CLK(clk_i_bF_buf101), .D(opcode_q_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_ra_i_4_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_245 ( .CLK(clk_i_bF_buf100), .D(opcode_q_21__FF_INPUT), .Q(opcode_q_21_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_246 ( .CLK(clk_i_bF_buf99), .D(opcode_q_22__FF_INPUT), .Q(opcode_q_22_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_247 ( .CLK(clk_i_bF_buf98), .D(opcode_q_23__FF_INPUT), .Q(opcode_q_23_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_248 ( .CLK(clk_i_bF_buf97), .D(opcode_q_24__FF_INPUT), .Q(opcode_q_24_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_249 ( .CLK(clk_i_bF_buf96), .D(opcode_q_25__FF_INPUT), .Q(opcode_q_25_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_25 ( .CLK(clk_i_bF_buf90), .D(pc_q_16__FF_INPUT), .Q(pc_q_16_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_250 ( .CLK(clk_i_bF_buf95), .D(opcode_q_26__FF_INPUT), .Q(inst_r_0_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_251 ( .CLK(clk_i_bF_buf94), .D(opcode_q_27__FF_INPUT), .Q(inst_r_1_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_252 ( .CLK(clk_i_bF_buf93), .D(opcode_q_28__FF_INPUT), .Q(inst_r_2_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_253 ( .CLK(clk_i_bF_buf92), .D(opcode_q_29__FF_INPUT), .Q(inst_r_3_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_254 ( .CLK(clk_i_bF_buf91), .D(opcode_q_30__FF_INPUT), .Q(inst_r_4_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_255 ( .CLK(clk_i_bF_buf90), .D(opcode_q_31__FF_INPUT), .Q(inst_r_5_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_256 ( .CLK(clk_i_bF_buf89), .D(mem_offset_q_0__FF_INPUT), .Q(mem_offset_q_0_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_257 ( .CLK(clk_i_bF_buf88), .D(mem_offset_q_1__FF_INPUT), .Q(mem_offset_q_1_), .R(_abc_43815_n4167_bF_buf15_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_258 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r1_sp_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_259 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r1_sp_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_26 ( .CLK(clk_i_bF_buf89), .D(pc_q_17__FF_INPUT), .Q(pc_q_17_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_260 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r1_sp_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_261 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r1_sp_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_262 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r1_sp_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_263 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r1_sp_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_264 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r1_sp_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_265 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r1_sp_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_266 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r1_sp_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_267 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r1_sp_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_268 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r1_sp_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_269 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r1_sp_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_27 ( .CLK(clk_i_bF_buf88), .D(pc_q_18__FF_INPUT), .Q(pc_q_18_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_270 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r1_sp_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_271 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r1_sp_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_272 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r1_sp_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_273 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r1_sp_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_274 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r1_sp_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_275 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r1_sp_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_276 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r1_sp_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_277 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r1_sp_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_278 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r1_sp_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_279 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r1_sp_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_28 ( .CLK(clk_i_bF_buf87), .D(pc_q_19__FF_INPUT), .Q(pc_q_19_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_280 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r1_sp_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_281 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r1_sp_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_282 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r1_sp_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_283 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r1_sp_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_284 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r1_sp_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_285 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r1_sp_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_286 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r1_sp_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_287 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r1_sp_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_288 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r1_sp_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_289 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r1_sp_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_29 ( .CLK(clk_i_bF_buf86), .D(pc_q_20__FF_INPUT), .Q(pc_q_20_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_290 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r2_fp_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_291 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r2_fp_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_292 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r2_fp_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_293 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r2_fp_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_294 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r2_fp_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_295 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r2_fp_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_296 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r2_fp_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_297 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r2_fp_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_298 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r2_fp_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_299 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r2_fp_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_3 ( .CLK(clk_i_bF_buf112), .D(_abc_27555_n343), .Q(state_q_2_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_30 ( .CLK(clk_i_bF_buf85), .D(pc_q_21__FF_INPUT), .Q(pc_q_21_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_300 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r2_fp_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_301 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r2_fp_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_302 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r2_fp_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_303 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r2_fp_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_304 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r2_fp_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_305 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r2_fp_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_306 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r2_fp_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_307 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r2_fp_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_308 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r2_fp_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_309 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r2_fp_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_31 ( .CLK(clk_i_bF_buf84), .D(pc_q_22__FF_INPUT), .Q(pc_q_22_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_310 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r2_fp_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_311 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r2_fp_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_312 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r2_fp_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_313 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r2_fp_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_314 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r2_fp_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_315 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r2_fp_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_316 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r2_fp_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_317 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r2_fp_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_318 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r2_fp_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_319 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r2_fp_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_32 ( .CLK(clk_i_bF_buf83), .D(pc_q_23__FF_INPUT), .Q(pc_q_23_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_320 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r2_fp_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_321 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r2_fp_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_322 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r3_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_323 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r3_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_324 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r3_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_325 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r3_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_326 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r3_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_327 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r3_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_328 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r3_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_329 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r3_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_33 ( .CLK(clk_i_bF_buf82), .D(pc_q_24__FF_INPUT), .Q(pc_q_24_), .R(_abc_43815_n4167_bF_buf15_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_330 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank_reg_r3_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_331 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank_reg_r3_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_332 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank_reg_r3_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_333 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank_reg_r3_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_334 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank_reg_r3_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_335 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank_reg_r3_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_336 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank_reg_r3_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_337 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank_reg_r3_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_338 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank_reg_r3_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_339 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank_reg_r3_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_34 ( .CLK(clk_i_bF_buf81), .D(pc_q_25__FF_INPUT), .Q(pc_q_25_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_340 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank_reg_r3_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_341 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank_reg_r3_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_342 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank_reg_r3_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_343 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank_reg_r3_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_344 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank_reg_r3_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_345 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank_reg_r3_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_346 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank_reg_r3_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_347 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank_reg_r3_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_348 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank_reg_r3_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_349 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank_reg_r3_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_35 ( .CLK(clk_i_bF_buf80), .D(pc_q_26__FF_INPUT), .Q(pc_q_26_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_350 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank_reg_r3_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_351 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank_reg_r3_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_352 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank_reg_r3_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_353 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank_reg_r3_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r3_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_354 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank_reg_r4_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_355 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank_reg_r4_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_356 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank_reg_r4_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_357 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank_reg_r4_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_358 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank_reg_r4_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_359 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank_reg_r4_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_36 ( .CLK(clk_i_bF_buf79), .D(pc_q_27__FF_INPUT), .Q(pc_q_27_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_360 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank_reg_r4_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_361 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank_reg_r4_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_362 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank_reg_r4_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_363 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank_reg_r4_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_364 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank_reg_r4_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_365 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank_reg_r4_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_366 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank_reg_r4_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_367 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank_reg_r4_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_368 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank_reg_r4_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_369 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank_reg_r4_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_37 ( .CLK(clk_i_bF_buf78), .D(pc_q_28__FF_INPUT), .Q(pc_q_28_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_370 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank_reg_r4_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_371 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank_reg_r4_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_372 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank_reg_r4_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_373 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r4_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_374 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r4_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_375 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r4_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_376 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r4_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_377 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r4_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_378 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r4_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_379 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r4_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_38 ( .CLK(clk_i_bF_buf77), .D(pc_q_29__FF_INPUT), .Q(pc_q_29_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_380 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r4_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_381 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r4_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_382 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r4_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_383 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r4_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_384 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r4_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_385 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r4_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r4_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_386 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r5_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_387 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r5_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_388 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r5_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_389 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r5_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_39 ( .CLK(clk_i_bF_buf76), .D(pc_q_30__FF_INPUT), .Q(pc_q_30_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_390 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r5_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_391 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r5_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_392 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r5_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_393 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r5_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_394 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r5_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_395 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r5_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_396 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r5_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_397 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r5_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_398 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r5_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_399 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r5_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_4 ( .CLK(clk_i_bF_buf111), .D(_abc_27555_n185), .Q(state_q_3_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_40 ( .CLK(clk_i_bF_buf75), .D(pc_q_31__FF_INPUT), .Q(pc_q_31_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_400 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r5_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_401 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r5_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_402 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r5_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_403 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r5_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_404 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r5_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_405 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r5_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_406 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r5_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_407 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r5_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_408 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r5_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_409 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r5_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_41 ( .CLK(clk_i_bF_buf74), .D(epc_q_0__FF_INPUT), .Q(epc_q_0_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_410 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r5_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_411 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r5_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_412 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r5_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_413 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r5_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_414 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r5_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_415 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r5_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_416 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r5_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_417 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r5_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r5_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_418 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r6_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_419 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r6_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_42 ( .CLK(clk_i_bF_buf73), .D(epc_q_1__FF_INPUT), .Q(epc_q_1_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_420 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r6_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_421 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r6_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_422 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r6_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_423 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r6_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_424 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r6_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_425 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r6_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_426 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r6_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_427 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r6_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_428 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r6_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_429 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r6_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_43 ( .CLK(clk_i_bF_buf72), .D(epc_q_2__FF_INPUT), .Q(epc_q_2_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_430 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r6_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_431 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r6_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_432 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r6_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_433 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r6_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_434 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r6_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_435 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r6_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_436 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r6_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_437 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r6_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_438 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r6_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_439 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r6_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_44 ( .CLK(clk_i_bF_buf71), .D(epc_q_3__FF_INPUT), .Q(epc_q_3_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_440 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r6_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_441 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r6_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_442 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r6_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_443 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r6_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_444 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r6_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_445 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank_reg_r6_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_446 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank_reg_r6_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_447 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank_reg_r6_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_448 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank_reg_r6_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_449 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank_reg_r6_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r6_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_45 ( .CLK(clk_i_bF_buf70), .D(epc_q_4__FF_INPUT), .Q(epc_q_4_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_450 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank_reg_r7_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_451 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank_reg_r7_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_452 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank_reg_r7_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_453 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank_reg_r7_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_454 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank_reg_r7_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_455 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank_reg_r7_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_456 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank_reg_r7_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_457 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank_reg_r7_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_458 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank_reg_r7_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_459 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank_reg_r7_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_46 ( .CLK(clk_i_bF_buf69), .D(epc_q_5__FF_INPUT), .Q(epc_q_5_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_460 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank_reg_r7_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_461 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank_reg_r7_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_462 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank_reg_r7_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_463 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank_reg_r7_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_464 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank_reg_r7_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_465 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank_reg_r7_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_466 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank_reg_r7_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_467 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank_reg_r7_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_468 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank_reg_r7_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_469 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank_reg_r7_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_47 ( .CLK(clk_i_bF_buf68), .D(epc_q_6__FF_INPUT), .Q(epc_q_6_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_470 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank_reg_r7_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_471 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank_reg_r7_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_472 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank_reg_r7_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_473 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank_reg_r7_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_474 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank_reg_r7_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_475 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank_reg_r7_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_476 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank_reg_r7_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_477 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank_reg_r7_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_478 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank_reg_r7_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_479 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank_reg_r7_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_48 ( .CLK(clk_i_bF_buf67), .D(epc_q_7__FF_INPUT), .Q(epc_q_7_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_480 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank_reg_r7_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_481 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank_reg_r7_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r7_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_482 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank_reg_r8_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_483 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank_reg_r8_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_484 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank_reg_r8_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_485 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank_reg_r8_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_486 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank_reg_r8_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_487 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank_reg_r8_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_488 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r8_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_489 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r8_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_49 ( .CLK(clk_i_bF_buf66), .D(epc_q_8__FF_INPUT), .Q(epc_q_8_), .R(_abc_43815_n4167_bF_buf15_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_490 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r8_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_491 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r8_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_492 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r8_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_493 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r8_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_494 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r8_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_495 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r8_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_496 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r8_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_497 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r8_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_498 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r8_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_499 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r8_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_5 ( .CLK(clk_i_bF_buf110), .D(_abc_27555_n288), .Q(state_q_4_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_50 ( .CLK(clk_i_bF_buf65), .D(epc_q_9__FF_INPUT), .Q(epc_q_9_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_500 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r8_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_501 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r8_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_502 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r8_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_503 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r8_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_504 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r8_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_505 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r8_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_506 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r8_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_507 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r8_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_508 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r8_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_509 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r8_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_51 ( .CLK(clk_i_bF_buf64), .D(epc_q_10__FF_INPUT), .Q(epc_q_10_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_510 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r8_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_511 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r8_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_512 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r8_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_513 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r8_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r8_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_514 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r9_lr_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_515 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r9_lr_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_516 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r9_lr_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_517 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r9_lr_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_518 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r9_lr_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_519 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r9_lr_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_52 ( .CLK(clk_i_bF_buf63), .D(epc_q_11__FF_INPUT), .Q(epc_q_11_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_520 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r9_lr_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_521 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r9_lr_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_522 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r9_lr_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_523 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r9_lr_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_524 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r9_lr_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_525 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r9_lr_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_526 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r9_lr_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_527 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r9_lr_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_528 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r9_lr_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_529 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r9_lr_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_53 ( .CLK(clk_i_bF_buf62), .D(epc_q_12__FF_INPUT), .Q(epc_q_12_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_530 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r9_lr_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_531 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r9_lr_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_532 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r9_lr_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_533 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r9_lr_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_534 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r9_lr_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_535 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r9_lr_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_536 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r9_lr_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_537 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r9_lr_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_538 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r9_lr_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_539 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r9_lr_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_54 ( .CLK(clk_i_bF_buf61), .D(epc_q_13__FF_INPUT), .Q(epc_q_13_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_540 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r9_lr_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_541 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r9_lr_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_542 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r9_lr_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_543 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r9_lr_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_544 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r9_lr_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_545 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r9_lr_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_546 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r10_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_547 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r10_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_548 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r10_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_549 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r10_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_55 ( .CLK(clk_i_bF_buf60), .D(epc_q_14__FF_INPUT), .Q(epc_q_14_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_550 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r10_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_551 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r10_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_552 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r10_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_553 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r10_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_554 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r10_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_555 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r10_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_556 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r10_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_557 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r10_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_558 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r10_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_559 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r10_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_56 ( .CLK(clk_i_bF_buf59), .D(epc_q_15__FF_INPUT), .Q(epc_q_15_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_560 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank_reg_r10_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_561 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank_reg_r10_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_562 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank_reg_r10_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_563 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank_reg_r10_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_564 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank_reg_r10_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_565 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank_reg_r10_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_566 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank_reg_r10_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_567 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank_reg_r10_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_568 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank_reg_r10_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_569 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank_reg_r10_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_57 ( .CLK(clk_i_bF_buf58), .D(epc_q_16__FF_INPUT), .Q(epc_q_16_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_570 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank_reg_r10_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_571 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank_reg_r10_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_572 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank_reg_r10_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_573 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank_reg_r10_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_574 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank_reg_r10_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_575 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank_reg_r10_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_576 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank_reg_r10_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_577 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank_reg_r10_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r10_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_578 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank_reg_r11_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_579 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank_reg_r11_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_58 ( .CLK(clk_i_bF_buf57), .D(epc_q_17__FF_INPUT), .Q(epc_q_17_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_580 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank_reg_r11_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_581 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank_reg_r11_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_582 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank_reg_r11_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_583 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank_reg_r11_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_584 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank_reg_r11_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_585 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank_reg_r11_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_586 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank_reg_r11_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_587 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank_reg_r11_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_588 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank_reg_r11_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_589 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank_reg_r11_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_59 ( .CLK(clk_i_bF_buf56), .D(epc_q_18__FF_INPUT), .Q(epc_q_18_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_590 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank_reg_r11_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_591 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank_reg_r11_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_592 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank_reg_r11_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_593 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank_reg_r11_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_594 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank_reg_r11_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_595 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank_reg_r11_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_596 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank_reg_r11_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_597 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank_reg_r11_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_598 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank_reg_r11_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_599 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank_reg_r11_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_6 ( .CLK(clk_i_bF_buf109), .D(_abc_27555_n4367_bF_buf7), .Q(state_q_5_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_60 ( .CLK(clk_i_bF_buf55), .D(epc_q_19__FF_INPUT), .Q(epc_q_19_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_600 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank_reg_r11_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_601 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank_reg_r11_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_602 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank_reg_r11_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_603 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r11_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_604 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r11_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_605 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r11_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_606 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r11_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_607 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r11_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_608 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r11_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_609 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r11_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r11_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_61 ( .CLK(clk_i_bF_buf54), .D(epc_q_20__FF_INPUT), .Q(epc_q_20_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_610 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r12_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_611 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r12_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_612 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r12_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_613 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r12_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_614 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r12_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_615 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r12_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_616 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r12_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_617 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r12_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_618 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r12_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_619 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r12_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_62 ( .CLK(clk_i_bF_buf53), .D(epc_q_21__FF_INPUT), .Q(epc_q_21_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_620 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r12_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_621 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r12_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_622 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r12_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_623 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r12_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_624 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r12_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_625 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r12_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_626 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r12_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_627 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r12_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_628 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r12_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_629 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r12_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_63 ( .CLK(clk_i_bF_buf52), .D(epc_q_22__FF_INPUT), .Q(epc_q_22_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_630 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r12_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_631 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r12_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_632 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r12_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_633 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r12_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_634 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r12_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_635 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r12_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_636 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r12_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_637 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r12_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_638 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r12_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_639 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r12_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_64 ( .CLK(clk_i_bF_buf51), .D(epc_q_23__FF_INPUT), .Q(epc_q_23_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_640 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r12_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_641 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r12_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r12_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_642 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r13_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_643 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r13_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_644 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r13_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_645 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r13_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_646 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r13_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_647 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r13_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_648 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r13_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_649 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r13_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_65 ( .CLK(clk_i_bF_buf50), .D(epc_q_24__FF_INPUT), .Q(epc_q_24_), .R(_abc_43815_n4167_bF_buf15_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_650 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r13_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_651 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r13_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_652 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r13_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_653 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r13_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_654 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r13_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_655 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r13_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_656 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r13_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_657 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r13_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_658 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r13_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_659 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r13_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_66 ( .CLK(clk_i_bF_buf49), .D(epc_q_25__FF_INPUT), .Q(epc_q_25_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_660 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r13_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_661 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r13_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_662 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r13_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_663 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r13_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_664 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r13_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_665 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r13_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_666 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r13_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_667 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r13_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_668 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r13_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_669 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r13_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_67 ( .CLK(clk_i_bF_buf48), .D(epc_q_26__FF_INPUT), .Q(epc_q_26_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_670 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r13_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_671 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r13_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_672 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r13_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_673 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r13_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r13_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_674 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r14_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_675 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank_reg_r14_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_676 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank_reg_r14_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_677 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank_reg_r14_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_678 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank_reg_r14_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_679 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank_reg_r14_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_68 ( .CLK(clk_i_bF_buf47), .D(epc_q_27__FF_INPUT), .Q(epc_q_27_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_680 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank_reg_r14_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_681 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank_reg_r14_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_682 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank_reg_r14_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_683 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank_reg_r14_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_684 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank_reg_r14_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_685 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank_reg_r14_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_686 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank_reg_r14_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_687 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank_reg_r14_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_688 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank_reg_r14_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_689 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank_reg_r14_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_69 ( .CLK(clk_i_bF_buf46), .D(epc_q_28__FF_INPUT), .Q(epc_q_28_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_690 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank_reg_r14_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_691 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank_reg_r14_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_692 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank_reg_r14_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_693 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank_reg_r14_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_694 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank_reg_r14_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_695 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank_reg_r14_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_696 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank_reg_r14_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_697 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank_reg_r14_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_698 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank_reg_r14_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_699 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank_reg_r14_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_7 ( .CLK(clk_i_bF_buf108), .D(inst_trap_w), .Q(_auto_iopadmap_cc_313_execute_47726), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_70 ( .CLK(clk_i_bF_buf45), .D(epc_q_29__FF_INPUT), .Q(epc_q_29_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_700 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank_reg_r14_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_701 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank_reg_r14_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_702 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank_reg_r14_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_703 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank_reg_r14_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_704 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank_reg_r14_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_705 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank_reg_r14_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r14_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_706 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank_reg_r15_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_707 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank_reg_r15_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_708 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank_reg_r15_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_709 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank_reg_r15_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_71 ( .CLK(clk_i_bF_buf44), .D(epc_q_30__FF_INPUT), .Q(epc_q_30_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_710 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank_reg_r15_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_711 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank_reg_r15_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_712 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank_reg_r15_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_713 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank_reg_r15_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_714 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank_reg_r15_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_715 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank_reg_r15_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_716 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank_reg_r15_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_717 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank_reg_r15_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_718 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r15_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_719 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r15_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_72 ( .CLK(clk_i_bF_buf43), .D(epc_q_31__FF_INPUT), .Q(epc_q_31_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_720 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r15_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_721 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r15_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_722 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r15_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_723 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r15_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_724 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r15_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_725 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r15_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_726 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r15_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_727 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r15_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_728 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r15_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_729 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r15_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_73 ( .CLK(clk_i_bF_buf42), .D(sr_q_2__FF_INPUT), .Q(sr_q_2_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_730 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r15_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_731 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r15_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_732 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r15_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_733 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r15_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_734 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r15_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_735 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r15_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_736 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r15_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_737 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r15_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r15_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_738 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r16_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_739 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r16_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_74 ( .CLK(clk_i_bF_buf41), .D(sr_q_9__FF_INPUT), .Q(sr_q_9_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_740 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r16_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_741 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r16_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_742 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r16_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_743 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r16_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_744 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r16_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_745 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r16_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_746 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r16_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_747 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r16_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_748 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r16_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_749 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r16_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_75 ( .CLK(clk_i_bF_buf40), .D(sr_q_10__FF_INPUT), .Q(alu_c_i), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_750 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r16_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_751 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r16_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_752 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r16_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_753 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r16_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_754 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r16_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_755 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r16_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_756 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r16_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_757 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r16_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_758 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r16_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_759 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r16_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_76 ( .CLK(clk_i_bF_buf39), .D(esr_q_2__FF_INPUT), .Q(esr_q_2_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_760 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r16_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_761 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r16_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_762 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r16_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_763 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r16_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_764 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r16_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_765 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r16_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_766 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r16_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_767 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r16_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_768 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r16_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_769 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r16_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r16_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_77 ( .CLK(clk_i_bF_buf38), .D(esr_q_9__FF_INPUT), .Q(esr_q_9_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_770 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r17_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_771 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r17_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_772 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r17_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_773 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r17_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_774 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r17_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_775 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r17_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_776 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r17_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_777 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r17_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_778 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r17_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_779 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r17_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_78 ( .CLK(clk_i_bF_buf37), .D(esr_q_10__FF_INPUT), .Q(esr_q_10_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_780 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r17_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_781 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r17_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_782 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r17_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_783 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r17_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_784 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r17_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_785 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r17_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_786 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r17_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_787 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r17_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_788 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r17_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_789 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r17_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_79 ( .CLK(clk_i_bF_buf36), .D(nmi_q_FF_INPUT), .Q(nmi_q), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_790 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank_reg_r17_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_791 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank_reg_r17_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_792 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank_reg_r17_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_793 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank_reg_r17_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_794 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank_reg_r17_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_795 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank_reg_r17_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_796 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank_reg_r17_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_797 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank_reg_r17_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_798 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank_reg_r17_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_799 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank_reg_r17_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_8 ( .CLK(clk_i_bF_buf107), .D(fault_o_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_47728), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_80 ( .CLK(clk_i_bF_buf35), .D(ex_rd_q_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rd_i_0_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_800 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank_reg_r17_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_801 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank_reg_r17_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r17_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_802 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank_reg_r18_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_803 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank_reg_r18_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_804 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank_reg_r18_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_805 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank_reg_r18_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_806 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank_reg_r18_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_807 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank_reg_r18_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_808 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank_reg_r18_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_809 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank_reg_r18_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_81 ( .CLK(clk_i_bF_buf34), .D(ex_rd_q_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rd_i_1_), .R(_abc_43815_n4167_bF_buf15_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_810 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank_reg_r18_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_811 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank_reg_r18_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_812 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank_reg_r18_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_813 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank_reg_r18_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_814 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank_reg_r18_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_815 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank_reg_r18_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_816 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank_reg_r18_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_817 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank_reg_r18_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_818 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank_reg_r18_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_819 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank_reg_r18_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_82 ( .CLK(clk_i_bF_buf33), .D(ex_rd_q_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rd_i_2_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_820 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank_reg_r18_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_821 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank_reg_r18_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_822 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank_reg_r18_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_823 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank_reg_r18_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_824 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank_reg_r18_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_825 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank_reg_r18_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_826 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank_reg_r18_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_827 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank_reg_r18_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_828 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank_reg_r18_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_829 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank_reg_r18_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_83 ( .CLK(clk_i_bF_buf32), .D(ex_rd_q_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rd_i_3_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_830 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank_reg_r18_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_831 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank_reg_r18_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_832 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank_reg_r18_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_833 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r18_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r18_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_834 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r19_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_835 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r19_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_836 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r19_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_837 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r19_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_838 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r19_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_839 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r19_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_84 ( .CLK(clk_i_bF_buf31), .D(ex_rd_q_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_rd_i_4_), .R(_abc_43815_n4167_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_840 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r19_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_841 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r19_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_842 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r19_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_843 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r19_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_844 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r19_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_845 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r19_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_846 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r19_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_847 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r19_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_848 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r19_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_849 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r19_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_85 ( .CLK(clk_i_bF_buf30), .D(alu_input_a_r_0_), .Q(alu_a_i_0_), .R(_abc_43815_n4167_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_850 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r19_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_851 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r19_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_852 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r19_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_853 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r19_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_854 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r19_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_855 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r19_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_856 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r19_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_857 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r19_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_858 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r19_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_859 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r19_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_86 ( .CLK(clk_i_bF_buf29), .D(alu_input_a_r_1_), .Q(alu_a_i_1_), .R(_abc_43815_n4167_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_860 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r19_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_861 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r19_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_862 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r19_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_863 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r19_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_864 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r19_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_865 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r19_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r19_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_866 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r20_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_867 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r20_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_868 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r20_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_869 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r20_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_87 ( .CLK(clk_i_bF_buf28), .D(alu_input_a_r_2_), .Q(alu_a_i_2_), .R(_abc_43815_n4167_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_870 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r20_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_871 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r20_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_872 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r20_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_873 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r20_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_874 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r20_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_875 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r20_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_876 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r20_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_877 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r20_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_878 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r20_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_879 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r20_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_88 ( .CLK(clk_i_bF_buf27), .D(alu_input_a_r_3_), .Q(alu_a_i_3_), .R(_abc_43815_n4167_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_880 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r20_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_881 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r20_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_882 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r20_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_883 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r20_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_884 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r20_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_885 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank_reg_r20_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_886 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank_reg_r20_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_887 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank_reg_r20_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_888 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank_reg_r20_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_889 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank_reg_r20_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_89 ( .CLK(clk_i_bF_buf26), .D(alu_input_a_r_4_), .Q(alu_a_i_4_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_890 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank_reg_r20_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_891 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank_reg_r20_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_892 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank_reg_r20_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_893 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank_reg_r20_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_894 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank_reg_r20_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_895 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank_reg_r20_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_896 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank_reg_r20_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_897 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank_reg_r20_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r20_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_898 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank_reg_r21_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_899 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank_reg_r21_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_9 ( .CLK(clk_i_bF_buf106), .D(pc_q_0__FF_INPUT), .Q(next_pc_r_0_), .R(_abc_43815_n4167_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_90 ( .CLK(clk_i_bF_buf25), .D(alu_input_a_r_5_), .Q(alu_a_i_5_), .R(_abc_43815_n4167_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_900 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank_reg_r21_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_901 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank_reg_r21_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_902 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank_reg_r21_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_903 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank_reg_r21_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_904 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank_reg_r21_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_905 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank_reg_r21_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_906 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank_reg_r21_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_907 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank_reg_r21_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_908 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank_reg_r21_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_909 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank_reg_r21_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_91 ( .CLK(clk_i_bF_buf24), .D(alu_input_a_r_6_), .Q(alu_a_i_6_), .R(_abc_43815_n4167_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_910 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank_reg_r21_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_911 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank_reg_r21_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_912 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank_reg_r21_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_913 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank_reg_r21_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_914 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank_reg_r21_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_915 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank_reg_r21_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_916 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank_reg_r21_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_917 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank_reg_r21_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_918 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank_reg_r21_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_919 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank_reg_r21_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_92 ( .CLK(clk_i_bF_buf23), .D(alu_input_a_r_7_), .Q(alu_a_i_7_), .R(_abc_43815_n4167_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_920 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank_reg_r21_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_921 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank_reg_r21_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_922 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank_reg_r21_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_923 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank_reg_r21_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_924 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank_reg_r21_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_925 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank_reg_r21_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_926 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank_reg_r21_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_927 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank_reg_r21_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_928 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank_reg_r21_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_929 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank_reg_r21_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r21_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_93 ( .CLK(clk_i_bF_buf22), .D(alu_input_a_r_8_), .Q(alu_a_i_8_), .R(_abc_43815_n4167_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_930 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank_reg_r22_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_931 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank_reg_r22_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_932 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank_reg_r22_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_933 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank_reg_r22_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_934 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank_reg_r22_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_935 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank_reg_r22_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_936 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank_reg_r22_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_937 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank_reg_r22_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_938 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank_reg_r22_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_939 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank_reg_r22_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_94 ( .CLK(clk_i_bF_buf21), .D(alu_input_a_r_9_), .Q(alu_a_i_9_), .R(_abc_43815_n4167_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_940 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank_reg_r22_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_941 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank_reg_r22_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_942 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank_reg_r22_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_943 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank_reg_r22_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_944 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank_reg_r22_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_945 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank_reg_r22_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_946 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank_reg_r22_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_947 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank_reg_r22_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_948 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank_reg_r22_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_949 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank_reg_r22_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_95 ( .CLK(clk_i_bF_buf20), .D(alu_input_a_r_10_), .Q(alu_a_i_10_), .R(_abc_43815_n4167_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_950 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank_reg_r22_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_951 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank_reg_r22_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf98), .S(1'b1) );
  DFFSR DFFSR_952 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank_reg_r22_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf97), .S(1'b1) );
  DFFSR DFFSR_953 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank_reg_r22_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf96), .S(1'b1) );
  DFFSR DFFSR_954 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank_reg_r22_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf95), .S(1'b1) );
  DFFSR DFFSR_955 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank_reg_r22_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf94), .S(1'b1) );
  DFFSR DFFSR_956 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank_reg_r22_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf93), .S(1'b1) );
  DFFSR DFFSR_957 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank_reg_r22_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf92), .S(1'b1) );
  DFFSR DFFSR_958 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank_reg_r22_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf91), .S(1'b1) );
  DFFSR DFFSR_959 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank_reg_r22_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf90), .S(1'b1) );
  DFFSR DFFSR_96 ( .CLK(clk_i_bF_buf19), .D(alu_input_a_r_11_), .Q(alu_a_i_11_), .R(_abc_43815_n4167_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_960 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank_reg_r22_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf89), .S(1'b1) );
  DFFSR DFFSR_961 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank_reg_r22_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r22_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_962 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank_reg_r23_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_963 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank_reg_r23_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_964 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank_reg_r23_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_965 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank_reg_r23_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_966 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank_reg_r23_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_967 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank_reg_r23_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_968 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank_reg_r23_6__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_6_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_969 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank_reg_r23_7__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_7_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_97 ( .CLK(clk_i_bF_buf18), .D(alu_input_a_r_12_), .Q(alu_a_i_12_), .R(_abc_43815_n4167_bF_buf15_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_970 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank_reg_r23_8__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_8_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_971 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank_reg_r23_9__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_9_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_972 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank_reg_r23_10__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_10_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_973 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank_reg_r23_11__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_11_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_974 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank_reg_r23_12__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_12_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_975 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank_reg_r23_13__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_13_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_976 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank_reg_r23_14__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_14_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_977 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank_reg_r23_15__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_15_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_978 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank_reg_r23_16__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_16_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_979 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank_reg_r23_17__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_17_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_98 ( .CLK(clk_i_bF_buf17), .D(alu_input_a_r_13_), .Q(alu_a_i_13_), .R(_abc_43815_n4167_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_980 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank_reg_r23_18__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_18_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_981 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank_reg_r23_19__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_19_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_982 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank_reg_r23_20__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_20_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_983 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank_reg_r23_21__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_21_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_984 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank_reg_r23_22__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_22_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_985 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank_reg_r23_23__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_23_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_986 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank_reg_r23_24__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_24_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_987 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank_reg_r23_25__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_25_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_988 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank_reg_r23_26__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_26_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_989 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank_reg_r23_27__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_27_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_99 ( .CLK(clk_i_bF_buf16), .D(alu_input_a_r_14_), .Q(alu_a_i_14_), .R(_abc_43815_n4167_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_990 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank_reg_r23_28__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_28_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_991 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank_reg_r23_29__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_29_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_992 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank_reg_r23_30__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_30_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_993 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank_reg_r23_31__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r23_31_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_994 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank_reg_r24_0__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_0_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_995 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank_reg_r24_1__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_1_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_996 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank_reg_r24_2__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_2_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_997 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank_reg_r24_3__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_3_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_998 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank_reg_r24_4__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_4_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_999 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank_reg_r24_5__FF_INPUT), .Q(REGFILE_SIM_reg_bank_reg_r24_5_), .R(REGFILE_SIM_reg_bank__abc_33898_n5245_bF_buf50), .S(1'b1) );
  INVX1 INVX1_1 ( .A(opcode_q_25_), .Y(_abc_43815_n621) );
  INVX1 INVX1_10 ( .A(_abc_43815_n653), .Y(_abc_43815_n664_1) );
  INVX1 INVX1_100 ( .A(_abc_43815_n1382), .Y(_abc_43815_n1383) );
  INVX1 INVX1_1000 ( .A(alu__abc_41358_n426), .Y(alu__abc_41358_n1347) );
  INVX1 INVX1_1001 ( .A(alu__abc_41358_n764), .Y(alu__abc_41358_n1350) );
  INVX1 INVX1_1002 ( .A(alu__abc_41358_n1387), .Y(alu__abc_41358_n1388) );
  INVX1 INVX1_1003 ( .A(alu__abc_41358_n407), .Y(alu__abc_41358_n1399) );
  INVX1 INVX1_1004 ( .A(alu__abc_41358_n765), .Y(alu__abc_41358_n1404) );
  INVX1 INVX1_1005 ( .A(alu__abc_41358_n1441), .Y(alu__abc_41358_n1442) );
  INVX1 INVX1_1006 ( .A(alu__abc_41358_n1452), .Y(alu__abc_41358_n1453) );
  INVX1 INVX1_1007 ( .A(alu__abc_41358_n766), .Y(alu__abc_41358_n1457) );
  INVX1 INVX1_1008 ( .A(alu__abc_41358_n1485), .Y(alu__abc_41358_n1486) );
  INVX1 INVX1_1009 ( .A(alu__abc_41358_n1496), .Y(alu__abc_41358_n1497) );
  INVX1 INVX1_101 ( .A(_abc_43815_n1389), .Y(_abc_43815_n1390) );
  INVX1 INVX1_1010 ( .A(alu__abc_41358_n1502), .Y(alu__abc_41358_n1503) );
  INVX1 INVX1_1011 ( .A(alu__abc_41358_n1530), .Y(alu__abc_41358_n1531) );
  INVX1 INVX1_1012 ( .A(alu__abc_41358_n1545), .Y(alu__abc_41358_n1546) );
  INVX1 INVX1_1013 ( .A(alu__abc_41358_n1549), .Y(alu__abc_41358_n1550) );
  INVX1 INVX1_1014 ( .A(alu__abc_41358_n1576), .Y(alu__abc_41358_n1577) );
  INVX1 INVX1_1015 ( .A(alu__abc_41358_n1588), .Y(alu__abc_41358_n1589) );
  INVX1 INVX1_1016 ( .A(alu__abc_41358_n1595), .Y(alu__abc_41358_n1596) );
  INVX1 INVX1_1017 ( .A(alu__abc_41358_n1599), .Y(alu__abc_41358_n1600) );
  INVX1 INVX1_1018 ( .A(alu__abc_41358_n1636), .Y(alu__abc_41358_n1637) );
  INVX1 INVX1_1019 ( .A(alu__abc_41358_n1640), .Y(alu__abc_41358_n1641) );
  INVX1 INVX1_102 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_43815_n1420) );
  INVX1 INVX1_1020 ( .A(alu__abc_41358_n1668), .Y(alu__abc_41358_n1669) );
  INVX1 INVX1_1021 ( .A(alu__abc_41358_n1679), .Y(alu__abc_41358_n1681) );
  INVX1 INVX1_1022 ( .A(alu__abc_41358_n1685), .Y(alu__abc_41358_n1686) );
  INVX1 INVX1_1023 ( .A(alu__abc_41358_n1713), .Y(alu__abc_41358_n1714) );
  INVX1 INVX1_1024 ( .A(alu__abc_41358_n1727), .Y(alu__abc_41358_n1728) );
  INVX1 INVX1_1025 ( .A(alu__abc_41358_n1734), .Y(alu__abc_41358_n1735) );
  INVX1 INVX1_1026 ( .A(alu__abc_41358_n1762), .Y(alu__abc_41358_n1763) );
  INVX1 INVX1_1027 ( .A(alu__abc_41358_n1772), .Y(alu__abc_41358_n1773) );
  INVX1 INVX1_1028 ( .A(alu__abc_41358_n1778), .Y(alu__abc_41358_n1779) );
  INVX1 INVX1_1029 ( .A(alu__abc_41358_n1783), .Y(alu__abc_41358_n1784) );
  INVX1 INVX1_103 ( .A(_abc_43815_n1421), .Y(_abc_43815_n1422) );
  INVX1 INVX1_1030 ( .A(alu__abc_41358_n1818), .Y(alu__abc_41358_n1819) );
  INVX1 INVX1_1031 ( .A(alu__abc_41358_n1823), .Y(alu__abc_41358_n1824) );
  INVX1 INVX1_1032 ( .A(alu__abc_41358_n1845), .Y(alu__abc_41358_n1846) );
  INVX1 INVX1_1033 ( .A(alu__abc_41358_n1859), .Y(alu__abc_41358_n1860) );
  INVX1 INVX1_1034 ( .A(alu__abc_41358_n811), .Y(alu__abc_41358_n1866) );
  INVX1 INVX1_1035 ( .A(alu__abc_41358_n1890), .Y(alu__abc_41358_n1891) );
  INVX1 INVX1_1036 ( .A(alu__abc_41358_n1902), .Y(alu__abc_41358_n1903) );
  INVX1 INVX1_1037 ( .A(alu__abc_41358_n1910), .Y(alu__abc_41358_n1911) );
  INVX1 INVX1_1038 ( .A(alu__abc_41358_n1934), .Y(alu__abc_41358_n1935) );
  INVX1 INVX1_1039 ( .A(alu__abc_41358_n1945), .Y(alu__abc_41358_n1947) );
  INVX1 INVX1_104 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_43815_n1442) );
  INVX1 INVX1_1040 ( .A(alu__abc_41358_n1952), .Y(alu__abc_41358_n1953) );
  INVX1 INVX1_1041 ( .A(alu__abc_41358_n1976), .Y(alu__abc_41358_n1977) );
  INVX1 INVX1_1042 ( .A(alu__abc_41358_n1988), .Y(alu__abc_41358_n1989) );
  INVX1 INVX1_1043 ( .A(alu__abc_41358_n1994), .Y(alu__abc_41358_n1995) );
  INVX1 INVX1_1044 ( .A(alu__abc_41358_n2015), .Y(alu__abc_41358_n2016) );
  INVX1 INVX1_1045 ( .A(alu__abc_41358_n2029), .Y(alu__abc_41358_n2030) );
  INVX1 INVX1_1046 ( .A(alu__abc_41358_n2033), .Y(alu__abc_41358_n2034) );
  INVX1 INVX1_1047 ( .A(alu__abc_41358_n2058), .Y(alu__abc_41358_n2059) );
  INVX1 INVX1_1048 ( .A(alu__abc_41358_n2071), .Y(alu__abc_41358_n2072) );
  INVX1 INVX1_1049 ( .A(alu__abc_41358_n2078), .Y(alu__abc_41358_n2079) );
  INVX1 INVX1_105 ( .A(_abc_43815_n1443_1), .Y(_abc_43815_n1444) );
  INVX1 INVX1_1050 ( .A(alu__abc_41358_n2101), .Y(alu__abc_41358_n2102) );
  INVX1 INVX1_1051 ( .A(alu__abc_41358_n2114), .Y(alu__abc_41358_n2115) );
  INVX1 INVX1_1052 ( .A(alu__abc_41358_n2118), .Y(alu__abc_41358_n2119) );
  INVX1 INVX1_1053 ( .A(alu__abc_41358_n2142), .Y(alu__abc_41358_n2143) );
  INVX1 INVX1_1054 ( .A(alu__abc_41358_n2155), .Y(alu__abc_41358_n2156) );
  INVX1 INVX1_1055 ( .A(alu__abc_41358_n2161), .Y(alu__abc_41358_n2162) );
  INVX1 INVX1_1056 ( .A(alu__abc_41358_n2180), .Y(alu__abc_41358_n2181) );
  INVX1 INVX1_1057 ( .A(alu__abc_41358_n2195), .Y(alu__abc_41358_n2196) );
  INVX1 INVX1_1058 ( .A(alu__abc_41358_n2199), .Y(alu__abc_41358_n2200) );
  INVX1 INVX1_1059 ( .A(alu__abc_41358_n2222), .Y(alu__abc_41358_n2223) );
  INVX1 INVX1_106 ( .A(sr_q_9_), .Y(_abc_43815_n1462) );
  INVX1 INVX1_1060 ( .A(alu__abc_41358_n2236), .Y(alu__abc_41358_n2237) );
  INVX1 INVX1_1061 ( .A(alu__abc_41358_n2241), .Y(alu__abc_41358_n2242) );
  INVX1 INVX1_1062 ( .A(alu__abc_41358_n2244), .Y(alu__abc_41358_n2245) );
  INVX1 INVX1_1063 ( .A(alu__abc_41358_n2266), .Y(alu__abc_41358_n2267) );
  INVX1 INVX1_1064 ( .A(alu__abc_41358_n2279), .Y(alu__abc_41358_n2280) );
  INVX1 INVX1_1065 ( .A(alu__abc_41358_n2283), .Y(alu__abc_41358_n2284) );
  INVX1 INVX1_1066 ( .A(alu__abc_41358_n2307), .Y(alu__abc_41358_n2308) );
  INVX1 INVX1_1067 ( .A(alu__abc_41358_n2321), .Y(alu__abc_41358_n2322) );
  INVX1 INVX1_1068 ( .A(alu__abc_41358_n2325), .Y(alu__abc_41358_n2326) );
  INVX1 INVX1_1069 ( .A(alu__abc_41358_n2344), .Y(alu__abc_41358_n2345) );
  INVX1 INVX1_107 ( .A(_abc_43815_n1463), .Y(_abc_43815_n1464) );
  INVX1 INVX1_1070 ( .A(alu__abc_41358_n2359), .Y(alu__abc_41358_n2360) );
  INVX1 INVX1_1071 ( .A(alu__abc_41358_n2363), .Y(alu__abc_41358_n2365) );
  INVX1 INVX1_1072 ( .A(alu__abc_41358_n2388), .Y(alu__abc_41358_n2389) );
  INVX1 INVX1_1073 ( .A(alu__abc_41358_n2401), .Y(alu__abc_41358_n2402) );
  INVX1 INVX1_1074 ( .A(alu__abc_41358_n2426), .Y(alu__abc_41358_n2427) );
  INVX1 INVX1_1075 ( .A(alu__abc_41358_n828), .Y(alu__abc_41358_n2440) );
  INVX1 INVX1_1076 ( .A(alu__abc_41358_n2464), .Y(alu__abc_41358_n2465) );
  INVX1 INVX1_1077 ( .A(alu__abc_41358_n2478), .Y(alu__abc_41358_n2479) );
  INVX1 INVX1_1078 ( .A(alu__abc_41358_n2560), .Y(alu_greater_than_o) );
  INVX1 INVX1_1079 ( .A(alu_equal_o), .Y(alu__abc_41358_n2562) );
  INVX1 INVX1_108 ( .A(_abc_43815_n1467), .Y(_abc_43815_n1468) );
  INVX1 INVX1_1080 ( .A(alu_less_than_signed_o), .Y(alu__abc_41358_n2563) );
  INVX1 INVX1_109 ( .A(_abc_43815_n1474), .Y(_abc_43815_n1475_1) );
  INVX1 INVX1_11 ( .A(_abc_43815_n640), .Y(_abc_43815_n665) );
  INVX1 INVX1_110 ( .A(pc_q_2_), .Y(_abc_43815_n1485) );
  INVX1 INVX1_111 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_43815_n1503) );
  INVX1 INVX1_112 ( .A(_abc_43815_n1504), .Y(_abc_43815_n1505) );
  INVX1 INVX1_113 ( .A(_abc_43815_n1510), .Y(_abc_43815_n1511) );
  INVX1 INVX1_114 ( .A(_abc_43815_n1513), .Y(_abc_43815_n1514) );
  INVX1 INVX1_115 ( .A(_abc_43815_n1524), .Y(_abc_43815_n1525) );
  INVX1 INVX1_116 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_43815_n1539) );
  INVX1 INVX1_117 ( .A(_abc_43815_n1540), .Y(_abc_43815_n1541) );
  INVX1 INVX1_118 ( .A(_abc_43815_n1547_1), .Y(_abc_43815_n1548) );
  INVX1 INVX1_119 ( .A(_abc_43815_n1551), .Y(_abc_43815_n1552) );
  INVX1 INVX1_12 ( .A(_abc_43815_n666), .Y(_abc_43815_n667) );
  INVX1 INVX1_120 ( .A(_abc_43815_n1561), .Y(_abc_43815_n1562) );
  INVX1 INVX1_121 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_43815_n1576) );
  INVX1 INVX1_122 ( .A(_abc_43815_n1577), .Y(_abc_43815_n1578) );
  INVX1 INVX1_123 ( .A(_abc_43815_n1582), .Y(_abc_43815_n1583_1) );
  INVX1 INVX1_124 ( .A(_abc_43815_n1585), .Y(_abc_43815_n1586_1) );
  INVX1 INVX1_125 ( .A(_abc_43815_n1590), .Y(_abc_43815_n1591) );
  INVX1 INVX1_126 ( .A(_abc_43815_n1601), .Y(_abc_43815_n1602_1) );
  INVX1 INVX1_127 ( .A(_abc_43815_n1618_1), .Y(_abc_43815_n1619) );
  INVX1 INVX1_128 ( .A(_abc_43815_n1622), .Y(_abc_43815_n1623) );
  INVX1 INVX1_129 ( .A(_abc_43815_n1633), .Y(_abc_43815_n1634_1) );
  INVX1 INVX1_13 ( .A(mem_ack_i), .Y(_abc_43815_n674_1) );
  INVX1 INVX1_130 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_43815_n1652) );
  INVX1 INVX1_131 ( .A(_abc_43815_n1653), .Y(_abc_43815_n1654) );
  INVX1 INVX1_132 ( .A(_abc_43815_n1658_1), .Y(_abc_43815_n1659) );
  INVX1 INVX1_133 ( .A(_abc_43815_n1664), .Y(_abc_43815_n1665) );
  INVX1 INVX1_134 ( .A(_abc_43815_n1666), .Y(_abc_43815_n1667) );
  INVX1 INVX1_135 ( .A(_abc_43815_n1678), .Y(_abc_43815_n1679) );
  INVX1 INVX1_136 ( .A(_abc_43815_n1694), .Y(_abc_43815_n1695) );
  INVX1 INVX1_137 ( .A(_abc_43815_n1701), .Y(_abc_43815_n1702) );
  INVX1 INVX1_138 ( .A(_abc_43815_n1705_1), .Y(_abc_43815_n1706_1) );
  INVX1 INVX1_139 ( .A(_abc_43815_n1709), .Y(_abc_43815_n1710) );
  INVX1 INVX1_14 ( .A(_abc_43815_n678), .Y(_abc_43815_n679_1) );
  INVX1 INVX1_140 ( .A(_abc_43815_n1731), .Y(_abc_43815_n1732) );
  INVX1 INVX1_141 ( .A(_abc_43815_n1096), .Y(_abc_43815_n1740) );
  INVX1 INVX1_142 ( .A(_abc_43815_n1742), .Y(_abc_43815_n1743) );
  INVX1 INVX1_143 ( .A(_abc_43815_n1745), .Y(_abc_43815_n1746) );
  INVX1 INVX1_144 ( .A(_abc_43815_n1747), .Y(_abc_43815_n1748) );
  INVX1 INVX1_145 ( .A(_abc_43815_n1770), .Y(_abc_43815_n1771) );
  INVX1 INVX1_146 ( .A(_abc_43815_n1425_1_bF_buf0), .Y(_abc_43815_n1779) );
  INVX1 INVX1_147 ( .A(_abc_43815_n1781_1), .Y(_abc_43815_n1782) );
  INVX1 INVX1_148 ( .A(_abc_43815_n1785_1), .Y(_abc_43815_n1786) );
  INVX1 INVX1_149 ( .A(_abc_43815_n1790), .Y(_abc_43815_n1791_1) );
  INVX1 INVX1_15 ( .A(mem_offset_q_0_), .Y(_abc_43815_n687) );
  INVX1 INVX1_150 ( .A(_abc_43815_n1811), .Y(_abc_43815_n1812) );
  INVX1 INVX1_151 ( .A(_abc_43815_n1818), .Y(_abc_43815_n1819) );
  INVX1 INVX1_152 ( .A(_abc_43815_n1821), .Y(_abc_43815_n1822) );
  INVX1 INVX1_153 ( .A(_abc_43815_n1823_1), .Y(_abc_43815_n1825) );
  INVX1 INVX1_154 ( .A(_abc_43815_n1847_1), .Y(_abc_43815_n1848) );
  INVX1 INVX1_155 ( .A(_abc_43815_n1860), .Y(_abc_43815_n1861) );
  INVX1 INVX1_156 ( .A(_abc_43815_n1864), .Y(_abc_43815_n1865_1) );
  INVX1 INVX1_157 ( .A(_abc_43815_n1868_1), .Y(_abc_43815_n1869) );
  INVX1 INVX1_158 ( .A(_abc_43815_n1871_1), .Y(_abc_43815_n1872) );
  INVX1 INVX1_159 ( .A(_abc_43815_n1891), .Y(_abc_43815_n1892) );
  INVX1 INVX1_16 ( .A(mem_offset_q_1_), .Y(_abc_43815_n688) );
  INVX1 INVX1_160 ( .A(_abc_43815_n1902), .Y(_abc_43815_n1903) );
  INVX1 INVX1_161 ( .A(_abc_43815_n1908), .Y(_abc_43815_n1909) );
  INVX1 INVX1_162 ( .A(_abc_43815_n1910), .Y(_abc_43815_n1911) );
  INVX1 INVX1_163 ( .A(_abc_43815_n1930), .Y(_abc_43815_n1931) );
  INVX1 INVX1_164 ( .A(_abc_43815_n1941), .Y(_abc_43815_n1942) );
  INVX1 INVX1_165 ( .A(_abc_43815_n1944), .Y(_abc_43815_n1945) );
  INVX1 INVX1_166 ( .A(_abc_43815_n1947), .Y(_abc_43815_n1948) );
  INVX1 INVX1_167 ( .A(_abc_43815_n1967), .Y(_abc_43815_n1968) );
  INVX1 INVX1_168 ( .A(_abc_43815_n1972), .Y(_abc_43815_n1973) );
  INVX1 INVX1_169 ( .A(_abc_43815_n1975), .Y(_abc_43815_n1976) );
  INVX1 INVX1_17 ( .A(_abc_43815_n644), .Y(_abc_43815_n690) );
  INVX1 INVX1_170 ( .A(_abc_43815_n1977), .Y(_abc_43815_n1979) );
  INVX1 INVX1_171 ( .A(_abc_43815_n2003), .Y(_abc_43815_n2004) );
  INVX1 INVX1_172 ( .A(_abc_43815_n2012), .Y(_abc_43815_n2013_1) );
  INVX1 INVX1_173 ( .A(_abc_43815_n2016), .Y(_abc_43815_n2017) );
  INVX1 INVX1_174 ( .A(_abc_43815_n2018), .Y(_abc_43815_n2019) );
  INVX1 INVX1_175 ( .A(_abc_43815_n2024), .Y(_abc_43815_n2025) );
  INVX1 INVX1_176 ( .A(_abc_43815_n2028), .Y(_abc_43815_n2029) );
  INVX1 INVX1_177 ( .A(_abc_43815_n2048), .Y(_abc_43815_n2049) );
  INVX1 INVX1_178 ( .A(_abc_43815_n2059), .Y(_abc_43815_n2060) );
  INVX1 INVX1_179 ( .A(_abc_43815_n2065), .Y(_abc_43815_n2066) );
  INVX1 INVX1_18 ( .A(opcode_q_21_), .Y(_abc_43815_n988) );
  INVX1 INVX1_180 ( .A(_abc_43815_n2067), .Y(_abc_43815_n2068) );
  INVX1 INVX1_181 ( .A(_abc_43815_n2087_1), .Y(_abc_43815_n2088) );
  INVX1 INVX1_182 ( .A(_abc_43815_n2094), .Y(_abc_43815_n2095) );
  INVX1 INVX1_183 ( .A(_abc_43815_n2097), .Y(_abc_43815_n2098) );
  INVX1 INVX1_184 ( .A(_abc_43815_n2100), .Y(_abc_43815_n2101_1) );
  INVX1 INVX1_185 ( .A(_abc_43815_n2124), .Y(_abc_43815_n2125) );
  INVX1 INVX1_186 ( .A(_abc_43815_n2129_1), .Y(_abc_43815_n2130) );
  INVX1 INVX1_187 ( .A(_abc_43815_n2132), .Y(_abc_43815_n2133) );
  INVX1 INVX1_188 ( .A(_abc_43815_n2134), .Y(_abc_43815_n2136) );
  INVX1 INVX1_189 ( .A(_abc_43815_n2160), .Y(_abc_43815_n2161) );
  INVX1 INVX1_19 ( .A(_abc_43815_n993_1), .Y(_abc_43815_n994_1) );
  INVX1 INVX1_190 ( .A(_abc_43815_n2093), .Y(_abc_43815_n2168) );
  INVX1 INVX1_191 ( .A(_abc_43815_n2175), .Y(_abc_43815_n2176) );
  INVX1 INVX1_192 ( .A(_abc_43815_n2179), .Y(_abc_43815_n2180) );
  INVX1 INVX1_193 ( .A(_abc_43815_n2203_1), .Y(_abc_43815_n2204) );
  INVX1 INVX1_194 ( .A(_abc_43815_n2210), .Y(_abc_43815_n2211) );
  INVX1 INVX1_195 ( .A(_abc_43815_n2218), .Y(_abc_43815_n2219) );
  INVX1 INVX1_196 ( .A(_abc_43815_n2241), .Y(_abc_43815_n2242_1) );
  INVX1 INVX1_197 ( .A(_abc_43815_n2247), .Y(_abc_43815_n2248) );
  INVX1 INVX1_198 ( .A(_abc_43815_n2250), .Y(_abc_43815_n2251) );
  INVX1 INVX1_199 ( .A(_abc_43815_n2253), .Y(_abc_43815_n2254) );
  INVX1 INVX1_2 ( .A(inst_r_4_), .Y(_abc_43815_n622) );
  INVX1 INVX1_20 ( .A(_abc_43815_n997), .Y(_abc_43815_n998) );
  INVX1 INVX1_200 ( .A(_abc_43815_n2277), .Y(_abc_43815_n2278) );
  INVX1 INVX1_201 ( .A(_abc_43815_n2282_1), .Y(_abc_43815_n2283) );
  INVX1 INVX1_202 ( .A(_abc_43815_n2285), .Y(_abc_43815_n2286) );
  INVX1 INVX1_203 ( .A(_abc_43815_n2287), .Y(_abc_43815_n2288) );
  INVX1 INVX1_204 ( .A(_abc_43815_n2313), .Y(_abc_43815_n2314) );
  INVX1 INVX1_205 ( .A(_abc_43815_n2328), .Y(_abc_43815_n2329) );
  INVX1 INVX1_206 ( .A(_abc_43815_n2331), .Y(_abc_43815_n2332_1) );
  INVX1 INVX1_207 ( .A(_abc_43815_n2356), .Y(_abc_43815_n2357) );
  INVX1 INVX1_208 ( .A(_abc_43815_n2362_1), .Y(_abc_43815_n2363) );
  INVX1 INVX1_209 ( .A(_abc_43815_n2368), .Y(_abc_43815_n2369) );
  INVX1 INVX1_21 ( .A(_abc_43815_n989), .Y(_abc_43815_n1001) );
  INVX1 INVX1_210 ( .A(_abc_43815_n2370), .Y(_abc_43815_n2371) );
  INVX1 INVX1_211 ( .A(_abc_43815_n2395), .Y(_abc_43815_n2396_1) );
  INVX1 INVX1_212 ( .A(_abc_43815_n2401), .Y(_abc_43815_n2402) );
  INVX1 INVX1_213 ( .A(_abc_43815_n2404), .Y(_abc_43815_n2405) );
  INVX1 INVX1_214 ( .A(_abc_43815_n2407), .Y(_abc_43815_n2408) );
  INVX1 INVX1_215 ( .A(_abc_43815_n2432), .Y(_abc_43815_n2433) );
  INVX1 INVX1_216 ( .A(_abc_43815_n2438), .Y(_abc_43815_n2439) );
  INVX1 INVX1_217 ( .A(_abc_43815_n2443), .Y(_abc_43815_n2444) );
  INVX1 INVX1_218 ( .A(_abc_43815_n2446), .Y(_abc_43815_n2447) );
  INVX1 INVX1_219 ( .A(_abc_43815_n2471), .Y(_abc_43815_n2472) );
  INVX1 INVX1_22 ( .A(opcode_q_23_), .Y(_abc_43815_n1002) );
  INVX1 INVX1_220 ( .A(_abc_43815_n2478), .Y(_abc_43815_n2479) );
  INVX1 INVX1_221 ( .A(_abc_43815_n2484), .Y(_abc_43815_n2485) );
  INVX1 INVX1_222 ( .A(_abc_43815_n2487), .Y(_abc_43815_n2488) );
  INVX1 INVX1_223 ( .A(_abc_43815_n2512), .Y(_abc_43815_n2513) );
  INVX1 INVX1_224 ( .A(_abc_43815_n2517_1), .Y(_abc_43815_n2518) );
  INVX1 INVX1_225 ( .A(_abc_43815_n2520), .Y(_abc_43815_n2521) );
  INVX1 INVX1_226 ( .A(_abc_43815_n2522), .Y(_abc_43815_n2523) );
  INVX1 INVX1_227 ( .A(_abc_43815_n2548), .Y(_abc_43815_n2549) );
  INVX1 INVX1_228 ( .A(_abc_43815_n2555), .Y(_abc_43815_n2556) );
  INVX1 INVX1_229 ( .A(_abc_43815_n2559), .Y(_abc_43815_n2560) );
  INVX1 INVX1_23 ( .A(_abc_43815_n1003), .Y(_abc_43815_n1004) );
  INVX1 INVX1_230 ( .A(_abc_43815_n2562), .Y(_abc_43815_n2563) );
  INVX1 INVX1_231 ( .A(_abc_43815_n2587), .Y(_abc_43815_n2588) );
  INVX1 INVX1_232 ( .A(_abc_43815_n2592), .Y(_abc_43815_n2593) );
  INVX1 INVX1_233 ( .A(pc_q_31_), .Y(_abc_43815_n2595) );
  INVX1 INVX1_234 ( .A(_abc_43815_n2597), .Y(_abc_43815_n2599) );
  INVX1 INVX1_235 ( .A(_abc_43815_n1190), .Y(_abc_43815_n2675) );
  INVX1 INVX1_236 ( .A(_abc_43815_n670_1), .Y(_abc_43815_n2762) );
  INVX1 INVX1_237 ( .A(_abc_43815_n984), .Y(_abc_43815_n2893) );
  INVX1 INVX1_238 ( .A(_abc_43815_n680_1_bF_buf2), .Y(_abc_43815_n3314) );
  INVX1 INVX1_239 ( .A(_abc_43815_n3315), .Y(_abc_43815_n3316_1) );
  INVX1 INVX1_24 ( .A(_abc_43815_n1009_1), .Y(_abc_43815_n1010) );
  INVX1 INVX1_240 ( .A(_abc_43815_n3321), .Y(_abc_43815_n3322) );
  INVX1 INVX1_241 ( .A(_abc_43815_n3323_1), .Y(_abc_43815_n3324_1) );
  INVX1 INVX1_242 ( .A(_abc_43815_n3327), .Y(_abc_43815_n3328) );
  INVX1 INVX1_243 ( .A(\mem_dat_i[0] ), .Y(_abc_43815_n3333) );
  INVX1 INVX1_244 ( .A(_abc_43815_n3334), .Y(_abc_43815_n3335) );
  INVX1 INVX1_245 ( .A(\mem_dat_i[1] ), .Y(_abc_43815_n3338) );
  INVX1 INVX1_246 ( .A(_abc_43815_n3339_1), .Y(_abc_43815_n3340_1) );
  INVX1 INVX1_247 ( .A(\mem_dat_i[2] ), .Y(_abc_43815_n3343) );
  INVX1 INVX1_248 ( .A(_abc_43815_n3344), .Y(_abc_43815_n3345) );
  INVX1 INVX1_249 ( .A(\mem_dat_i[3] ), .Y(_abc_43815_n3348_1) );
  INVX1 INVX1_25 ( .A(_abc_43815_n1014), .Y(_abc_43815_n1015) );
  INVX1 INVX1_250 ( .A(_abc_43815_n3349), .Y(_abc_43815_n3350) );
  INVX1 INVX1_251 ( .A(\mem_dat_i[4] ), .Y(_abc_43815_n3353) );
  INVX1 INVX1_252 ( .A(_abc_43815_n3354), .Y(_abc_43815_n3355) );
  INVX1 INVX1_253 ( .A(\mem_dat_i[5] ), .Y(_abc_43815_n3358) );
  INVX1 INVX1_254 ( .A(_abc_43815_n3359_1), .Y(_abc_43815_n3360_1) );
  INVX1 INVX1_255 ( .A(\mem_dat_i[6] ), .Y(_abc_43815_n3363) );
  INVX1 INVX1_256 ( .A(_abc_43815_n3364), .Y(_abc_43815_n3365) );
  INVX1 INVX1_257 ( .A(\mem_dat_i[7] ), .Y(_abc_43815_n3368) );
  INVX1 INVX1_258 ( .A(_abc_43815_n3369_1), .Y(_abc_43815_n3370_1) );
  INVX1 INVX1_259 ( .A(\mem_dat_i[8] ), .Y(_abc_43815_n3373) );
  INVX1 INVX1_26 ( .A(opcode_q_24_), .Y(_abc_43815_n1016) );
  INVX1 INVX1_260 ( .A(_abc_43815_n3374), .Y(_abc_43815_n3375) );
  INVX1 INVX1_261 ( .A(\mem_dat_i[9] ), .Y(_abc_43815_n3378) );
  INVX1 INVX1_262 ( .A(_abc_43815_n3379_1), .Y(_abc_43815_n3380_1) );
  INVX1 INVX1_263 ( .A(\mem_dat_i[10] ), .Y(_abc_43815_n3383) );
  INVX1 INVX1_264 ( .A(_abc_43815_n3384), .Y(_abc_43815_n3385) );
  INVX1 INVX1_265 ( .A(\mem_dat_i[11] ), .Y(_abc_43815_n3388) );
  INVX1 INVX1_266 ( .A(_abc_43815_n3389_1), .Y(_abc_43815_n3390_1) );
  INVX1 INVX1_267 ( .A(\mem_dat_i[12] ), .Y(_abc_43815_n3393) );
  INVX1 INVX1_268 ( .A(_abc_43815_n3394), .Y(_abc_43815_n3395) );
  INVX1 INVX1_269 ( .A(\mem_dat_i[13] ), .Y(_abc_43815_n3398) );
  INVX1 INVX1_27 ( .A(_abc_43815_n1020), .Y(_abc_43815_n1021) );
  INVX1 INVX1_270 ( .A(_abc_43815_n3399_1), .Y(_abc_43815_n3400_1) );
  INVX1 INVX1_271 ( .A(\mem_dat_i[14] ), .Y(_abc_43815_n3403) );
  INVX1 INVX1_272 ( .A(_abc_43815_n3404), .Y(_abc_43815_n3405) );
  INVX1 INVX1_273 ( .A(\mem_dat_i[15] ), .Y(_abc_43815_n3408) );
  INVX1 INVX1_274 ( .A(_abc_43815_n3409_1), .Y(_abc_43815_n3410_1) );
  INVX1 INVX1_275 ( .A(\mem_dat_i[16] ), .Y(_abc_43815_n3413) );
  INVX1 INVX1_276 ( .A(_abc_43815_n3414), .Y(_abc_43815_n3415) );
  INVX1 INVX1_277 ( .A(\mem_dat_i[17] ), .Y(_abc_43815_n3418) );
  INVX1 INVX1_278 ( .A(_abc_43815_n3419_1), .Y(_abc_43815_n3420_1) );
  INVX1 INVX1_279 ( .A(\mem_dat_i[18] ), .Y(_abc_43815_n3423) );
  INVX1 INVX1_28 ( .A(_abc_43815_n1024), .Y(_abc_43815_n1025) );
  INVX1 INVX1_280 ( .A(_abc_43815_n3424), .Y(_abc_43815_n3425) );
  INVX1 INVX1_281 ( .A(\mem_dat_i[19] ), .Y(_abc_43815_n3428) );
  INVX1 INVX1_282 ( .A(_abc_43815_n3429_1), .Y(_abc_43815_n3430_1) );
  INVX1 INVX1_283 ( .A(\mem_dat_i[20] ), .Y(_abc_43815_n3433) );
  INVX1 INVX1_284 ( .A(_abc_43815_n3434), .Y(_abc_43815_n3435) );
  INVX1 INVX1_285 ( .A(\mem_dat_i[21] ), .Y(_abc_43815_n3438_1) );
  INVX1 INVX1_286 ( .A(_abc_43815_n3439_1), .Y(_abc_43815_n3440) );
  INVX1 INVX1_287 ( .A(\mem_dat_i[22] ), .Y(_abc_43815_n3443) );
  INVX1 INVX1_288 ( .A(_abc_43815_n3444), .Y(_abc_43815_n3445) );
  INVX1 INVX1_289 ( .A(\mem_dat_i[23] ), .Y(_abc_43815_n3448_1) );
  INVX1 INVX1_29 ( .A(opcode_q_22_), .Y(_abc_43815_n1033) );
  INVX1 INVX1_290 ( .A(_abc_43815_n3449), .Y(_abc_43815_n3450) );
  INVX1 INVX1_291 ( .A(\mem_dat_i[24] ), .Y(_abc_43815_n3453) );
  INVX1 INVX1_292 ( .A(_abc_43815_n3454), .Y(_abc_43815_n3455) );
  INVX1 INVX1_293 ( .A(\mem_dat_i[25] ), .Y(_abc_43815_n3458) );
  INVX1 INVX1_294 ( .A(_abc_43815_n3459), .Y(_abc_43815_n3460) );
  INVX1 INVX1_295 ( .A(\mem_dat_i[26] ), .Y(_abc_43815_n3463) );
  INVX1 INVX1_296 ( .A(_abc_43815_n3464), .Y(_abc_43815_n3465_1) );
  INVX1 INVX1_297 ( .A(\mem_dat_i[27] ), .Y(_abc_43815_n3468) );
  INVX1 INVX1_298 ( .A(_abc_43815_n3469), .Y(_abc_43815_n3470) );
  INVX1 INVX1_299 ( .A(\mem_dat_i[28] ), .Y(_abc_43815_n3473) );
  INVX1 INVX1_3 ( .A(inst_r_5_), .Y(_abc_43815_n623) );
  INVX1 INVX1_30 ( .A(_abc_43815_n1034), .Y(_abc_43815_n1035) );
  INVX1 INVX1_300 ( .A(_abc_43815_n3474_1), .Y(_abc_43815_n3475_1) );
  INVX1 INVX1_301 ( .A(\mem_dat_i[29] ), .Y(_abc_43815_n3478) );
  INVX1 INVX1_302 ( .A(_abc_43815_n3479), .Y(_abc_43815_n3480) );
  INVX1 INVX1_303 ( .A(\mem_dat_i[30] ), .Y(_abc_43815_n3483_1) );
  INVX1 INVX1_304 ( .A(_abc_43815_n3484_1), .Y(_abc_43815_n3485) );
  INVX1 INVX1_305 ( .A(\mem_dat_i[31] ), .Y(_abc_43815_n3488) );
  INVX1 INVX1_306 ( .A(_abc_43815_n3489), .Y(_abc_43815_n3490) );
  INVX1 INVX1_307 ( .A(_abc_43815_n651_1), .Y(_abc_43815_n3493_1) );
  INVX1 INVX1_308 ( .A(_abc_43815_n3317_bF_buf2), .Y(_abc_43815_n3495) );
  INVX1 INVX1_309 ( .A(_abc_43815_n3540), .Y(_abc_43815_n3964) );
  INVX1 INVX1_31 ( .A(_abc_43815_n624_1), .Y(_abc_43815_n1041) );
  INVX1 INVX1_310 ( .A(state_q_3_bF_buf4), .Y(_abc_43815_n3967) );
  INVX1 INVX1_311 ( .A(state_q_2_), .Y(_abc_43815_n3977) );
  INVX1 INVX1_312 ( .A(_abc_43815_n3992), .Y(_abc_43815_n3993) );
  INVX1 INVX1_313 ( .A(_abc_43815_n3995_1), .Y(_abc_43815_n3996) );
  INVX1 INVX1_314 ( .A(_abc_43815_n4010), .Y(_abc_43815_n4011) );
  INVX1 INVX1_315 ( .A(_abc_43815_n4009), .Y(_abc_43815_n4014) );
  INVX1 INVX1_316 ( .A(_abc_43815_n4012), .Y(_abc_43815_n4015_1) );
  INVX1 INVX1_317 ( .A(_abc_43815_n4021), .Y(_abc_43815_n4022_1) );
  INVX1 INVX1_318 ( .A(_abc_43815_n4026), .Y(_abc_43815_n4027) );
  INVX1 INVX1_319 ( .A(_abc_43815_n4039), .Y(_abc_43815_n4040) );
  INVX1 INVX1_32 ( .A(_abc_43815_n1044), .Y(_abc_43815_n1045) );
  INVX1 INVX1_320 ( .A(_abc_43815_n4041_1), .Y(_abc_43815_n4042) );
  INVX1 INVX1_321 ( .A(_abc_43815_n4038), .Y(_abc_43815_n4044) );
  INVX1 INVX1_322 ( .A(_abc_43815_n4052), .Y(_abc_43815_n4053) );
  INVX1 INVX1_323 ( .A(_abc_43815_n4058), .Y(_abc_43815_n4059) );
  INVX1 INVX1_324 ( .A(_abc_43815_n4067), .Y(_abc_43815_n4068_1) );
  INVX1 INVX1_325 ( .A(_abc_43815_n4069), .Y(_abc_43815_n4070) );
  INVX1 INVX1_326 ( .A(_abc_43815_n4066), .Y(_abc_43815_n4072) );
  INVX1 INVX1_327 ( .A(_abc_43815_n4082_1), .Y(_abc_43815_n4083) );
  INVX1 INVX1_328 ( .A(_abc_43815_n4084), .Y(_abc_43815_n4085) );
  INVX1 INVX1_329 ( .A(_abc_43815_n4089_1), .Y(_abc_43815_n4090) );
  INVX1 INVX1_33 ( .A(_abc_43815_n1048), .Y(_abc_43815_n1049) );
  INVX1 INVX1_330 ( .A(_abc_43815_n4081), .Y(_abc_43815_n4097) );
  INVX1 INVX1_331 ( .A(_abc_43815_n4099), .Y(_abc_43815_n4100) );
  INVX1 INVX1_332 ( .A(_abc_43815_n4101_1), .Y(_abc_43815_n4102) );
  INVX1 INVX1_333 ( .A(_abc_43815_n4098), .Y(_abc_43815_n4104) );
  INVX1 INVX1_334 ( .A(_abc_43815_n4115), .Y(_abc_43815_n4116) );
  INVX1 INVX1_335 ( .A(_abc_43815_n4120), .Y(_abc_43815_n4121) );
  INVX1 INVX1_336 ( .A(_abc_43815_n4123), .Y(_abc_43815_n4124_1) );
  INVX1 INVX1_337 ( .A(_abc_43815_n4119_1), .Y(_abc_43815_n4131_1) );
  INVX1 INVX1_338 ( .A(_abc_43815_n4136), .Y(_abc_43815_n4137) );
  INVX1 INVX1_339 ( .A(_abc_43815_n4139), .Y(_abc_43815_n4140) );
  INVX1 INVX1_34 ( .A(_abc_43815_n1050), .Y(_abc_43815_n1051) );
  INVX1 INVX1_340 ( .A(_abc_43815_n4132), .Y(_abc_43815_n4142) );
  INVX1 INVX1_341 ( .A(_abc_43815_n4153), .Y(_abc_43815_n4154) );
  INVX1 INVX1_342 ( .A(_abc_43815_n4166_1), .Y(_abc_43815_n4167_1) );
  INVX1 INVX1_343 ( .A(_abc_43815_n4177), .Y(_abc_43815_n4178) );
  INVX1 INVX1_344 ( .A(_abc_43815_n4184), .Y(_abc_43815_n4185) );
  INVX1 INVX1_345 ( .A(_abc_43815_n4186), .Y(_abc_43815_n4187) );
  INVX1 INVX1_346 ( .A(_abc_43815_n4196), .Y(_abc_43815_n4197) );
  INVX1 INVX1_347 ( .A(_abc_43815_n4201), .Y(_abc_43815_n4202) );
  INVX1 INVX1_348 ( .A(_abc_43815_n4205), .Y(_abc_43815_n4206) );
  INVX1 INVX1_349 ( .A(_abc_43815_n4218), .Y(_abc_43815_n4219) );
  INVX1 INVX1_35 ( .A(_abc_43815_n1058), .Y(_abc_43815_n1059) );
  INVX1 INVX1_350 ( .A(_abc_43815_n4221), .Y(_abc_43815_n4222) );
  INVX1 INVX1_351 ( .A(_abc_43815_n4223), .Y(_abc_43815_n4224) );
  INVX1 INVX1_352 ( .A(_abc_43815_n4214), .Y(_abc_43815_n4226) );
  INVX1 INVX1_353 ( .A(_abc_43815_n4234), .Y(_abc_43815_n4235) );
  INVX1 INVX1_354 ( .A(_abc_43815_n4238), .Y(_abc_43815_n4239) );
  INVX1 INVX1_355 ( .A(_abc_43815_n4240), .Y(_abc_43815_n4241) );
  INVX1 INVX1_356 ( .A(_abc_43815_n4245), .Y(_abc_43815_n4246) );
  INVX1 INVX1_357 ( .A(_abc_43815_n4250), .Y(_abc_43815_n4251) );
  INVX1 INVX1_358 ( .A(_abc_43815_n4259), .Y(_abc_43815_n4260) );
  INVX1 INVX1_359 ( .A(_abc_43815_n4262), .Y(_abc_43815_n4263) );
  INVX1 INVX1_36 ( .A(_abc_43815_n1060_bF_buf3), .Y(_abc_43815_n1061) );
  INVX1 INVX1_360 ( .A(_abc_43815_n4258), .Y(_abc_43815_n4265) );
  INVX1 INVX1_361 ( .A(_abc_43815_n4273), .Y(_abc_43815_n4274) );
  INVX1 INVX1_362 ( .A(_abc_43815_n4277), .Y(_abc_43815_n4278) );
  INVX1 INVX1_363 ( .A(_abc_43815_n4283), .Y(_abc_43815_n4284) );
  INVX1 INVX1_364 ( .A(_abc_43815_n4292), .Y(_abc_43815_n4293) );
  INVX1 INVX1_365 ( .A(_abc_43815_n4295), .Y(_abc_43815_n4296) );
  INVX1 INVX1_366 ( .A(_abc_43815_n4291), .Y(_abc_43815_n4298) );
  INVX1 INVX1_367 ( .A(_abc_43815_n4309), .Y(_abc_43815_n4310) );
  INVX1 INVX1_368 ( .A(_abc_43815_n4312), .Y(_abc_43815_n4313) );
  INVX1 INVX1_369 ( .A(_abc_43815_n4315), .Y(_abc_43815_n4316) );
  INVX1 INVX1_37 ( .A(_abc_43815_n1069), .Y(_abc_43815_n1070) );
  INVX1 INVX1_370 ( .A(_abc_43815_n4320), .Y(_abc_43815_n4321) );
  INVX1 INVX1_371 ( .A(_abc_43815_n4329), .Y(_abc_43815_n4330) );
  INVX1 INVX1_372 ( .A(_abc_43815_n4332), .Y(_abc_43815_n4333) );
  INVX1 INVX1_373 ( .A(_abc_43815_n4328), .Y(_abc_43815_n4335) );
  INVX1 INVX1_374 ( .A(_abc_43815_n4347), .Y(_abc_43815_n4348) );
  INVX1 INVX1_375 ( .A(_abc_43815_n4352), .Y(_abc_43815_n4353) );
  INVX1 INVX1_376 ( .A(_abc_43815_n4360), .Y(_abc_43815_n4361) );
  INVX1 INVX1_377 ( .A(_abc_43815_n4362), .Y(_abc_43815_n4363) );
  INVX1 INVX1_378 ( .A(_abc_43815_n4365), .Y(_abc_43815_n4367) );
  INVX1 INVX1_379 ( .A(_abc_43815_n4376), .Y(_abc_43815_n4377) );
  INVX1 INVX1_38 ( .A(_abc_43815_n1073), .Y(_abc_43815_n1074) );
  INVX1 INVX1_380 ( .A(_abc_43815_n4379), .Y(_abc_43815_n4380) );
  INVX1 INVX1_381 ( .A(_abc_43815_n4384), .Y(_abc_43815_n4385) );
  INVX1 INVX1_382 ( .A(_abc_43815_n4389), .Y(_abc_43815_n4390) );
  INVX1 INVX1_383 ( .A(_abc_43815_n4398), .Y(_abc_43815_n4399) );
  INVX1 INVX1_384 ( .A(_abc_43815_n4401), .Y(_abc_43815_n4402) );
  INVX1 INVX1_385 ( .A(_abc_43815_n4397), .Y(_abc_43815_n4404) );
  INVX1 INVX1_386 ( .A(_abc_43815_n4414), .Y(_abc_43815_n4415) );
  INVX1 INVX1_387 ( .A(_abc_43815_n4417), .Y(_abc_43815_n4418) );
  INVX1 INVX1_388 ( .A(_abc_43815_n4422), .Y(_abc_43815_n4423) );
  INVX1 INVX1_389 ( .A(_abc_43815_n4431), .Y(_abc_43815_n4432) );
  INVX1 INVX1_39 ( .A(_abc_43815_n1075), .Y(_abc_43815_n1076) );
  INVX1 INVX1_390 ( .A(_abc_43815_n4434), .Y(_abc_43815_n4435) );
  INVX1 INVX1_391 ( .A(_abc_43815_n4430), .Y(_abc_43815_n4437) );
  INVX1 INVX1_392 ( .A(_abc_43815_n4383), .Y(_abc_43815_n4445) );
  INVX1 INVX1_393 ( .A(_abc_43815_n4412), .Y(_abc_43815_n4446) );
  INVX1 INVX1_394 ( .A(_abc_43815_n4447), .Y(_abc_43815_n4448) );
  INVX1 INVX1_395 ( .A(_abc_43815_n4451), .Y(_abc_43815_n4452) );
  INVX1 INVX1_396 ( .A(_abc_43815_n4455), .Y(_abc_43815_n4456) );
  INVX1 INVX1_397 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_43815_n4458) );
  INVX1 INVX1_398 ( .A(_abc_43815_n4460), .Y(_abc_43815_n4461) );
  INVX1 INVX1_399 ( .A(_abc_43815_n4463), .Y(_abc_43815_n4464) );
  INVX1 INVX1_4 ( .A(inst_r_2_), .Y(_abc_43815_n625) );
  INVX1 INVX1_40 ( .A(_abc_43815_n1080), .Y(_abc_43815_n1081) );
  INVX1 INVX1_400 ( .A(_abc_43815_n4471), .Y(_abc_43815_n4472) );
  INVX1 INVX1_401 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_43815_n4474) );
  INVX1 INVX1_402 ( .A(_abc_43815_n4476), .Y(_abc_43815_n4478) );
  INVX1 INVX1_403 ( .A(_abc_43815_n4486), .Y(_abc_43815_n4487) );
  INVX1 INVX1_404 ( .A(_abc_43815_n4492), .Y(_abc_43815_n4493) );
  INVX1 INVX1_405 ( .A(_abc_43815_n4495), .Y(_abc_43815_n4496) );
  INVX1 INVX1_406 ( .A(_abc_43815_n4489), .Y(_abc_43815_n4498) );
  INVX1 INVX1_407 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_43815_n4507) );
  INVX1 INVX1_408 ( .A(_abc_43815_n4510), .Y(_abc_43815_n4511) );
  INVX1 INVX1_409 ( .A(_abc_43815_n4506), .Y(_abc_43815_n4513) );
  INVX1 INVX1_41 ( .A(_abc_43815_n1011), .Y(_abc_43815_n1086_1) );
  INVX1 INVX1_410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2106_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2107) );
  INVX1 INVX1_411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2111_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2112_1) );
  INVX1 INVX1_412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2116), .Y(REGFILE_SIM_reg_bank__abc_33898_n2117_1) );
  INVX1 INVX1_413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2121_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2122) );
  INVX1 INVX1_414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2126_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2127_1) );
  INVX1 INVX1_415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2131), .Y(REGFILE_SIM_reg_bank__abc_33898_n2132_1) );
  INVX1 INVX1_416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2136_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2137) );
  INVX1 INVX1_417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2141_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2142_1) );
  INVX1 INVX1_418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2146), .Y(REGFILE_SIM_reg_bank__abc_33898_n2147_1) );
  INVX1 INVX1_419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2151_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2152) );
  INVX1 INVX1_42 ( .A(_abc_43815_n1017), .Y(_abc_43815_n1090) );
  INVX1 INVX1_420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2156_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2157_1) );
  INVX1 INVX1_421 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2161), .Y(REGFILE_SIM_reg_bank__abc_33898_n2162_1) );
  INVX1 INVX1_422 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2166_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2167) );
  INVX1 INVX1_423 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2171_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2172_1) );
  INVX1 INVX1_424 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2176), .Y(REGFILE_SIM_reg_bank__abc_33898_n2177_1) );
  INVX1 INVX1_425 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2181_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2182) );
  INVX1 INVX1_426 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2186_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2187_1) );
  INVX1 INVX1_427 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2191), .Y(REGFILE_SIM_reg_bank__abc_33898_n2192_1) );
  INVX1 INVX1_428 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2196_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2197) );
  INVX1 INVX1_429 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2201), .Y(REGFILE_SIM_reg_bank__abc_33898_n2202_1) );
  INVX1 INVX1_43 ( .A(alu_op_r_7_), .Y(_abc_43815_n1107) );
  INVX1 INVX1_430 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2206_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2207) );
  INVX1 INVX1_431 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2211_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2212_1) );
  INVX1 INVX1_432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2216), .Y(REGFILE_SIM_reg_bank__abc_33898_n2217_1) );
  INVX1 INVX1_433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2221_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2222) );
  INVX1 INVX1_434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2226_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2227_1) );
  INVX1 INVX1_435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2231), .Y(REGFILE_SIM_reg_bank__abc_33898_n2232_1) );
  INVX1 INVX1_436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2236_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2237) );
  INVX1 INVX1_437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2241_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2242_1) );
  INVX1 INVX1_438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2246), .Y(REGFILE_SIM_reg_bank__abc_33898_n2247_1) );
  INVX1 INVX1_439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2251_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2252) );
  INVX1 INVX1_44 ( .A(alu_op_r_6_), .Y(_abc_43815_n1108_1) );
  INVX1 INVX1_440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2256_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2257_1) );
  INVX1 INVX1_441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2261), .Y(REGFILE_SIM_reg_bank__abc_33898_n2262_1) );
  INVX1 INVX1_442 ( .A(REGFILE_SIM_reg_bank_rd_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2264) );
  INVX1 INVX1_443 ( .A(REGFILE_SIM_reg_bank_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2365_1) );
  INVX1 INVX1_444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2470), .Y(REGFILE_SIM_reg_bank__abc_33898_n2471_1) );
  INVX1 INVX1_445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2474_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2475_1) );
  INVX1 INVX1_446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2478_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2479) );
  INVX1 INVX1_447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2482), .Y(REGFILE_SIM_reg_bank__abc_33898_n2483_1) );
  INVX1 INVX1_448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2486_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2487_1) );
  INVX1 INVX1_449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2490), .Y(REGFILE_SIM_reg_bank__abc_33898_n2491_1) );
  INVX1 INVX1_45 ( .A(alu_op_r_4_), .Y(_abc_43815_n1110) );
  INVX1 INVX1_450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2494_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2495) );
  INVX1 INVX1_451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2498), .Y(REGFILE_SIM_reg_bank__abc_33898_n2499_1) );
  INVX1 INVX1_452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2502_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2503_1) );
  INVX1 INVX1_453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2506_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2507) );
  INVX1 INVX1_454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2510), .Y(REGFILE_SIM_reg_bank__abc_33898_n2511_1) );
  INVX1 INVX1_455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2514_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2515_1) );
  INVX1 INVX1_456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2518_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2519) );
  INVX1 INVX1_457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2522), .Y(REGFILE_SIM_reg_bank__abc_33898_n2523_1) );
  INVX1 INVX1_458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2526_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2527_1) );
  INVX1 INVX1_459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2530_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2531) );
  INVX1 INVX1_46 ( .A(alu_op_r_5_), .Y(_abc_43815_n1111) );
  INVX1 INVX1_460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2534), .Y(REGFILE_SIM_reg_bank__abc_33898_n2535_1) );
  INVX1 INVX1_461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2538_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2539_1) );
  INVX1 INVX1_462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2542_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2543) );
  INVX1 INVX1_463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2546), .Y(REGFILE_SIM_reg_bank__abc_33898_n2547_1) );
  INVX1 INVX1_464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2550_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2551_1) );
  INVX1 INVX1_465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2554_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2555) );
  INVX1 INVX1_466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2558), .Y(REGFILE_SIM_reg_bank__abc_33898_n2559_1) );
  INVX1 INVX1_467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2562_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2563_1) );
  INVX1 INVX1_468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2566_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2567) );
  INVX1 INVX1_469 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2570), .Y(REGFILE_SIM_reg_bank__abc_33898_n2571_1) );
  INVX1 INVX1_47 ( .A(alu_op_r_2_), .Y(_abc_43815_n1114) );
  INVX1 INVX1_470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2574_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2575_1) );
  INVX1 INVX1_471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2578_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2579) );
  INVX1 INVX1_472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2582), .Y(REGFILE_SIM_reg_bank__abc_33898_n2583_1) );
  INVX1 INVX1_473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2586_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2587) );
  INVX1 INVX1_474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2590_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2591_1) );
  INVX1 INVX1_475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2594_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2595) );
  INVX1 INVX1_476 ( .A(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2597_1) );
  INVX1 INVX1_477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2701), .Y(REGFILE_SIM_reg_bank__abc_33898_n2702_1) );
  INVX1 INVX1_478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2705_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2706_1) );
  INVX1 INVX1_479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2709_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2710) );
  INVX1 INVX1_48 ( .A(alu_op_r_1_), .Y(_abc_43815_n1116_1) );
  INVX1 INVX1_480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2713), .Y(REGFILE_SIM_reg_bank__abc_33898_n2714_1) );
  INVX1 INVX1_481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2717_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2718_1) );
  INVX1 INVX1_482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2721_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2722) );
  INVX1 INVX1_483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2725), .Y(REGFILE_SIM_reg_bank__abc_33898_n2726_1) );
  INVX1 INVX1_484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2729_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2730_1) );
  INVX1 INVX1_485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2733_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2734) );
  INVX1 INVX1_486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2737), .Y(REGFILE_SIM_reg_bank__abc_33898_n2738_1) );
  INVX1 INVX1_487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2741_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2742_1) );
  INVX1 INVX1_488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2745_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2746) );
  INVX1 INVX1_489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2749), .Y(REGFILE_SIM_reg_bank__abc_33898_n2750_1) );
  INVX1 INVX1_49 ( .A(alu_op_r_0_), .Y(_abc_43815_n1117) );
  INVX1 INVX1_490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2753_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2754_1) );
  INVX1 INVX1_491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2757_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2758) );
  INVX1 INVX1_492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2761), .Y(REGFILE_SIM_reg_bank__abc_33898_n2762_1) );
  INVX1 INVX1_493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2765_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2766_1) );
  INVX1 INVX1_494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2769_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2770) );
  INVX1 INVX1_495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2773), .Y(REGFILE_SIM_reg_bank__abc_33898_n2774_1) );
  INVX1 INVX1_496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2777_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2778_1) );
  INVX1 INVX1_497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2781), .Y(REGFILE_SIM_reg_bank__abc_33898_n2782_1) );
  INVX1 INVX1_498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2785_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2786) );
  INVX1 INVX1_499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2789), .Y(REGFILE_SIM_reg_bank__abc_33898_n2790_1) );
  INVX1 INVX1_5 ( .A(inst_r_1_), .Y(_abc_43815_n629) );
  INVX1 INVX1_50 ( .A(_abc_43815_n1121), .Y(_abc_43815_n1122) );
  INVX1 INVX1_500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2793_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2794_1) );
  INVX1 INVX1_501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2797_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2798) );
  INVX1 INVX1_502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2801), .Y(REGFILE_SIM_reg_bank__abc_33898_n2802_1) );
  INVX1 INVX1_503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2805_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2806_1) );
  INVX1 INVX1_504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2809_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2810) );
  INVX1 INVX1_505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2813), .Y(REGFILE_SIM_reg_bank__abc_33898_n2814_1) );
  INVX1 INVX1_506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2817_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2818_1) );
  INVX1 INVX1_507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2821_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2822) );
  INVX1 INVX1_508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2825), .Y(REGFILE_SIM_reg_bank__abc_33898_n2826_1) );
  INVX1 INVX1_509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2831), .Y(REGFILE_SIM_reg_bank__abc_33898_n2832_1) );
  INVX1 INVX1_51 ( .A(_abc_43815_n1126), .Y(_abc_43815_n1127) );
  INVX1 INVX1_510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2835_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2836_1) );
  INVX1 INVX1_511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2839_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2840) );
  INVX1 INVX1_512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2843), .Y(REGFILE_SIM_reg_bank__abc_33898_n2844_1) );
  INVX1 INVX1_513 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2847_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2848_1) );
  INVX1 INVX1_514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2851_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2852) );
  INVX1 INVX1_515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2855), .Y(REGFILE_SIM_reg_bank__abc_33898_n2856_1) );
  INVX1 INVX1_516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2859_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2860_1) );
  INVX1 INVX1_517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2863_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2864) );
  INVX1 INVX1_518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2867), .Y(REGFILE_SIM_reg_bank__abc_33898_n2868_1) );
  INVX1 INVX1_519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2871_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2872_1) );
  INVX1 INVX1_52 ( .A(alu_op_r_3_), .Y(_abc_43815_n1129) );
  INVX1 INVX1_520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2875_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2876) );
  INVX1 INVX1_521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2879_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2880) );
  INVX1 INVX1_522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2883), .Y(REGFILE_SIM_reg_bank__abc_33898_n2884_1) );
  INVX1 INVX1_523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2887_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2888_1) );
  INVX1 INVX1_524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2891_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2892) );
  INVX1 INVX1_525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2895), .Y(REGFILE_SIM_reg_bank__abc_33898_n2896_1) );
  INVX1 INVX1_526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2899_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2900_1) );
  INVX1 INVX1_527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2903_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2904) );
  INVX1 INVX1_528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2907), .Y(REGFILE_SIM_reg_bank__abc_33898_n2908_1) );
  INVX1 INVX1_529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2911_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2912_1) );
  INVX1 INVX1_53 ( .A(_abc_43815_n1134), .Y(_abc_43815_n1135_1) );
  INVX1 INVX1_530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2915_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2916) );
  INVX1 INVX1_531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2919), .Y(REGFILE_SIM_reg_bank__abc_33898_n2920_1) );
  INVX1 INVX1_532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2923_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2924_1) );
  INVX1 INVX1_533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2927_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2928) );
  INVX1 INVX1_534 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2931), .Y(REGFILE_SIM_reg_bank__abc_33898_n2932_1) );
  INVX1 INVX1_535 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2935_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2936_1) );
  INVX1 INVX1_536 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2939_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2940) );
  INVX1 INVX1_537 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2943), .Y(REGFILE_SIM_reg_bank__abc_33898_n2944_1) );
  INVX1 INVX1_538 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2947_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2948_1) );
  INVX1 INVX1_539 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2951_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2952) );
  INVX1 INVX1_54 ( .A(_abc_43815_n1106), .Y(_abc_43815_n1136_1) );
  INVX1 INVX1_540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2955), .Y(REGFILE_SIM_reg_bank__abc_33898_n2956_1) );
  INVX1 INVX1_541 ( .A(REGFILE_SIM_reg_bank_rd_i_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3056_1) );
  INVX1 INVX1_542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3160), .Y(REGFILE_SIM_reg_bank__abc_33898_n3161) );
  INVX1 INVX1_543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3164), .Y(REGFILE_SIM_reg_bank__abc_33898_n3165) );
  INVX1 INVX1_544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3168), .Y(REGFILE_SIM_reg_bank__abc_33898_n3169) );
  INVX1 INVX1_545 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3172), .Y(REGFILE_SIM_reg_bank__abc_33898_n3173) );
  INVX1 INVX1_546 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3176), .Y(REGFILE_SIM_reg_bank__abc_33898_n3177) );
  INVX1 INVX1_547 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3180), .Y(REGFILE_SIM_reg_bank__abc_33898_n3181) );
  INVX1 INVX1_548 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3184), .Y(REGFILE_SIM_reg_bank__abc_33898_n3185) );
  INVX1 INVX1_549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3188), .Y(REGFILE_SIM_reg_bank__abc_33898_n3189) );
  INVX1 INVX1_55 ( .A(_abc_43815_n1139), .Y(_abc_43815_n1140) );
  INVX1 INVX1_550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3192), .Y(REGFILE_SIM_reg_bank__abc_33898_n3193) );
  INVX1 INVX1_551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3196), .Y(REGFILE_SIM_reg_bank__abc_33898_n3197_1) );
  INVX1 INVX1_552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3200), .Y(REGFILE_SIM_reg_bank__abc_33898_n3201) );
  INVX1 INVX1_553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3204), .Y(REGFILE_SIM_reg_bank__abc_33898_n3205) );
  INVX1 INVX1_554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3208), .Y(REGFILE_SIM_reg_bank__abc_33898_n3209) );
  INVX1 INVX1_555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3212), .Y(REGFILE_SIM_reg_bank__abc_33898_n3213) );
  INVX1 INVX1_556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3216), .Y(REGFILE_SIM_reg_bank__abc_33898_n3217) );
  INVX1 INVX1_557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3220), .Y(REGFILE_SIM_reg_bank__abc_33898_n3221) );
  INVX1 INVX1_558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3224), .Y(REGFILE_SIM_reg_bank__abc_33898_n3225) );
  INVX1 INVX1_559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3228), .Y(REGFILE_SIM_reg_bank__abc_33898_n3229_1) );
  INVX1 INVX1_56 ( .A(_abc_43815_n1113), .Y(_abc_43815_n1144) );
  INVX1 INVX1_560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3232), .Y(REGFILE_SIM_reg_bank__abc_33898_n3233) );
  INVX1 INVX1_561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3236), .Y(REGFILE_SIM_reg_bank__abc_33898_n3237) );
  INVX1 INVX1_562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3240), .Y(REGFILE_SIM_reg_bank__abc_33898_n3241) );
  INVX1 INVX1_563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3244), .Y(REGFILE_SIM_reg_bank__abc_33898_n3245) );
  INVX1 INVX1_564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3248), .Y(REGFILE_SIM_reg_bank__abc_33898_n3249) );
  INVX1 INVX1_565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3252), .Y(REGFILE_SIM_reg_bank__abc_33898_n3253) );
  INVX1 INVX1_566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3256), .Y(REGFILE_SIM_reg_bank__abc_33898_n3257) );
  INVX1 INVX1_567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3260), .Y(REGFILE_SIM_reg_bank__abc_33898_n3261_1) );
  INVX1 INVX1_568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3264), .Y(REGFILE_SIM_reg_bank__abc_33898_n3265) );
  INVX1 INVX1_569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3268), .Y(REGFILE_SIM_reg_bank__abc_33898_n3269) );
  INVX1 INVX1_57 ( .A(_abc_43815_n1130), .Y(_abc_43815_n1145) );
  INVX1 INVX1_570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3272), .Y(REGFILE_SIM_reg_bank__abc_33898_n3273) );
  INVX1 INVX1_571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3276), .Y(REGFILE_SIM_reg_bank__abc_33898_n3277) );
  INVX1 INVX1_572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3280), .Y(REGFILE_SIM_reg_bank__abc_33898_n3281) );
  INVX1 INVX1_573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3284), .Y(REGFILE_SIM_reg_bank__abc_33898_n3285) );
  INVX1 INVX1_574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3290), .Y(REGFILE_SIM_reg_bank__abc_33898_n3291) );
  INVX1 INVX1_575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3294), .Y(REGFILE_SIM_reg_bank__abc_33898_n3295) );
  INVX1 INVX1_576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3298), .Y(REGFILE_SIM_reg_bank__abc_33898_n3299) );
  INVX1 INVX1_577 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3302), .Y(REGFILE_SIM_reg_bank__abc_33898_n3303) );
  INVX1 INVX1_578 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3306), .Y(REGFILE_SIM_reg_bank__abc_33898_n3307) );
  INVX1 INVX1_579 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3310), .Y(REGFILE_SIM_reg_bank__abc_33898_n3311) );
  INVX1 INVX1_58 ( .A(_abc_43815_n1118), .Y(_abc_43815_n1146) );
  INVX1 INVX1_580 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3314), .Y(REGFILE_SIM_reg_bank__abc_33898_n3315) );
  INVX1 INVX1_581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3318), .Y(REGFILE_SIM_reg_bank__abc_33898_n3319) );
  INVX1 INVX1_582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3322), .Y(REGFILE_SIM_reg_bank__abc_33898_n3323) );
  INVX1 INVX1_583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3326), .Y(REGFILE_SIM_reg_bank__abc_33898_n3327) );
  INVX1 INVX1_584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3330), .Y(REGFILE_SIM_reg_bank__abc_33898_n3331) );
  INVX1 INVX1_585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3334), .Y(REGFILE_SIM_reg_bank__abc_33898_n3335) );
  INVX1 INVX1_586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3338), .Y(REGFILE_SIM_reg_bank__abc_33898_n3339) );
  INVX1 INVX1_587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3342), .Y(REGFILE_SIM_reg_bank__abc_33898_n3343) );
  INVX1 INVX1_588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3346), .Y(REGFILE_SIM_reg_bank__abc_33898_n3347) );
  INVX1 INVX1_589 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3350), .Y(REGFILE_SIM_reg_bank__abc_33898_n3351) );
  INVX1 INVX1_59 ( .A(_abc_43815_n1153_1), .Y(_abc_43815_n1154) );
  INVX1 INVX1_590 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3354), .Y(REGFILE_SIM_reg_bank__abc_33898_n3355) );
  INVX1 INVX1_591 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3358), .Y(REGFILE_SIM_reg_bank__abc_33898_n3359) );
  INVX1 INVX1_592 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3362), .Y(REGFILE_SIM_reg_bank__abc_33898_n3363) );
  INVX1 INVX1_593 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3366), .Y(REGFILE_SIM_reg_bank__abc_33898_n3367) );
  INVX1 INVX1_594 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3370), .Y(REGFILE_SIM_reg_bank__abc_33898_n3371) );
  INVX1 INVX1_595 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3374), .Y(REGFILE_SIM_reg_bank__abc_33898_n3375) );
  INVX1 INVX1_596 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3378), .Y(REGFILE_SIM_reg_bank__abc_33898_n3379) );
  INVX1 INVX1_597 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3382), .Y(REGFILE_SIM_reg_bank__abc_33898_n3383) );
  INVX1 INVX1_598 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3386), .Y(REGFILE_SIM_reg_bank__abc_33898_n3387) );
  INVX1 INVX1_599 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3390), .Y(REGFILE_SIM_reg_bank__abc_33898_n3391) );
  INVX1 INVX1_6 ( .A(inst_r_0_), .Y(_abc_43815_n630) );
  INVX1 INVX1_60 ( .A(_abc_43815_n1159), .Y(_abc_43815_n1160) );
  INVX1 INVX1_600 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3394), .Y(REGFILE_SIM_reg_bank__abc_33898_n3395) );
  INVX1 INVX1_601 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3398), .Y(REGFILE_SIM_reg_bank__abc_33898_n3399) );
  INVX1 INVX1_602 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3402), .Y(REGFILE_SIM_reg_bank__abc_33898_n3403) );
  INVX1 INVX1_603 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3406), .Y(REGFILE_SIM_reg_bank__abc_33898_n3407) );
  INVX1 INVX1_604 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3410), .Y(REGFILE_SIM_reg_bank__abc_33898_n3411) );
  INVX1 INVX1_605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3414), .Y(REGFILE_SIM_reg_bank__abc_33898_n3415) );
  INVX1 INVX1_606 ( .A(REGFILE_SIM_reg_bank_rd_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3911) );
  INVX1 INVX1_607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3915), .Y(REGFILE_SIM_reg_bank__abc_33898_n3916) );
  INVX1 INVX1_608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3919), .Y(REGFILE_SIM_reg_bank__abc_33898_n3920) );
  INVX1 INVX1_609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3923), .Y(REGFILE_SIM_reg_bank__abc_33898_n3924) );
  INVX1 INVX1_61 ( .A(_abc_43815_n1164), .Y(_abc_43815_n1165) );
  INVX1 INVX1_610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3927), .Y(REGFILE_SIM_reg_bank__abc_33898_n3928) );
  INVX1 INVX1_611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3931), .Y(REGFILE_SIM_reg_bank__abc_33898_n3932) );
  INVX1 INVX1_612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3935), .Y(REGFILE_SIM_reg_bank__abc_33898_n3936) );
  INVX1 INVX1_613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3939), .Y(REGFILE_SIM_reg_bank__abc_33898_n3940) );
  INVX1 INVX1_614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3943), .Y(REGFILE_SIM_reg_bank__abc_33898_n3944) );
  INVX1 INVX1_615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3947), .Y(REGFILE_SIM_reg_bank__abc_33898_n3948) );
  INVX1 INVX1_616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3951), .Y(REGFILE_SIM_reg_bank__abc_33898_n3952) );
  INVX1 INVX1_617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3955), .Y(REGFILE_SIM_reg_bank__abc_33898_n3956) );
  INVX1 INVX1_618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3959), .Y(REGFILE_SIM_reg_bank__abc_33898_n3960) );
  INVX1 INVX1_619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3963), .Y(REGFILE_SIM_reg_bank__abc_33898_n3964) );
  INVX1 INVX1_62 ( .A(_abc_43815_n1177), .Y(_abc_43815_n1178_1) );
  INVX1 INVX1_620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3967), .Y(REGFILE_SIM_reg_bank__abc_33898_n3968) );
  INVX1 INVX1_621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3971), .Y(REGFILE_SIM_reg_bank__abc_33898_n3972) );
  INVX1 INVX1_622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3975), .Y(REGFILE_SIM_reg_bank__abc_33898_n3976) );
  INVX1 INVX1_623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3979), .Y(REGFILE_SIM_reg_bank__abc_33898_n3980) );
  INVX1 INVX1_624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3983), .Y(REGFILE_SIM_reg_bank__abc_33898_n3984) );
  INVX1 INVX1_625 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3987), .Y(REGFILE_SIM_reg_bank__abc_33898_n3988) );
  INVX1 INVX1_626 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3991), .Y(REGFILE_SIM_reg_bank__abc_33898_n3992) );
  INVX1 INVX1_627 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3995), .Y(REGFILE_SIM_reg_bank__abc_33898_n3996) );
  INVX1 INVX1_628 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3999), .Y(REGFILE_SIM_reg_bank__abc_33898_n4000) );
  INVX1 INVX1_629 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4003), .Y(REGFILE_SIM_reg_bank__abc_33898_n4004) );
  INVX1 INVX1_63 ( .A(_abc_43815_n1180), .Y(_abc_43815_n1181) );
  INVX1 INVX1_630 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4007), .Y(REGFILE_SIM_reg_bank__abc_33898_n4008) );
  INVX1 INVX1_631 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4011), .Y(REGFILE_SIM_reg_bank__abc_33898_n4012) );
  INVX1 INVX1_632 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4015), .Y(REGFILE_SIM_reg_bank__abc_33898_n4016) );
  INVX1 INVX1_633 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4019), .Y(REGFILE_SIM_reg_bank__abc_33898_n4020) );
  INVX1 INVX1_634 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4023), .Y(REGFILE_SIM_reg_bank__abc_33898_n4024) );
  INVX1 INVX1_635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4027), .Y(REGFILE_SIM_reg_bank__abc_33898_n4028) );
  INVX1 INVX1_636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4031), .Y(REGFILE_SIM_reg_bank__abc_33898_n4032) );
  INVX1 INVX1_637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4035), .Y(REGFILE_SIM_reg_bank__abc_33898_n4036) );
  INVX1 INVX1_638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4039), .Y(REGFILE_SIM_reg_bank__abc_33898_n4040) );
  INVX1 INVX1_639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4437), .Y(REGFILE_SIM_reg_bank__abc_33898_n4438) );
  INVX1 INVX1_64 ( .A(_abc_43815_n1185), .Y(_abc_43815_n1186_1) );
  INVX1 INVX1_640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4441), .Y(REGFILE_SIM_reg_bank__abc_33898_n4442) );
  INVX1 INVX1_641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4445), .Y(REGFILE_SIM_reg_bank__abc_33898_n4446) );
  INVX1 INVX1_642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4449), .Y(REGFILE_SIM_reg_bank__abc_33898_n4450) );
  INVX1 INVX1_643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4453), .Y(REGFILE_SIM_reg_bank__abc_33898_n4454) );
  INVX1 INVX1_644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4457), .Y(REGFILE_SIM_reg_bank__abc_33898_n4458) );
  INVX1 INVX1_645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4461), .Y(REGFILE_SIM_reg_bank__abc_33898_n4462) );
  INVX1 INVX1_646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4465), .Y(REGFILE_SIM_reg_bank__abc_33898_n4466) );
  INVX1 INVX1_647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4469), .Y(REGFILE_SIM_reg_bank__abc_33898_n4470) );
  INVX1 INVX1_648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4473), .Y(REGFILE_SIM_reg_bank__abc_33898_n4474) );
  INVX1 INVX1_649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4477), .Y(REGFILE_SIM_reg_bank__abc_33898_n4478) );
  INVX1 INVX1_65 ( .A(_abc_43815_n1192), .Y(_abc_43815_n1193) );
  INVX1 INVX1_650 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4481), .Y(REGFILE_SIM_reg_bank__abc_33898_n4482) );
  INVX1 INVX1_651 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4485), .Y(REGFILE_SIM_reg_bank__abc_33898_n4486) );
  INVX1 INVX1_652 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4489), .Y(REGFILE_SIM_reg_bank__abc_33898_n4490) );
  INVX1 INVX1_653 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4493_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4494) );
  INVX1 INVX1_654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4497), .Y(REGFILE_SIM_reg_bank__abc_33898_n4498) );
  INVX1 INVX1_655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4501), .Y(REGFILE_SIM_reg_bank__abc_33898_n4502) );
  INVX1 INVX1_656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4505), .Y(REGFILE_SIM_reg_bank__abc_33898_n4506) );
  INVX1 INVX1_657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4509), .Y(REGFILE_SIM_reg_bank__abc_33898_n4510) );
  INVX1 INVX1_658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4513), .Y(REGFILE_SIM_reg_bank__abc_33898_n4514) );
  INVX1 INVX1_659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4517), .Y(REGFILE_SIM_reg_bank__abc_33898_n4518) );
  INVX1 INVX1_66 ( .A(_abc_43815_n1195), .Y(_abc_43815_n1196) );
  INVX1 INVX1_660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4521), .Y(REGFILE_SIM_reg_bank__abc_33898_n4522) );
  INVX1 INVX1_661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4525), .Y(REGFILE_SIM_reg_bank__abc_33898_n4526) );
  INVX1 INVX1_662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4529), .Y(REGFILE_SIM_reg_bank__abc_33898_n4530) );
  INVX1 INVX1_663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4533), .Y(REGFILE_SIM_reg_bank__abc_33898_n4534) );
  INVX1 INVX1_664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4537), .Y(REGFILE_SIM_reg_bank__abc_33898_n4538) );
  INVX1 INVX1_665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4541), .Y(REGFILE_SIM_reg_bank__abc_33898_n4542) );
  INVX1 INVX1_666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4545), .Y(REGFILE_SIM_reg_bank__abc_33898_n4546) );
  INVX1 INVX1_667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4549), .Y(REGFILE_SIM_reg_bank__abc_33898_n4550) );
  INVX1 INVX1_668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4553_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4554) );
  INVX1 INVX1_669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4557), .Y(REGFILE_SIM_reg_bank__abc_33898_n4558) );
  INVX1 INVX1_67 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_8_), .Y(_abc_43815_n1198) );
  INVX1 INVX1_670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4561), .Y(REGFILE_SIM_reg_bank__abc_33898_n4562) );
  INVX1 INVX1_671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4566), .Y(REGFILE_SIM_reg_bank__abc_33898_n4567) );
  INVX1 INVX1_672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4570), .Y(REGFILE_SIM_reg_bank__abc_33898_n4571) );
  INVX1 INVX1_673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4574), .Y(REGFILE_SIM_reg_bank__abc_33898_n4575) );
  INVX1 INVX1_674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4578), .Y(REGFILE_SIM_reg_bank__abc_33898_n4579) );
  INVX1 INVX1_675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4582), .Y(REGFILE_SIM_reg_bank__abc_33898_n4583_1) );
  INVX1 INVX1_676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4586), .Y(REGFILE_SIM_reg_bank__abc_33898_n4587) );
  INVX1 INVX1_677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4590), .Y(REGFILE_SIM_reg_bank__abc_33898_n4591) );
  INVX1 INVX1_678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4594), .Y(REGFILE_SIM_reg_bank__abc_33898_n4595) );
  INVX1 INVX1_679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4598), .Y(REGFILE_SIM_reg_bank__abc_33898_n4599) );
  INVX1 INVX1_68 ( .A(int32_r_10_), .Y(_abc_43815_n1199) );
  INVX1 INVX1_680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4602), .Y(REGFILE_SIM_reg_bank__abc_33898_n4603) );
  INVX1 INVX1_681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4606), .Y(REGFILE_SIM_reg_bank__abc_33898_n4607) );
  INVX1 INVX1_682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4610), .Y(REGFILE_SIM_reg_bank__abc_33898_n4611) );
  INVX1 INVX1_683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4614), .Y(REGFILE_SIM_reg_bank__abc_33898_n4615) );
  INVX1 INVX1_684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4618), .Y(REGFILE_SIM_reg_bank__abc_33898_n4619) );
  INVX1 INVX1_685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4622), .Y(REGFILE_SIM_reg_bank__abc_33898_n4623) );
  INVX1 INVX1_686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4626), .Y(REGFILE_SIM_reg_bank__abc_33898_n4627) );
  INVX1 INVX1_687 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4630), .Y(REGFILE_SIM_reg_bank__abc_33898_n4631) );
  INVX1 INVX1_688 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4634), .Y(REGFILE_SIM_reg_bank__abc_33898_n4635) );
  INVX1 INVX1_689 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4638), .Y(REGFILE_SIM_reg_bank__abc_33898_n4639) );
  INVX1 INVX1_69 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_10_), .Y(_abc_43815_n1201) );
  INVX1 INVX1_690 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4642), .Y(REGFILE_SIM_reg_bank__abc_33898_n4643_1) );
  INVX1 INVX1_691 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4646), .Y(REGFILE_SIM_reg_bank__abc_33898_n4647) );
  INVX1 INVX1_692 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4650), .Y(REGFILE_SIM_reg_bank__abc_33898_n4651) );
  INVX1 INVX1_693 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4654), .Y(REGFILE_SIM_reg_bank__abc_33898_n4655) );
  INVX1 INVX1_694 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4658), .Y(REGFILE_SIM_reg_bank__abc_33898_n4659) );
  INVX1 INVX1_695 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4662), .Y(REGFILE_SIM_reg_bank__abc_33898_n4663) );
  INVX1 INVX1_696 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4666), .Y(REGFILE_SIM_reg_bank__abc_33898_n4667) );
  INVX1 INVX1_697 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4670), .Y(REGFILE_SIM_reg_bank__abc_33898_n4671) );
  INVX1 INVX1_698 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4674), .Y(REGFILE_SIM_reg_bank__abc_33898_n4675) );
  INVX1 INVX1_699 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4678), .Y(REGFILE_SIM_reg_bank__abc_33898_n4679) );
  INVX1 INVX1_7 ( .A(enable_i_bF_buf6), .Y(_abc_43815_n634) );
  INVX1 INVX1_70 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_43815_n1204) );
  INVX1 INVX1_700 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4682), .Y(REGFILE_SIM_reg_bank__abc_33898_n4683) );
  INVX1 INVX1_701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4686), .Y(REGFILE_SIM_reg_bank__abc_33898_n4687) );
  INVX1 INVX1_702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4690), .Y(REGFILE_SIM_reg_bank__abc_33898_n4691) );
  INVX1 INVX1_703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4891), .Y(REGFILE_SIM_reg_bank__abc_33898_n4892) );
  INVX1 INVX1_704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4895), .Y(REGFILE_SIM_reg_bank__abc_33898_n4896) );
  INVX1 INVX1_705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4899), .Y(REGFILE_SIM_reg_bank__abc_33898_n4900) );
  INVX1 INVX1_706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4903), .Y(REGFILE_SIM_reg_bank__abc_33898_n4904) );
  INVX1 INVX1_707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4907), .Y(REGFILE_SIM_reg_bank__abc_33898_n4908) );
  INVX1 INVX1_708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4911), .Y(REGFILE_SIM_reg_bank__abc_33898_n4912) );
  INVX1 INVX1_709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4915), .Y(REGFILE_SIM_reg_bank__abc_33898_n4916) );
  INVX1 INVX1_71 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_43815_n1205_1) );
  INVX1 INVX1_710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4919), .Y(REGFILE_SIM_reg_bank__abc_33898_n4920) );
  INVX1 INVX1_711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4923), .Y(REGFILE_SIM_reg_bank__abc_33898_n4924) );
  INVX1 INVX1_712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4927), .Y(REGFILE_SIM_reg_bank__abc_33898_n4928) );
  INVX1 INVX1_713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4931), .Y(REGFILE_SIM_reg_bank__abc_33898_n4932) );
  INVX1 INVX1_714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4935), .Y(REGFILE_SIM_reg_bank__abc_33898_n4936) );
  INVX1 INVX1_715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4939), .Y(REGFILE_SIM_reg_bank__abc_33898_n4940) );
  INVX1 INVX1_716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4943_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4944) );
  INVX1 INVX1_717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4947), .Y(REGFILE_SIM_reg_bank__abc_33898_n4948) );
  INVX1 INVX1_718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4951), .Y(REGFILE_SIM_reg_bank__abc_33898_n4952) );
  INVX1 INVX1_719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4955), .Y(REGFILE_SIM_reg_bank__abc_33898_n4956) );
  INVX1 INVX1_72 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_43815_n1206_1) );
  INVX1 INVX1_720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4959), .Y(REGFILE_SIM_reg_bank__abc_33898_n4960) );
  INVX1 INVX1_721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4963), .Y(REGFILE_SIM_reg_bank__abc_33898_n4964) );
  INVX1 INVX1_722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4967), .Y(REGFILE_SIM_reg_bank__abc_33898_n4968) );
  INVX1 INVX1_723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4971), .Y(REGFILE_SIM_reg_bank__abc_33898_n4972) );
  INVX1 INVX1_724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4975), .Y(REGFILE_SIM_reg_bank__abc_33898_n4976) );
  INVX1 INVX1_725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4979), .Y(REGFILE_SIM_reg_bank__abc_33898_n4980) );
  INVX1 INVX1_726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4983), .Y(REGFILE_SIM_reg_bank__abc_33898_n4984) );
  INVX1 INVX1_727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4987), .Y(REGFILE_SIM_reg_bank__abc_33898_n4988) );
  INVX1 INVX1_728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4991), .Y(REGFILE_SIM_reg_bank__abc_33898_n4992) );
  INVX1 INVX1_729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4995), .Y(REGFILE_SIM_reg_bank__abc_33898_n4996) );
  INVX1 INVX1_73 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_43815_n1209) );
  INVX1 INVX1_730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4999), .Y(REGFILE_SIM_reg_bank__abc_33898_n5000) );
  INVX1 INVX1_731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5003_1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5004) );
  INVX1 INVX1_732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5007), .Y(REGFILE_SIM_reg_bank__abc_33898_n5008) );
  INVX1 INVX1_733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5011), .Y(REGFILE_SIM_reg_bank__abc_33898_n5012) );
  INVX1 INVX1_734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5015), .Y(REGFILE_SIM_reg_bank__abc_33898_n5016) );
  INVX1 INVX1_735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5020), .Y(REGFILE_SIM_reg_bank__abc_33898_n5021) );
  INVX1 INVX1_736 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5024), .Y(REGFILE_SIM_reg_bank__abc_33898_n5025) );
  INVX1 INVX1_737 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5028), .Y(REGFILE_SIM_reg_bank__abc_33898_n5029) );
  INVX1 INVX1_738 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5032), .Y(REGFILE_SIM_reg_bank__abc_33898_n5033_1) );
  INVX1 INVX1_739 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5036), .Y(REGFILE_SIM_reg_bank__abc_33898_n5037) );
  INVX1 INVX1_74 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_43815_n1210) );
  INVX1 INVX1_740 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5040), .Y(REGFILE_SIM_reg_bank__abc_33898_n5041) );
  INVX1 INVX1_741 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5044), .Y(REGFILE_SIM_reg_bank__abc_33898_n5045) );
  INVX1 INVX1_742 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5048), .Y(REGFILE_SIM_reg_bank__abc_33898_n5049) );
  INVX1 INVX1_743 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5052), .Y(REGFILE_SIM_reg_bank__abc_33898_n5053) );
  INVX1 INVX1_744 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5056), .Y(REGFILE_SIM_reg_bank__abc_33898_n5057) );
  INVX1 INVX1_745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5060), .Y(REGFILE_SIM_reg_bank__abc_33898_n5061) );
  INVX1 INVX1_746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5064), .Y(REGFILE_SIM_reg_bank__abc_33898_n5065) );
  INVX1 INVX1_747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5068), .Y(REGFILE_SIM_reg_bank__abc_33898_n5069) );
  INVX1 INVX1_748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5072), .Y(REGFILE_SIM_reg_bank__abc_33898_n5073) );
  INVX1 INVX1_749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5076), .Y(REGFILE_SIM_reg_bank__abc_33898_n5077) );
  INVX1 INVX1_75 ( .A(_abc_43815_n1212), .Y(_abc_43815_n1213) );
  INVX1 INVX1_750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5080), .Y(REGFILE_SIM_reg_bank__abc_33898_n5081) );
  INVX1 INVX1_751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5084), .Y(REGFILE_SIM_reg_bank__abc_33898_n5085) );
  INVX1 INVX1_752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5088), .Y(REGFILE_SIM_reg_bank__abc_33898_n5089) );
  INVX1 INVX1_753 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5092), .Y(REGFILE_SIM_reg_bank__abc_33898_n5093_1) );
  INVX1 INVX1_754 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5096), .Y(REGFILE_SIM_reg_bank__abc_33898_n5097) );
  INVX1 INVX1_755 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5100), .Y(REGFILE_SIM_reg_bank__abc_33898_n5101) );
  INVX1 INVX1_756 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5104), .Y(REGFILE_SIM_reg_bank__abc_33898_n5105) );
  INVX1 INVX1_757 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5108), .Y(REGFILE_SIM_reg_bank__abc_33898_n5109) );
  INVX1 INVX1_758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5112), .Y(REGFILE_SIM_reg_bank__abc_33898_n5113) );
  INVX1 INVX1_759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5116), .Y(REGFILE_SIM_reg_bank__abc_33898_n5117) );
  INVX1 INVX1_76 ( .A(_abc_43815_n1217), .Y(_abc_43815_n1218) );
  INVX1 INVX1_760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5120), .Y(REGFILE_SIM_reg_bank__abc_33898_n5121) );
  INVX1 INVX1_761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5124), .Y(REGFILE_SIM_reg_bank__abc_33898_n5125) );
  INVX1 INVX1_762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5128), .Y(REGFILE_SIM_reg_bank__abc_33898_n5129) );
  INVX1 INVX1_763 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5132), .Y(REGFILE_SIM_reg_bank__abc_33898_n5133) );
  INVX1 INVX1_764 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5136), .Y(REGFILE_SIM_reg_bank__abc_33898_n5137) );
  INVX1 INVX1_765 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5140), .Y(REGFILE_SIM_reg_bank__abc_33898_n5141) );
  INVX1 INVX1_766 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5144), .Y(REGFILE_SIM_reg_bank__abc_33898_n5145) );
  INVX1 INVX1_767 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5540) );
  INVX1 INVX1_768 ( .A(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5543) );
  INVX1 INVX1_769 ( .A(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5551) );
  INVX1 INVX1_77 ( .A(_abc_43815_n1219), .Y(_abc_43815_n1220) );
  INVX1 INVX1_770 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5561) );
  INVX1 INVX1_771 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7549) );
  INVX1 INVX1_772 ( .A(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7552) );
  INVX1 INVX1_773 ( .A(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7560) );
  INVX1 INVX1_774 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7570) );
  INVX1 INVX1_775 ( .A(alu__abc_41358_n110), .Y(alu__abc_41358_n111) );
  INVX1 INVX1_776 ( .A(alu_b_i_25_), .Y(alu__abc_41358_n112_1) );
  INVX1 INVX1_777 ( .A(alu_a_i_25_), .Y(alu__abc_41358_n113_1) );
  INVX1 INVX1_778 ( .A(alu__abc_41358_n114), .Y(alu__abc_41358_n115) );
  INVX1 INVX1_779 ( .A(alu__abc_41358_n116), .Y(alu__abc_41358_n117) );
  INVX1 INVX1_78 ( .A(_abc_43815_n1222), .Y(_abc_43815_n1223) );
  INVX1 INVX1_780 ( .A(alu__abc_41358_n118), .Y(alu__abc_41358_n119_1) );
  INVX1 INVX1_781 ( .A(alu_b_i_24_), .Y(alu__abc_41358_n120_1) );
  INVX1 INVX1_782 ( .A(alu_a_i_24_), .Y(alu__abc_41358_n121) );
  INVX1 INVX1_783 ( .A(alu__abc_41358_n122), .Y(alu__abc_41358_n123) );
  INVX1 INVX1_784 ( .A(alu__abc_41358_n124_1), .Y(alu__abc_41358_n125_1) );
  INVX1 INVX1_785 ( .A(alu__abc_41358_n127), .Y(alu__abc_41358_n128) );
  INVX1 INVX1_786 ( .A(alu_b_i_26_), .Y(alu__abc_41358_n129) );
  INVX1 INVX1_787 ( .A(alu_a_i_26_), .Y(alu__abc_41358_n130_1) );
  INVX1 INVX1_788 ( .A(alu__abc_41358_n131_1), .Y(alu__abc_41358_n132) );
  INVX1 INVX1_789 ( .A(alu__abc_41358_n133), .Y(alu__abc_41358_n134) );
  INVX1 INVX1_79 ( .A(_abc_43815_n1224), .Y(_abc_43815_n1225) );
  INVX1 INVX1_790 ( .A(alu__abc_41358_n135_1), .Y(alu__abc_41358_n136_1) );
  INVX1 INVX1_791 ( .A(alu_b_i_27_), .Y(alu__abc_41358_n137) );
  INVX1 INVX1_792 ( .A(alu_a_i_27_), .Y(alu__abc_41358_n138) );
  INVX1 INVX1_793 ( .A(alu__abc_41358_n139), .Y(alu__abc_41358_n140) );
  INVX1 INVX1_794 ( .A(alu__abc_41358_n145), .Y(alu__abc_41358_n146) );
  INVX1 INVX1_795 ( .A(alu_b_i_28_), .Y(alu__abc_41358_n147) );
  INVX1 INVX1_796 ( .A(alu_a_i_28_), .Y(alu__abc_41358_n148_1) );
  INVX1 INVX1_797 ( .A(alu__abc_41358_n149_1), .Y(alu__abc_41358_n150) );
  INVX1 INVX1_798 ( .A(alu__abc_41358_n151), .Y(alu__abc_41358_n152) );
  INVX1 INVX1_799 ( .A(alu__abc_41358_n153), .Y(alu__abc_41358_n154_1) );
  INVX1 INVX1_8 ( .A(inst_r_3_), .Y(_abc_43815_n637) );
  INVX1 INVX1_80 ( .A(_abc_43815_n1228), .Y(_abc_43815_n1229) );
  INVX1 INVX1_800 ( .A(alu_b_i_29_), .Y(alu__abc_41358_n155_1) );
  INVX1 INVX1_801 ( .A(alu_a_i_29_), .Y(alu__abc_41358_n156) );
  INVX1 INVX1_802 ( .A(alu__abc_41358_n157), .Y(alu__abc_41358_n158) );
  INVX1 INVX1_803 ( .A(alu__abc_41358_n159_1), .Y(alu__abc_41358_n160_1) );
  INVX1 INVX1_804 ( .A(alu__abc_41358_n162), .Y(alu__abc_41358_n163) );
  INVX1 INVX1_805 ( .A(alu_b_i_30_), .Y(alu__abc_41358_n164) );
  INVX1 INVX1_806 ( .A(alu_a_i_30_), .Y(alu__abc_41358_n165) );
  INVX1 INVX1_807 ( .A(alu__abc_41358_n166_1), .Y(alu__abc_41358_n167_1) );
  INVX1 INVX1_808 ( .A(alu__abc_41358_n168), .Y(alu__abc_41358_n169) );
  INVX1 INVX1_809 ( .A(alu_b_i_31_), .Y(alu__abc_41358_n171_1) );
  INVX1 INVX1_81 ( .A(_abc_43815_n1230_1), .Y(_abc_43815_n1231) );
  INVX1 INVX1_810 ( .A(alu_a_i_31_), .Y(alu__abc_41358_n172_1) );
  INVX1 INVX1_811 ( .A(alu__abc_41358_n178_1), .Y(alu__abc_41358_n179) );
  INVX1 INVX1_812 ( .A(alu_b_i_22_), .Y(alu__abc_41358_n180) );
  INVX1 INVX1_813 ( .A(alu_a_i_22_), .Y(alu__abc_41358_n181) );
  INVX1 INVX1_814 ( .A(alu__abc_41358_n182_1), .Y(alu__abc_41358_n183_1) );
  INVX1 INVX1_815 ( .A(alu__abc_41358_n184), .Y(alu__abc_41358_n185) );
  INVX1 INVX1_816 ( .A(alu__abc_41358_n186), .Y(alu__abc_41358_n187) );
  INVX1 INVX1_817 ( .A(alu_b_i_23_), .Y(alu__abc_41358_n188) );
  INVX1 INVX1_818 ( .A(alu_a_i_23_), .Y(alu__abc_41358_n189) );
  INVX1 INVX1_819 ( .A(alu__abc_41358_n190), .Y(alu__abc_41358_n191_1) );
  INVX1 INVX1_82 ( .A(_abc_43815_n1234), .Y(_abc_43815_n1235) );
  INVX1 INVX1_820 ( .A(alu__abc_41358_n195), .Y(alu__abc_41358_n196_1) );
  INVX1 INVX1_821 ( .A(alu_b_i_20_), .Y(alu__abc_41358_n197) );
  INVX1 INVX1_822 ( .A(alu_a_i_20_), .Y(alu__abc_41358_n198_1) );
  INVX1 INVX1_823 ( .A(alu__abc_41358_n199), .Y(alu__abc_41358_n200) );
  INVX1 INVX1_824 ( .A(alu__abc_41358_n201), .Y(alu__abc_41358_n202) );
  INVX1 INVX1_825 ( .A(alu__abc_41358_n203_1), .Y(alu__abc_41358_n204) );
  INVX1 INVX1_826 ( .A(alu_b_i_21_), .Y(alu__abc_41358_n205) );
  INVX1 INVX1_827 ( .A(alu_a_i_21_), .Y(alu__abc_41358_n206_1) );
  INVX1 INVX1_828 ( .A(alu__abc_41358_n207), .Y(alu__abc_41358_n208) );
  INVX1 INVX1_829 ( .A(alu__abc_41358_n209), .Y(alu__abc_41358_n210) );
  INVX1 INVX1_83 ( .A(_abc_43815_n1240), .Y(_abc_43815_n1241) );
  INVX1 INVX1_830 ( .A(alu__abc_41358_n213), .Y(alu__abc_41358_n214) );
  INVX1 INVX1_831 ( .A(alu_b_i_18_), .Y(alu__abc_41358_n215) );
  INVX1 INVX1_832 ( .A(alu_a_i_18_), .Y(alu__abc_41358_n216) );
  INVX1 INVX1_833 ( .A(alu__abc_41358_n217), .Y(alu__abc_41358_n218) );
  INVX1 INVX1_834 ( .A(alu__abc_41358_n219), .Y(alu__abc_41358_n220) );
  INVX1 INVX1_835 ( .A(alu__abc_41358_n221), .Y(alu__abc_41358_n222) );
  INVX1 INVX1_836 ( .A(alu_b_i_19_), .Y(alu__abc_41358_n223) );
  INVX1 INVX1_837 ( .A(alu_a_i_19_), .Y(alu__abc_41358_n224) );
  INVX1 INVX1_838 ( .A(alu__abc_41358_n225), .Y(alu__abc_41358_n226) );
  INVX1 INVX1_839 ( .A(alu__abc_41358_n230), .Y(alu__abc_41358_n231) );
  INVX1 INVX1_84 ( .A(_abc_43815_n1246), .Y(_abc_43815_n1247) );
  INVX1 INVX1_840 ( .A(alu_b_i_16_), .Y(alu__abc_41358_n232) );
  INVX1 INVX1_841 ( .A(alu_a_i_16_), .Y(alu__abc_41358_n233) );
  INVX1 INVX1_842 ( .A(alu__abc_41358_n234), .Y(alu__abc_41358_n235) );
  INVX1 INVX1_843 ( .A(alu__abc_41358_n236), .Y(alu__abc_41358_n237) );
  INVX1 INVX1_844 ( .A(alu__abc_41358_n238), .Y(alu__abc_41358_n239) );
  INVX1 INVX1_845 ( .A(alu_b_i_17_), .Y(alu__abc_41358_n240) );
  INVX1 INVX1_846 ( .A(alu_a_i_17_), .Y(alu__abc_41358_n241) );
  INVX1 INVX1_847 ( .A(alu__abc_41358_n242), .Y(alu__abc_41358_n243) );
  INVX1 INVX1_848 ( .A(alu__abc_41358_n244), .Y(alu__abc_41358_n245) );
  INVX1 INVX1_849 ( .A(alu_a_i_1_), .Y(alu__abc_41358_n251) );
  INVX1 INVX1_85 ( .A(_abc_43815_n1221), .Y(_abc_43815_n1248) );
  INVX1 INVX1_850 ( .A(alu_a_i_0_), .Y(alu__abc_41358_n255) );
  INVX1 INVX1_851 ( .A(alu__abc_41358_n256), .Y(alu__abc_41358_n257) );
  INVX1 INVX1_852 ( .A(alu__abc_41358_n260), .Y(alu__abc_41358_n261) );
  INVX1 INVX1_853 ( .A(alu__abc_41358_n263), .Y(alu__abc_41358_n264) );
  INVX1 INVX1_854 ( .A(alu_b_i_6_), .Y(alu__abc_41358_n265) );
  INVX1 INVX1_855 ( .A(alu_a_i_6_), .Y(alu__abc_41358_n266) );
  INVX1 INVX1_856 ( .A(alu__abc_41358_n267), .Y(alu__abc_41358_n268) );
  INVX1 INVX1_857 ( .A(alu__abc_41358_n269), .Y(alu__abc_41358_n270) );
  INVX1 INVX1_858 ( .A(alu_b_i_7_), .Y(alu__abc_41358_n272) );
  INVX1 INVX1_859 ( .A(alu_a_i_7_), .Y(alu__abc_41358_n273) );
  INVX1 INVX1_86 ( .A(_abc_43815_n1216), .Y(_abc_43815_n1250_1) );
  INVX1 INVX1_860 ( .A(alu__abc_41358_n277), .Y(alu__abc_41358_n278) );
  INVX1 INVX1_861 ( .A(alu_a_i_4_), .Y(alu__abc_41358_n280) );
  INVX1 INVX1_862 ( .A(alu__abc_41358_n281), .Y(alu__abc_41358_n282) );
  INVX1 INVX1_863 ( .A(alu__abc_41358_n283), .Y(alu__abc_41358_n284) );
  INVX1 INVX1_864 ( .A(alu_b_i_5_), .Y(alu__abc_41358_n286) );
  INVX1 INVX1_865 ( .A(alu_a_i_5_), .Y(alu__abc_41358_n287) );
  INVX1 INVX1_866 ( .A(alu_a_i_3_), .Y(alu__abc_41358_n293) );
  INVX1 INVX1_867 ( .A(alu_a_i_2_), .Y(alu__abc_41358_n298) );
  INVX1 INVX1_868 ( .A(alu__abc_41358_n305), .Y(alu__abc_41358_n306) );
  INVX1 INVX1_869 ( .A(alu_b_i_12_), .Y(alu__abc_41358_n307) );
  INVX1 INVX1_87 ( .A(_abc_43815_n1233_1), .Y(_abc_43815_n1251) );
  INVX1 INVX1_870 ( .A(alu_a_i_12_), .Y(alu__abc_41358_n308) );
  INVX1 INVX1_871 ( .A(alu__abc_41358_n309), .Y(alu__abc_41358_n310) );
  INVX1 INVX1_872 ( .A(alu__abc_41358_n311), .Y(alu__abc_41358_n312) );
  INVX1 INVX1_873 ( .A(alu__abc_41358_n313), .Y(alu__abc_41358_n314) );
  INVX1 INVX1_874 ( .A(alu_b_i_13_), .Y(alu__abc_41358_n315) );
  INVX1 INVX1_875 ( .A(alu_a_i_13_), .Y(alu__abc_41358_n316) );
  INVX1 INVX1_876 ( .A(alu__abc_41358_n317), .Y(alu__abc_41358_n318) );
  INVX1 INVX1_877 ( .A(alu__abc_41358_n319), .Y(alu__abc_41358_n320) );
  INVX1 INVX1_878 ( .A(alu__abc_41358_n322), .Y(alu__abc_41358_n323) );
  INVX1 INVX1_879 ( .A(alu_b_i_14_), .Y(alu__abc_41358_n324) );
  INVX1 INVX1_88 ( .A(_abc_43815_n1252), .Y(_abc_43815_n1253) );
  INVX1 INVX1_880 ( .A(alu_a_i_14_), .Y(alu__abc_41358_n325) );
  INVX1 INVX1_881 ( .A(alu__abc_41358_n326), .Y(alu__abc_41358_n327) );
  INVX1 INVX1_882 ( .A(alu__abc_41358_n328), .Y(alu__abc_41358_n329_1) );
  INVX1 INVX1_883 ( .A(alu__abc_41358_n330), .Y(alu__abc_41358_n331) );
  INVX1 INVX1_884 ( .A(alu_b_i_15_), .Y(alu__abc_41358_n332) );
  INVX1 INVX1_885 ( .A(alu_a_i_15_), .Y(alu__abc_41358_n333) );
  INVX1 INVX1_886 ( .A(alu__abc_41358_n334), .Y(alu__abc_41358_n335) );
  INVX1 INVX1_887 ( .A(alu__abc_41358_n340), .Y(alu__abc_41358_n341) );
  INVX1 INVX1_888 ( .A(alu_b_i_10_), .Y(alu__abc_41358_n342) );
  INVX1 INVX1_889 ( .A(alu_a_i_10_), .Y(alu__abc_41358_n343) );
  INVX1 INVX1_89 ( .A(_abc_43815_n1197), .Y(_abc_43815_n1273) );
  INVX1 INVX1_890 ( .A(alu__abc_41358_n344), .Y(alu__abc_41358_n345) );
  INVX1 INVX1_891 ( .A(alu__abc_41358_n346), .Y(alu__abc_41358_n347) );
  INVX1 INVX1_892 ( .A(alu__abc_41358_n348), .Y(alu__abc_41358_n349) );
  INVX1 INVX1_893 ( .A(alu_b_i_11_), .Y(alu__abc_41358_n350) );
  INVX1 INVX1_894 ( .A(alu_a_i_11_), .Y(alu__abc_41358_n351) );
  INVX1 INVX1_895 ( .A(alu__abc_41358_n352), .Y(alu__abc_41358_n353) );
  INVX1 INVX1_896 ( .A(alu__abc_41358_n357), .Y(alu__abc_41358_n358) );
  INVX1 INVX1_897 ( .A(alu_b_i_8_), .Y(alu__abc_41358_n359) );
  INVX1 INVX1_898 ( .A(alu_a_i_8_), .Y(alu__abc_41358_n360) );
  INVX1 INVX1_899 ( .A(alu__abc_41358_n361), .Y(alu__abc_41358_n362) );
  INVX1 INVX1_9 ( .A(_abc_43815_n662), .Y(_abc_43815_n663) );
  INVX1 INVX1_90 ( .A(alu_flag_update_o), .Y(_abc_43815_n1286) );
  INVX1 INVX1_900 ( .A(alu__abc_41358_n365), .Y(alu__abc_41358_n366) );
  INVX1 INVX1_901 ( .A(alu_b_i_9_), .Y(alu__abc_41358_n367) );
  INVX1 INVX1_902 ( .A(alu_a_i_9_), .Y(alu__abc_41358_n368) );
  INVX1 INVX1_903 ( .A(alu__abc_41358_n369), .Y(alu__abc_41358_n370) );
  INVX1 INVX1_904 ( .A(alu__abc_41358_n371), .Y(alu__abc_41358_n372) );
  INVX1 INVX1_905 ( .A(alu_op_i_1_), .Y(alu__abc_41358_n378) );
  INVX1 INVX1_906 ( .A(alu_op_i_3_), .Y(alu__abc_41358_n379) );
  INVX1 INVX1_907 ( .A(alu_op_i_2_), .Y(alu__abc_41358_n382) );
  INVX1 INVX1_908 ( .A(alu_op_i_0_bF_buf5), .Y(alu__abc_41358_n384) );
  INVX1 INVX1_909 ( .A(alu__abc_41358_n391), .Y(alu__abc_41358_n392) );
  INVX1 INVX1_91 ( .A(_abc_43815_n1291), .Y(_abc_43815_n1292) );
  INVX1 INVX1_910 ( .A(alu__abc_41358_n143_1), .Y(alu__abc_41358_n393) );
  INVX1 INVX1_911 ( .A(alu__abc_41358_n395), .Y(alu__abc_41358_n396) );
  INVX1 INVX1_912 ( .A(alu__abc_41358_n397), .Y(alu__abc_41358_n398) );
  INVX1 INVX1_913 ( .A(alu__abc_41358_n402), .Y(alu__abc_41358_n403) );
  INVX1 INVX1_914 ( .A(alu__abc_41358_n405), .Y(alu__abc_41358_n406) );
  INVX1 INVX1_915 ( .A(alu__abc_41358_n409), .Y(alu__abc_41358_n410) );
  INVX1 INVX1_916 ( .A(alu__abc_41358_n413), .Y(alu__abc_41358_n414) );
  INVX1 INVX1_917 ( .A(alu__abc_41358_n431), .Y(alu__abc_41358_n432) );
  INVX1 INVX1_918 ( .A(alu__abc_41358_n433), .Y(alu__abc_41358_n434) );
  INVX1 INVX1_919 ( .A(alu__abc_41358_n437), .Y(alu__abc_41358_n438) );
  INVX1 INVX1_92 ( .A(_abc_43815_n1295), .Y(_abc_43815_n1296) );
  INVX1 INVX1_920 ( .A(alu__abc_41358_n446), .Y(alu__abc_41358_n447) );
  INVX1 INVX1_921 ( .A(alu__abc_41358_n448), .Y(alu__abc_41358_n449) );
  INVX1 INVX1_922 ( .A(alu__abc_41358_n452), .Y(alu__abc_41358_n453) );
  INVX1 INVX1_923 ( .A(alu__abc_41358_n463), .Y(alu__abc_41358_n464) );
  INVX1 INVX1_924 ( .A(alu__abc_41358_n465), .Y(alu__abc_41358_n466) );
  INVX1 INVX1_925 ( .A(alu__abc_41358_n469), .Y(alu__abc_41358_n470) );
  INVX1 INVX1_926 ( .A(alu__abc_41358_n478), .Y(alu__abc_41358_n479) );
  INVX1 INVX1_927 ( .A(alu__abc_41358_n480), .Y(alu__abc_41358_n481) );
  INVX1 INVX1_928 ( .A(alu__abc_41358_n484), .Y(alu__abc_41358_n485) );
  INVX1 INVX1_929 ( .A(alu__abc_41358_n498), .Y(alu__abc_41358_n499) );
  INVX1 INVX1_93 ( .A(alu_equal_o), .Y(_abc_43815_n1300_1) );
  INVX1 INVX1_930 ( .A(alu__abc_41358_n500), .Y(alu__abc_41358_n501) );
  INVX1 INVX1_931 ( .A(alu__abc_41358_n503), .Y(alu__abc_41358_n504) );
  INVX1 INVX1_932 ( .A(alu__abc_41358_n506), .Y(alu__abc_41358_n507) );
  INVX1 INVX1_933 ( .A(alu__abc_41358_n508), .Y(alu__abc_41358_n509) );
  INVX1 INVX1_934 ( .A(alu__abc_41358_n515), .Y(alu__abc_41358_n516) );
  INVX1 INVX1_935 ( .A(alu__abc_41358_n174), .Y(alu__abc_41358_n522) );
  INVX1 INVX1_936 ( .A(alu__abc_41358_n527), .Y(alu__abc_41358_n528) );
  INVX1 INVX1_937 ( .A(alu__abc_41358_n173), .Y(alu__abc_41358_n530) );
  INVX1 INVX1_938 ( .A(alu__abc_41358_n540), .Y(alu__abc_41358_n541) );
  INVX1 INVX1_939 ( .A(alu__abc_41358_n544), .Y(alu__abc_41358_n545) );
  INVX1 INVX1_94 ( .A(_abc_43815_n1348), .Y(_abc_43815_n1349) );
  INVX1 INVX1_940 ( .A(alu__abc_41358_n549), .Y(alu__abc_41358_n550) );
  INVX1 INVX1_941 ( .A(alu__abc_41358_n565_1), .Y(alu__abc_41358_n566) );
  INVX1 INVX1_942 ( .A(alu__abc_41358_n250), .Y(alu__abc_41358_n575) );
  INVX1 INVX1_943 ( .A(alu__abc_41358_n581), .Y(alu__abc_41358_n582) );
  INVX1 INVX1_944 ( .A(alu__abc_41358_n295), .Y(alu__abc_41358_n584) );
  INVX1 INVX1_945 ( .A(alu__abc_41358_n275), .Y(alu__abc_41358_n588) );
  INVX1 INVX1_946 ( .A(alu__abc_41358_n289), .Y(alu__abc_41358_n590) );
  INVX1 INVX1_947 ( .A(alu__abc_41358_n288), .Y(alu__abc_41358_n594) );
  INVX1 INVX1_948 ( .A(alu__abc_41358_n274), .Y(alu__abc_41358_n598) );
  INVX1 INVX1_949 ( .A(alu__abc_41358_n621), .Y(alu__abc_41358_n622) );
  INVX1 INVX1_95 ( .A(_abc_43815_n1352_1), .Y(_abc_43815_n1353_1) );
  INVX1 INVX1_950 ( .A(alu__abc_41358_n623), .Y(alu__abc_41358_n624) );
  INVX1 INVX1_951 ( .A(alu__abc_41358_n630), .Y(alu__abc_41358_n631) );
  INVX1 INVX1_952 ( .A(alu__abc_41358_n632), .Y(alu__abc_41358_n633) );
  INVX1 INVX1_953 ( .A(alu__abc_41358_n643), .Y(alu__abc_41358_n644) );
  INVX1 INVX1_954 ( .A(alu__abc_41358_n645), .Y(alu__abc_41358_n646) );
  INVX1 INVX1_955 ( .A(alu__abc_41358_n651), .Y(alu__abc_41358_n652) );
  INVX1 INVX1_956 ( .A(alu__abc_41358_n653), .Y(alu__abc_41358_n654) );
  INVX1 INVX1_957 ( .A(alu__abc_41358_n613), .Y(alu__abc_41358_n660) );
  INVX1 INVX1_958 ( .A(alu__abc_41358_n661), .Y(alu__abc_41358_n662) );
  INVX1 INVX1_959 ( .A(alu__abc_41358_n673), .Y(alu__abc_41358_n674) );
  INVX1 INVX1_96 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n1356) );
  INVX1 INVX1_960 ( .A(alu__abc_41358_n677), .Y(alu__abc_41358_n678) );
  INVX1 INVX1_961 ( .A(alu__abc_41358_n679), .Y(alu__abc_41358_n680) );
  INVX1 INVX1_962 ( .A(alu__abc_41358_n686), .Y(alu__abc_41358_n687) );
  INVX1 INVX1_963 ( .A(alu__abc_41358_n688), .Y(alu__abc_41358_n690) );
  INVX1 INVX1_964 ( .A(alu__abc_41358_n700), .Y(alu__abc_41358_n701) );
  INVX1 INVX1_965 ( .A(alu__abc_41358_n578), .Y(alu__abc_41358_n706) );
  INVX1 INVX1_966 ( .A(alu__abc_41358_n586), .Y(alu__abc_41358_n710) );
  INVX1 INVX1_967 ( .A(alu__abc_41358_n592), .Y(alu__abc_41358_n712) );
  INVX1 INVX1_968 ( .A(alu__abc_41358_n601), .Y(alu__abc_41358_n714) );
  INVX1 INVX1_969 ( .A(alu__abc_41358_n717), .Y(alu__abc_41358_n718) );
  INVX1 INVX1_97 ( .A(_abc_43815_n1357), .Y(_abc_43815_n1358) );
  INVX1 INVX1_970 ( .A(alu__abc_41358_n596), .Y(alu__abc_41358_n724) );
  INVX1 INVX1_971 ( .A(alu__abc_41358_n591), .Y(alu__abc_41358_n725) );
  INVX1 INVX1_972 ( .A(alu__abc_41358_n741), .Y(alu__abc_41358_n742) );
  INVX1 INVX1_973 ( .A(alu__abc_41358_n301), .Y(alu__abc_41358_n747) );
  INVX1 INVX1_974 ( .A(alu__abc_41358_n296), .Y(alu__abc_41358_n751) );
  INVX1 INVX1_975 ( .A(alu__abc_41358_n297), .Y(alu__abc_41358_n752) );
  INVX1 INVX1_976 ( .A(alu__abc_41358_n570), .Y(alu__abc_41358_n767) );
  INVX1 INVX1_977 ( .A(alu__abc_41358_n604), .Y(alu__abc_41358_n768) );
  INVX1 INVX1_978 ( .A(alu__abc_41358_n603), .Y(alu__abc_41358_n774) );
  INVX1 INVX1_979 ( .A(alu__abc_41358_n699), .Y(alu__abc_41358_n797) );
  INVX1 INVX1_98 ( .A(alu_c_update_o), .Y(_abc_43815_n1367) );
  INVX1 INVX1_980 ( .A(alu__abc_41358_n816), .Y(alu__abc_41358_n818_1) );
  INVX1 INVX1_981 ( .A(alu__abc_41358_n927_bF_buf4), .Y(alu__abc_41358_n928) );
  INVX1 INVX1_982 ( .A(alu__abc_41358_n744), .Y(alu__abc_41358_n943) );
  INVX1 INVX1_983 ( .A(alu__abc_41358_n258), .Y(alu__abc_41358_n1056) );
  INVX1 INVX1_984 ( .A(alu__abc_41358_n1065), .Y(alu__abc_41358_n1066) );
  INVX1 INVX1_985 ( .A(alu__abc_41358_n745), .Y(alu__abc_41358_n1072) );
  INVX1 INVX1_986 ( .A(alu__abc_41358_n1132), .Y(alu__abc_41358_n1133) );
  INVX1 INVX1_987 ( .A(alu__abc_41358_n300), .Y(alu__abc_41358_n1134) );
  INVX1 INVX1_988 ( .A(alu__abc_41358_n418), .Y(alu__abc_41358_n1137_1) );
  INVX1 INVX1_989 ( .A(alu__abc_41358_n1143), .Y(alu__abc_41358_n1144) );
  INVX1 INVX1_99 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_43815_n1381) );
  INVX1 INVX1_990 ( .A(alu__abc_41358_n750), .Y(alu__abc_41358_n1151) );
  INVX1 INVX1_991 ( .A(alu__abc_41358_n759), .Y(alu__abc_41358_n1208) );
  INVX1 INVX1_992 ( .A(alu__abc_41358_n415), .Y(alu__abc_41358_n1211) );
  INVX1 INVX1_993 ( .A(alu__abc_41358_n1226), .Y(alu__abc_41358_n1227) );
  INVX1 INVX1_994 ( .A(alu__abc_41358_n762), .Y(alu__abc_41358_n1239) );
  INVX1 INVX1_995 ( .A(alu__abc_41358_n422), .Y(alu__abc_41358_n1265) );
  INVX1 INVX1_996 ( .A(alu__abc_41358_n1281), .Y(alu__abc_41358_n1282) );
  INVX1 INVX1_997 ( .A(alu__abc_41358_n763), .Y(alu__abc_41358_n1292) );
  INVX1 INVX1_998 ( .A(alu__abc_41358_n1296), .Y(alu__abc_41358_n1297) );
  INVX1 INVX1_999 ( .A(alu__abc_41358_n411), .Y(alu__abc_41358_n1318) );
  INVX2 INVX2_1 ( .A(_abc_43815_n992), .Y(_abc_43815_n1000) );
  INVX2 INVX2_10 ( .A(alu__abc_41358_n227), .Y(alu__abc_41358_n228) );
  INVX2 INVX2_11 ( .A(alu__abc_41358_n336), .Y(alu__abc_41358_n337) );
  INVX2 INVX2_12 ( .A(alu__abc_41358_n354), .Y(alu__abc_41358_n355) );
  INVX2 INVX2_13 ( .A(alu__abc_41358_n363), .Y(alu__abc_41358_n364) );
  INVX2 INVX2_2 ( .A(_abc_43815_n1056), .Y(_abc_43815_n1057) );
  INVX2 INVX2_3 ( .A(_abc_43815_n1065_1_bF_buf4), .Y(_abc_43815_n1066) );
  INVX2 INVX2_4 ( .A(_abc_43815_n1097), .Y(_abc_43815_n1098) );
  INVX2 INVX2_5 ( .A(_abc_43815_n671_bF_buf3), .Y(_abc_43815_n3502_1) );
  INVX2 INVX2_6 ( .A(_abc_43815_n652), .Y(_abc_43815_n3509) );
  INVX2 INVX2_7 ( .A(_abc_43815_n4217_bF_buf3), .Y(_abc_43815_n4220) );
  INVX2 INVX2_8 ( .A(alu__abc_41358_n141), .Y(alu__abc_41358_n142) );
  INVX2 INVX2_9 ( .A(alu__abc_41358_n192_1), .Y(alu__abc_41358_n193) );
  INVX4 INVX4_1 ( .A(_abc_43815_n645_1_bF_buf4), .Y(_abc_43815_n646_1) );
  INVX4 INVX4_10 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2125) );
  INVX4 INVX4_11 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2130_1) );
  INVX4 INVX4_12 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2135_1) );
  INVX4 INVX4_13 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2140) );
  INVX4 INVX4_14 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2145_1) );
  INVX4 INVX4_15 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2150_1) );
  INVX4 INVX4_16 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2155) );
  INVX4 INVX4_17 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2160_1) );
  INVX4 INVX4_18 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2165_1) );
  INVX4 INVX4_19 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2170) );
  INVX4 INVX4_2 ( .A(state_q_1_bF_buf2), .Y(_abc_43815_n682) );
  INVX4 INVX4_20 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2175_1) );
  INVX4 INVX4_21 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2180_1) );
  INVX4 INVX4_22 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2185) );
  INVX4 INVX4_23 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2190_1) );
  INVX4 INVX4_24 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2195_1) );
  INVX4 INVX4_25 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2200_1) );
  INVX4 INVX4_26 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2205_1) );
  INVX4 INVX4_27 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2210) );
  INVX4 INVX4_28 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2215_1) );
  INVX4 INVX4_29 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2220_1) );
  INVX4 INVX4_3 ( .A(_abc_43815_n692_bF_buf3), .Y(_abc_43815_n693) );
  INVX4 INVX4_30 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2225) );
  INVX4 INVX4_31 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2230_1) );
  INVX4 INVX4_32 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2235_1) );
  INVX4 INVX4_33 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2240) );
  INVX4 INVX4_34 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2245_1) );
  INVX4 INVX4_35 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2250_1) );
  INVX4 INVX4_36 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2255) );
  INVX4 INVX4_37 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2260_1) );
  INVX4 INVX4_38 ( .A(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5539) );
  INVX4 INVX4_39 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n7548) );
  INVX4 INVX4_4 ( .A(_abc_43815_n987), .Y(_abc_43815_n999) );
  INVX4 INVX4_5 ( .A(_abc_43815_n1398), .Y(_abc_43815_n1692) );
  INVX4 INVX4_6 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2105_1) );
  INVX4 INVX4_7 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2110) );
  INVX4 INVX4_8 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2115_1) );
  INVX4 INVX4_9 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2120_1) );
  INVX8 INVX8_1 ( .A(_abc_43815_n641_bF_buf3), .Y(_abc_43815_n642_1) );
  INVX8 INVX8_10 ( .A(_abc_43815_n1418_bF_buf1), .Y(_abc_43815_n1489) );
  INVX8 INVX8_11 ( .A(state_q_5_), .Y(_abc_43815_n3549) );
  INVX8 INVX8_12 ( .A(rst_i), .Y(_abc_43815_n4167) );
  INVX8 INVX8_13 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2269_1) );
  INVX8 INVX8_14 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2370) );
  INVX8 INVX8_15 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2602_1) );
  INVX8 INVX8_16 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2960_1) );
  INVX8 INVX8_17 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3061) );
  INVX8 INVX8_18 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3419) );
  INVX8 INVX8_19 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3519) );
  INVX8 INVX8_2 ( .A(_abc_43815_n649_bF_buf4), .Y(_abc_43815_n650) );
  INVX8 INVX8_20 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3618) );
  INVX8 INVX8_21 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3717) );
  INVX8 INVX8_22 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3815) );
  INVX8 INVX8_23 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4044) );
  INVX8 INVX8_24 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4142) );
  INVX8 INVX8_25 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4241) );
  INVX8 INVX8_26 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4339) );
  INVX8 INVX8_27 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4695) );
  INVX8 INVX8_28 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4793_1) );
  INVX8 INVX8_29 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5149) );
  INVX8 INVX8_3 ( .A(_abc_43815_n685), .Y(_abc_43815_n686_1) );
  INVX8 INVX8_30 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5247) );
  INVX8 INVX8_31 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5345) );
  INVX8 INVX8_32 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5443) );
  INVX8 INVX8_33 ( .A(rst_i), .Y(REGFILE_SIM_reg_bank__abc_33898_n5245) );
  INVX8 INVX8_34 ( .A(alu_b_i_1_bF_buf6), .Y(alu__abc_41358_n252) );
  INVX8 INVX8_35 ( .A(alu_b_i_0_bF_buf3), .Y(alu__abc_41358_n259) );
  INVX8 INVX8_36 ( .A(alu_b_i_4_bF_buf3), .Y(alu__abc_41358_n279) );
  INVX8 INVX8_37 ( .A(alu_b_i_3_bF_buf5), .Y(alu__abc_41358_n294) );
  INVX8 INVX8_38 ( .A(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n299) );
  INVX8 INVX8_4 ( .A(_abc_43815_n1171_bF_buf5), .Y(_abc_43815_n1172_1) );
  INVX8 INVX8_5 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .Y(_abc_43815_n1278) );
  INVX8 INVX8_6 ( .A(_abc_43815_n1350_bF_buf2), .Y(_abc_43815_n1413) );
  INVX8 INVX8_7 ( .A(_abc_43815_n1428_bF_buf3), .Y(_abc_43815_n1431_1) );
  INVX8 INVX8_8 ( .A(_abc_43815_n1351_bF_buf0), .Y(_abc_43815_n1461) );
  INVX8 INVX8_9 ( .A(_abc_43815_n1472_1_bF_buf4), .Y(_abc_43815_n1473) );
  OR2X2 OR2X2_1 ( .A(state_q_0_), .B(state_q_4_), .Y(_abc_43815_n618) );
  OR2X2 OR2X2_10 ( .A(_abc_43815_n691), .B(_abc_43815_n664_1), .Y(_abc_43815_n692) );
  OR2X2 OR2X2_100 ( .A(state_q_1_bF_buf4), .B(alu_p_o_17_), .Y(_abc_43815_n896) );
  OR2X2 OR2X2_1000 ( .A(_abc_43815_n3266_1), .B(_abc_43815_n3267), .Y(alu_input_a_r_28_) );
  OR2X2 OR2X2_1001 ( .A(_abc_43815_n2514), .B(_abc_43815_n1172_1_bF_buf2), .Y(_abc_43815_n3269) );
  OR2X2 OR2X2_1002 ( .A(_abc_43815_n1171_bF_buf2), .B(_abc_43815_n3272_1), .Y(_abc_43815_n3273) );
  OR2X2 OR2X2_1003 ( .A(_abc_43815_n3271), .B(_abc_43815_n3273), .Y(_abc_43815_n3274_1) );
  OR2X2 OR2X2_1004 ( .A(_abc_43815_n3274_1), .B(_abc_43815_n3270_1), .Y(_abc_43815_n3275) );
  OR2X2 OR2X2_1005 ( .A(_abc_43815_n3276_1), .B(_abc_43815_n3277), .Y(alu_input_a_r_29_) );
  OR2X2 OR2X2_1006 ( .A(_abc_43815_n2550), .B(_abc_43815_n1172_1_bF_buf1), .Y(_abc_43815_n3279) );
  OR2X2 OR2X2_1007 ( .A(_abc_43815_n1171_bF_buf1), .B(_abc_43815_n3282_1), .Y(_abc_43815_n3283) );
  OR2X2 OR2X2_1008 ( .A(_abc_43815_n3281), .B(_abc_43815_n3283), .Y(_abc_43815_n3284_1) );
  OR2X2 OR2X2_1009 ( .A(_abc_43815_n3284_1), .B(_abc_43815_n3280_1), .Y(_abc_43815_n3285) );
  OR2X2 OR2X2_101 ( .A(_abc_43815_n898), .B(_abc_43815_n885_1), .Y(_abc_43815_n899) );
  OR2X2 OR2X2_1010 ( .A(_abc_43815_n3286_1), .B(_abc_43815_n3287), .Y(alu_input_a_r_30_) );
  OR2X2 OR2X2_1011 ( .A(_abc_43815_n2589_1), .B(_abc_43815_n1172_1_bF_buf0), .Y(_abc_43815_n3289) );
  OR2X2 OR2X2_1012 ( .A(_abc_43815_n1171_bF_buf0), .B(_abc_43815_n3292_1), .Y(_abc_43815_n3293) );
  OR2X2 OR2X2_1013 ( .A(_abc_43815_n3291), .B(_abc_43815_n3293), .Y(_abc_43815_n3294_1) );
  OR2X2 OR2X2_1014 ( .A(_abc_43815_n3294_1), .B(_abc_43815_n3290_1), .Y(_abc_43815_n3295) );
  OR2X2 OR2X2_1015 ( .A(_abc_43815_n3296_1), .B(_abc_43815_n3297), .Y(alu_input_a_r_31_) );
  OR2X2 OR2X2_1016 ( .A(_abc_43815_n2788), .B(_abc_43815_n1055), .Y(_abc_43815_n3299) );
  OR2X2 OR2X2_1017 ( .A(_abc_43815_n1153_1), .B(_abc_43815_n2775), .Y(_abc_43815_n3300_1) );
  OR2X2 OR2X2_1018 ( .A(_abc_43815_n3300_1), .B(_abc_43815_n1164), .Y(_abc_43815_n3301) );
  OR2X2 OR2X2_1019 ( .A(_abc_43815_n1126), .B(_abc_43815_n1050), .Y(_abc_43815_n3302_1) );
  OR2X2 OR2X2_102 ( .A(_abc_43815_n900_1), .B(_abc_43815_n832_1_bF_buf1), .Y(_abc_43815_n901) );
  OR2X2 OR2X2_1020 ( .A(_abc_43815_n3302_1), .B(_abc_43815_n1177), .Y(_abc_43815_n3303) );
  OR2X2 OR2X2_1021 ( .A(_abc_43815_n3301), .B(_abc_43815_n3303), .Y(_abc_43815_n3304_1) );
  OR2X2 OR2X2_1022 ( .A(_abc_43815_n3304_1), .B(_abc_43815_n3299), .Y(alu_func_r_0_) );
  OR2X2 OR2X2_1023 ( .A(_abc_43815_n2815), .B(_abc_43815_n2790), .Y(_abc_43815_n3306_1) );
  OR2X2 OR2X2_1024 ( .A(_abc_43815_n987), .B(_abc_43815_n1164), .Y(_abc_43815_n3307) );
  OR2X2 OR2X2_1025 ( .A(_abc_43815_n3307), .B(_abc_43815_n1055), .Y(_abc_43815_n3308_1) );
  OR2X2 OR2X2_1026 ( .A(_abc_43815_n3308_1), .B(_abc_43815_n3306_1), .Y(_abc_43815_n3309) );
  OR2X2 OR2X2_1027 ( .A(_abc_43815_n3309), .B(_abc_43815_n1185), .Y(alu_func_r_1_) );
  OR2X2 OR2X2_1028 ( .A(_abc_43815_n1177), .B(_abc_43815_n1159), .Y(_abc_43815_n3311) );
  OR2X2 OR2X2_1029 ( .A(_abc_43815_n2990), .B(_abc_43815_n3311), .Y(alu_func_r_3_) );
  OR2X2 OR2X2_103 ( .A(state_q_1_bF_buf3), .B(alu_p_o_18_), .Y(_abc_43815_n902) );
  OR2X2 OR2X2_1030 ( .A(_abc_43815_n680_1_bF_buf3), .B(mem_offset_q_0_), .Y(_abc_43815_n3313) );
  OR2X2 OR2X2_1031 ( .A(_abc_43815_n3314), .B(_abc_43815_n3317_bF_buf3), .Y(_abc_43815_n3318) );
  OR2X2 OR2X2_1032 ( .A(_abc_43815_n680_1_bF_buf1), .B(mem_offset_q_1_), .Y(_abc_43815_n3320) );
  OR2X2 OR2X2_1033 ( .A(_abc_43815_n3325), .B(_abc_43815_n3326), .Y(_abc_43815_n3327) );
  OR2X2 OR2X2_1034 ( .A(_abc_43815_n3314), .B(_abc_43815_n3328), .Y(_abc_43815_n3329) );
  OR2X2 OR2X2_1035 ( .A(_abc_27555_n4367_bF_buf7), .B(alu_op_r_0_), .Y(_abc_43815_n3332_1) );
  OR2X2 OR2X2_1036 ( .A(_abc_27555_n4367_bF_buf5), .B(alu_op_r_1_), .Y(_abc_43815_n3337) );
  OR2X2 OR2X2_1037 ( .A(_abc_27555_n4367_bF_buf3), .B(alu_op_r_2_), .Y(_abc_43815_n3342) );
  OR2X2 OR2X2_1038 ( .A(_abc_27555_n4367_bF_buf1), .B(alu_op_r_3_), .Y(_abc_43815_n3347_1) );
  OR2X2 OR2X2_1039 ( .A(_abc_27555_n4367_bF_buf7), .B(int32_r_4_), .Y(_abc_43815_n3352) );
  OR2X2 OR2X2_104 ( .A(_abc_43815_n904), .B(_abc_43815_n885_1), .Y(_abc_43815_n905) );
  OR2X2 OR2X2_1040 ( .A(_abc_27555_n4367_bF_buf5), .B(int32_r_5_), .Y(_abc_43815_n3357) );
  OR2X2 OR2X2_1041 ( .A(_abc_27555_n4367_bF_buf3), .B(alu_op_r_4_), .Y(_abc_43815_n3362) );
  OR2X2 OR2X2_1042 ( .A(_abc_27555_n4367_bF_buf1), .B(alu_op_r_5_), .Y(_abc_43815_n3367) );
  OR2X2 OR2X2_1043 ( .A(_abc_27555_n4367_bF_buf7), .B(alu_op_r_6_), .Y(_abc_43815_n3372) );
  OR2X2 OR2X2_1044 ( .A(_abc_27555_n4367_bF_buf5), .B(alu_op_r_7_), .Y(_abc_43815_n3377) );
  OR2X2 OR2X2_1045 ( .A(_abc_27555_n4367_bF_buf3), .B(int32_r_10_), .Y(_abc_43815_n3382) );
  OR2X2 OR2X2_1046 ( .A(_abc_27555_n4367_bF_buf1), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_43815_n3387) );
  OR2X2 OR2X2_1047 ( .A(_abc_27555_n4367_bF_buf7), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_43815_n3392) );
  OR2X2 OR2X2_1048 ( .A(_abc_27555_n4367_bF_buf5), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_43815_n3397) );
  OR2X2 OR2X2_1049 ( .A(_abc_27555_n4367_bF_buf3), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_43815_n3402) );
  OR2X2 OR2X2_105 ( .A(_abc_43815_n906), .B(_abc_43815_n832_1_bF_buf0), .Y(_abc_43815_n907) );
  OR2X2 OR2X2_1050 ( .A(_abc_27555_n4367_bF_buf1), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0), .Y(_abc_43815_n3407) );
  OR2X2 OR2X2_1051 ( .A(_abc_27555_n4367_bF_buf7), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(_abc_43815_n3412) );
  OR2X2 OR2X2_1052 ( .A(_abc_27555_n4367_bF_buf5), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(_abc_43815_n3417) );
  OR2X2 OR2X2_1053 ( .A(_abc_27555_n4367_bF_buf3), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(_abc_43815_n3422) );
  OR2X2 OR2X2_1054 ( .A(_abc_27555_n4367_bF_buf1), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(_abc_43815_n3427) );
  OR2X2 OR2X2_1055 ( .A(_abc_27555_n4367_bF_buf7), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(_abc_43815_n3432) );
  OR2X2 OR2X2_1056 ( .A(_abc_27555_n4367_bF_buf5), .B(opcode_q_21_), .Y(_abc_43815_n3437) );
  OR2X2 OR2X2_1057 ( .A(_abc_27555_n4367_bF_buf3), .B(opcode_q_22_), .Y(_abc_43815_n3442) );
  OR2X2 OR2X2_1058 ( .A(_abc_27555_n4367_bF_buf1), .B(opcode_q_23_), .Y(_abc_43815_n3447_1) );
  OR2X2 OR2X2_1059 ( .A(_abc_27555_n4367_bF_buf7), .B(opcode_q_24_), .Y(_abc_43815_n3452) );
  OR2X2 OR2X2_106 ( .A(state_q_1_bF_buf2), .B(alu_p_o_19_), .Y(_abc_43815_n908) );
  OR2X2 OR2X2_1060 ( .A(_abc_27555_n4367_bF_buf5), .B(opcode_q_25_), .Y(_abc_43815_n3457_1) );
  OR2X2 OR2X2_1061 ( .A(_abc_27555_n4367_bF_buf3), .B(inst_r_0_), .Y(_abc_43815_n3462) );
  OR2X2 OR2X2_1062 ( .A(_abc_27555_n4367_bF_buf1), .B(inst_r_1_), .Y(_abc_43815_n3467) );
  OR2X2 OR2X2_1063 ( .A(_abc_27555_n4367_bF_buf7), .B(inst_r_2_), .Y(_abc_43815_n3472) );
  OR2X2 OR2X2_1064 ( .A(_abc_27555_n4367_bF_buf5), .B(inst_r_3_), .Y(_abc_43815_n3477) );
  OR2X2 OR2X2_1065 ( .A(_abc_27555_n4367_bF_buf3), .B(inst_r_4_), .Y(_abc_43815_n3482) );
  OR2X2 OR2X2_1066 ( .A(_abc_27555_n4367_bF_buf1), .B(inst_r_5_), .Y(_abc_43815_n3487) );
  OR2X2 OR2X2_1067 ( .A(state_q_5_), .B(_auto_iopadmap_cc_313_execute_47802_0_), .Y(_abc_43815_n3492_1) );
  OR2X2 OR2X2_1068 ( .A(_abc_43815_n3493_1), .B(_auto_iopadmap_cc_313_execute_47802_0_), .Y(_abc_43815_n3494) );
  OR2X2 OR2X2_1069 ( .A(_abc_43815_n650_bF_buf2), .B(_abc_43815_n3497), .Y(_abc_43815_n3498) );
  OR2X2 OR2X2_107 ( .A(_abc_43815_n910), .B(_abc_43815_n885_1), .Y(_abc_43815_n911) );
  OR2X2 OR2X2_1070 ( .A(_abc_43815_n3496_bF_buf3), .B(_abc_43815_n3498), .Y(_abc_43815_n3499) );
  OR2X2 OR2X2_1071 ( .A(_abc_43815_n3502_1), .B(_abc_43815_n3504), .Y(_abc_43815_n3505) );
  OR2X2 OR2X2_1072 ( .A(_abc_43815_n3505), .B(_abc_43815_n3501_1), .Y(_abc_43815_n3506) );
  OR2X2 OR2X2_1073 ( .A(state_q_5_), .B(_auto_iopadmap_cc_313_execute_47802_1_), .Y(_abc_43815_n3508) );
  OR2X2 OR2X2_1074 ( .A(_abc_43815_n3509), .B(_auto_iopadmap_cc_313_execute_47802_1_), .Y(_abc_43815_n3510) );
  OR2X2 OR2X2_1075 ( .A(_abc_43815_n3496_bF_buf2), .B(_abc_43815_n1079), .Y(_abc_43815_n3513) );
  OR2X2 OR2X2_1076 ( .A(_abc_43815_n3513), .B(_abc_43815_n3512_1), .Y(_abc_43815_n3514) );
  OR2X2 OR2X2_1077 ( .A(_abc_43815_n3515), .B(_abc_43815_n3502_1), .Y(_abc_43815_n3516) );
  OR2X2 OR2X2_1078 ( .A(state_q_5_), .B(_auto_iopadmap_cc_313_execute_47802_2_), .Y(_abc_43815_n3518) );
  OR2X2 OR2X2_1079 ( .A(_abc_43815_n3493_1), .B(_auto_iopadmap_cc_313_execute_47802_2_), .Y(_abc_43815_n3519) );
  OR2X2 OR2X2_108 ( .A(_abc_43815_n912), .B(_abc_43815_n832_1_bF_buf3), .Y(_abc_43815_n913) );
  OR2X2 OR2X2_1080 ( .A(_abc_43815_n650_bF_buf1), .B(_abc_43815_n3522_1), .Y(_abc_43815_n3523) );
  OR2X2 OR2X2_1081 ( .A(_abc_43815_n3521_1_bF_buf3), .B(_abc_43815_n3523), .Y(_abc_43815_n3524) );
  OR2X2 OR2X2_1082 ( .A(_abc_43815_n3502_1), .B(_abc_43815_n3526), .Y(_abc_43815_n3527) );
  OR2X2 OR2X2_1083 ( .A(_abc_43815_n3527), .B(_abc_43815_n3525), .Y(_abc_43815_n3528) );
  OR2X2 OR2X2_1084 ( .A(state_q_5_), .B(_auto_iopadmap_cc_313_execute_47802_3_), .Y(_abc_43815_n3530) );
  OR2X2 OR2X2_1085 ( .A(_abc_43815_n3509), .B(_auto_iopadmap_cc_313_execute_47802_3_), .Y(_abc_43815_n3531_1) );
  OR2X2 OR2X2_1086 ( .A(_abc_43815_n3521_1_bF_buf2), .B(_abc_43815_n1079), .Y(_abc_43815_n3533) );
  OR2X2 OR2X2_1087 ( .A(_abc_43815_n3533), .B(_abc_43815_n3532_1), .Y(_abc_43815_n3534) );
  OR2X2 OR2X2_1088 ( .A(_abc_43815_n3535), .B(_abc_43815_n3502_1), .Y(_abc_43815_n3536) );
  OR2X2 OR2X2_1089 ( .A(_abc_43815_n3504), .B(_abc_43815_n645_1_bF_buf3), .Y(_abc_43815_n3538) );
  OR2X2 OR2X2_109 ( .A(state_q_1_bF_buf1), .B(alu_p_o_20_), .Y(_abc_43815_n914) );
  OR2X2 OR2X2_1090 ( .A(_abc_43815_n651_1), .B(_abc_43815_n3540), .Y(_abc_43815_n3541_1) );
  OR2X2 OR2X2_1091 ( .A(_abc_43815_n3544), .B(_abc_43815_n3542_1), .Y(_abc_43815_n3545) );
  OR2X2 OR2X2_1092 ( .A(_abc_43815_n3546), .B(_abc_43815_n3539), .Y(_abc_43815_n3547) );
  OR2X2 OR2X2_1093 ( .A(_abc_43815_n3548), .B(_abc_43815_n3550), .Y(mem_dat_o_0__FF_INPUT) );
  OR2X2 OR2X2_1094 ( .A(_abc_43815_n3555), .B(_abc_43815_n3553), .Y(_abc_43815_n3556) );
  OR2X2 OR2X2_1095 ( .A(_abc_43815_n3557), .B(_abc_43815_n3552_1), .Y(_abc_43815_n3558) );
  OR2X2 OR2X2_1096 ( .A(_abc_43815_n3559), .B(_abc_43815_n3560), .Y(mem_dat_o_1__FF_INPUT) );
  OR2X2 OR2X2_1097 ( .A(_abc_43815_n3565), .B(_abc_43815_n3563), .Y(_abc_43815_n3566) );
  OR2X2 OR2X2_1098 ( .A(_abc_43815_n3567), .B(_abc_43815_n3562_1), .Y(_abc_43815_n3568) );
  OR2X2 OR2X2_1099 ( .A(_abc_43815_n3569), .B(_abc_43815_n3570), .Y(mem_dat_o_2__FF_INPUT) );
  OR2X2 OR2X2_11 ( .A(_abc_43815_n692_bF_buf2), .B(_abc_43815_n696), .Y(_abc_43815_n697) );
  OR2X2 OR2X2_110 ( .A(_abc_43815_n916_1), .B(_abc_43815_n885_1), .Y(_abc_43815_n917_1) );
  OR2X2 OR2X2_1100 ( .A(_abc_43815_n3575), .B(_abc_43815_n3573), .Y(_abc_43815_n3576) );
  OR2X2 OR2X2_1101 ( .A(_abc_43815_n3577), .B(_abc_43815_n3572_1), .Y(_abc_43815_n3578) );
  OR2X2 OR2X2_1102 ( .A(_abc_43815_n3579), .B(_abc_43815_n3580), .Y(mem_dat_o_3__FF_INPUT) );
  OR2X2 OR2X2_1103 ( .A(_abc_43815_n3585), .B(_abc_43815_n3583), .Y(_abc_43815_n3586) );
  OR2X2 OR2X2_1104 ( .A(_abc_43815_n3587), .B(_abc_43815_n3582_1), .Y(_abc_43815_n3588) );
  OR2X2 OR2X2_1105 ( .A(_abc_43815_n3589), .B(_abc_43815_n3590_1), .Y(mem_dat_o_4__FF_INPUT) );
  OR2X2 OR2X2_1106 ( .A(_abc_43815_n3595), .B(_abc_43815_n3593), .Y(_abc_43815_n3596) );
  OR2X2 OR2X2_1107 ( .A(_abc_43815_n3597), .B(_abc_43815_n3592), .Y(_abc_43815_n3598) );
  OR2X2 OR2X2_1108 ( .A(_abc_43815_n3599_1), .B(_abc_43815_n3600_1), .Y(mem_dat_o_5__FF_INPUT) );
  OR2X2 OR2X2_1109 ( .A(_abc_43815_n3605), .B(_abc_43815_n3603), .Y(_abc_43815_n3606) );
  OR2X2 OR2X2_111 ( .A(_abc_43815_n918), .B(_abc_43815_n832_1_bF_buf2), .Y(_abc_43815_n919) );
  OR2X2 OR2X2_1110 ( .A(_abc_43815_n3607), .B(_abc_43815_n3602), .Y(_abc_43815_n3608_1) );
  OR2X2 OR2X2_1111 ( .A(_abc_43815_n3609_1), .B(_abc_43815_n3610), .Y(mem_dat_o_6__FF_INPUT) );
  OR2X2 OR2X2_1112 ( .A(_abc_43815_n3615), .B(_abc_43815_n3613), .Y(_abc_43815_n3616) );
  OR2X2 OR2X2_1113 ( .A(_abc_43815_n3617_1), .B(_abc_43815_n3612), .Y(_abc_43815_n3618_1) );
  OR2X2 OR2X2_1114 ( .A(_abc_43815_n3619), .B(_abc_43815_n3620), .Y(mem_dat_o_7__FF_INPUT) );
  OR2X2 OR2X2_1115 ( .A(_abc_43815_n650_bF_buf0), .B(_abc_43815_n3624), .Y(_abc_43815_n3625) );
  OR2X2 OR2X2_1116 ( .A(_abc_43815_n3623), .B(_abc_43815_n3625), .Y(_abc_43815_n3626_1) );
  OR2X2 OR2X2_1117 ( .A(_abc_43815_n3628), .B(_abc_43815_n649_bF_buf4), .Y(_abc_43815_n3629) );
  OR2X2 OR2X2_1118 ( .A(_abc_43815_n3629), .B(_abc_43815_n3627_1), .Y(_abc_43815_n3630) );
  OR2X2 OR2X2_1119 ( .A(_abc_43815_n3631), .B(_abc_43815_n641_bF_buf1), .Y(_abc_43815_n3632) );
  OR2X2 OR2X2_112 ( .A(state_q_1_bF_buf0), .B(alu_p_o_21_), .Y(_abc_43815_n920) );
  OR2X2 OR2X2_1120 ( .A(_abc_43815_n3543), .B(_abc_43815_n642_1_bF_buf4), .Y(_abc_43815_n3633) );
  OR2X2 OR2X2_1121 ( .A(_abc_43815_n3635_1), .B(_abc_43815_n3622), .Y(mem_dat_o_8__FF_INPUT) );
  OR2X2 OR2X2_1122 ( .A(_abc_43815_n650_bF_buf4), .B(_abc_43815_n3639), .Y(_abc_43815_n3640) );
  OR2X2 OR2X2_1123 ( .A(_abc_43815_n3638), .B(_abc_43815_n3640), .Y(_abc_43815_n3641) );
  OR2X2 OR2X2_1124 ( .A(_abc_43815_n3643), .B(_abc_43815_n649_bF_buf3), .Y(_abc_43815_n3644_1) );
  OR2X2 OR2X2_1125 ( .A(_abc_43815_n3644_1), .B(_abc_43815_n3642), .Y(_abc_43815_n3645_1) );
  OR2X2 OR2X2_1126 ( .A(_abc_43815_n3646), .B(_abc_43815_n641_bF_buf0), .Y(_abc_43815_n3647) );
  OR2X2 OR2X2_1127 ( .A(_abc_43815_n3554), .B(_abc_43815_n642_1_bF_buf3), .Y(_abc_43815_n3648) );
  OR2X2 OR2X2_1128 ( .A(_abc_43815_n3650), .B(_abc_43815_n3637), .Y(mem_dat_o_9__FF_INPUT) );
  OR2X2 OR2X2_1129 ( .A(_abc_43815_n650_bF_buf3), .B(_abc_43815_n3654), .Y(_abc_43815_n3655_1) );
  OR2X2 OR2X2_113 ( .A(_abc_43815_n922), .B(_abc_43815_n885_1), .Y(_abc_43815_n923) );
  OR2X2 OR2X2_1130 ( .A(_abc_43815_n3653_1), .B(_abc_43815_n3655_1), .Y(_abc_43815_n3656) );
  OR2X2 OR2X2_1131 ( .A(_abc_43815_n3658), .B(_abc_43815_n649_bF_buf2), .Y(_abc_43815_n3659) );
  OR2X2 OR2X2_1132 ( .A(_abc_43815_n3659), .B(_abc_43815_n3657), .Y(_abc_43815_n3660) );
  OR2X2 OR2X2_1133 ( .A(_abc_43815_n3661), .B(_abc_43815_n641_bF_buf3), .Y(_abc_43815_n3662) );
  OR2X2 OR2X2_1134 ( .A(_abc_43815_n3564), .B(_abc_43815_n642_1_bF_buf2), .Y(_abc_43815_n3663) );
  OR2X2 OR2X2_1135 ( .A(_abc_43815_n3665), .B(_abc_43815_n3652), .Y(mem_dat_o_10__FF_INPUT) );
  OR2X2 OR2X2_1136 ( .A(_abc_43815_n650_bF_buf2), .B(_abc_43815_n3669_1), .Y(_abc_43815_n3670) );
  OR2X2 OR2X2_1137 ( .A(_abc_43815_n3668_1), .B(_abc_43815_n3670), .Y(_abc_43815_n3671) );
  OR2X2 OR2X2_1138 ( .A(_abc_43815_n3673), .B(_abc_43815_n649_bF_buf1), .Y(_abc_43815_n3674) );
  OR2X2 OR2X2_1139 ( .A(_abc_43815_n3674), .B(_abc_43815_n3672), .Y(_abc_43815_n3675) );
  OR2X2 OR2X2_114 ( .A(_abc_43815_n924), .B(_abc_43815_n832_1_bF_buf1), .Y(_abc_43815_n925) );
  OR2X2 OR2X2_1140 ( .A(_abc_43815_n3676), .B(_abc_43815_n641_bF_buf2), .Y(_abc_43815_n3677) );
  OR2X2 OR2X2_1141 ( .A(_abc_43815_n3574), .B(_abc_43815_n642_1_bF_buf1), .Y(_abc_43815_n3678) );
  OR2X2 OR2X2_1142 ( .A(_abc_43815_n3680_1), .B(_abc_43815_n3667_1), .Y(mem_dat_o_11__FF_INPUT) );
  OR2X2 OR2X2_1143 ( .A(_abc_43815_n650_bF_buf1), .B(_abc_43815_n3684), .Y(_abc_43815_n3685) );
  OR2X2 OR2X2_1144 ( .A(_abc_43815_n3683_1), .B(_abc_43815_n3685), .Y(_abc_43815_n3686) );
  OR2X2 OR2X2_1145 ( .A(_abc_43815_n3688), .B(_abc_43815_n649_bF_buf0), .Y(_abc_43815_n3689) );
  OR2X2 OR2X2_1146 ( .A(_abc_43815_n3689), .B(_abc_43815_n3687), .Y(_abc_43815_n3690) );
  OR2X2 OR2X2_1147 ( .A(_abc_43815_n3691), .B(_abc_43815_n641_bF_buf1), .Y(_abc_43815_n3692) );
  OR2X2 OR2X2_1148 ( .A(_abc_43815_n3584), .B(_abc_43815_n642_1_bF_buf0), .Y(_abc_43815_n3693) );
  OR2X2 OR2X2_1149 ( .A(_abc_43815_n3695_1), .B(_abc_43815_n3682), .Y(mem_dat_o_12__FF_INPUT) );
  OR2X2 OR2X2_115 ( .A(state_q_1_bF_buf4), .B(alu_p_o_22_), .Y(_abc_43815_n926) );
  OR2X2 OR2X2_1150 ( .A(_abc_43815_n650_bF_buf0), .B(_abc_43815_n3699), .Y(_abc_43815_n3700) );
  OR2X2 OR2X2_1151 ( .A(_abc_43815_n3698), .B(_abc_43815_n3700), .Y(_abc_43815_n3701_1) );
  OR2X2 OR2X2_1152 ( .A(_abc_43815_n3703), .B(_abc_43815_n649_bF_buf4), .Y(_abc_43815_n3704) );
  OR2X2 OR2X2_1153 ( .A(_abc_43815_n3704), .B(_abc_43815_n3702_1), .Y(_abc_43815_n3705) );
  OR2X2 OR2X2_1154 ( .A(_abc_43815_n3706), .B(_abc_43815_n641_bF_buf0), .Y(_abc_43815_n3707_1) );
  OR2X2 OR2X2_1155 ( .A(_abc_43815_n3594), .B(_abc_43815_n642_1_bF_buf5), .Y(_abc_43815_n3708) );
  OR2X2 OR2X2_1156 ( .A(_abc_43815_n3710), .B(_abc_43815_n3697), .Y(mem_dat_o_13__FF_INPUT) );
  OR2X2 OR2X2_1157 ( .A(_abc_43815_n650_bF_buf4), .B(_abc_43815_n3714), .Y(_abc_43815_n3715) );
  OR2X2 OR2X2_1158 ( .A(_abc_43815_n3713_1), .B(_abc_43815_n3715), .Y(_abc_43815_n3716) );
  OR2X2 OR2X2_1159 ( .A(_abc_43815_n3718), .B(_abc_43815_n649_bF_buf3), .Y(_abc_43815_n3719) );
  OR2X2 OR2X2_116 ( .A(_abc_43815_n928), .B(_abc_43815_n885_1), .Y(_abc_43815_n929) );
  OR2X2 OR2X2_1160 ( .A(_abc_43815_n3719), .B(_abc_43815_n3717), .Y(_abc_43815_n3720_1) );
  OR2X2 OR2X2_1161 ( .A(_abc_43815_n3721), .B(_abc_43815_n641_bF_buf3), .Y(_abc_43815_n3722) );
  OR2X2 OR2X2_1162 ( .A(_abc_43815_n3604), .B(_abc_43815_n642_1_bF_buf4), .Y(_abc_43815_n3723) );
  OR2X2 OR2X2_1163 ( .A(_abc_43815_n3725), .B(_abc_43815_n3712), .Y(mem_dat_o_14__FF_INPUT) );
  OR2X2 OR2X2_1164 ( .A(_abc_43815_n650_bF_buf3), .B(_abc_43815_n3729), .Y(_abc_43815_n3730) );
  OR2X2 OR2X2_1165 ( .A(_abc_43815_n3728), .B(_abc_43815_n3730), .Y(_abc_43815_n3731) );
  OR2X2 OR2X2_1166 ( .A(_abc_43815_n3733_1), .B(_abc_43815_n649_bF_buf2), .Y(_abc_43815_n3734) );
  OR2X2 OR2X2_1167 ( .A(_abc_43815_n3734), .B(_abc_43815_n3732), .Y(_abc_43815_n3735) );
  OR2X2 OR2X2_1168 ( .A(_abc_43815_n3736), .B(_abc_43815_n641_bF_buf2), .Y(_abc_43815_n3737) );
  OR2X2 OR2X2_1169 ( .A(_abc_43815_n3614), .B(_abc_43815_n642_1_bF_buf3), .Y(_abc_43815_n3738) );
  OR2X2 OR2X2_117 ( .A(_abc_43815_n930), .B(_abc_43815_n832_1_bF_buf0), .Y(_abc_43815_n931) );
  OR2X2 OR2X2_1170 ( .A(_abc_43815_n3740), .B(_abc_43815_n3727), .Y(mem_dat_o_15__FF_INPUT) );
  OR2X2 OR2X2_1171 ( .A(_abc_43815_n3746), .B(_abc_43815_n3748), .Y(_abc_43815_n3749) );
  OR2X2 OR2X2_1172 ( .A(_abc_43815_n3749), .B(_abc_43815_n3745), .Y(_abc_43815_n3750_1) );
  OR2X2 OR2X2_1173 ( .A(_abc_43815_n3751), .B(_abc_43815_n3743_1), .Y(_abc_43815_n3752) );
  OR2X2 OR2X2_1174 ( .A(_abc_43815_n3753), .B(_abc_43815_n3742), .Y(mem_dat_o_16__FF_INPUT) );
  OR2X2 OR2X2_1175 ( .A(_abc_43815_n3759), .B(_abc_43815_n3761), .Y(_abc_43815_n3762) );
  OR2X2 OR2X2_1176 ( .A(_abc_43815_n3762), .B(_abc_43815_n3758), .Y(_abc_43815_n3763_1) );
  OR2X2 OR2X2_1177 ( .A(_abc_43815_n3764), .B(_abc_43815_n3756_1), .Y(_abc_43815_n3765) );
  OR2X2 OR2X2_1178 ( .A(_abc_43815_n3766), .B(_abc_43815_n3755), .Y(mem_dat_o_17__FF_INPUT) );
  OR2X2 OR2X2_1179 ( .A(_abc_43815_n3772), .B(_abc_43815_n3774), .Y(_abc_43815_n3775) );
  OR2X2 OR2X2_118 ( .A(state_q_1_bF_buf3), .B(alu_p_o_23_), .Y(_abc_43815_n932) );
  OR2X2 OR2X2_1180 ( .A(_abc_43815_n3775), .B(_abc_43815_n3771), .Y(_abc_43815_n3776) );
  OR2X2 OR2X2_1181 ( .A(_abc_43815_n3777), .B(_abc_43815_n3769), .Y(_abc_43815_n3778) );
  OR2X2 OR2X2_1182 ( .A(_abc_43815_n3779), .B(_abc_43815_n3768), .Y(mem_dat_o_18__FF_INPUT) );
  OR2X2 OR2X2_1183 ( .A(_abc_43815_n3786_1), .B(_abc_43815_n3785), .Y(_abc_43815_n3787) );
  OR2X2 OR2X2_1184 ( .A(_abc_43815_n3787), .B(_abc_43815_n3784), .Y(_abc_43815_n3788) );
  OR2X2 OR2X2_1185 ( .A(_abc_43815_n3789), .B(_abc_43815_n3782), .Y(_abc_43815_n3790) );
  OR2X2 OR2X2_1186 ( .A(_abc_43815_n3791), .B(_abc_43815_n3781), .Y(mem_dat_o_19__FF_INPUT) );
  OR2X2 OR2X2_1187 ( .A(_abc_43815_n3797), .B(_abc_43815_n3799), .Y(_abc_43815_n3800) );
  OR2X2 OR2X2_1188 ( .A(_abc_43815_n3800), .B(_abc_43815_n3796), .Y(_abc_43815_n3801) );
  OR2X2 OR2X2_1189 ( .A(_abc_43815_n3802), .B(_abc_43815_n3794), .Y(_abc_43815_n3803) );
  OR2X2 OR2X2_119 ( .A(_abc_43815_n934_1), .B(_abc_43815_n885_1), .Y(_abc_43815_n935) );
  OR2X2 OR2X2_1190 ( .A(_abc_43815_n3804), .B(_abc_43815_n3793_1), .Y(mem_dat_o_20__FF_INPUT) );
  OR2X2 OR2X2_1191 ( .A(_abc_43815_n3810), .B(_abc_43815_n3812_1), .Y(_abc_43815_n3813) );
  OR2X2 OR2X2_1192 ( .A(_abc_43815_n3813), .B(_abc_43815_n3809), .Y(_abc_43815_n3814) );
  OR2X2 OR2X2_1193 ( .A(_abc_43815_n3815), .B(_abc_43815_n3807), .Y(_abc_43815_n3816) );
  OR2X2 OR2X2_1194 ( .A(_abc_43815_n3817), .B(_abc_43815_n3806), .Y(mem_dat_o_21__FF_INPUT) );
  OR2X2 OR2X2_1195 ( .A(_abc_43815_n3823), .B(_abc_43815_n3825_1), .Y(_abc_43815_n3826) );
  OR2X2 OR2X2_1196 ( .A(_abc_43815_n3826), .B(_abc_43815_n3822), .Y(_abc_43815_n3827) );
  OR2X2 OR2X2_1197 ( .A(_abc_43815_n3828), .B(_abc_43815_n3820), .Y(_abc_43815_n3829) );
  OR2X2 OR2X2_1198 ( .A(_abc_43815_n3830), .B(_abc_43815_n3819), .Y(mem_dat_o_22__FF_INPUT) );
  OR2X2 OR2X2_1199 ( .A(_abc_43815_n3837), .B(_abc_43815_n3836), .Y(_abc_43815_n3838) );
  OR2X2 OR2X2_12 ( .A(_abc_43815_n695), .B(_abc_43815_n698), .Y(_abc_43815_n699) );
  OR2X2 OR2X2_120 ( .A(_abc_43815_n936), .B(_abc_43815_n832_1_bF_buf3), .Y(_abc_43815_n937_1) );
  OR2X2 OR2X2_1200 ( .A(_abc_43815_n3838), .B(_abc_43815_n3835_1), .Y(_abc_43815_n3839) );
  OR2X2 OR2X2_1201 ( .A(_abc_43815_n3840), .B(_abc_43815_n3833), .Y(_abc_43815_n3841) );
  OR2X2 OR2X2_1202 ( .A(_abc_43815_n3842_1), .B(_abc_43815_n3832), .Y(mem_dat_o_23__FF_INPUT) );
  OR2X2 OR2X2_1203 ( .A(_abc_43815_n3744), .B(_abc_43815_n642_1_bF_buf0), .Y(_abc_43815_n3845) );
  OR2X2 OR2X2_1204 ( .A(_abc_43815_n3846), .B(_abc_43815_n3847), .Y(_abc_43815_n3848) );
  OR2X2 OR2X2_1205 ( .A(_abc_43815_n3848), .B(_abc_43815_n649_bF_buf3), .Y(_abc_43815_n3849_1) );
  OR2X2 OR2X2_1206 ( .A(_abc_43815_n650_bF_buf1), .B(_abc_43815_n3851), .Y(_abc_43815_n3852) );
  OR2X2 OR2X2_1207 ( .A(_abc_43815_n3850), .B(_abc_43815_n3852), .Y(_abc_43815_n3853) );
  OR2X2 OR2X2_1208 ( .A(_abc_43815_n3854), .B(_abc_43815_n641_bF_buf1), .Y(_abc_43815_n3855) );
  OR2X2 OR2X2_1209 ( .A(_abc_43815_n3857), .B(_abc_43815_n3844), .Y(mem_dat_o_24__FF_INPUT) );
  OR2X2 OR2X2_121 ( .A(state_q_1_bF_buf2), .B(alu_p_o_24_), .Y(_abc_43815_n938) );
  OR2X2 OR2X2_1210 ( .A(_abc_43815_n3757), .B(_abc_43815_n642_1_bF_buf5), .Y(_abc_43815_n3860) );
  OR2X2 OR2X2_1211 ( .A(_abc_43815_n3861), .B(_abc_43815_n3862), .Y(_abc_43815_n3863) );
  OR2X2 OR2X2_1212 ( .A(_abc_43815_n3863), .B(_abc_43815_n649_bF_buf2), .Y(_abc_43815_n3864) );
  OR2X2 OR2X2_1213 ( .A(_abc_43815_n650_bF_buf0), .B(_abc_43815_n3866), .Y(_abc_43815_n3867) );
  OR2X2 OR2X2_1214 ( .A(_abc_43815_n3865), .B(_abc_43815_n3867), .Y(_abc_43815_n3868) );
  OR2X2 OR2X2_1215 ( .A(_abc_43815_n3869), .B(_abc_43815_n641_bF_buf0), .Y(_abc_43815_n3870_1) );
  OR2X2 OR2X2_1216 ( .A(_abc_43815_n3872), .B(_abc_43815_n3859), .Y(mem_dat_o_25__FF_INPUT) );
  OR2X2 OR2X2_1217 ( .A(_abc_43815_n3770), .B(_abc_43815_n642_1_bF_buf4), .Y(_abc_43815_n3875) );
  OR2X2 OR2X2_1218 ( .A(_abc_43815_n3876), .B(_abc_43815_n3877_1), .Y(_abc_43815_n3878) );
  OR2X2 OR2X2_1219 ( .A(_abc_43815_n3878), .B(_abc_43815_n649_bF_buf1), .Y(_abc_43815_n3879) );
  OR2X2 OR2X2_122 ( .A(_abc_43815_n940), .B(_abc_43815_n885_1), .Y(_abc_43815_n941) );
  OR2X2 OR2X2_1220 ( .A(_abc_43815_n650_bF_buf4), .B(_abc_43815_n3881), .Y(_abc_43815_n3882) );
  OR2X2 OR2X2_1221 ( .A(_abc_43815_n3880), .B(_abc_43815_n3882), .Y(_abc_43815_n3883) );
  OR2X2 OR2X2_1222 ( .A(_abc_43815_n3884_1), .B(_abc_43815_n641_bF_buf3), .Y(_abc_43815_n3885) );
  OR2X2 OR2X2_1223 ( .A(_abc_43815_n3887), .B(_abc_43815_n3874), .Y(mem_dat_o_26__FF_INPUT) );
  OR2X2 OR2X2_1224 ( .A(_abc_43815_n3783), .B(_abc_43815_n642_1_bF_buf3), .Y(_abc_43815_n3890) );
  OR2X2 OR2X2_1225 ( .A(_abc_43815_n3891_1), .B(_abc_43815_n3892), .Y(_abc_43815_n3893) );
  OR2X2 OR2X2_1226 ( .A(_abc_43815_n3893), .B(_abc_43815_n649_bF_buf0), .Y(_abc_43815_n3894) );
  OR2X2 OR2X2_1227 ( .A(_abc_43815_n650_bF_buf3), .B(_abc_43815_n3896), .Y(_abc_43815_n3897) );
  OR2X2 OR2X2_1228 ( .A(_abc_43815_n3895), .B(_abc_43815_n3897), .Y(_abc_43815_n3898) );
  OR2X2 OR2X2_1229 ( .A(_abc_43815_n3899), .B(_abc_43815_n641_bF_buf2), .Y(_abc_43815_n3900) );
  OR2X2 OR2X2_123 ( .A(_abc_43815_n942), .B(_abc_43815_n832_1_bF_buf2), .Y(_abc_43815_n943) );
  OR2X2 OR2X2_1230 ( .A(_abc_43815_n3902), .B(_abc_43815_n3889), .Y(mem_dat_o_27__FF_INPUT) );
  OR2X2 OR2X2_1231 ( .A(_abc_43815_n3795), .B(_abc_43815_n642_1_bF_buf2), .Y(_abc_43815_n3905) );
  OR2X2 OR2X2_1232 ( .A(_abc_43815_n3906), .B(_abc_43815_n3907), .Y(_abc_43815_n3908_1) );
  OR2X2 OR2X2_1233 ( .A(_abc_43815_n3908_1), .B(_abc_43815_n649_bF_buf4), .Y(_abc_43815_n3909) );
  OR2X2 OR2X2_1234 ( .A(_abc_43815_n650_bF_buf2), .B(_abc_43815_n3911), .Y(_abc_43815_n3912) );
  OR2X2 OR2X2_1235 ( .A(_abc_43815_n3910), .B(_abc_43815_n3912), .Y(_abc_43815_n3913) );
  OR2X2 OR2X2_1236 ( .A(_abc_43815_n3914), .B(_abc_43815_n641_bF_buf1), .Y(_abc_43815_n3915) );
  OR2X2 OR2X2_1237 ( .A(_abc_43815_n3917), .B(_abc_43815_n3904), .Y(mem_dat_o_28__FF_INPUT) );
  OR2X2 OR2X2_1238 ( .A(_abc_43815_n3808), .B(_abc_43815_n642_1_bF_buf1), .Y(_abc_43815_n3920) );
  OR2X2 OR2X2_1239 ( .A(_abc_43815_n3921), .B(_abc_43815_n3922), .Y(_abc_43815_n3923_1) );
  OR2X2 OR2X2_124 ( .A(state_q_1_bF_buf1), .B(alu_p_o_25_), .Y(_abc_43815_n944) );
  OR2X2 OR2X2_1240 ( .A(_abc_43815_n3923_1), .B(_abc_43815_n649_bF_buf3), .Y(_abc_43815_n3924) );
  OR2X2 OR2X2_1241 ( .A(_abc_43815_n650_bF_buf1), .B(_abc_43815_n3926), .Y(_abc_43815_n3927) );
  OR2X2 OR2X2_1242 ( .A(_abc_43815_n3925), .B(_abc_43815_n3927), .Y(_abc_43815_n3928) );
  OR2X2 OR2X2_1243 ( .A(_abc_43815_n3929), .B(_abc_43815_n641_bF_buf0), .Y(_abc_43815_n3930) );
  OR2X2 OR2X2_1244 ( .A(_abc_43815_n3932), .B(_abc_43815_n3919), .Y(mem_dat_o_29__FF_INPUT) );
  OR2X2 OR2X2_1245 ( .A(_abc_43815_n3821), .B(_abc_43815_n642_1_bF_buf0), .Y(_abc_43815_n3935) );
  OR2X2 OR2X2_1246 ( .A(_abc_43815_n3936), .B(_abc_43815_n3937), .Y(_abc_43815_n3938_1) );
  OR2X2 OR2X2_1247 ( .A(_abc_43815_n3938_1), .B(_abc_43815_n649_bF_buf2), .Y(_abc_43815_n3939) );
  OR2X2 OR2X2_1248 ( .A(_abc_43815_n650_bF_buf0), .B(_abc_43815_n3941), .Y(_abc_43815_n3942) );
  OR2X2 OR2X2_1249 ( .A(_abc_43815_n3940), .B(_abc_43815_n3942), .Y(_abc_43815_n3943) );
  OR2X2 OR2X2_125 ( .A(_abc_43815_n946), .B(_abc_43815_n885_1), .Y(_abc_43815_n947) );
  OR2X2 OR2X2_1250 ( .A(_abc_43815_n3944), .B(_abc_43815_n641_bF_buf3), .Y(_abc_43815_n3945_1) );
  OR2X2 OR2X2_1251 ( .A(_abc_43815_n3947), .B(_abc_43815_n3934), .Y(mem_dat_o_30__FF_INPUT) );
  OR2X2 OR2X2_1252 ( .A(_abc_43815_n3834), .B(_abc_43815_n642_1_bF_buf5), .Y(_abc_43815_n3950) );
  OR2X2 OR2X2_1253 ( .A(_abc_43815_n3951_1), .B(_abc_43815_n3952), .Y(_abc_43815_n3953) );
  OR2X2 OR2X2_1254 ( .A(_abc_43815_n3953), .B(_abc_43815_n649_bF_buf1), .Y(_abc_43815_n3954) );
  OR2X2 OR2X2_1255 ( .A(_abc_43815_n650_bF_buf4), .B(_abc_43815_n3956), .Y(_abc_43815_n3957) );
  OR2X2 OR2X2_1256 ( .A(_abc_43815_n3955), .B(_abc_43815_n3957), .Y(_abc_43815_n3958_1) );
  OR2X2 OR2X2_1257 ( .A(_abc_43815_n3959), .B(_abc_43815_n641_bF_buf2), .Y(_abc_43815_n3960) );
  OR2X2 OR2X2_1258 ( .A(_abc_43815_n3962), .B(_abc_43815_n3949), .Y(mem_dat_o_31__FF_INPUT) );
  OR2X2 OR2X2_1259 ( .A(_abc_43815_n3965), .B(_auto_iopadmap_cc_313_execute_47809), .Y(_abc_43815_n3966_1) );
  OR2X2 OR2X2_126 ( .A(_abc_43815_n948), .B(_abc_43815_n832_1_bF_buf1), .Y(_abc_43815_n949) );
  OR2X2 OR2X2_1260 ( .A(_abc_43815_n671_bF_buf0), .B(_abc_43815_n3969), .Y(_abc_43815_n3970) );
  OR2X2 OR2X2_1261 ( .A(_abc_43815_n2762), .B(_abc_43815_n3965), .Y(_abc_43815_n3972) );
  OR2X2 OR2X2_1262 ( .A(_abc_43815_n3974), .B(state_q_3_bF_buf3), .Y(_abc_43815_n3975) );
  OR2X2 OR2X2_1263 ( .A(_abc_43815_n3973_1), .B(_abc_43815_n3975), .Y(mem_stb_o_FF_INPUT) );
  OR2X2 OR2X2_1264 ( .A(_abc_43815_n674_1), .B(state_q_5_), .Y(_abc_43815_n3979) );
  OR2X2 OR2X2_1265 ( .A(_abc_43815_n3979), .B(_abc_43815_n3978_1), .Y(_abc_43815_n3980) );
  OR2X2 OR2X2_1266 ( .A(_abc_43815_n3981), .B(state_q_3_bF_buf2), .Y(_abc_43815_n3982) );
  OR2X2 OR2X2_1267 ( .A(_abc_43815_n3973_1), .B(_abc_43815_n3982), .Y(mem_cyc_o_FF_INPUT) );
  OR2X2 OR2X2_1268 ( .A(_abc_43815_n672), .B(_abc_43815_n3968), .Y(_abc_43815_n3985_1) );
  OR2X2 OR2X2_1269 ( .A(_abc_43815_n3986), .B(_abc_43815_n3984), .Y(mem_addr_o_0__FF_INPUT) );
  OR2X2 OR2X2_127 ( .A(state_q_1_bF_buf0), .B(alu_p_o_26_), .Y(_abc_43815_n950) );
  OR2X2 OR2X2_1270 ( .A(_abc_43815_n3989), .B(_abc_43815_n3988), .Y(mem_addr_o_1__FF_INPUT) );
  OR2X2 OR2X2_1271 ( .A(_abc_43815_n3326), .B(_abc_43815_n3321), .Y(_abc_43815_n3991) );
  OR2X2 OR2X2_1272 ( .A(_abc_43815_n3991), .B(_abc_43815_n3994), .Y(_abc_43815_n3997) );
  OR2X2 OR2X2_1273 ( .A(_abc_43815_n3999), .B(_abc_43815_n4000), .Y(_abc_43815_n4001) );
  OR2X2 OR2X2_1274 ( .A(_abc_43815_n4003), .B(_abc_43815_n4004), .Y(_abc_43815_n4005) );
  OR2X2 OR2X2_1275 ( .A(_abc_43815_n4002_1), .B(_abc_43815_n4005), .Y(mem_addr_o_2__FF_INPUT) );
  OR2X2 OR2X2_1276 ( .A(_abc_43815_n3995_1), .B(_abc_43815_n3992), .Y(_abc_43815_n4009) );
  OR2X2 OR2X2_1277 ( .A(_abc_43815_n4009), .B(_abc_43815_n4012), .Y(_abc_43815_n4013) );
  OR2X2 OR2X2_1278 ( .A(_abc_43815_n4014), .B(_abc_43815_n4015_1), .Y(_abc_43815_n4016) );
  OR2X2 OR2X2_1279 ( .A(_abc_43815_n4018), .B(_abc_43815_n4008_1), .Y(_abc_43815_n4019) );
  OR2X2 OR2X2_128 ( .A(_abc_43815_n952), .B(_abc_43815_n885_1), .Y(_abc_43815_n953) );
  OR2X2 OR2X2_1280 ( .A(_abc_43815_n4019), .B(_abc_43815_n4007), .Y(mem_addr_o_3__FF_INPUT) );
  OR2X2 OR2X2_1281 ( .A(_abc_43815_n4024), .B(_abc_43815_n4010), .Y(_abc_43815_n4025) );
  OR2X2 OR2X2_1282 ( .A(_abc_43815_n4025), .B(_abc_43815_n4023), .Y(_abc_43815_n4028) );
  OR2X2 OR2X2_1283 ( .A(_abc_43815_n4030), .B(_abc_43815_n4031), .Y(_abc_43815_n4032) );
  OR2X2 OR2X2_1284 ( .A(_abc_43815_n4034_1), .B(_abc_43815_n4035), .Y(_abc_43815_n4036) );
  OR2X2 OR2X2_1285 ( .A(_abc_43815_n4033), .B(_abc_43815_n4036), .Y(mem_addr_o_4__FF_INPUT) );
  OR2X2 OR2X2_1286 ( .A(_abc_43815_n4026), .B(_abc_43815_n4021), .Y(_abc_43815_n4038) );
  OR2X2 OR2X2_1287 ( .A(_abc_43815_n4045), .B(_abc_43815_n4043), .Y(_abc_43815_n4046) );
  OR2X2 OR2X2_1288 ( .A(_abc_43815_n4049), .B(_abc_43815_n4048), .Y(_abc_43815_n4050) );
  OR2X2 OR2X2_1289 ( .A(_abc_43815_n4047), .B(_abc_43815_n4050), .Y(mem_addr_o_5__FF_INPUT) );
  OR2X2 OR2X2_129 ( .A(_abc_43815_n954), .B(_abc_43815_n832_1_bF_buf0), .Y(_abc_43815_n955_1) );
  OR2X2 OR2X2_1290 ( .A(_abc_43815_n4055_1), .B(_abc_43815_n4039), .Y(_abc_43815_n4056) );
  OR2X2 OR2X2_1291 ( .A(_abc_43815_n4056), .B(_abc_43815_n4054), .Y(_abc_43815_n4057) );
  OR2X2 OR2X2_1292 ( .A(_abc_43815_n4063), .B(_abc_43815_n4062_1), .Y(_abc_43815_n4064) );
  OR2X2 OR2X2_1293 ( .A(_abc_43815_n4061), .B(_abc_43815_n4064), .Y(mem_addr_o_6__FF_INPUT) );
  OR2X2 OR2X2_1294 ( .A(_abc_43815_n4066), .B(_abc_43815_n4070), .Y(_abc_43815_n4071) );
  OR2X2 OR2X2_1295 ( .A(_abc_43815_n4072), .B(_abc_43815_n4069), .Y(_abc_43815_n4073) );
  OR2X2 OR2X2_1296 ( .A(_abc_43815_n4077), .B(_abc_43815_n4076), .Y(_abc_43815_n4078) );
  OR2X2 OR2X2_1297 ( .A(_abc_43815_n4075_1), .B(_abc_43815_n4078), .Y(mem_addr_o_7__FF_INPUT) );
  OR2X2 OR2X2_1298 ( .A(_abc_43815_n4080), .B(_abc_43815_n4081), .Y(_abc_43815_n4082_1) );
  OR2X2 OR2X2_1299 ( .A(_abc_43815_n4058), .B(_abc_43815_n4085), .Y(_abc_43815_n4086) );
  OR2X2 OR2X2_13 ( .A(_abc_43815_n701), .B(_abc_43815_n702), .Y(_abc_43815_n703) );
  OR2X2 OR2X2_130 ( .A(state_q_1_bF_buf4), .B(alu_p_o_27_), .Y(_abc_43815_n956_1) );
  OR2X2 OR2X2_1300 ( .A(_abc_43815_n4087), .B(_abc_43815_n4083), .Y(_abc_43815_n4088) );
  OR2X2 OR2X2_1301 ( .A(_abc_43815_n4094_1), .B(_abc_43815_n4093), .Y(_abc_43815_n4095) );
  OR2X2 OR2X2_1302 ( .A(_abc_43815_n4092), .B(_abc_43815_n4095), .Y(mem_addr_o_8__FF_INPUT) );
  OR2X2 OR2X2_1303 ( .A(_abc_43815_n4098), .B(_abc_43815_n4102), .Y(_abc_43815_n4103) );
  OR2X2 OR2X2_1304 ( .A(_abc_43815_n4104), .B(_abc_43815_n4101_1), .Y(_abc_43815_n4105) );
  OR2X2 OR2X2_1305 ( .A(_abc_43815_n4109), .B(_abc_43815_n4108), .Y(_abc_43815_n4110) );
  OR2X2 OR2X2_1306 ( .A(_abc_43815_n4107), .B(_abc_43815_n4110), .Y(mem_addr_o_9__FF_INPUT) );
  OR2X2 OR2X2_1307 ( .A(_abc_43815_n4114), .B(_abc_43815_n1213), .Y(_abc_43815_n4115) );
  OR2X2 OR2X2_1308 ( .A(_abc_43815_n4113), .B(_abc_43815_n4116), .Y(_abc_43815_n4117) );
  OR2X2 OR2X2_1309 ( .A(_abc_43815_n4118), .B(_abc_43815_n4119_1), .Y(_abc_43815_n4120) );
  OR2X2 OR2X2_131 ( .A(_abc_43815_n958), .B(_abc_43815_n885_1), .Y(_abc_43815_n959) );
  OR2X2 OR2X2_1310 ( .A(_abc_43815_n4117), .B(_abc_43815_n4121), .Y(_abc_43815_n4122) );
  OR2X2 OR2X2_1311 ( .A(_abc_43815_n4128), .B(_abc_43815_n4127), .Y(_abc_43815_n4129) );
  OR2X2 OR2X2_1312 ( .A(_abc_43815_n4126), .B(_abc_43815_n4129), .Y(mem_addr_o_10__FF_INPUT) );
  OR2X2 OR2X2_1313 ( .A(_abc_43815_n4134), .B(_abc_43815_n4133), .Y(_abc_43815_n4135) );
  OR2X2 OR2X2_1314 ( .A(_abc_43815_n4135), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_43815_n4138_1) );
  OR2X2 OR2X2_1315 ( .A(_abc_43815_n4132), .B(_abc_43815_n4140), .Y(_abc_43815_n4141) );
  OR2X2 OR2X2_1316 ( .A(_abc_43815_n4142), .B(_abc_43815_n4139), .Y(_abc_43815_n4143) );
  OR2X2 OR2X2_1317 ( .A(_abc_43815_n4147), .B(_abc_43815_n4146), .Y(_abc_43815_n4148) );
  OR2X2 OR2X2_1318 ( .A(_abc_43815_n4145_1), .B(_abc_43815_n4148), .Y(mem_addr_o_11__FF_INPUT) );
  OR2X2 OR2X2_1319 ( .A(_abc_43815_n4151), .B(_abc_43815_n4150_1), .Y(_abc_43815_n4152) );
  OR2X2 OR2X2_132 ( .A(_abc_43815_n960), .B(_abc_43815_n832_1_bF_buf3), .Y(_abc_43815_n961) );
  OR2X2 OR2X2_1320 ( .A(_abc_43815_n4152), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_43815_n4155) );
  OR2X2 OR2X2_1321 ( .A(_abc_43815_n4160), .B(_abc_43815_n4136), .Y(_abc_43815_n4161_1) );
  OR2X2 OR2X2_1322 ( .A(_abc_43815_n4162_1), .B(_abc_43815_n4161_1), .Y(_abc_43815_n4163) );
  OR2X2 OR2X2_1323 ( .A(_abc_43815_n4159), .B(_abc_43815_n4163), .Y(_abc_43815_n4164_1) );
  OR2X2 OR2X2_1324 ( .A(_abc_43815_n4164_1), .B(_abc_43815_n4156), .Y(_abc_43815_n4165_1) );
  OR2X2 OR2X2_1325 ( .A(_abc_43815_n4171), .B(_abc_43815_n4170), .Y(_abc_43815_n4172) );
  OR2X2 OR2X2_1326 ( .A(_abc_43815_n4169), .B(_abc_43815_n4172), .Y(mem_addr_o_12__FF_INPUT) );
  OR2X2 OR2X2_1327 ( .A(_abc_43815_n4175), .B(_abc_43815_n4174), .Y(_abc_43815_n4176) );
  OR2X2 OR2X2_1328 ( .A(_abc_43815_n4176), .B(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_43815_n4179) );
  OR2X2 OR2X2_1329 ( .A(_abc_43815_n4180), .B(_abc_43815_n4153), .Y(_abc_43815_n4181) );
  OR2X2 OR2X2_133 ( .A(state_q_1_bF_buf3), .B(alu_p_o_28_), .Y(_abc_43815_n962) );
  OR2X2 OR2X2_1330 ( .A(_abc_43815_n4166_1), .B(_abc_43815_n4181), .Y(_abc_43815_n4182) );
  OR2X2 OR2X2_1331 ( .A(_abc_43815_n4192), .B(_abc_43815_n4191), .Y(_abc_43815_n4193) );
  OR2X2 OR2X2_1332 ( .A(_abc_43815_n4190), .B(_abc_43815_n4193), .Y(mem_addr_o_13__FF_INPUT) );
  OR2X2 OR2X2_1333 ( .A(_abc_43815_n4199), .B(_abc_43815_n4198), .Y(_abc_43815_n4200) );
  OR2X2 OR2X2_1334 ( .A(_abc_43815_n4200), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_43815_n4203) );
  OR2X2 OR2X2_1335 ( .A(_abc_43815_n4197), .B(_abc_43815_n4204), .Y(_abc_43815_n4207) );
  OR2X2 OR2X2_1336 ( .A(_abc_43815_n4211), .B(_abc_43815_n4210), .Y(_abc_43815_n4212) );
  OR2X2 OR2X2_1337 ( .A(_abc_43815_n4209), .B(_abc_43815_n4212), .Y(mem_addr_o_14__FF_INPUT) );
  OR2X2 OR2X2_1338 ( .A(_abc_43815_n4216), .B(_abc_43815_n4215), .Y(_abc_43815_n4217) );
  OR2X2 OR2X2_1339 ( .A(_abc_43815_n4214), .B(_abc_43815_n4224), .Y(_abc_43815_n4225) );
  OR2X2 OR2X2_134 ( .A(_abc_43815_n964_1), .B(_abc_43815_n885_1), .Y(_abc_43815_n965) );
  OR2X2 OR2X2_1340 ( .A(_abc_43815_n4226), .B(_abc_43815_n4223), .Y(_abc_43815_n4227) );
  OR2X2 OR2X2_1341 ( .A(_abc_43815_n4231), .B(_abc_43815_n4230), .Y(_abc_43815_n4232) );
  OR2X2 OR2X2_1342 ( .A(_abc_43815_n4229), .B(_abc_43815_n4232), .Y(mem_addr_o_15__FF_INPUT) );
  OR2X2 OR2X2_1343 ( .A(_abc_43815_n4195), .B(_abc_43815_n4235), .Y(_abc_43815_n4236) );
  OR2X2 OR2X2_1344 ( .A(_abc_43815_n4237), .B(_abc_43815_n4218), .Y(_abc_43815_n4238) );
  OR2X2 OR2X2_1345 ( .A(_abc_43815_n4243), .B(_abc_43815_n4241), .Y(_abc_43815_n4244) );
  OR2X2 OR2X2_1346 ( .A(_abc_43815_n4217_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_43815_n4247) );
  OR2X2 OR2X2_1347 ( .A(_abc_43815_n4244), .B(_abc_43815_n4248), .Y(_abc_43815_n4249) );
  OR2X2 OR2X2_1348 ( .A(_abc_43815_n4255), .B(_abc_43815_n4254), .Y(_abc_43815_n4256) );
  OR2X2 OR2X2_1349 ( .A(_abc_43815_n4253), .B(_abc_43815_n4256), .Y(mem_addr_o_16__FF_INPUT) );
  OR2X2 OR2X2_135 ( .A(_abc_43815_n966), .B(_abc_43815_n832_1_bF_buf2), .Y(_abc_43815_n967) );
  OR2X2 OR2X2_1350 ( .A(_abc_43815_n4217_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_43815_n4261) );
  OR2X2 OR2X2_1351 ( .A(_abc_43815_n4258), .B(_abc_43815_n4263), .Y(_abc_43815_n4264) );
  OR2X2 OR2X2_1352 ( .A(_abc_43815_n4265), .B(_abc_43815_n4262), .Y(_abc_43815_n4266) );
  OR2X2 OR2X2_1353 ( .A(_abc_43815_n4270), .B(_abc_43815_n4269), .Y(_abc_43815_n4271) );
  OR2X2 OR2X2_1354 ( .A(_abc_43815_n4268), .B(_abc_43815_n4271), .Y(mem_addr_o_17__FF_INPUT) );
  OR2X2 OR2X2_1355 ( .A(_abc_43815_n4217_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_43815_n4275) );
  OR2X2 OR2X2_1356 ( .A(_abc_43815_n4280), .B(_abc_43815_n4278), .Y(_abc_43815_n4281) );
  OR2X2 OR2X2_1357 ( .A(_abc_43815_n4281), .B(_abc_43815_n4276), .Y(_abc_43815_n4282) );
  OR2X2 OR2X2_1358 ( .A(_abc_43815_n4288), .B(_abc_43815_n4287), .Y(_abc_43815_n4289) );
  OR2X2 OR2X2_1359 ( .A(_abc_43815_n4286), .B(_abc_43815_n4289), .Y(mem_addr_o_18__FF_INPUT) );
  OR2X2 OR2X2_136 ( .A(state_q_1_bF_buf2), .B(alu_p_o_29_), .Y(_abc_43815_n968) );
  OR2X2 OR2X2_1360 ( .A(_abc_43815_n4217_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_43815_n4294) );
  OR2X2 OR2X2_1361 ( .A(_abc_43815_n4291), .B(_abc_43815_n4296), .Y(_abc_43815_n4297) );
  OR2X2 OR2X2_1362 ( .A(_abc_43815_n4298), .B(_abc_43815_n4295), .Y(_abc_43815_n4299) );
  OR2X2 OR2X2_1363 ( .A(_abc_43815_n4303), .B(_abc_43815_n4302), .Y(_abc_43815_n4304) );
  OR2X2 OR2X2_1364 ( .A(_abc_43815_n4301), .B(_abc_43815_n4304), .Y(mem_addr_o_19__FF_INPUT) );
  OR2X2 OR2X2_1365 ( .A(_abc_43815_n4308), .B(_abc_43815_n4313), .Y(_abc_43815_n4314) );
  OR2X2 OR2X2_1366 ( .A(_abc_43815_n4217_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_43815_n4317) );
  OR2X2 OR2X2_1367 ( .A(_abc_43815_n4314), .B(_abc_43815_n4318), .Y(_abc_43815_n4319) );
  OR2X2 OR2X2_1368 ( .A(_abc_43815_n4325), .B(_abc_43815_n4324), .Y(_abc_43815_n4326) );
  OR2X2 OR2X2_1369 ( .A(_abc_43815_n4323), .B(_abc_43815_n4326), .Y(mem_addr_o_20__FF_INPUT) );
  OR2X2 OR2X2_137 ( .A(_abc_43815_n970), .B(_abc_43815_n885_1), .Y(_abc_43815_n971) );
  OR2X2 OR2X2_1370 ( .A(_abc_43815_n4217_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_43815_n4331) );
  OR2X2 OR2X2_1371 ( .A(_abc_43815_n4328), .B(_abc_43815_n4333), .Y(_abc_43815_n4334) );
  OR2X2 OR2X2_1372 ( .A(_abc_43815_n4335), .B(_abc_43815_n4332), .Y(_abc_43815_n4336) );
  OR2X2 OR2X2_1373 ( .A(_abc_43815_n4340), .B(_abc_43815_n4339), .Y(_abc_43815_n4341) );
  OR2X2 OR2X2_1374 ( .A(_abc_43815_n4338), .B(_abc_43815_n4341), .Y(mem_addr_o_21__FF_INPUT) );
  OR2X2 OR2X2_1375 ( .A(_abc_43815_n4315), .B(_abc_43815_n4329), .Y(_abc_43815_n4343) );
  OR2X2 OR2X2_1376 ( .A(_abc_43815_n4345), .B(_abc_43815_n4343), .Y(_abc_43815_n4346) );
  OR2X2 OR2X2_1377 ( .A(_abc_43815_n4217_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_43815_n4349) );
  OR2X2 OR2X2_1378 ( .A(_abc_43815_n4346), .B(_abc_43815_n4350), .Y(_abc_43815_n4351) );
  OR2X2 OR2X2_1379 ( .A(_abc_43815_n4357), .B(_abc_43815_n4356), .Y(_abc_43815_n4358) );
  OR2X2 OR2X2_138 ( .A(_abc_43815_n972), .B(_abc_43815_n832_1_bF_buf1), .Y(_abc_43815_n973) );
  OR2X2 OR2X2_1380 ( .A(_abc_43815_n4355), .B(_abc_43815_n4358), .Y(mem_addr_o_22__FF_INPUT) );
  OR2X2 OR2X2_1381 ( .A(_abc_43815_n4217_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_43815_n4364) );
  OR2X2 OR2X2_1382 ( .A(_abc_43815_n4361), .B(_abc_43815_n4365), .Y(_abc_43815_n4366) );
  OR2X2 OR2X2_1383 ( .A(_abc_43815_n4360), .B(_abc_43815_n4367), .Y(_abc_43815_n4368) );
  OR2X2 OR2X2_1384 ( .A(_abc_43815_n4372), .B(_abc_43815_n4371), .Y(_abc_43815_n4373) );
  OR2X2 OR2X2_1385 ( .A(_abc_43815_n4370), .B(_abc_43815_n4373), .Y(mem_addr_o_23__FF_INPUT) );
  OR2X2 OR2X2_1386 ( .A(_abc_43815_n4382), .B(_abc_43815_n4380), .Y(_abc_43815_n4383) );
  OR2X2 OR2X2_1387 ( .A(_abc_43815_n4217_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_43815_n4386) );
  OR2X2 OR2X2_1388 ( .A(_abc_43815_n4383), .B(_abc_43815_n4387), .Y(_abc_43815_n4388) );
  OR2X2 OR2X2_1389 ( .A(_abc_43815_n4394), .B(_abc_43815_n4393), .Y(_abc_43815_n4395) );
  OR2X2 OR2X2_139 ( .A(state_q_1_bF_buf1), .B(alu_p_o_30_), .Y(_abc_43815_n974) );
  OR2X2 OR2X2_1390 ( .A(_abc_43815_n4392), .B(_abc_43815_n4395), .Y(mem_addr_o_24__FF_INPUT) );
  OR2X2 OR2X2_1391 ( .A(_abc_43815_n4217_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_43815_n4400) );
  OR2X2 OR2X2_1392 ( .A(_abc_43815_n4397), .B(_abc_43815_n4402), .Y(_abc_43815_n4403) );
  OR2X2 OR2X2_1393 ( .A(_abc_43815_n4404), .B(_abc_43815_n4401), .Y(_abc_43815_n4405) );
  OR2X2 OR2X2_1394 ( .A(_abc_43815_n4409), .B(_abc_43815_n4408), .Y(_abc_43815_n4410) );
  OR2X2 OR2X2_1395 ( .A(_abc_43815_n4407), .B(_abc_43815_n4410), .Y(mem_addr_o_25__FF_INPUT) );
  OR2X2 OR2X2_1396 ( .A(_abc_43815_n4413), .B(_abc_43815_n4415), .Y(_abc_43815_n4416) );
  OR2X2 OR2X2_1397 ( .A(_abc_43815_n4217_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_43815_n4419) );
  OR2X2 OR2X2_1398 ( .A(_abc_43815_n4416), .B(_abc_43815_n4420), .Y(_abc_43815_n4421) );
  OR2X2 OR2X2_1399 ( .A(_abc_43815_n4427), .B(_abc_43815_n4426), .Y(_abc_43815_n4428) );
  OR2X2 OR2X2_14 ( .A(_abc_43815_n705), .B(_abc_43815_n707_1), .Y(_abc_43815_n708) );
  OR2X2 OR2X2_140 ( .A(_abc_43815_n976), .B(_abc_43815_n885_1), .Y(_abc_43815_n977) );
  OR2X2 OR2X2_1400 ( .A(_abc_43815_n4425), .B(_abc_43815_n4428), .Y(mem_addr_o_26__FF_INPUT) );
  OR2X2 OR2X2_1401 ( .A(_abc_43815_n4217_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_43815_n4433) );
  OR2X2 OR2X2_1402 ( .A(_abc_43815_n4430), .B(_abc_43815_n4435), .Y(_abc_43815_n4436) );
  OR2X2 OR2X2_1403 ( .A(_abc_43815_n4437), .B(_abc_43815_n4434), .Y(_abc_43815_n4438) );
  OR2X2 OR2X2_1404 ( .A(_abc_43815_n4442), .B(_abc_43815_n4441), .Y(_abc_43815_n4443) );
  OR2X2 OR2X2_1405 ( .A(_abc_43815_n4440), .B(_abc_43815_n4443), .Y(mem_addr_o_27__FF_INPUT) );
  OR2X2 OR2X2_1406 ( .A(_abc_43815_n4446), .B(_abc_43815_n4448), .Y(_abc_43815_n4449) );
  OR2X2 OR2X2_1407 ( .A(_abc_43815_n4445), .B(_abc_43815_n4449), .Y(_abc_43815_n4450) );
  OR2X2 OR2X2_1408 ( .A(_abc_43815_n4459), .B(_abc_43815_n4457), .Y(_abc_43815_n4460) );
  OR2X2 OR2X2_1409 ( .A(_abc_43815_n4456), .B(_abc_43815_n4461), .Y(_abc_43815_n4462) );
  OR2X2 OR2X2_141 ( .A(_abc_43815_n978), .B(_abc_43815_n832_1_bF_buf0), .Y(_abc_43815_n979) );
  OR2X2 OR2X2_1410 ( .A(_abc_43815_n4468), .B(_abc_43815_n4467), .Y(_abc_43815_n4469) );
  OR2X2 OR2X2_1411 ( .A(_abc_43815_n4466), .B(_abc_43815_n4469), .Y(mem_addr_o_28__FF_INPUT) );
  OR2X2 OR2X2_1412 ( .A(_abc_43815_n4463), .B(_abc_43815_n4457), .Y(_abc_43815_n4471) );
  OR2X2 OR2X2_1413 ( .A(_abc_43815_n4475), .B(_abc_43815_n4473), .Y(_abc_43815_n4476) );
  OR2X2 OR2X2_1414 ( .A(_abc_43815_n4472), .B(_abc_43815_n4476), .Y(_abc_43815_n4477) );
  OR2X2 OR2X2_1415 ( .A(_abc_43815_n4471), .B(_abc_43815_n4478), .Y(_abc_43815_n4479) );
  OR2X2 OR2X2_1416 ( .A(_abc_43815_n4483), .B(_abc_43815_n4482), .Y(_abc_43815_n4484) );
  OR2X2 OR2X2_1417 ( .A(_abc_43815_n4481), .B(_abc_43815_n4484), .Y(mem_addr_o_29__FF_INPUT) );
  OR2X2 OR2X2_1418 ( .A(_abc_43815_n4217_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_43815_n4488) );
  OR2X2 OR2X2_1419 ( .A(_abc_43815_n4220), .B(_abc_43815_n4490), .Y(_abc_43815_n4491) );
  OR2X2 OR2X2_142 ( .A(state_q_1_bF_buf0), .B(alu_p_o_31_), .Y(_abc_43815_n980) );
  OR2X2 OR2X2_1420 ( .A(_abc_43815_n4455), .B(_abc_43815_n4493), .Y(_abc_43815_n4494) );
  OR2X2 OR2X2_1421 ( .A(_abc_43815_n4496), .B(_abc_43815_n4489), .Y(_abc_43815_n4497) );
  OR2X2 OR2X2_1422 ( .A(_abc_43815_n4495), .B(_abc_43815_n4498), .Y(_abc_43815_n4499) );
  OR2X2 OR2X2_1423 ( .A(_abc_43815_n4503), .B(_abc_43815_n4502), .Y(_abc_43815_n4504) );
  OR2X2 OR2X2_1424 ( .A(_abc_43815_n4501), .B(_abc_43815_n4504), .Y(mem_addr_o_30__FF_INPUT) );
  OR2X2 OR2X2_1425 ( .A(_abc_43815_n4220), .B(_abc_43815_n4507), .Y(_abc_43815_n4508) );
  OR2X2 OR2X2_1426 ( .A(_abc_43815_n4217_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_43815_n4509) );
  OR2X2 OR2X2_1427 ( .A(_abc_43815_n4506), .B(_abc_43815_n4511), .Y(_abc_43815_n4512) );
  OR2X2 OR2X2_1428 ( .A(_abc_43815_n4513), .B(_abc_43815_n4510), .Y(_abc_43815_n4514) );
  OR2X2 OR2X2_1429 ( .A(_abc_43815_n4518), .B(_abc_43815_n4517), .Y(_abc_43815_n4519) );
  OR2X2 OR2X2_143 ( .A(_abc_43815_n617), .B(state_q_4_), .Y(REGFILE_SIM_reg_bank_wr_i) );
  OR2X2 OR2X2_1430 ( .A(_abc_43815_n4516), .B(_abc_43815_n4519), .Y(mem_addr_o_31__FF_INPUT) );
  OR2X2 OR2X2_1431 ( .A(_abc_43815_n1280), .B(_auto_iopadmap_cc_313_execute_47728), .Y(_abc_43815_n4524) );
  OR2X2 OR2X2_1432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2104) );
  OR2X2 OR2X2_1433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2109_1) );
  OR2X2 OR2X2_1434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2114_1) );
  OR2X2 OR2X2_1435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2119) );
  OR2X2 OR2X2_1436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2124_1) );
  OR2X2 OR2X2_1437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2129_1) );
  OR2X2 OR2X2_1438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2134) );
  OR2X2 OR2X2_1439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2139_1) );
  OR2X2 OR2X2_144 ( .A(_abc_43815_n984), .B(_abc_43815_n986_bF_buf4), .Y(_abc_43815_n987) );
  OR2X2 OR2X2_1440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2144_1) );
  OR2X2 OR2X2_1441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2149) );
  OR2X2 OR2X2_1442 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2154_1) );
  OR2X2 OR2X2_1443 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2159_1) );
  OR2X2 OR2X2_1444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2164) );
  OR2X2 OR2X2_1445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2169_1) );
  OR2X2 OR2X2_1446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2174_1) );
  OR2X2 OR2X2_1447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2179) );
  OR2X2 OR2X2_1448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2184_1) );
  OR2X2 OR2X2_1449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2189_1) );
  OR2X2 OR2X2_145 ( .A(opcode_q_24_), .B(opcode_q_23_), .Y(_abc_43815_n993_1) );
  OR2X2 OR2X2_1450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2194) );
  OR2X2 OR2X2_1451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2199) );
  OR2X2 OR2X2_1452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2204) );
  OR2X2 OR2X2_1453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2209_1) );
  OR2X2 OR2X2_1454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2214_1) );
  OR2X2 OR2X2_1455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2219) );
  OR2X2 OR2X2_1456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2224_1) );
  OR2X2 OR2X2_1457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2229_1) );
  OR2X2 OR2X2_1458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2234) );
  OR2X2 OR2X2_1459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2239_1) );
  OR2X2 OR2X2_146 ( .A(_abc_43815_n1001), .B(_abc_43815_n1004), .Y(_abc_43815_n1005) );
  OR2X2 OR2X2_1460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2244_1) );
  OR2X2 OR2X2_1461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2249) );
  OR2X2 OR2X2_1462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2254_1) );
  OR2X2 OR2X2_1463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2103_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2259_1) );
  OR2X2 OR2X2_1464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2268_1) );
  OR2X2 OR2X2_1465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2270) );
  OR2X2 OR2X2_1466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2272_1) );
  OR2X2 OR2X2_1467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2273) );
  OR2X2 OR2X2_1468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2275_1) );
  OR2X2 OR2X2_1469 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2276) );
  OR2X2 OR2X2_147 ( .A(_abc_43815_n1005), .B(_abc_43815_n1000), .Y(_abc_43815_n1006) );
  OR2X2 OR2X2_1470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2278_1) );
  OR2X2 OR2X2_1471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2279) );
  OR2X2 OR2X2_1472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2281_1) );
  OR2X2 OR2X2_1473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2282) );
  OR2X2 OR2X2_1474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2284_1) );
  OR2X2 OR2X2_1475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2285) );
  OR2X2 OR2X2_1476 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2287_1) );
  OR2X2 OR2X2_1477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2288) );
  OR2X2 OR2X2_1478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2290_1) );
  OR2X2 OR2X2_1479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2291) );
  OR2X2 OR2X2_148 ( .A(_abc_43815_n999), .B(_abc_43815_n1006), .Y(_abc_43815_n1007) );
  OR2X2 OR2X2_1480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2293_1) );
  OR2X2 OR2X2_1481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2294) );
  OR2X2 OR2X2_1482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2296) );
  OR2X2 OR2X2_1483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2297_1) );
  OR2X2 OR2X2_1484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2299_1) );
  OR2X2 OR2X2_1485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2300_1) );
  OR2X2 OR2X2_1486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2302_1) );
  OR2X2 OR2X2_1487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2303_1) );
  OR2X2 OR2X2_1488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2305_1) );
  OR2X2 OR2X2_1489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2306_1) );
  OR2X2 OR2X2_149 ( .A(_abc_43815_n988), .B(opcode_q_22_), .Y(_abc_43815_n1009_1) );
  OR2X2 OR2X2_1490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2308_1) );
  OR2X2 OR2X2_1491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2309_1) );
  OR2X2 OR2X2_1492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2311_1) );
  OR2X2 OR2X2_1493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2312_1) );
  OR2X2 OR2X2_1494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2314_1) );
  OR2X2 OR2X2_1495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2315_1) );
  OR2X2 OR2X2_1496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2317_1) );
  OR2X2 OR2X2_1497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2318_1) );
  OR2X2 OR2X2_1498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2320_1) );
  OR2X2 OR2X2_1499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2321_1) );
  OR2X2 OR2X2_15 ( .A(_abc_43815_n703), .B(_abc_43815_n708), .Y(_abc_43815_n709) );
  OR2X2 OR2X2_150 ( .A(_abc_43815_n1004), .B(_abc_43815_n1025), .Y(_abc_43815_n1026) );
  OR2X2 OR2X2_1500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2323_1) );
  OR2X2 OR2X2_1501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2324_1) );
  OR2X2 OR2X2_1502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2326_1) );
  OR2X2 OR2X2_1503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2327_1) );
  OR2X2 OR2X2_1504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2329_1) );
  OR2X2 OR2X2_1505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2330_1) );
  OR2X2 OR2X2_1506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2332_1) );
  OR2X2 OR2X2_1507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2333_1) );
  OR2X2 OR2X2_1508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2335_1) );
  OR2X2 OR2X2_1509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2336_1) );
  OR2X2 OR2X2_151 ( .A(_abc_43815_n1026), .B(_abc_43815_n1000), .Y(_abc_43815_n1027) );
  OR2X2 OR2X2_1510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2338_1) );
  OR2X2 OR2X2_1511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2339_1) );
  OR2X2 OR2X2_1512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2341_1) );
  OR2X2 OR2X2_1513 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2342_1) );
  OR2X2 OR2X2_1514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2344_1) );
  OR2X2 OR2X2_1515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2345_1) );
  OR2X2 OR2X2_1516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2347_1) );
  OR2X2 OR2X2_1517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2348_1) );
  OR2X2 OR2X2_1518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2350_1) );
  OR2X2 OR2X2_1519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2351_1) );
  OR2X2 OR2X2_152 ( .A(_abc_43815_n999), .B(_abc_43815_n1027), .Y(_abc_43815_n1028) );
  OR2X2 OR2X2_1520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2353_1) );
  OR2X2 OR2X2_1521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2354_1) );
  OR2X2 OR2X2_1522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2356_1) );
  OR2X2 OR2X2_1523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2357_1) );
  OR2X2 OR2X2_1524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2359_1) );
  OR2X2 OR2X2_1525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2360_1) );
  OR2X2 OR2X2_1526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2267_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2362_1) );
  OR2X2 OR2X2_1527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2269_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n2363_1) );
  OR2X2 OR2X2_1528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2369_1) );
  OR2X2 OR2X2_1529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2371_1) );
  OR2X2 OR2X2_153 ( .A(_abc_43815_n1025), .B(_abc_43815_n993_1), .Y(_abc_43815_n1029) );
  OR2X2 OR2X2_1530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2373) );
  OR2X2 OR2X2_1531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2374_1) );
  OR2X2 OR2X2_1532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2376) );
  OR2X2 OR2X2_1533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2377_1) );
  OR2X2 OR2X2_1534 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2379) );
  OR2X2 OR2X2_1535 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2380_1) );
  OR2X2 OR2X2_1536 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2382) );
  OR2X2 OR2X2_1537 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2383_1) );
  OR2X2 OR2X2_1538 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2385) );
  OR2X2 OR2X2_1539 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2386_1) );
  OR2X2 OR2X2_154 ( .A(_abc_43815_n1000), .B(_abc_43815_n1029), .Y(_abc_43815_n1030) );
  OR2X2 OR2X2_1540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2388) );
  OR2X2 OR2X2_1541 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2389_1) );
  OR2X2 OR2X2_1542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2391) );
  OR2X2 OR2X2_1543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2392_1) );
  OR2X2 OR2X2_1544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2394_1) );
  OR2X2 OR2X2_1545 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2395) );
  OR2X2 OR2X2_1546 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2397_1) );
  OR2X2 OR2X2_1547 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2398) );
  OR2X2 OR2X2_1548 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2400_1) );
  OR2X2 OR2X2_1549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2401) );
  OR2X2 OR2X2_155 ( .A(_abc_43815_n999), .B(_abc_43815_n1030), .Y(_abc_43815_n1031_1) );
  OR2X2 OR2X2_1550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2403_1) );
  OR2X2 OR2X2_1551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2404) );
  OR2X2 OR2X2_1552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2406_1) );
  OR2X2 OR2X2_1553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2407) );
  OR2X2 OR2X2_1554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2409_1) );
  OR2X2 OR2X2_1555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2410) );
  OR2X2 OR2X2_1556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2412_1) );
  OR2X2 OR2X2_1557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2413) );
  OR2X2 OR2X2_1558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2415_1) );
  OR2X2 OR2X2_1559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2416) );
  OR2X2 OR2X2_156 ( .A(_abc_43815_n1035), .B(_abc_43815_n993_1), .Y(_abc_43815_n1036) );
  OR2X2 OR2X2_1560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2418_1) );
  OR2X2 OR2X2_1561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2419) );
  OR2X2 OR2X2_1562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2421_1) );
  OR2X2 OR2X2_1563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2422) );
  OR2X2 OR2X2_1564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2424_1) );
  OR2X2 OR2X2_1565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2425) );
  OR2X2 OR2X2_1566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2427_1) );
  OR2X2 OR2X2_1567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2428) );
  OR2X2 OR2X2_1568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2430_1) );
  OR2X2 OR2X2_1569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2431) );
  OR2X2 OR2X2_157 ( .A(_abc_43815_n1036), .B(_abc_43815_n1000), .Y(_abc_43815_n1037) );
  OR2X2 OR2X2_1570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2433_1) );
  OR2X2 OR2X2_1571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2434) );
  OR2X2 OR2X2_1572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2436_1) );
  OR2X2 OR2X2_1573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2437) );
  OR2X2 OR2X2_1574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2439_1) );
  OR2X2 OR2X2_1575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2440) );
  OR2X2 OR2X2_1576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2442_1) );
  OR2X2 OR2X2_1577 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2443) );
  OR2X2 OR2X2_1578 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2445_1) );
  OR2X2 OR2X2_1579 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2446) );
  OR2X2 OR2X2_158 ( .A(_abc_43815_n999), .B(_abc_43815_n1037), .Y(_abc_43815_n1038) );
  OR2X2 OR2X2_1580 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2448_1) );
  OR2X2 OR2X2_1581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2449) );
  OR2X2 OR2X2_1582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2451_1) );
  OR2X2 OR2X2_1583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2452) );
  OR2X2 OR2X2_1584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2454_1) );
  OR2X2 OR2X2_1585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2455) );
  OR2X2 OR2X2_1586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2457_1) );
  OR2X2 OR2X2_1587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2458) );
  OR2X2 OR2X2_1588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2460_1) );
  OR2X2 OR2X2_1589 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2461) );
  OR2X2 OR2X2_159 ( .A(_abc_43815_n690), .B(_abc_43815_n1041), .Y(_abc_43815_n1042) );
  OR2X2 OR2X2_1590 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2368_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2463_1) );
  OR2X2 OR2X2_1591 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2370_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n2464) );
  OR2X2 OR2X2_1592 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2469_1) );
  OR2X2 OR2X2_1593 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2473) );
  OR2X2 OR2X2_1594 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2477_1) );
  OR2X2 OR2X2_1595 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2481_1) );
  OR2X2 OR2X2_1596 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2485) );
  OR2X2 OR2X2_1597 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2489_1) );
  OR2X2 OR2X2_1598 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2493_1) );
  OR2X2 OR2X2_1599 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2497_1) );
  OR2X2 OR2X2_16 ( .A(_abc_43815_n700), .B(_abc_43815_n710), .Y(_abc_43815_n711) );
  OR2X2 OR2X2_160 ( .A(_abc_43815_n1055), .B(_abc_43815_n1054), .Y(_abc_43815_n1056) );
  OR2X2 OR2X2_1600 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2501) );
  OR2X2 OR2X2_1601 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2505_1) );
  OR2X2 OR2X2_1602 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2509_1) );
  OR2X2 OR2X2_1603 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2513) );
  OR2X2 OR2X2_1604 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2517_1) );
  OR2X2 OR2X2_1605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2521_1) );
  OR2X2 OR2X2_1606 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2525) );
  OR2X2 OR2X2_1607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2529_1) );
  OR2X2 OR2X2_1608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2533_1) );
  OR2X2 OR2X2_1609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2537) );
  OR2X2 OR2X2_161 ( .A(_abc_43815_n1035), .B(_abc_43815_n1086_1), .Y(_abc_43815_n1087) );
  OR2X2 OR2X2_1610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2541_1) );
  OR2X2 OR2X2_1611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2545_1) );
  OR2X2 OR2X2_1612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2549) );
  OR2X2 OR2X2_1613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2553_1) );
  OR2X2 OR2X2_1614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2557_1) );
  OR2X2 OR2X2_1615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2561) );
  OR2X2 OR2X2_1616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2565_1) );
  OR2X2 OR2X2_1617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2569_1) );
  OR2X2 OR2X2_1618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2573) );
  OR2X2 OR2X2_1619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2577_1) );
  OR2X2 OR2X2_162 ( .A(_abc_43815_n1087), .B(_abc_43815_n1000), .Y(_abc_43815_n1088) );
  OR2X2 OR2X2_1620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2581_1) );
  OR2X2 OR2X2_1621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2585) );
  OR2X2 OR2X2_1622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2589) );
  OR2X2 OR2X2_1623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2468_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2593_1) );
  OR2X2 OR2X2_1624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2601) );
  OR2X2 OR2X2_1625 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2603_1) );
  OR2X2 OR2X2_1626 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2605_1) );
  OR2X2 OR2X2_1627 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2606_1) );
  OR2X2 OR2X2_1628 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2608_1) );
  OR2X2 OR2X2_1629 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2609_1) );
  OR2X2 OR2X2_163 ( .A(_abc_43815_n999), .B(_abc_43815_n1088), .Y(_abc_43815_n1089) );
  OR2X2 OR2X2_1630 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2611_1) );
  OR2X2 OR2X2_1631 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2612_1) );
  OR2X2 OR2X2_1632 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2614_1) );
  OR2X2 OR2X2_1633 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2615_1) );
  OR2X2 OR2X2_1634 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2617_1) );
  OR2X2 OR2X2_1635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2618_1) );
  OR2X2 OR2X2_1636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2620_1) );
  OR2X2 OR2X2_1637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2621_1) );
  OR2X2 OR2X2_1638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2623_1) );
  OR2X2 OR2X2_1639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2624_1) );
  OR2X2 OR2X2_164 ( .A(_abc_43815_n1035), .B(_abc_43815_n1090), .Y(_abc_43815_n1091) );
  OR2X2 OR2X2_1640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2626_1) );
  OR2X2 OR2X2_1641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2627_1) );
  OR2X2 OR2X2_1642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2629_1) );
  OR2X2 OR2X2_1643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2630_1) );
  OR2X2 OR2X2_1644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2632_1) );
  OR2X2 OR2X2_1645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2633_1) );
  OR2X2 OR2X2_1646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2635_1) );
  OR2X2 OR2X2_1647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2636_1) );
  OR2X2 OR2X2_1648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2638_1) );
  OR2X2 OR2X2_1649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2639_1) );
  OR2X2 OR2X2_165 ( .A(_abc_43815_n1091), .B(_abc_43815_n1000), .Y(_abc_43815_n1092) );
  OR2X2 OR2X2_1650 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2641_1) );
  OR2X2 OR2X2_1651 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2642_1) );
  OR2X2 OR2X2_1652 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2644_1) );
  OR2X2 OR2X2_1653 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2645_1) );
  OR2X2 OR2X2_1654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2647_1) );
  OR2X2 OR2X2_1655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2648_1) );
  OR2X2 OR2X2_1656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2650_1) );
  OR2X2 OR2X2_1657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2651_1) );
  OR2X2 OR2X2_1658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2653_1) );
  OR2X2 OR2X2_1659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2654_1) );
  OR2X2 OR2X2_166 ( .A(_abc_43815_n999), .B(_abc_43815_n1092), .Y(_abc_43815_n1093) );
  OR2X2 OR2X2_1660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2656_1) );
  OR2X2 OR2X2_1661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2657_1) );
  OR2X2 OR2X2_1662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2659_1) );
  OR2X2 OR2X2_1663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2660_1) );
  OR2X2 OR2X2_1664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2662_1) );
  OR2X2 OR2X2_1665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2663_1) );
  OR2X2 OR2X2_1666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2665_1) );
  OR2X2 OR2X2_1667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2666_1) );
  OR2X2 OR2X2_1668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2668_1) );
  OR2X2 OR2X2_1669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2669_1) );
  OR2X2 OR2X2_167 ( .A(inst_trap_w), .B(_abc_43815_n1096), .Y(_abc_43815_n1097) );
  OR2X2 OR2X2_1670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2671_1) );
  OR2X2 OR2X2_1671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2672_1) );
  OR2X2 OR2X2_1672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2674_1) );
  OR2X2 OR2X2_1673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2675_1) );
  OR2X2 OR2X2_1674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2677_1) );
  OR2X2 OR2X2_1675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2678_1) );
  OR2X2 OR2X2_1676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2680_1) );
  OR2X2 OR2X2_1677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2681_1) );
  OR2X2 OR2X2_1678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2683_1) );
  OR2X2 OR2X2_1679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2684) );
  OR2X2 OR2X2_168 ( .A(_abc_43815_n1009_1), .B(_abc_43815_n993_1), .Y(_abc_43815_n1099) );
  OR2X2 OR2X2_1680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2686) );
  OR2X2 OR2X2_1681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2687_1) );
  OR2X2 OR2X2_1682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2689) );
  OR2X2 OR2X2_1683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2690_1) );
  OR2X2 OR2X2_1684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2692) );
  OR2X2 OR2X2_1685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2693_1) );
  OR2X2 OR2X2_1686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2600_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2695) );
  OR2X2 OR2X2_1687 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2602_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n2696_1) );
  OR2X2 OR2X2_1688 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2700_1) );
  OR2X2 OR2X2_1689 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2704) );
  OR2X2 OR2X2_169 ( .A(_abc_43815_n1000), .B(_abc_43815_n1099), .Y(_abc_43815_n1100) );
  OR2X2 OR2X2_1690 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2708_1) );
  OR2X2 OR2X2_1691 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2712_1) );
  OR2X2 OR2X2_1692 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2716) );
  OR2X2 OR2X2_1693 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2720_1) );
  OR2X2 OR2X2_1694 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2724_1) );
  OR2X2 OR2X2_1695 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2728) );
  OR2X2 OR2X2_1696 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2732_1) );
  OR2X2 OR2X2_1697 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2736_1) );
  OR2X2 OR2X2_1698 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2740) );
  OR2X2 OR2X2_1699 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2744_1) );
  OR2X2 OR2X2_17 ( .A(_abc_43815_n712), .B(_abc_43815_n683), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_) );
  OR2X2 OR2X2_170 ( .A(_abc_43815_n999), .B(_abc_43815_n1100), .Y(_abc_43815_n1101) );
  OR2X2 OR2X2_1700 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2748_1) );
  OR2X2 OR2X2_1701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2752) );
  OR2X2 OR2X2_1702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2756_1) );
  OR2X2 OR2X2_1703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2760_1) );
  OR2X2 OR2X2_1704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2764) );
  OR2X2 OR2X2_1705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2768_1) );
  OR2X2 OR2X2_1706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2772_1) );
  OR2X2 OR2X2_1707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2776) );
  OR2X2 OR2X2_1708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2780_1) );
  OR2X2 OR2X2_1709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2784_1) );
  OR2X2 OR2X2_171 ( .A(_abc_43815_n1140), .B(_abc_43815_n1136_1), .Y(_abc_43815_n1141) );
  OR2X2 OR2X2_1710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2788_1) );
  OR2X2 OR2X2_1711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2792) );
  OR2X2 OR2X2_1712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2796_1) );
  OR2X2 OR2X2_1713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2800_1) );
  OR2X2 OR2X2_1714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2804) );
  OR2X2 OR2X2_1715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2808_1) );
  OR2X2 OR2X2_1716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2812_1) );
  OR2X2 OR2X2_1717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2816) );
  OR2X2 OR2X2_1718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2820_1) );
  OR2X2 OR2X2_1719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2699_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2824_1) );
  OR2X2 OR2X2_172 ( .A(_abc_43815_n1145), .B(_abc_43815_n1146), .Y(_abc_43815_n1147) );
  OR2X2 OR2X2_1720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2830_1) );
  OR2X2 OR2X2_1721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2834) );
  OR2X2 OR2X2_1722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2838_1) );
  OR2X2 OR2X2_1723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2842_1) );
  OR2X2 OR2X2_1724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2846) );
  OR2X2 OR2X2_1725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2850_1) );
  OR2X2 OR2X2_1726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2854_1) );
  OR2X2 OR2X2_1727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2858) );
  OR2X2 OR2X2_1728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2862_1) );
  OR2X2 OR2X2_1729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2866_1) );
  OR2X2 OR2X2_173 ( .A(_abc_43815_n1147), .B(_abc_43815_n1144), .Y(_abc_43815_n1148) );
  OR2X2 OR2X2_1730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2870) );
  OR2X2 OR2X2_1731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2874_1) );
  OR2X2 OR2X2_1732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2878) );
  OR2X2 OR2X2_1733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2882_1) );
  OR2X2 OR2X2_1734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2886) );
  OR2X2 OR2X2_1735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2890_1) );
  OR2X2 OR2X2_1736 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2894_1) );
  OR2X2 OR2X2_1737 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2898) );
  OR2X2 OR2X2_1738 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2902_1) );
  OR2X2 OR2X2_1739 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2906_1) );
  OR2X2 OR2X2_174 ( .A(_abc_43815_n1148), .B(_abc_43815_n1136_1), .Y(_abc_43815_n1149) );
  OR2X2 OR2X2_1740 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2910) );
  OR2X2 OR2X2_1741 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2914_1) );
  OR2X2 OR2X2_1742 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2918_1) );
  OR2X2 OR2X2_1743 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2922) );
  OR2X2 OR2X2_1744 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2926_1) );
  OR2X2 OR2X2_1745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2930_1) );
  OR2X2 OR2X2_1746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2934) );
  OR2X2 OR2X2_1747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2938_1) );
  OR2X2 OR2X2_1748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2942_1) );
  OR2X2 OR2X2_1749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2946) );
  OR2X2 OR2X2_175 ( .A(_abc_43815_n1169), .B(_abc_43815_n1170), .Y(_abc_43815_n1171) );
  OR2X2 OR2X2_1750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2950_1) );
  OR2X2 OR2X2_1751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2829_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2954_1) );
  OR2X2 OR2X2_1752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2959_1) );
  OR2X2 OR2X2_1753 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2961) );
  OR2X2 OR2X2_1754 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2963_1) );
  OR2X2 OR2X2_1755 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2964) );
  OR2X2 OR2X2_1756 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2966_1) );
  OR2X2 OR2X2_1757 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2967) );
  OR2X2 OR2X2_1758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2969_1) );
  OR2X2 OR2X2_1759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2970) );
  OR2X2 OR2X2_176 ( .A(_abc_43815_n1183), .B(_abc_43815_n1184), .Y(_abc_43815_n1185) );
  OR2X2 OR2X2_1760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2972_1) );
  OR2X2 OR2X2_1761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2973) );
  OR2X2 OR2X2_1762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2975) );
  OR2X2 OR2X2_1763 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2976_1) );
  OR2X2 OR2X2_1764 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2978_1) );
  OR2X2 OR2X2_1765 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2979_1) );
  OR2X2 OR2X2_1766 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2981_1) );
  OR2X2 OR2X2_1767 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2982_1) );
  OR2X2 OR2X2_1768 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2984_1) );
  OR2X2 OR2X2_1769 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2985_1) );
  OR2X2 OR2X2_177 ( .A(_abc_43815_n1190), .B(next_pc_r_1_), .Y(_abc_43815_n1191) );
  OR2X2 OR2X2_1770 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2987_1) );
  OR2X2 OR2X2_1771 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2988_1) );
  OR2X2 OR2X2_1772 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2990_1) );
  OR2X2 OR2X2_1773 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2991_1) );
  OR2X2 OR2X2_1774 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2993_1) );
  OR2X2 OR2X2_1775 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2994_1) );
  OR2X2 OR2X2_1776 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2996_1) );
  OR2X2 OR2X2_1777 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n2997_1) );
  OR2X2 OR2X2_1778 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n2999_1) );
  OR2X2 OR2X2_1779 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3000_1) );
  OR2X2 OR2X2_178 ( .A(_abc_43815_n1191), .B(next_pc_r_0_), .Y(_abc_43815_n1192) );
  OR2X2 OR2X2_1780 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3002_1) );
  OR2X2 OR2X2_1781 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3003_1) );
  OR2X2 OR2X2_1782 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3005_1) );
  OR2X2 OR2X2_1783 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3006_1) );
  OR2X2 OR2X2_1784 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3008_1) );
  OR2X2 OR2X2_1785 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3009_1) );
  OR2X2 OR2X2_1786 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3011_1) );
  OR2X2 OR2X2_1787 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3012_1) );
  OR2X2 OR2X2_1788 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3014_1) );
  OR2X2 OR2X2_1789 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3015_1) );
  OR2X2 OR2X2_179 ( .A(nmi_q), .B(nmi_i), .Y(_abc_43815_n1195) );
  OR2X2 OR2X2_1790 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3017_1) );
  OR2X2 OR2X2_1791 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3018_1) );
  OR2X2 OR2X2_1792 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3020_1) );
  OR2X2 OR2X2_1793 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3021_1) );
  OR2X2 OR2X2_1794 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3023_1) );
  OR2X2 OR2X2_1795 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3024_1) );
  OR2X2 OR2X2_1796 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3026_1) );
  OR2X2 OR2X2_1797 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3027_1) );
  OR2X2 OR2X2_1798 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3029_1) );
  OR2X2 OR2X2_1799 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3030_1) );
  OR2X2 OR2X2_18 ( .A(_abc_43815_n716), .B(_abc_43815_n685), .Y(_abc_43815_n717) );
  OR2X2 OR2X2_180 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_9_), .B(alu_op_r_7_), .Y(_abc_43815_n1212) );
  OR2X2 OR2X2_1800 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3032_1) );
  OR2X2 OR2X2_1801 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3033_1) );
  OR2X2 OR2X2_1802 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3035_1) );
  OR2X2 OR2X2_1803 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3036_1) );
  OR2X2 OR2X2_1804 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3038_1) );
  OR2X2 OR2X2_1805 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3039_1) );
  OR2X2 OR2X2_1806 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3041_1) );
  OR2X2 OR2X2_1807 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3042_1) );
  OR2X2 OR2X2_1808 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3044_1) );
  OR2X2 OR2X2_1809 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3045_1) );
  OR2X2 OR2X2_181 ( .A(alu_op_r_2_), .B(REGFILE_SIM_reg_bank_reg_ra_o_2_), .Y(_abc_43815_n1217) );
  OR2X2 OR2X2_1810 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3047_1) );
  OR2X2 OR2X2_1811 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3048_1) );
  OR2X2 OR2X2_1812 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3050_1) );
  OR2X2 OR2X2_1813 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3051_1) );
  OR2X2 OR2X2_1814 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2958_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3053_1) );
  OR2X2 OR2X2_1815 ( .A(REGFILE_SIM_reg_bank__abc_33898_n2960_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3054_1) );
  OR2X2 OR2X2_1816 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3060_1) );
  OR2X2 OR2X2_1817 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3062_1) );
  OR2X2 OR2X2_1818 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3064) );
  OR2X2 OR2X2_1819 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3065_1) );
  OR2X2 OR2X2_182 ( .A(alu_op_r_3_), .B(REGFILE_SIM_reg_bank_reg_ra_o_3_), .Y(_abc_43815_n1219) );
  OR2X2 OR2X2_1820 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3067) );
  OR2X2 OR2X2_1821 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3068_1) );
  OR2X2 OR2X2_1822 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3070) );
  OR2X2 OR2X2_1823 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3071_1) );
  OR2X2 OR2X2_1824 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3073) );
  OR2X2 OR2X2_1825 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3074_1) );
  OR2X2 OR2X2_1826 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3076) );
  OR2X2 OR2X2_1827 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3077_1) );
  OR2X2 OR2X2_1828 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3079_1) );
  OR2X2 OR2X2_1829 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3080) );
  OR2X2 OR2X2_183 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_0_), .B(alu_op_r_0_), .Y(_abc_43815_n1222) );
  OR2X2 OR2X2_1830 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3082) );
  OR2X2 OR2X2_1831 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3083) );
  OR2X2 OR2X2_1832 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3085) );
  OR2X2 OR2X2_1833 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3086) );
  OR2X2 OR2X2_1834 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3088) );
  OR2X2 OR2X2_1835 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3089) );
  OR2X2 OR2X2_1836 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3091) );
  OR2X2 OR2X2_1837 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3092) );
  OR2X2 OR2X2_1838 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3094) );
  OR2X2 OR2X2_1839 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3095) );
  OR2X2 OR2X2_184 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_1_), .B(alu_op_r_1_), .Y(_abc_43815_n1224) );
  OR2X2 OR2X2_1840 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3097) );
  OR2X2 OR2X2_1841 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3098) );
  OR2X2 OR2X2_1842 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3100) );
  OR2X2 OR2X2_1843 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3101) );
  OR2X2 OR2X2_1844 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3103) );
  OR2X2 OR2X2_1845 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3104) );
  OR2X2 OR2X2_1846 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3106) );
  OR2X2 OR2X2_1847 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3107) );
  OR2X2 OR2X2_1848 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3109) );
  OR2X2 OR2X2_1849 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3110) );
  OR2X2 OR2X2_185 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_4_), .B(int32_r_4_), .Y(_abc_43815_n1228) );
  OR2X2 OR2X2_1850 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3112) );
  OR2X2 OR2X2_1851 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3113) );
  OR2X2 OR2X2_1852 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3115) );
  OR2X2 OR2X2_1853 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3116) );
  OR2X2 OR2X2_1854 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3118) );
  OR2X2 OR2X2_1855 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3119) );
  OR2X2 OR2X2_1856 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3121) );
  OR2X2 OR2X2_1857 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3122) );
  OR2X2 OR2X2_1858 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3124) );
  OR2X2 OR2X2_1859 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3125) );
  OR2X2 OR2X2_186 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_7_), .B(alu_op_r_5_), .Y(_abc_43815_n1230_1) );
  OR2X2 OR2X2_1860 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3127) );
  OR2X2 OR2X2_1861 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3128) );
  OR2X2 OR2X2_1862 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3130) );
  OR2X2 OR2X2_1863 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3131) );
  OR2X2 OR2X2_1864 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3133) );
  OR2X2 OR2X2_1865 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3134) );
  OR2X2 OR2X2_1866 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3136) );
  OR2X2 OR2X2_1867 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3137) );
  OR2X2 OR2X2_1868 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3139) );
  OR2X2 OR2X2_1869 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3140) );
  OR2X2 OR2X2_187 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_6_), .B(alu_op_r_4_), .Y(_abc_43815_n1233_1) );
  OR2X2 OR2X2_1870 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3142) );
  OR2X2 OR2X2_1871 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3143) );
  OR2X2 OR2X2_1872 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3145) );
  OR2X2 OR2X2_1873 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3146) );
  OR2X2 OR2X2_1874 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3148) );
  OR2X2 OR2X2_1875 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3149) );
  OR2X2 OR2X2_1876 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3151) );
  OR2X2 OR2X2_1877 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3152) );
  OR2X2 OR2X2_1878 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3059_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3154) );
  OR2X2 OR2X2_1879 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3061_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3155) );
  OR2X2 OR2X2_188 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_5_), .B(int32_r_5_), .Y(_abc_43815_n1234) );
  OR2X2 OR2X2_1880 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3159) );
  OR2X2 OR2X2_1881 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3163) );
  OR2X2 OR2X2_1882 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3167) );
  OR2X2 OR2X2_1883 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3171) );
  OR2X2 OR2X2_1884 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3175) );
  OR2X2 OR2X2_1885 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3179) );
  OR2X2 OR2X2_1886 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3183) );
  OR2X2 OR2X2_1887 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3187) );
  OR2X2 OR2X2_1888 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3191) );
  OR2X2 OR2X2_1889 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3195) );
  OR2X2 OR2X2_189 ( .A(_abc_43815_n1242), .B(_abc_43815_n1243), .Y(_abc_43815_n1244) );
  OR2X2 OR2X2_1890 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3199) );
  OR2X2 OR2X2_1891 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3203) );
  OR2X2 OR2X2_1892 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3207) );
  OR2X2 OR2X2_1893 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3211) );
  OR2X2 OR2X2_1894 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3215) );
  OR2X2 OR2X2_1895 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3219) );
  OR2X2 OR2X2_1896 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3223) );
  OR2X2 OR2X2_1897 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3227) );
  OR2X2 OR2X2_1898 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3231) );
  OR2X2 OR2X2_1899 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3235) );
  OR2X2 OR2X2_19 ( .A(_abc_43815_n717), .B(_abc_43815_n715), .Y(_abc_43815_n718) );
  OR2X2 OR2X2_190 ( .A(_abc_43815_n1248), .B(_abc_43815_n1247), .Y(_abc_43815_n1249_1) );
  OR2X2 OR2X2_1900 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3239) );
  OR2X2 OR2X2_1901 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3243) );
  OR2X2 OR2X2_1902 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3247) );
  OR2X2 OR2X2_1903 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3251) );
  OR2X2 OR2X2_1904 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3255) );
  OR2X2 OR2X2_1905 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3259) );
  OR2X2 OR2X2_1906 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3263) );
  OR2X2 OR2X2_1907 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3267) );
  OR2X2 OR2X2_1908 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3271) );
  OR2X2 OR2X2_1909 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3275) );
  OR2X2 OR2X2_191 ( .A(_abc_43815_n1224), .B(_abc_43815_n1234), .Y(_abc_43815_n1254) );
  OR2X2 OR2X2_1910 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3279) );
  OR2X2 OR2X2_1911 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3158_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3283) );
  OR2X2 OR2X2_1912 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3289) );
  OR2X2 OR2X2_1913 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3293_1) );
  OR2X2 OR2X2_1914 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3297) );
  OR2X2 OR2X2_1915 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3301) );
  OR2X2 OR2X2_1916 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3305) );
  OR2X2 OR2X2_1917 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3309) );
  OR2X2 OR2X2_1918 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3313) );
  OR2X2 OR2X2_1919 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3317) );
  OR2X2 OR2X2_192 ( .A(_abc_43815_n1253), .B(_abc_43815_n1254), .Y(_abc_43815_n1255_1) );
  OR2X2 OR2X2_1920 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3321) );
  OR2X2 OR2X2_1921 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3325_1) );
  OR2X2 OR2X2_1922 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3329) );
  OR2X2 OR2X2_1923 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3333) );
  OR2X2 OR2X2_1924 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3337) );
  OR2X2 OR2X2_1925 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3341) );
  OR2X2 OR2X2_1926 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3345) );
  OR2X2 OR2X2_1927 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3349) );
  OR2X2 OR2X2_1928 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3353) );
  OR2X2 OR2X2_1929 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3357_1) );
  OR2X2 OR2X2_193 ( .A(_abc_43815_n1250_1), .B(_abc_43815_n1255_1), .Y(_abc_43815_n1256) );
  OR2X2 OR2X2_1930 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3361) );
  OR2X2 OR2X2_1931 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3365) );
  OR2X2 OR2X2_1932 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3369) );
  OR2X2 OR2X2_1933 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3373) );
  OR2X2 OR2X2_1934 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3377) );
  OR2X2 OR2X2_1935 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3381) );
  OR2X2 OR2X2_1936 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3385) );
  OR2X2 OR2X2_1937 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3389_1) );
  OR2X2 OR2X2_1938 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3393) );
  OR2X2 OR2X2_1939 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3397) );
  OR2X2 OR2X2_194 ( .A(_abc_43815_n1256), .B(_abc_43815_n1249_1), .Y(_abc_43815_n1257) );
  OR2X2 OR2X2_1940 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3401) );
  OR2X2 OR2X2_1941 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3405) );
  OR2X2 OR2X2_1942 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3409) );
  OR2X2 OR2X2_1943 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3288_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3413) );
  OR2X2 OR2X2_1944 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3418) );
  OR2X2 OR2X2_1945 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3420) );
  OR2X2 OR2X2_1946 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3422) );
  OR2X2 OR2X2_1947 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3423) );
  OR2X2 OR2X2_1948 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3425) );
  OR2X2 OR2X2_1949 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3426) );
  OR2X2 OR2X2_195 ( .A(_abc_43815_n1258), .B(_abc_43815_n1265), .Y(_abc_43815_n1266_1) );
  OR2X2 OR2X2_1950 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3428) );
  OR2X2 OR2X2_1951 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3429) );
  OR2X2 OR2X2_1952 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3431) );
  OR2X2 OR2X2_1953 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3432) );
  OR2X2 OR2X2_1954 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3434) );
  OR2X2 OR2X2_1955 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3435) );
  OR2X2 OR2X2_1956 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3437) );
  OR2X2 OR2X2_1957 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3438) );
  OR2X2 OR2X2_1958 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3440) );
  OR2X2 OR2X2_1959 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3441) );
  OR2X2 OR2X2_196 ( .A(_abc_43815_n1268), .B(_abc_43815_n1269), .Y(_abc_43815_n1270) );
  OR2X2 OR2X2_1960 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3443) );
  OR2X2 OR2X2_1961 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3444) );
  OR2X2 OR2X2_1962 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3446) );
  OR2X2 OR2X2_1963 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3447) );
  OR2X2 OR2X2_1964 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3449) );
  OR2X2 OR2X2_1965 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3450) );
  OR2X2 OR2X2_1966 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3452) );
  OR2X2 OR2X2_1967 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3453_1) );
  OR2X2 OR2X2_1968 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3455) );
  OR2X2 OR2X2_1969 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3456) );
  OR2X2 OR2X2_197 ( .A(_abc_43815_n1267), .B(_abc_43815_n1271), .Y(_abc_43815_n1272) );
  OR2X2 OR2X2_1970 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3458) );
  OR2X2 OR2X2_1971 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3459) );
  OR2X2 OR2X2_1972 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3461) );
  OR2X2 OR2X2_1973 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3462) );
  OR2X2 OR2X2_1974 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3464) );
  OR2X2 OR2X2_1975 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3465) );
  OR2X2 OR2X2_1976 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3467) );
  OR2X2 OR2X2_1977 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3468) );
  OR2X2 OR2X2_1978 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3470) );
  OR2X2 OR2X2_1979 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3471) );
  OR2X2 OR2X2_198 ( .A(_abc_43815_n1273), .B(intr_i), .Y(_abc_43815_n1274) );
  OR2X2 OR2X2_1980 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3473) );
  OR2X2 OR2X2_1981 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3474) );
  OR2X2 OR2X2_1982 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3476) );
  OR2X2 OR2X2_1983 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3477) );
  OR2X2 OR2X2_1984 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3479) );
  OR2X2 OR2X2_1985 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3480) );
  OR2X2 OR2X2_1986 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3482) );
  OR2X2 OR2X2_1987 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3483) );
  OR2X2 OR2X2_1988 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3485_1) );
  OR2X2 OR2X2_1989 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3486) );
  OR2X2 OR2X2_199 ( .A(_abc_43815_n1275), .B(_abc_43815_n1245), .Y(_abc_43815_n1276) );
  OR2X2 OR2X2_1990 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3488) );
  OR2X2 OR2X2_1991 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3489) );
  OR2X2 OR2X2_1992 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3491) );
  OR2X2 OR2X2_1993 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3492) );
  OR2X2 OR2X2_1994 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3494) );
  OR2X2 OR2X2_1995 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3495) );
  OR2X2 OR2X2_1996 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3497) );
  OR2X2 OR2X2_1997 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3498) );
  OR2X2 OR2X2_1998 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3500) );
  OR2X2 OR2X2_1999 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3501) );
  OR2X2 OR2X2_2 ( .A(_abc_43815_n619), .B(_abc_43815_n617), .Y(_abc_27555_n185) );
  OR2X2 OR2X2_20 ( .A(_abc_43815_n720), .B(_abc_43815_n719), .Y(_abc_43815_n721) );
  OR2X2 OR2X2_200 ( .A(_abc_43815_n1281), .B(_abc_43815_n1279), .Y(_abc_43815_n1282_1) );
  OR2X2 OR2X2_2000 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3503) );
  OR2X2 OR2X2_2001 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3504) );
  OR2X2 OR2X2_2002 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3506) );
  OR2X2 OR2X2_2003 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3507) );
  OR2X2 OR2X2_2004 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3509) );
  OR2X2 OR2X2_2005 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3510) );
  OR2X2 OR2X2_2006 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3417_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3512) );
  OR2X2 OR2X2_2007 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3419_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3513) );
  OR2X2 OR2X2_2008 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3518) );
  OR2X2 OR2X2_2009 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3520) );
  OR2X2 OR2X2_201 ( .A(_abc_43815_n1282_1), .B(_abc_43815_n1277), .Y(_abc_43815_n1283_1) );
  OR2X2 OR2X2_2010 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3522) );
  OR2X2 OR2X2_2011 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3523) );
  OR2X2 OR2X2_2012 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3525) );
  OR2X2 OR2X2_2013 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3526) );
  OR2X2 OR2X2_2014 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3528) );
  OR2X2 OR2X2_2015 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3529) );
  OR2X2 OR2X2_2016 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3531) );
  OR2X2 OR2X2_2017 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3532) );
  OR2X2 OR2X2_2018 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3534) );
  OR2X2 OR2X2_2019 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3535) );
  OR2X2 OR2X2_202 ( .A(sr_q_9_), .B(alu_flag_update_o), .Y(_abc_43815_n1285) );
  OR2X2 OR2X2_2020 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3537) );
  OR2X2 OR2X2_2021 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3538) );
  OR2X2 OR2X2_2022 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3540) );
  OR2X2 OR2X2_2023 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3541) );
  OR2X2 OR2X2_2024 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3543) );
  OR2X2 OR2X2_2025 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3544) );
  OR2X2 OR2X2_2026 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3546) );
  OR2X2 OR2X2_2027 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3547) );
  OR2X2 OR2X2_2028 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3549_1) );
  OR2X2 OR2X2_2029 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3550) );
  OR2X2 OR2X2_203 ( .A(_abc_43815_n1298), .B(alu_equal_o), .Y(_abc_43815_n1299) );
  OR2X2 OR2X2_2030 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3552) );
  OR2X2 OR2X2_2031 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3553) );
  OR2X2 OR2X2_2032 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3555) );
  OR2X2 OR2X2_2033 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3556) );
  OR2X2 OR2X2_2034 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3558) );
  OR2X2 OR2X2_2035 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3559) );
  OR2X2 OR2X2_2036 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3561) );
  OR2X2 OR2X2_2037 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3562) );
  OR2X2 OR2X2_2038 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3564) );
  OR2X2 OR2X2_2039 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3565) );
  OR2X2 OR2X2_204 ( .A(_abc_43815_n1101), .B(_abc_43815_n1300_1), .Y(_abc_43815_n1301) );
  OR2X2 OR2X2_2040 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3567) );
  OR2X2 OR2X2_2041 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3568) );
  OR2X2 OR2X2_2042 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3570) );
  OR2X2 OR2X2_2043 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3571) );
  OR2X2 OR2X2_2044 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3573) );
  OR2X2 OR2X2_2045 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3574) );
  OR2X2 OR2X2_2046 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3576) );
  OR2X2 OR2X2_2047 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3577) );
  OR2X2 OR2X2_2048 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3579) );
  OR2X2 OR2X2_2049 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3580) );
  OR2X2 OR2X2_205 ( .A(_abc_43815_n1306), .B(_abc_43815_n1305), .Y(_abc_43815_n1307) );
  OR2X2 OR2X2_2050 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3582) );
  OR2X2 OR2X2_2051 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3583) );
  OR2X2 OR2X2_2052 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3585) );
  OR2X2 OR2X2_2053 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3586) );
  OR2X2 OR2X2_2054 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3588) );
  OR2X2 OR2X2_2055 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3589) );
  OR2X2 OR2X2_2056 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3591) );
  OR2X2 OR2X2_2057 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3592) );
  OR2X2 OR2X2_2058 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3594) );
  OR2X2 OR2X2_2059 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3595) );
  OR2X2 OR2X2_206 ( .A(_abc_43815_n1303_1), .B(_abc_43815_n1307), .Y(_abc_43815_n1308) );
  OR2X2 OR2X2_2060 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3597) );
  OR2X2 OR2X2_2061 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3598) );
  OR2X2 OR2X2_2062 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3600) );
  OR2X2 OR2X2_2063 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3601) );
  OR2X2 OR2X2_2064 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3603) );
  OR2X2 OR2X2_2065 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3604) );
  OR2X2 OR2X2_2066 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3606) );
  OR2X2 OR2X2_2067 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3607) );
  OR2X2 OR2X2_2068 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3609) );
  OR2X2 OR2X2_2069 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3610) );
  OR2X2 OR2X2_207 ( .A(_abc_43815_n1089), .B(alu_less_than_signed_o), .Y(_abc_43815_n1309) );
  OR2X2 OR2X2_2070 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3517_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3612) );
  OR2X2 OR2X2_2071 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3519_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n3613_1) );
  OR2X2 OR2X2_2072 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3617) );
  OR2X2 OR2X2_2073 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3619) );
  OR2X2 OR2X2_2074 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3621) );
  OR2X2 OR2X2_2075 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3622) );
  OR2X2 OR2X2_2076 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3624) );
  OR2X2 OR2X2_2077 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3625) );
  OR2X2 OR2X2_2078 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3627) );
  OR2X2 OR2X2_2079 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3628) );
  OR2X2 OR2X2_208 ( .A(_abc_43815_n1310), .B(_abc_43815_n1020), .Y(_abc_43815_n1311) );
  OR2X2 OR2X2_2080 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3630) );
  OR2X2 OR2X2_2081 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3631) );
  OR2X2 OR2X2_2082 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3633) );
  OR2X2 OR2X2_2083 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3634) );
  OR2X2 OR2X2_2084 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3636) );
  OR2X2 OR2X2_2085 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3637) );
  OR2X2 OR2X2_2086 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3639) );
  OR2X2 OR2X2_2087 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3640) );
  OR2X2 OR2X2_2088 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3642) );
  OR2X2 OR2X2_2089 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3643) );
  OR2X2 OR2X2_209 ( .A(alu_less_than_o), .B(alu_equal_o), .Y(_abc_43815_n1312) );
  OR2X2 OR2X2_2090 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3645_1) );
  OR2X2 OR2X2_2091 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3646) );
  OR2X2 OR2X2_2092 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3648) );
  OR2X2 OR2X2_2093 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3649) );
  OR2X2 OR2X2_2094 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3651) );
  OR2X2 OR2X2_2095 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3652) );
  OR2X2 OR2X2_2096 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3654) );
  OR2X2 OR2X2_2097 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3655) );
  OR2X2 OR2X2_2098 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3657) );
  OR2X2 OR2X2_2099 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3658) );
  OR2X2 OR2X2_21 ( .A(_abc_43815_n722), .B(_abc_43815_n723), .Y(_abc_43815_n724) );
  OR2X2 OR2X2_210 ( .A(_abc_43815_n1021), .B(_abc_43815_n1312), .Y(_abc_43815_n1313) );
  OR2X2 OR2X2_2100 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3660) );
  OR2X2 OR2X2_2101 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3661) );
  OR2X2 OR2X2_2102 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3663) );
  OR2X2 OR2X2_2103 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3664) );
  OR2X2 OR2X2_2104 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3666) );
  OR2X2 OR2X2_2105 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3667) );
  OR2X2 OR2X2_2106 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3669) );
  OR2X2 OR2X2_2107 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3670) );
  OR2X2 OR2X2_2108 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3672) );
  OR2X2 OR2X2_2109 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3673) );
  OR2X2 OR2X2_211 ( .A(_abc_43815_n1314), .B(_abc_43815_n1014), .Y(_abc_43815_n1315) );
  OR2X2 OR2X2_2110 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3675) );
  OR2X2 OR2X2_2111 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3676) );
  OR2X2 OR2X2_2112 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3678) );
  OR2X2 OR2X2_2113 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3679) );
  OR2X2 OR2X2_2114 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3681) );
  OR2X2 OR2X2_2115 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3682) );
  OR2X2 OR2X2_2116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3684) );
  OR2X2 OR2X2_2117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3685) );
  OR2X2 OR2X2_2118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3687) );
  OR2X2 OR2X2_2119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3688) );
  OR2X2 OR2X2_212 ( .A(alu_less_than_signed_o), .B(alu_equal_o), .Y(_abc_43815_n1316) );
  OR2X2 OR2X2_2120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3690) );
  OR2X2 OR2X2_2121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3691) );
  OR2X2 OR2X2_2122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3693) );
  OR2X2 OR2X2_2123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3694) );
  OR2X2 OR2X2_2124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3696) );
  OR2X2 OR2X2_2125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3697) );
  OR2X2 OR2X2_2126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3699) );
  OR2X2 OR2X2_2127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3700) );
  OR2X2 OR2X2_2128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3702) );
  OR2X2 OR2X2_2129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3703) );
  OR2X2 OR2X2_213 ( .A(_abc_43815_n1015), .B(_abc_43815_n1316), .Y(_abc_43815_n1317) );
  OR2X2 OR2X2_2130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3705) );
  OR2X2 OR2X2_2131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3706) );
  OR2X2 OR2X2_2132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3708) );
  OR2X2 OR2X2_2133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3709_1) );
  OR2X2 OR2X2_2134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3616_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3711) );
  OR2X2 OR2X2_2135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3618_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n3712) );
  OR2X2 OR2X2_2136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3716) );
  OR2X2 OR2X2_2137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3718) );
  OR2X2 OR2X2_2138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3720) );
  OR2X2 OR2X2_2139 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3721) );
  OR2X2 OR2X2_214 ( .A(_abc_43815_n1318), .B(_abc_43815_n997), .Y(_abc_43815_n1319_1) );
  OR2X2 OR2X2_2140 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3723) );
  OR2X2 OR2X2_2141 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3724) );
  OR2X2 OR2X2_2142 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3726) );
  OR2X2 OR2X2_2143 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3727) );
  OR2X2 OR2X2_2144 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3729) );
  OR2X2 OR2X2_2145 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3730) );
  OR2X2 OR2X2_2146 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3732) );
  OR2X2 OR2X2_2147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3733) );
  OR2X2 OR2X2_2148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3735) );
  OR2X2 OR2X2_2149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3736) );
  OR2X2 OR2X2_215 ( .A(_abc_43815_n998), .B(alu_greater_than_o), .Y(_abc_43815_n1320_1) );
  OR2X2 OR2X2_2150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3738) );
  OR2X2 OR2X2_2151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3739) );
  OR2X2 OR2X2_2152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3741_1) );
  OR2X2 OR2X2_2153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3742) );
  OR2X2 OR2X2_2154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3744) );
  OR2X2 OR2X2_2155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3745) );
  OR2X2 OR2X2_2156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3747) );
  OR2X2 OR2X2_2157 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3748) );
  OR2X2 OR2X2_2158 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3750) );
  OR2X2 OR2X2_2159 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3751) );
  OR2X2 OR2X2_216 ( .A(_abc_43815_n1324), .B(_abc_43815_n1323), .Y(_abc_43815_n1325_1) );
  OR2X2 OR2X2_2160 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3753) );
  OR2X2 OR2X2_2161 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3754) );
  OR2X2 OR2X2_2162 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3756) );
  OR2X2 OR2X2_2163 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3757) );
  OR2X2 OR2X2_2164 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3759) );
  OR2X2 OR2X2_2165 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3760) );
  OR2X2 OR2X2_2166 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3762) );
  OR2X2 OR2X2_2167 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3763) );
  OR2X2 OR2X2_2168 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3765) );
  OR2X2 OR2X2_2169 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3766) );
  OR2X2 OR2X2_217 ( .A(_abc_43815_n1322), .B(_abc_43815_n1325_1), .Y(_abc_43815_n1326) );
  OR2X2 OR2X2_2170 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3768) );
  OR2X2 OR2X2_2171 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3769) );
  OR2X2 OR2X2_2172 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3771) );
  OR2X2 OR2X2_2173 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3772) );
  OR2X2 OR2X2_2174 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3774) );
  OR2X2 OR2X2_2175 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3775) );
  OR2X2 OR2X2_2176 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3777) );
  OR2X2 OR2X2_2177 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3778) );
  OR2X2 OR2X2_2178 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3780) );
  OR2X2 OR2X2_2179 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3781) );
  OR2X2 OR2X2_218 ( .A(alu_greater_than_o), .B(alu_equal_o), .Y(_abc_43815_n1327) );
  OR2X2 OR2X2_2180 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3783) );
  OR2X2 OR2X2_2181 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3784) );
  OR2X2 OR2X2_2182 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3786) );
  OR2X2 OR2X2_2183 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3787) );
  OR2X2 OR2X2_2184 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3789) );
  OR2X2 OR2X2_2185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3790) );
  OR2X2 OR2X2_2186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3792) );
  OR2X2 OR2X2_2187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3793) );
  OR2X2 OR2X2_2188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3795) );
  OR2X2 OR2X2_2189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3796) );
  OR2X2 OR2X2_219 ( .A(_abc_43815_n1031_1), .B(_abc_43815_n1327), .Y(_abc_43815_n1328) );
  OR2X2 OR2X2_2190 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3798) );
  OR2X2 OR2X2_2191 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3799) );
  OR2X2 OR2X2_2192 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3801) );
  OR2X2 OR2X2_2193 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3802) );
  OR2X2 OR2X2_2194 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3804) );
  OR2X2 OR2X2_2195 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3805_1) );
  OR2X2 OR2X2_2196 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3807) );
  OR2X2 OR2X2_2197 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3808) );
  OR2X2 OR2X2_2198 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3715_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3810) );
  OR2X2 OR2X2_2199 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3717_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n3811) );
  OR2X2 OR2X2_22 ( .A(_abc_43815_n724), .B(_abc_43815_n721), .Y(_abc_43815_n725) );
  OR2X2 OR2X2_220 ( .A(_abc_43815_n1329), .B(_abc_43815_n1289_1), .Y(_abc_43815_n1330) );
  OR2X2 OR2X2_2200 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3814) );
  OR2X2 OR2X2_2201 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3816) );
  OR2X2 OR2X2_2202 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3818) );
  OR2X2 OR2X2_2203 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3819) );
  OR2X2 OR2X2_2204 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3821) );
  OR2X2 OR2X2_2205 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3822) );
  OR2X2 OR2X2_2206 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3824) );
  OR2X2 OR2X2_2207 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3825) );
  OR2X2 OR2X2_2208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3827) );
  OR2X2 OR2X2_2209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3828) );
  OR2X2 OR2X2_221 ( .A(alu_greater_than_signed_o), .B(alu_equal_o), .Y(_abc_43815_n1331) );
  OR2X2 OR2X2_2210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3830) );
  OR2X2 OR2X2_2211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3831) );
  OR2X2 OR2X2_2212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3833) );
  OR2X2 OR2X2_2213 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3834) );
  OR2X2 OR2X2_2214 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3836) );
  OR2X2 OR2X2_2215 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3837_1) );
  OR2X2 OR2X2_2216 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3839) );
  OR2X2 OR2X2_2217 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3840) );
  OR2X2 OR2X2_2218 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3842) );
  OR2X2 OR2X2_2219 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3843) );
  OR2X2 OR2X2_222 ( .A(_abc_43815_n1028), .B(_abc_43815_n1331), .Y(_abc_43815_n1332) );
  OR2X2 OR2X2_2220 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3845) );
  OR2X2 OR2X2_2221 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3846) );
  OR2X2 OR2X2_2222 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3848) );
  OR2X2 OR2X2_2223 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3849) );
  OR2X2 OR2X2_2224 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3851) );
  OR2X2 OR2X2_2225 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3852) );
  OR2X2 OR2X2_2226 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3854) );
  OR2X2 OR2X2_2227 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3855) );
  OR2X2 OR2X2_2228 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3857) );
  OR2X2 OR2X2_2229 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3858) );
  OR2X2 OR2X2_223 ( .A(_abc_43815_n1333_1), .B(_abc_43815_n1286), .Y(_abc_43815_n1334) );
  OR2X2 OR2X2_2230 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3860) );
  OR2X2 OR2X2_2231 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3861) );
  OR2X2 OR2X2_2232 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3863) );
  OR2X2 OR2X2_2233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3864) );
  OR2X2 OR2X2_2234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3866) );
  OR2X2 OR2X2_2235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3867) );
  OR2X2 OR2X2_2236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3869_1) );
  OR2X2 OR2X2_2237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3870) );
  OR2X2 OR2X2_2238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3872) );
  OR2X2 OR2X2_2239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3873) );
  OR2X2 OR2X2_224 ( .A(_abc_43815_n1337), .B(_abc_43815_n1081), .Y(_abc_43815_n1338) );
  OR2X2 OR2X2_2240 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3875) );
  OR2X2 OR2X2_2241 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3876) );
  OR2X2 OR2X2_2242 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3878) );
  OR2X2 OR2X2_2243 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3879) );
  OR2X2 OR2X2_2244 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3881) );
  OR2X2 OR2X2_2245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3882) );
  OR2X2 OR2X2_2246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3884) );
  OR2X2 OR2X2_2247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3885) );
  OR2X2 OR2X2_2248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3887) );
  OR2X2 OR2X2_2249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3888) );
  OR2X2 OR2X2_225 ( .A(_abc_43815_n1336_1), .B(_abc_43815_n1338), .Y(_abc_43815_n1339) );
  OR2X2 OR2X2_2250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3890) );
  OR2X2 OR2X2_2251 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3891) );
  OR2X2 OR2X2_2252 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3893) );
  OR2X2 OR2X2_2253 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3894) );
  OR2X2 OR2X2_2254 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3896) );
  OR2X2 OR2X2_2255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3897) );
  OR2X2 OR2X2_2256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3899) );
  OR2X2 OR2X2_2257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3900) );
  OR2X2 OR2X2_2258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3902) );
  OR2X2 OR2X2_2259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3903) );
  OR2X2 OR2X2_226 ( .A(_abc_43815_n1335), .B(_abc_43815_n987), .Y(_abc_43815_n1340) );
  OR2X2 OR2X2_2260 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3905) );
  OR2X2 OR2X2_2261 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3906) );
  OR2X2 OR2X2_2262 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3813_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3908) );
  OR2X2 OR2X2_2263 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3815_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n3909) );
  OR2X2 OR2X2_2264 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3914) );
  OR2X2 OR2X2_2265 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3918) );
  OR2X2 OR2X2_2266 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3922) );
  OR2X2 OR2X2_2267 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3926) );
  OR2X2 OR2X2_2268 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3930) );
  OR2X2 OR2X2_2269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3934) );
  OR2X2 OR2X2_227 ( .A(_abc_43815_n1333_1), .B(_abc_43815_n999), .Y(_abc_43815_n1341) );
  OR2X2 OR2X2_2270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3938) );
  OR2X2 OR2X2_2271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3942) );
  OR2X2 OR2X2_2272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3946) );
  OR2X2 OR2X2_2273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3950) );
  OR2X2 OR2X2_2274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3954) );
  OR2X2 OR2X2_2275 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3958) );
  OR2X2 OR2X2_2276 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3962) );
  OR2X2 OR2X2_2277 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3966) );
  OR2X2 OR2X2_2278 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3970) );
  OR2X2 OR2X2_2279 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3974) );
  OR2X2 OR2X2_228 ( .A(_abc_43815_n1344), .B(_abc_43815_n1080), .Y(_abc_43815_n1345) );
  OR2X2 OR2X2_2280 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3978) );
  OR2X2 OR2X2_2281 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3982) );
  OR2X2 OR2X2_2282 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3986) );
  OR2X2 OR2X2_2283 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3990) );
  OR2X2 OR2X2_2284 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3994) );
  OR2X2 OR2X2_2285 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n3998) );
  OR2X2 OR2X2_2286 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4002) );
  OR2X2 OR2X2_2287 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4006) );
  OR2X2 OR2X2_2288 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4010) );
  OR2X2 OR2X2_2289 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4014) );
  OR2X2 OR2X2_229 ( .A(_abc_43815_n1343), .B(_abc_43815_n1345), .Y(_abc_43815_n1346) );
  OR2X2 OR2X2_2290 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4018) );
  OR2X2 OR2X2_2291 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4022) );
  OR2X2 OR2X2_2292 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4026) );
  OR2X2 OR2X2_2293 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4030) );
  OR2X2 OR2X2_2294 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4034) );
  OR2X2 OR2X2_2295 ( .A(REGFILE_SIM_reg_bank__abc_33898_n3913_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4038) );
  OR2X2 OR2X2_2296 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4043) );
  OR2X2 OR2X2_2297 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4045) );
  OR2X2 OR2X2_2298 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4047) );
  OR2X2 OR2X2_2299 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4048) );
  OR2X2 OR2X2_23 ( .A(_abc_43815_n686_1_bF_buf3), .B(_abc_43815_n725), .Y(_abc_43815_n726) );
  OR2X2 OR2X2_230 ( .A(_abc_43815_n1240), .B(esr_q_9_), .Y(_abc_43815_n1355) );
  OR2X2 OR2X2_2300 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4050) );
  OR2X2 OR2X2_2301 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4051) );
  OR2X2 OR2X2_2302 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4053) );
  OR2X2 OR2X2_2303 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4054) );
  OR2X2 OR2X2_2304 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4056) );
  OR2X2 OR2X2_2305 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4057) );
  OR2X2 OR2X2_2306 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4059) );
  OR2X2 OR2X2_2307 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4060) );
  OR2X2 OR2X2_2308 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4062) );
  OR2X2 OR2X2_2309 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4063) );
  OR2X2 OR2X2_231 ( .A(_abc_43815_n1360_1), .B(_abc_43815_n1278_bF_buf6), .Y(_abc_43815_n1361) );
  OR2X2 OR2X2_2310 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4065) );
  OR2X2 OR2X2_2311 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4066) );
  OR2X2 OR2X2_2312 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4068) );
  OR2X2 OR2X2_2313 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4069) );
  OR2X2 OR2X2_2314 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4071) );
  OR2X2 OR2X2_2315 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4072) );
  OR2X2 OR2X2_2316 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4074) );
  OR2X2 OR2X2_2317 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4075) );
  OR2X2 OR2X2_2318 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4077) );
  OR2X2 OR2X2_2319 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4078) );
  OR2X2 OR2X2_232 ( .A(_abc_43815_n1354), .B(_abc_43815_n1361), .Y(_abc_43815_n1362) );
  OR2X2 OR2X2_2320 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4080) );
  OR2X2 OR2X2_2321 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4081) );
  OR2X2 OR2X2_2322 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4083) );
  OR2X2 OR2X2_2323 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4084) );
  OR2X2 OR2X2_2324 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4086) );
  OR2X2 OR2X2_2325 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4087) );
  OR2X2 OR2X2_2326 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4089) );
  OR2X2 OR2X2_2327 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4090) );
  OR2X2 OR2X2_2328 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4092) );
  OR2X2 OR2X2_2329 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4093_1) );
  OR2X2 OR2X2_233 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(esr_q_9_), .Y(_abc_43815_n1363) );
  OR2X2 OR2X2_2330 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4095) );
  OR2X2 OR2X2_2331 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4096) );
  OR2X2 OR2X2_2332 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4098) );
  OR2X2 OR2X2_2333 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4099) );
  OR2X2 OR2X2_2334 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4101) );
  OR2X2 OR2X2_2335 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4102) );
  OR2X2 OR2X2_2336 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4104) );
  OR2X2 OR2X2_2337 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4105) );
  OR2X2 OR2X2_2338 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4107) );
  OR2X2 OR2X2_2339 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4108) );
  OR2X2 OR2X2_234 ( .A(alu_c_i), .B(alu_c_update_o), .Y(_abc_43815_n1366) );
  OR2X2 OR2X2_2340 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4110) );
  OR2X2 OR2X2_2341 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4111) );
  OR2X2 OR2X2_2342 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4113) );
  OR2X2 OR2X2_2343 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4114) );
  OR2X2 OR2X2_2344 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4116) );
  OR2X2 OR2X2_2345 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4117) );
  OR2X2 OR2X2_2346 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4119) );
  OR2X2 OR2X2_2347 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4120) );
  OR2X2 OR2X2_2348 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4122) );
  OR2X2 OR2X2_2349 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4123) );
  OR2X2 OR2X2_235 ( .A(_abc_43815_n1367), .B(alu_c_o), .Y(_abc_43815_n1368) );
  OR2X2 OR2X2_2350 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4125_1) );
  OR2X2 OR2X2_2351 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4126) );
  OR2X2 OR2X2_2352 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4128) );
  OR2X2 OR2X2_2353 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4129) );
  OR2X2 OR2X2_2354 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4131) );
  OR2X2 OR2X2_2355 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4132) );
  OR2X2 OR2X2_2356 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4134) );
  OR2X2 OR2X2_2357 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4135) );
  OR2X2 OR2X2_2358 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4042_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4137) );
  OR2X2 OR2X2_2359 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4044_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4138) );
  OR2X2 OR2X2_236 ( .A(_abc_43815_n1371), .B(_abc_43815_n1080), .Y(_abc_43815_n1372_1) );
  OR2X2 OR2X2_2360 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4141) );
  OR2X2 OR2X2_2361 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4143) );
  OR2X2 OR2X2_2362 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4145) );
  OR2X2 OR2X2_2363 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4146) );
  OR2X2 OR2X2_2364 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4148) );
  OR2X2 OR2X2_2365 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4149) );
  OR2X2 OR2X2_2366 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4151) );
  OR2X2 OR2X2_2367 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4152) );
  OR2X2 OR2X2_2368 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4154) );
  OR2X2 OR2X2_2369 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4155) );
  OR2X2 OR2X2_237 ( .A(_abc_43815_n1372_1), .B(_abc_43815_n1370), .Y(_abc_43815_n1373) );
  OR2X2 OR2X2_2370 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4157_1) );
  OR2X2 OR2X2_2371 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4158) );
  OR2X2 OR2X2_2372 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4160) );
  OR2X2 OR2X2_2373 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4161) );
  OR2X2 OR2X2_2374 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4163) );
  OR2X2 OR2X2_2375 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4164) );
  OR2X2 OR2X2_2376 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4166) );
  OR2X2 OR2X2_2377 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4167) );
  OR2X2 OR2X2_2378 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4169) );
  OR2X2 OR2X2_2379 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4170) );
  OR2X2 OR2X2_238 ( .A(_abc_43815_n1379), .B(_abc_43815_n1369), .Y(_abc_43815_n1380) );
  OR2X2 OR2X2_2380 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4172) );
  OR2X2 OR2X2_2381 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4173) );
  OR2X2 OR2X2_2382 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4175) );
  OR2X2 OR2X2_2383 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4176) );
  OR2X2 OR2X2_2384 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4178) );
  OR2X2 OR2X2_2385 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4179) );
  OR2X2 OR2X2_2386 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4181) );
  OR2X2 OR2X2_2387 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4182) );
  OR2X2 OR2X2_2388 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4184) );
  OR2X2 OR2X2_2389 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4185) );
  OR2X2 OR2X2_239 ( .A(_abc_43815_n1384), .B(_abc_43815_n1081), .Y(_abc_43815_n1385) );
  OR2X2 OR2X2_2390 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4187) );
  OR2X2 OR2X2_2391 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4188) );
  OR2X2 OR2X2_2392 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4190_1) );
  OR2X2 OR2X2_2393 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4191) );
  OR2X2 OR2X2_2394 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4193_1) );
  OR2X2 OR2X2_2395 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4194) );
  OR2X2 OR2X2_2396 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4196) );
  OR2X2 OR2X2_2397 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4197_1) );
  OR2X2 OR2X2_2398 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4199) );
  OR2X2 OR2X2_2399 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4200) );
  OR2X2 OR2X2_24 ( .A(_abc_43815_n728), .B(_abc_43815_n714), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_) );
  OR2X2 OR2X2_240 ( .A(_abc_43815_n1240), .B(esr_q_10_), .Y(_abc_43815_n1388) );
  OR2X2 OR2X2_2400 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4202) );
  OR2X2 OR2X2_2401 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4203) );
  OR2X2 OR2X2_2402 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4205) );
  OR2X2 OR2X2_2403 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4206) );
  OR2X2 OR2X2_2404 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4208) );
  OR2X2 OR2X2_2405 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4209) );
  OR2X2 OR2X2_2406 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4211) );
  OR2X2 OR2X2_2407 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4212) );
  OR2X2 OR2X2_2408 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4214) );
  OR2X2 OR2X2_2409 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4215) );
  OR2X2 OR2X2_241 ( .A(_abc_43815_n1392_1), .B(_abc_43815_n1278_bF_buf5), .Y(_abc_43815_n1393) );
  OR2X2 OR2X2_2410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4217) );
  OR2X2 OR2X2_2411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4218) );
  OR2X2 OR2X2_2412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4220) );
  OR2X2 OR2X2_2413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4221) );
  OR2X2 OR2X2_2414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4223) );
  OR2X2 OR2X2_2415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4224) );
  OR2X2 OR2X2_2416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4226) );
  OR2X2 OR2X2_2417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4227) );
  OR2X2 OR2X2_2418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4229) );
  OR2X2 OR2X2_2419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4230) );
  OR2X2 OR2X2_242 ( .A(_abc_43815_n1393), .B(_abc_43815_n1387), .Y(_abc_43815_n1394) );
  OR2X2 OR2X2_2420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4232) );
  OR2X2 OR2X2_2421 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4233) );
  OR2X2 OR2X2_2422 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4140_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4235) );
  OR2X2 OR2X2_2423 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4142_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4236) );
  OR2X2 OR2X2_2424 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4240) );
  OR2X2 OR2X2_2425 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4242) );
  OR2X2 OR2X2_2426 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4244) );
  OR2X2 OR2X2_2427 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4245) );
  OR2X2 OR2X2_2428 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4247) );
  OR2X2 OR2X2_2429 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4248) );
  OR2X2 OR2X2_243 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(esr_q_10_), .Y(_abc_43815_n1395) );
  OR2X2 OR2X2_2430 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4250) );
  OR2X2 OR2X2_2431 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4251) );
  OR2X2 OR2X2_2432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4253) );
  OR2X2 OR2X2_2433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4254) );
  OR2X2 OR2X2_2434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4256) );
  OR2X2 OR2X2_2435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4257) );
  OR2X2 OR2X2_2436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4259) );
  OR2X2 OR2X2_2437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4260) );
  OR2X2 OR2X2_2438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4262) );
  OR2X2 OR2X2_2439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4263) );
  OR2X2 OR2X2_244 ( .A(_abc_43815_n1400), .B(_abc_43815_n1401), .Y(_abc_43815_n1402) );
  OR2X2 OR2X2_2440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4265) );
  OR2X2 OR2X2_2441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4266) );
  OR2X2 OR2X2_2442 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4268) );
  OR2X2 OR2X2_2443 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4269) );
  OR2X2 OR2X2_2444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4271) );
  OR2X2 OR2X2_2445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4272) );
  OR2X2 OR2X2_2446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4274) );
  OR2X2 OR2X2_2447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4275) );
  OR2X2 OR2X2_2448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4277) );
  OR2X2 OR2X2_2449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4278) );
  OR2X2 OR2X2_245 ( .A(_abc_43815_n1404), .B(_abc_43815_n1405_1), .Y(_abc_43815_n1406) );
  OR2X2 OR2X2_2450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4280) );
  OR2X2 OR2X2_2451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4281) );
  OR2X2 OR2X2_2452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4283) );
  OR2X2 OR2X2_2453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4284) );
  OR2X2 OR2X2_2454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4286) );
  OR2X2 OR2X2_2455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4287) );
  OR2X2 OR2X2_2456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4289) );
  OR2X2 OR2X2_2457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4290) );
  OR2X2 OR2X2_2458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4292) );
  OR2X2 OR2X2_2459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4293) );
  OR2X2 OR2X2_246 ( .A(_abc_43815_n1409), .B(_abc_43815_n1408_1), .Y(_abc_43815_n1410) );
  OR2X2 OR2X2_2460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4295) );
  OR2X2 OR2X2_2461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4296) );
  OR2X2 OR2X2_2462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4298) );
  OR2X2 OR2X2_2463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4299) );
  OR2X2 OR2X2_2464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4301) );
  OR2X2 OR2X2_2465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4302) );
  OR2X2 OR2X2_2466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4304) );
  OR2X2 OR2X2_2467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4305) );
  OR2X2 OR2X2_2468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4307) );
  OR2X2 OR2X2_2469 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4308) );
  OR2X2 OR2X2_247 ( .A(_abc_43815_n1278_bF_buf1), .B(next_pc_r_0_), .Y(_abc_43815_n1412) );
  OR2X2 OR2X2_2470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4310) );
  OR2X2 OR2X2_2471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4311) );
  OR2X2 OR2X2_2472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4313_1) );
  OR2X2 OR2X2_2473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4314) );
  OR2X2 OR2X2_2474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4316) );
  OR2X2 OR2X2_2475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4317) );
  OR2X2 OR2X2_2476 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4319) );
  OR2X2 OR2X2_2477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4320) );
  OR2X2 OR2X2_2478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4322) );
  OR2X2 OR2X2_2479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4323) );
  OR2X2 OR2X2_248 ( .A(_abc_43815_n1418_bF_buf5), .B(epc_q_0_), .Y(_abc_43815_n1419) );
  OR2X2 OR2X2_2480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4325) );
  OR2X2 OR2X2_2481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4326) );
  OR2X2 OR2X2_2482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4328) );
  OR2X2 OR2X2_2483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4329) );
  OR2X2 OR2X2_2484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4331) );
  OR2X2 OR2X2_2485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4332) );
  OR2X2 OR2X2_2486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4239_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4334) );
  OR2X2 OR2X2_2487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4241_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n4335) );
  OR2X2 OR2X2_2488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4338) );
  OR2X2 OR2X2_2489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4340) );
  OR2X2 OR2X2_249 ( .A(_abc_43815_n1413_bF_buf4), .B(_abc_43815_n1423), .Y(_abc_43815_n1424_1) );
  OR2X2 OR2X2_2490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4342) );
  OR2X2 OR2X2_2491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4343_1) );
  OR2X2 OR2X2_2492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4345) );
  OR2X2 OR2X2_2493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4346) );
  OR2X2 OR2X2_2494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4348) );
  OR2X2 OR2X2_2495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4349) );
  OR2X2 OR2X2_2496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4351) );
  OR2X2 OR2X2_2497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4352) );
  OR2X2 OR2X2_2498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4354) );
  OR2X2 OR2X2_2499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4355) );
  OR2X2 OR2X2_25 ( .A(_abc_43815_n731), .B(_abc_43815_n732), .Y(_abc_43815_n733_1) );
  OR2X2 OR2X2_250 ( .A(_abc_43815_n1169), .B(_abc_43815_n1069), .Y(_abc_43815_n1428) );
  OR2X2 OR2X2_2500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4357) );
  OR2X2 OR2X2_2501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4358) );
  OR2X2 OR2X2_2502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4360) );
  OR2X2 OR2X2_2503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4361) );
  OR2X2 OR2X2_2504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4363) );
  OR2X2 OR2X2_2505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4364) );
  OR2X2 OR2X2_2506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4366) );
  OR2X2 OR2X2_2507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4367) );
  OR2X2 OR2X2_2508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4369) );
  OR2X2 OR2X2_2509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4370) );
  OR2X2 OR2X2_251 ( .A(_abc_43815_n1428_bF_buf4), .B(_abc_43815_n1427), .Y(_abc_43815_n1429) );
  OR2X2 OR2X2_2510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4372) );
  OR2X2 OR2X2_2511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4373_1) );
  OR2X2 OR2X2_2512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4375) );
  OR2X2 OR2X2_2513 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4376) );
  OR2X2 OR2X2_2514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4378) );
  OR2X2 OR2X2_2515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4379) );
  OR2X2 OR2X2_2516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4381) );
  OR2X2 OR2X2_2517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4382) );
  OR2X2 OR2X2_2518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4384) );
  OR2X2 OR2X2_2519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4385) );
  OR2X2 OR2X2_252 ( .A(_abc_43815_n1426), .B(_abc_43815_n1429), .Y(_abc_43815_n1430) );
  OR2X2 OR2X2_2520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4387) );
  OR2X2 OR2X2_2521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4388) );
  OR2X2 OR2X2_2522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4390) );
  OR2X2 OR2X2_2523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4391) );
  OR2X2 OR2X2_2524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4393) );
  OR2X2 OR2X2_2525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4394) );
  OR2X2 OR2X2_2526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4396) );
  OR2X2 OR2X2_2527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4397) );
  OR2X2 OR2X2_2528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4399) );
  OR2X2 OR2X2_2529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4400) );
  OR2X2 OR2X2_253 ( .A(_abc_43815_n1431_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_43815_n1432) );
  OR2X2 OR2X2_2530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4402) );
  OR2X2 OR2X2_2531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4403_1) );
  OR2X2 OR2X2_2532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4405) );
  OR2X2 OR2X2_2533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4406) );
  OR2X2 OR2X2_2534 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4408) );
  OR2X2 OR2X2_2535 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4409) );
  OR2X2 OR2X2_2536 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4411) );
  OR2X2 OR2X2_2537 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4412) );
  OR2X2 OR2X2_2538 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4414) );
  OR2X2 OR2X2_2539 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4415) );
  OR2X2 OR2X2_254 ( .A(_abc_43815_n1350_bF_buf1), .B(_abc_43815_n1433), .Y(_abc_43815_n1434) );
  OR2X2 OR2X2_2540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4417) );
  OR2X2 OR2X2_2541 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4418) );
  OR2X2 OR2X2_2542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4420) );
  OR2X2 OR2X2_2543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4421) );
  OR2X2 OR2X2_2544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4423) );
  OR2X2 OR2X2_2545 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4424) );
  OR2X2 OR2X2_2546 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4426) );
  OR2X2 OR2X2_2547 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4427) );
  OR2X2 OR2X2_2548 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4429) );
  OR2X2 OR2X2_2549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4430) );
  OR2X2 OR2X2_255 ( .A(_abc_43815_n1436), .B(_abc_43815_n1412), .Y(_abc_43815_n1437) );
  OR2X2 OR2X2_2550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4337_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4432) );
  OR2X2 OR2X2_2551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4339_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n4433_1) );
  OR2X2 OR2X2_2552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4436) );
  OR2X2 OR2X2_2553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4440) );
  OR2X2 OR2X2_2554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4444) );
  OR2X2 OR2X2_2555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4448) );
  OR2X2 OR2X2_2556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4452) );
  OR2X2 OR2X2_2557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4456) );
  OR2X2 OR2X2_2558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4460) );
  OR2X2 OR2X2_2559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4464) );
  OR2X2 OR2X2_256 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_0_), .Y(_abc_43815_n1438) );
  OR2X2 OR2X2_2560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4468) );
  OR2X2 OR2X2_2561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4472) );
  OR2X2 OR2X2_2562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4476) );
  OR2X2 OR2X2_2563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4480) );
  OR2X2 OR2X2_2564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4484) );
  OR2X2 OR2X2_2565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4488) );
  OR2X2 OR2X2_2566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4492) );
  OR2X2 OR2X2_2567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4496) );
  OR2X2 OR2X2_2568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4500) );
  OR2X2 OR2X2_2569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4504) );
  OR2X2 OR2X2_257 ( .A(_abc_43815_n1418_bF_buf3), .B(epc_q_1_), .Y(_abc_43815_n1441) );
  OR2X2 OR2X2_2570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4508) );
  OR2X2 OR2X2_2571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4512) );
  OR2X2 OR2X2_2572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4516) );
  OR2X2 OR2X2_2573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4520) );
  OR2X2 OR2X2_2574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4524) );
  OR2X2 OR2X2_2575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4528) );
  OR2X2 OR2X2_2576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4532) );
  OR2X2 OR2X2_2577 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4536) );
  OR2X2 OR2X2_2578 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4540) );
  OR2X2 OR2X2_2579 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4544) );
  OR2X2 OR2X2_258 ( .A(_abc_43815_n1413_bF_buf3), .B(_abc_43815_n1445), .Y(_abc_43815_n1446) );
  OR2X2 OR2X2_2580 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4548) );
  OR2X2 OR2X2_2581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4552) );
  OR2X2 OR2X2_2582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4556) );
  OR2X2 OR2X2_2583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4435_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4560) );
  OR2X2 OR2X2_2584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4565) );
  OR2X2 OR2X2_2585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4569) );
  OR2X2 OR2X2_2586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4573) );
  OR2X2 OR2X2_2587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4577) );
  OR2X2 OR2X2_2588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4581) );
  OR2X2 OR2X2_2589 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4585) );
  OR2X2 OR2X2_259 ( .A(_abc_43815_n1428_bF_buf2), .B(_abc_43815_n1448), .Y(_abc_43815_n1449) );
  OR2X2 OR2X2_2590 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4589) );
  OR2X2 OR2X2_2591 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4593) );
  OR2X2 OR2X2_2592 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4597) );
  OR2X2 OR2X2_2593 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4601) );
  OR2X2 OR2X2_2594 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4605) );
  OR2X2 OR2X2_2595 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4609) );
  OR2X2 OR2X2_2596 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4613_1) );
  OR2X2 OR2X2_2597 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4617) );
  OR2X2 OR2X2_2598 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4621) );
  OR2X2 OR2X2_2599 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4625) );
  OR2X2 OR2X2_26 ( .A(_abc_43815_n735), .B(_abc_43815_n736), .Y(_abc_43815_n737) );
  OR2X2 OR2X2_260 ( .A(_abc_43815_n1447), .B(_abc_43815_n1449), .Y(_abc_43815_n1450) );
  OR2X2 OR2X2_2600 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4629) );
  OR2X2 OR2X2_2601 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4633) );
  OR2X2 OR2X2_2602 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4637) );
  OR2X2 OR2X2_2603 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4641) );
  OR2X2 OR2X2_2604 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4645) );
  OR2X2 OR2X2_2605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4649) );
  OR2X2 OR2X2_2606 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4653) );
  OR2X2 OR2X2_2607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4657) );
  OR2X2 OR2X2_2608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4661) );
  OR2X2 OR2X2_2609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4665) );
  OR2X2 OR2X2_261 ( .A(_abc_43815_n1431_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_43815_n1451) );
  OR2X2 OR2X2_2610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4669) );
  OR2X2 OR2X2_2611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4673_1) );
  OR2X2 OR2X2_2612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4677) );
  OR2X2 OR2X2_2613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4681) );
  OR2X2 OR2X2_2614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4685) );
  OR2X2 OR2X2_2615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4564_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4689) );
  OR2X2 OR2X2_2616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4694) );
  OR2X2 OR2X2_2617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4696) );
  OR2X2 OR2X2_2618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4698) );
  OR2X2 OR2X2_2619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4699) );
  OR2X2 OR2X2_262 ( .A(_abc_43815_n1350_bF_buf0), .B(_abc_43815_n1452), .Y(_abc_43815_n1453) );
  OR2X2 OR2X2_2620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4701) );
  OR2X2 OR2X2_2621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4702) );
  OR2X2 OR2X2_2622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4704) );
  OR2X2 OR2X2_2623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4705) );
  OR2X2 OR2X2_2624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4707) );
  OR2X2 OR2X2_2625 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4708) );
  OR2X2 OR2X2_2626 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4710) );
  OR2X2 OR2X2_2627 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4711) );
  OR2X2 OR2X2_2628 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4713) );
  OR2X2 OR2X2_2629 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4714) );
  OR2X2 OR2X2_263 ( .A(_abc_43815_n1278_bF_buf0), .B(next_pc_r_1_), .Y(_abc_43815_n1456) );
  OR2X2 OR2X2_2630 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4716) );
  OR2X2 OR2X2_2631 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4717) );
  OR2X2 OR2X2_2632 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4719) );
  OR2X2 OR2X2_2633 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4720) );
  OR2X2 OR2X2_2634 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4722) );
  OR2X2 OR2X2_2635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4723) );
  OR2X2 OR2X2_2636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4725) );
  OR2X2 OR2X2_2637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4726) );
  OR2X2 OR2X2_2638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4728) );
  OR2X2 OR2X2_2639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4729) );
  OR2X2 OR2X2_264 ( .A(_abc_43815_n1455), .B(_abc_43815_n1456), .Y(_abc_43815_n1457) );
  OR2X2 OR2X2_2640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4731) );
  OR2X2 OR2X2_2641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4732) );
  OR2X2 OR2X2_2642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4734) );
  OR2X2 OR2X2_2643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4735) );
  OR2X2 OR2X2_2644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4737) );
  OR2X2 OR2X2_2645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4738) );
  OR2X2 OR2X2_2646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4740) );
  OR2X2 OR2X2_2647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4741) );
  OR2X2 OR2X2_2648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4743) );
  OR2X2 OR2X2_2649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4744) );
  OR2X2 OR2X2_265 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_1_), .Y(_abc_43815_n1458) );
  OR2X2 OR2X2_2650 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4746) );
  OR2X2 OR2X2_2651 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4747) );
  OR2X2 OR2X2_2652 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4749) );
  OR2X2 OR2X2_2653 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4750) );
  OR2X2 OR2X2_2654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4752) );
  OR2X2 OR2X2_2655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4753) );
  OR2X2 OR2X2_2656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4755) );
  OR2X2 OR2X2_2657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4756) );
  OR2X2 OR2X2_2658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4758) );
  OR2X2 OR2X2_2659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4759) );
  OR2X2 OR2X2_266 ( .A(_abc_43815_n1468), .B(_abc_43815_n1469), .Y(_abc_43815_n1470) );
  OR2X2 OR2X2_2660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4761) );
  OR2X2 OR2X2_2661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4762) );
  OR2X2 OR2X2_2662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4764) );
  OR2X2 OR2X2_2663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4765) );
  OR2X2 OR2X2_2664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4767) );
  OR2X2 OR2X2_2665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4768) );
  OR2X2 OR2X2_2666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4770) );
  OR2X2 OR2X2_2667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4771) );
  OR2X2 OR2X2_2668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4773) );
  OR2X2 OR2X2_2669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4774) );
  OR2X2 OR2X2_267 ( .A(_abc_43815_n1470), .B(_abc_43815_n1075), .Y(_abc_43815_n1471) );
  OR2X2 OR2X2_2670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4776) );
  OR2X2 OR2X2_2671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4777) );
  OR2X2 OR2X2_2672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4779) );
  OR2X2 OR2X2_2673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4780) );
  OR2X2 OR2X2_2674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4782) );
  OR2X2 OR2X2_2675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4783) );
  OR2X2 OR2X2_2676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4785) );
  OR2X2 OR2X2_2677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4786) );
  OR2X2 OR2X2_2678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4693_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4788) );
  OR2X2 OR2X2_2679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4695_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n4789) );
  OR2X2 OR2X2_268 ( .A(alu_op_r_0_), .B(pc_q_2_), .Y(_abc_43815_n1476) );
  OR2X2 OR2X2_2680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4792) );
  OR2X2 OR2X2_2681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4794) );
  OR2X2 OR2X2_2682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4796) );
  OR2X2 OR2X2_2683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4797) );
  OR2X2 OR2X2_2684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4799) );
  OR2X2 OR2X2_2685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4800) );
  OR2X2 OR2X2_2686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4802) );
  OR2X2 OR2X2_2687 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4803) );
  OR2X2 OR2X2_2688 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4805) );
  OR2X2 OR2X2_2689 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4806) );
  OR2X2 OR2X2_269 ( .A(_abc_43815_n1428_bF_buf1), .B(_abc_43815_n1479), .Y(_abc_43815_n1480) );
  OR2X2 OR2X2_2690 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4808) );
  OR2X2 OR2X2_2691 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4809) );
  OR2X2 OR2X2_2692 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4811) );
  OR2X2 OR2X2_2693 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4812) );
  OR2X2 OR2X2_2694 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4814) );
  OR2X2 OR2X2_2695 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4815) );
  OR2X2 OR2X2_2696 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4817) );
  OR2X2 OR2X2_2697 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4818) );
  OR2X2 OR2X2_2698 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4820) );
  OR2X2 OR2X2_2699 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4821) );
  OR2X2 OR2X2_27 ( .A(_abc_43815_n738), .B(_abc_43815_n739), .Y(_abc_43815_n740) );
  OR2X2 OR2X2_270 ( .A(_abc_43815_n1478), .B(_abc_43815_n1480), .Y(_abc_43815_n1481) );
  OR2X2 OR2X2_2700 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4823_1) );
  OR2X2 OR2X2_2701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4824) );
  OR2X2 OR2X2_2702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4826) );
  OR2X2 OR2X2_2703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4827) );
  OR2X2 OR2X2_2704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4829) );
  OR2X2 OR2X2_2705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4830) );
  OR2X2 OR2X2_2706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4832) );
  OR2X2 OR2X2_2707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4833) );
  OR2X2 OR2X2_2708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4835) );
  OR2X2 OR2X2_2709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4836) );
  OR2X2 OR2X2_271 ( .A(_abc_43815_n1431_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_43815_n1482) );
  OR2X2 OR2X2_2710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4838) );
  OR2X2 OR2X2_2711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4839) );
  OR2X2 OR2X2_2712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4841) );
  OR2X2 OR2X2_2713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4842) );
  OR2X2 OR2X2_2714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4844) );
  OR2X2 OR2X2_2715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4845) );
  OR2X2 OR2X2_2716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4847) );
  OR2X2 OR2X2_2717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4848) );
  OR2X2 OR2X2_2718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4850) );
  OR2X2 OR2X2_2719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4851) );
  OR2X2 OR2X2_272 ( .A(_abc_43815_n1473_bF_buf4), .B(_abc_43815_n1483), .Y(_abc_43815_n1484) );
  OR2X2 OR2X2_2720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4853_1) );
  OR2X2 OR2X2_2721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4854) );
  OR2X2 OR2X2_2722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4856) );
  OR2X2 OR2X2_2723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4857) );
  OR2X2 OR2X2_2724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4859) );
  OR2X2 OR2X2_2725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4860) );
  OR2X2 OR2X2_2726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4862) );
  OR2X2 OR2X2_2727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4863) );
  OR2X2 OR2X2_2728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4865) );
  OR2X2 OR2X2_2729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4866) );
  OR2X2 OR2X2_273 ( .A(_abc_43815_n1472_1_bF_buf3), .B(_abc_43815_n1485), .Y(_abc_43815_n1486) );
  OR2X2 OR2X2_2730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4868) );
  OR2X2 OR2X2_2731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4869) );
  OR2X2 OR2X2_2732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4871) );
  OR2X2 OR2X2_2733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4872) );
  OR2X2 OR2X2_2734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4874) );
  OR2X2 OR2X2_2735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4875) );
  OR2X2 OR2X2_2736 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4877) );
  OR2X2 OR2X2_2737 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4878) );
  OR2X2 OR2X2_2738 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4880) );
  OR2X2 OR2X2_2739 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4881) );
  OR2X2 OR2X2_274 ( .A(_abc_43815_n1487), .B(_abc_43815_n1350_bF_buf4), .Y(_abc_43815_n1488) );
  OR2X2 OR2X2_2740 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4883_1) );
  OR2X2 OR2X2_2741 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4884) );
  OR2X2 OR2X2_2742 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4791_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4886) );
  OR2X2 OR2X2_2743 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4793_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n4887) );
  OR2X2 OR2X2_2744 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4890) );
  OR2X2 OR2X2_2745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4894) );
  OR2X2 OR2X2_2746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4898) );
  OR2X2 OR2X2_2747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4902) );
  OR2X2 OR2X2_2748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4906) );
  OR2X2 OR2X2_2749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4910) );
  OR2X2 OR2X2_275 ( .A(_abc_43815_n1490), .B(_abc_43815_n1491_1), .Y(_abc_43815_n1492_1) );
  OR2X2 OR2X2_2750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4914) );
  OR2X2 OR2X2_2751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4918) );
  OR2X2 OR2X2_2752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4922) );
  OR2X2 OR2X2_2753 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4926) );
  OR2X2 OR2X2_2754 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4930) );
  OR2X2 OR2X2_2755 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4934) );
  OR2X2 OR2X2_2756 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4938) );
  OR2X2 OR2X2_2757 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4942) );
  OR2X2 OR2X2_2758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4946) );
  OR2X2 OR2X2_2759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4950) );
  OR2X2 OR2X2_276 ( .A(_abc_43815_n1413_bF_buf2), .B(_abc_43815_n1492_1), .Y(_abc_43815_n1493) );
  OR2X2 OR2X2_2760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4954) );
  OR2X2 OR2X2_2761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4958) );
  OR2X2 OR2X2_2762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4962) );
  OR2X2 OR2X2_2763 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4966) );
  OR2X2 OR2X2_2764 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4970) );
  OR2X2 OR2X2_2765 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4974) );
  OR2X2 OR2X2_2766 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4978) );
  OR2X2 OR2X2_2767 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4982) );
  OR2X2 OR2X2_2768 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4986) );
  OR2X2 OR2X2_2769 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4990) );
  OR2X2 OR2X2_277 ( .A(_abc_43815_n1494), .B(_abc_43815_n1461_bF_buf3), .Y(_abc_43815_n1495) );
  OR2X2 OR2X2_2770 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4994) );
  OR2X2 OR2X2_2771 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n4998) );
  OR2X2 OR2X2_2772 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5002) );
  OR2X2 OR2X2_2773 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5006) );
  OR2X2 OR2X2_2774 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5010) );
  OR2X2 OR2X2_2775 ( .A(REGFILE_SIM_reg_bank__abc_33898_n4889_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5014) );
  OR2X2 OR2X2_2776 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5019) );
  OR2X2 OR2X2_2777 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5023) );
  OR2X2 OR2X2_2778 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5027) );
  OR2X2 OR2X2_2779 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5031) );
  OR2X2 OR2X2_278 ( .A(_abc_43815_n1351_bF_buf4), .B(_abc_43815_n1485), .Y(_abc_43815_n1496) );
  OR2X2 OR2X2_2780 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5035) );
  OR2X2 OR2X2_2781 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5039) );
  OR2X2 OR2X2_2782 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5043) );
  OR2X2 OR2X2_2783 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5047) );
  OR2X2 OR2X2_2784 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5051) );
  OR2X2 OR2X2_2785 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5055) );
  OR2X2 OR2X2_2786 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5059) );
  OR2X2 OR2X2_2787 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5063_1) );
  OR2X2 OR2X2_2788 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5067) );
  OR2X2 OR2X2_2789 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5071) );
  OR2X2 OR2X2_279 ( .A(_abc_43815_n1497), .B(_abc_43815_n1278_bF_buf7), .Y(_abc_43815_n1498) );
  OR2X2 OR2X2_2790 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5075) );
  OR2X2 OR2X2_2791 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5079) );
  OR2X2 OR2X2_2792 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5083) );
  OR2X2 OR2X2_2793 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5087) );
  OR2X2 OR2X2_2794 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5091) );
  OR2X2 OR2X2_2795 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5095) );
  OR2X2 OR2X2_2796 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5099) );
  OR2X2 OR2X2_2797 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5103) );
  OR2X2 OR2X2_2798 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5107) );
  OR2X2 OR2X2_2799 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5111) );
  OR2X2 OR2X2_28 ( .A(_abc_43815_n737), .B(_abc_43815_n740), .Y(_abc_43815_n741) );
  OR2X2 OR2X2_280 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_2_), .Y(_abc_43815_n1499) );
  OR2X2 OR2X2_2800 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5115) );
  OR2X2 OR2X2_2801 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5119) );
  OR2X2 OR2X2_2802 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5123_1) );
  OR2X2 OR2X2_2803 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5127) );
  OR2X2 OR2X2_2804 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5131) );
  OR2X2 OR2X2_2805 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5135) );
  OR2X2 OR2X2_2806 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5139) );
  OR2X2 OR2X2_2807 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5018_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5143) );
  OR2X2 OR2X2_2808 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5148) );
  OR2X2 OR2X2_2809 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5150) );
  OR2X2 OR2X2_281 ( .A(_abc_43815_n1418_bF_buf5), .B(epc_q_3_), .Y(_abc_43815_n1502) );
  OR2X2 OR2X2_2810 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5152) );
  OR2X2 OR2X2_2811 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5153_1) );
  OR2X2 OR2X2_2812 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5155) );
  OR2X2 OR2X2_2813 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5156) );
  OR2X2 OR2X2_2814 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5158) );
  OR2X2 OR2X2_2815 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5159) );
  OR2X2 OR2X2_2816 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5161) );
  OR2X2 OR2X2_2817 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5162) );
  OR2X2 OR2X2_2818 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5164) );
  OR2X2 OR2X2_2819 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5165) );
  OR2X2 OR2X2_282 ( .A(_abc_43815_n1413_bF_buf1), .B(_abc_43815_n1506), .Y(_abc_43815_n1507) );
  OR2X2 OR2X2_2820 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5167) );
  OR2X2 OR2X2_2821 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5168) );
  OR2X2 OR2X2_2822 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5170) );
  OR2X2 OR2X2_2823 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5171) );
  OR2X2 OR2X2_2824 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5173) );
  OR2X2 OR2X2_2825 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5174) );
  OR2X2 OR2X2_2826 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5176) );
  OR2X2 OR2X2_2827 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5177) );
  OR2X2 OR2X2_2828 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5179) );
  OR2X2 OR2X2_2829 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5180) );
  OR2X2 OR2X2_283 ( .A(_abc_43815_n1431_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_43815_n1508) );
  OR2X2 OR2X2_2830 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5182) );
  OR2X2 OR2X2_2831 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5183_1) );
  OR2X2 OR2X2_2832 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5185) );
  OR2X2 OR2X2_2833 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5186) );
  OR2X2 OR2X2_2834 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5188) );
  OR2X2 OR2X2_2835 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5189) );
  OR2X2 OR2X2_2836 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5191) );
  OR2X2 OR2X2_2837 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5192) );
  OR2X2 OR2X2_2838 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5194) );
  OR2X2 OR2X2_2839 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5195) );
  OR2X2 OR2X2_284 ( .A(alu_op_r_1_), .B(pc_q_3_), .Y(_abc_43815_n1509) );
  OR2X2 OR2X2_2840 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5197) );
  OR2X2 OR2X2_2841 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5198) );
  OR2X2 OR2X2_2842 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5200) );
  OR2X2 OR2X2_2843 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5201) );
  OR2X2 OR2X2_2844 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5203) );
  OR2X2 OR2X2_2845 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5204) );
  OR2X2 OR2X2_2846 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5206) );
  OR2X2 OR2X2_2847 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5207) );
  OR2X2 OR2X2_2848 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5209) );
  OR2X2 OR2X2_2849 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5210) );
  OR2X2 OR2X2_285 ( .A(_abc_43815_n1512), .B(_abc_43815_n1474), .Y(_abc_43815_n1515_1) );
  OR2X2 OR2X2_2850 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5212) );
  OR2X2 OR2X2_2851 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5213_1) );
  OR2X2 OR2X2_2852 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5215) );
  OR2X2 OR2X2_2853 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5216) );
  OR2X2 OR2X2_2854 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5218) );
  OR2X2 OR2X2_2855 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5219) );
  OR2X2 OR2X2_2856 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5221) );
  OR2X2 OR2X2_2857 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5222) );
  OR2X2 OR2X2_2858 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5224) );
  OR2X2 OR2X2_2859 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5225) );
  OR2X2 OR2X2_286 ( .A(_abc_43815_n1428_bF_buf0), .B(_abc_43815_n1518_1), .Y(_abc_43815_n1519) );
  OR2X2 OR2X2_2860 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5227) );
  OR2X2 OR2X2_2861 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5228) );
  OR2X2 OR2X2_2862 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5230) );
  OR2X2 OR2X2_2863 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5231) );
  OR2X2 OR2X2_2864 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5233) );
  OR2X2 OR2X2_2865 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5234) );
  OR2X2 OR2X2_2866 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5236) );
  OR2X2 OR2X2_2867 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5237) );
  OR2X2 OR2X2_2868 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5239) );
  OR2X2 OR2X2_2869 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5240) );
  OR2X2 OR2X2_287 ( .A(_abc_43815_n1517), .B(_abc_43815_n1519), .Y(_abc_43815_n1520) );
  OR2X2 OR2X2_2870 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5147_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5242) );
  OR2X2 OR2X2_2871 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5149_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_33898_n5243_1) );
  OR2X2 OR2X2_2872 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5246) );
  OR2X2 OR2X2_2873 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5248) );
  OR2X2 OR2X2_2874 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5250) );
  OR2X2 OR2X2_2875 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5251) );
  OR2X2 OR2X2_2876 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5253) );
  OR2X2 OR2X2_2877 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5254) );
  OR2X2 OR2X2_2878 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5256) );
  OR2X2 OR2X2_2879 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5257) );
  OR2X2 OR2X2_288 ( .A(_abc_43815_n1473_bF_buf3), .B(_abc_43815_n1521), .Y(_abc_43815_n1522) );
  OR2X2 OR2X2_2880 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5259) );
  OR2X2 OR2X2_2881 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5260) );
  OR2X2 OR2X2_2882 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5262) );
  OR2X2 OR2X2_2883 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5263) );
  OR2X2 OR2X2_2884 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5265) );
  OR2X2 OR2X2_2885 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5266) );
  OR2X2 OR2X2_2886 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5268) );
  OR2X2 OR2X2_2887 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5269) );
  OR2X2 OR2X2_2888 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5271) );
  OR2X2 OR2X2_2889 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5272) );
  OR2X2 OR2X2_289 ( .A(pc_q_2_), .B(pc_q_3_), .Y(_abc_43815_n1523) );
  OR2X2 OR2X2_2890 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5274) );
  OR2X2 OR2X2_2891 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5275) );
  OR2X2 OR2X2_2892 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5277) );
  OR2X2 OR2X2_2893 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5278) );
  OR2X2 OR2X2_2894 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5280) );
  OR2X2 OR2X2_2895 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5281) );
  OR2X2 OR2X2_2896 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5283) );
  OR2X2 OR2X2_2897 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5284) );
  OR2X2 OR2X2_2898 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5286) );
  OR2X2 OR2X2_2899 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5287) );
  OR2X2 OR2X2_29 ( .A(_abc_43815_n734), .B(_abc_43815_n742), .Y(_abc_43815_n743) );
  OR2X2 OR2X2_290 ( .A(_abc_43815_n1472_1_bF_buf2), .B(_abc_43815_n1526), .Y(_abc_43815_n1527) );
  OR2X2 OR2X2_2900 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5289) );
  OR2X2 OR2X2_2901 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5290) );
  OR2X2 OR2X2_2902 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5292) );
  OR2X2 OR2X2_2903 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5293) );
  OR2X2 OR2X2_2904 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5295) );
  OR2X2 OR2X2_2905 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5296) );
  OR2X2 OR2X2_2906 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5298) );
  OR2X2 OR2X2_2907 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5299) );
  OR2X2 OR2X2_2908 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5301) );
  OR2X2 OR2X2_2909 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5302) );
  OR2X2 OR2X2_291 ( .A(_abc_43815_n1528), .B(_abc_43815_n1350_bF_buf3), .Y(_abc_43815_n1529) );
  OR2X2 OR2X2_2910 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5304) );
  OR2X2 OR2X2_2911 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5305) );
  OR2X2 OR2X2_2912 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5307) );
  OR2X2 OR2X2_2913 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5308) );
  OR2X2 OR2X2_2914 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5310) );
  OR2X2 OR2X2_2915 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5311) );
  OR2X2 OR2X2_2916 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5313) );
  OR2X2 OR2X2_2917 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5314) );
  OR2X2 OR2X2_2918 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5316) );
  OR2X2 OR2X2_2919 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5317) );
  OR2X2 OR2X2_292 ( .A(_abc_43815_n1530), .B(_abc_43815_n1461_bF_buf2), .Y(_abc_43815_n1531) );
  OR2X2 OR2X2_2920 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5319) );
  OR2X2 OR2X2_2921 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5320) );
  OR2X2 OR2X2_2922 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5322) );
  OR2X2 OR2X2_2923 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5323) );
  OR2X2 OR2X2_2924 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5325) );
  OR2X2 OR2X2_2925 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5326) );
  OR2X2 OR2X2_2926 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5328) );
  OR2X2 OR2X2_2927 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5329) );
  OR2X2 OR2X2_2928 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5331) );
  OR2X2 OR2X2_2929 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5332) );
  OR2X2 OR2X2_293 ( .A(_abc_43815_n1351_bF_buf3), .B(_abc_43815_n1526), .Y(_abc_43815_n1532) );
  OR2X2 OR2X2_2930 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5334) );
  OR2X2 OR2X2_2931 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5335) );
  OR2X2 OR2X2_2932 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5337) );
  OR2X2 OR2X2_2933 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5338) );
  OR2X2 OR2X2_2934 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5245_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5340) );
  OR2X2 OR2X2_2935 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5247_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_33898_n5341) );
  OR2X2 OR2X2_2936 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5344) );
  OR2X2 OR2X2_2937 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5346) );
  OR2X2 OR2X2_2938 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5348) );
  OR2X2 OR2X2_2939 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5349) );
  OR2X2 OR2X2_294 ( .A(_abc_43815_n1533), .B(_abc_43815_n1278_bF_buf6), .Y(_abc_43815_n1534_1) );
  OR2X2 OR2X2_2940 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5351) );
  OR2X2 OR2X2_2941 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5352) );
  OR2X2 OR2X2_2942 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5354) );
  OR2X2 OR2X2_2943 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5355) );
  OR2X2 OR2X2_2944 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5357) );
  OR2X2 OR2X2_2945 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5358) );
  OR2X2 OR2X2_2946 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5360) );
  OR2X2 OR2X2_2947 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5361) );
  OR2X2 OR2X2_2948 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5363) );
  OR2X2 OR2X2_2949 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5364) );
  OR2X2 OR2X2_295 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_3_), .Y(_abc_43815_n1535_1) );
  OR2X2 OR2X2_2950 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5366) );
  OR2X2 OR2X2_2951 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5367) );
  OR2X2 OR2X2_2952 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5369) );
  OR2X2 OR2X2_2953 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5370) );
  OR2X2 OR2X2_2954 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5372) );
  OR2X2 OR2X2_2955 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5373) );
  OR2X2 OR2X2_2956 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5375) );
  OR2X2 OR2X2_2957 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5376) );
  OR2X2 OR2X2_2958 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5378) );
  OR2X2 OR2X2_2959 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5379) );
  OR2X2 OR2X2_296 ( .A(_abc_43815_n1418_bF_buf3), .B(epc_q_4_), .Y(_abc_43815_n1538) );
  OR2X2 OR2X2_2960 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5381) );
  OR2X2 OR2X2_2961 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5382) );
  OR2X2 OR2X2_2962 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5384) );
  OR2X2 OR2X2_2963 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5385) );
  OR2X2 OR2X2_2964 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5387) );
  OR2X2 OR2X2_2965 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5388) );
  OR2X2 OR2X2_2966 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5390) );
  OR2X2 OR2X2_2967 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5391) );
  OR2X2 OR2X2_2968 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5393) );
  OR2X2 OR2X2_2969 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5394) );
  OR2X2 OR2X2_297 ( .A(_abc_43815_n1413_bF_buf0), .B(_abc_43815_n1542), .Y(_abc_43815_n1543) );
  OR2X2 OR2X2_2970 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5396) );
  OR2X2 OR2X2_2971 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5397) );
  OR2X2 OR2X2_2972 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5399) );
  OR2X2 OR2X2_2973 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5400) );
  OR2X2 OR2X2_2974 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5402) );
  OR2X2 OR2X2_2975 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5403) );
  OR2X2 OR2X2_2976 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5405) );
  OR2X2 OR2X2_2977 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5406) );
  OR2X2 OR2X2_2978 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5408) );
  OR2X2 OR2X2_2979 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5409) );
  OR2X2 OR2X2_298 ( .A(_abc_43815_n1431_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_43815_n1544) );
  OR2X2 OR2X2_2980 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5411) );
  OR2X2 OR2X2_2981 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5412) );
  OR2X2 OR2X2_2982 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5414) );
  OR2X2 OR2X2_2983 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5415) );
  OR2X2 OR2X2_2984 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5417) );
  OR2X2 OR2X2_2985 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5418) );
  OR2X2 OR2X2_2986 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5420) );
  OR2X2 OR2X2_2987 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5421) );
  OR2X2 OR2X2_2988 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5423) );
  OR2X2 OR2X2_2989 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5424) );
  OR2X2 OR2X2_299 ( .A(_abc_43815_n1513), .B(_abc_43815_n1510), .Y(_abc_43815_n1545) );
  OR2X2 OR2X2_2990 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5426) );
  OR2X2 OR2X2_2991 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5427) );
  OR2X2 OR2X2_2992 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5429) );
  OR2X2 OR2X2_2993 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5430) );
  OR2X2 OR2X2_2994 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5432) );
  OR2X2 OR2X2_2995 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5433) );
  OR2X2 OR2X2_2996 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5435) );
  OR2X2 OR2X2_2997 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5436) );
  OR2X2 OR2X2_2998 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5343_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5438) );
  OR2X2 OR2X2_2999 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5345_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_33898_n5439) );
  OR2X2 OR2X2_3 ( .A(_abc_43815_n658), .B(_abc_43815_n660), .Y(_abc_43815_n661) );
  OR2X2 OR2X2_30 ( .A(_abc_43815_n744), .B(_abc_43815_n730_1), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_) );
  OR2X2 OR2X2_300 ( .A(alu_op_r_2_), .B(pc_q_4_), .Y(_abc_43815_n1546) );
  OR2X2 OR2X2_3000 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5442) );
  OR2X2 OR2X2_3001 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5444) );
  OR2X2 OR2X2_3002 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5446) );
  OR2X2 OR2X2_3003 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5447) );
  OR2X2 OR2X2_3004 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5449) );
  OR2X2 OR2X2_3005 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5450) );
  OR2X2 OR2X2_3006 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5452) );
  OR2X2 OR2X2_3007 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5453) );
  OR2X2 OR2X2_3008 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5455) );
  OR2X2 OR2X2_3009 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5456) );
  OR2X2 OR2X2_301 ( .A(_abc_43815_n1545), .B(_abc_43815_n1549), .Y(_abc_43815_n1550_1) );
  OR2X2 OR2X2_3010 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5458) );
  OR2X2 OR2X2_3011 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5459) );
  OR2X2 OR2X2_3012 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5461) );
  OR2X2 OR2X2_3013 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5462) );
  OR2X2 OR2X2_3014 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5464) );
  OR2X2 OR2X2_3015 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5465) );
  OR2X2 OR2X2_3016 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5467) );
  OR2X2 OR2X2_3017 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5468) );
  OR2X2 OR2X2_3018 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5470) );
  OR2X2 OR2X2_3019 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5471) );
  OR2X2 OR2X2_302 ( .A(_abc_43815_n1428_bF_buf4), .B(_abc_43815_n1555), .Y(_abc_43815_n1556) );
  OR2X2 OR2X2_3020 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5473) );
  OR2X2 OR2X2_3021 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5474) );
  OR2X2 OR2X2_3022 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5476) );
  OR2X2 OR2X2_3023 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5477) );
  OR2X2 OR2X2_3024 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5479) );
  OR2X2 OR2X2_3025 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5480) );
  OR2X2 OR2X2_3026 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5482) );
  OR2X2 OR2X2_3027 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5483) );
  OR2X2 OR2X2_3028 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5485) );
  OR2X2 OR2X2_3029 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5486) );
  OR2X2 OR2X2_303 ( .A(_abc_43815_n1554), .B(_abc_43815_n1556), .Y(_abc_43815_n1557) );
  OR2X2 OR2X2_3030 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5488) );
  OR2X2 OR2X2_3031 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5489) );
  OR2X2 OR2X2_3032 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5491) );
  OR2X2 OR2X2_3033 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5492) );
  OR2X2 OR2X2_3034 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5494) );
  OR2X2 OR2X2_3035 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5495) );
  OR2X2 OR2X2_3036 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5497) );
  OR2X2 OR2X2_3037 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5498) );
  OR2X2 OR2X2_3038 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5500) );
  OR2X2 OR2X2_3039 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5501) );
  OR2X2 OR2X2_304 ( .A(_abc_43815_n1473_bF_buf2), .B(_abc_43815_n1558), .Y(_abc_43815_n1559) );
  OR2X2 OR2X2_3040 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5503) );
  OR2X2 OR2X2_3041 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5504) );
  OR2X2 OR2X2_3042 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5506) );
  OR2X2 OR2X2_3043 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5507) );
  OR2X2 OR2X2_3044 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5509) );
  OR2X2 OR2X2_3045 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5510) );
  OR2X2 OR2X2_3046 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5512) );
  OR2X2 OR2X2_3047 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5513) );
  OR2X2 OR2X2_3048 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5515) );
  OR2X2 OR2X2_3049 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5516) );
  OR2X2 OR2X2_305 ( .A(_abc_43815_n1524), .B(pc_q_4_), .Y(_abc_43815_n1560) );
  OR2X2 OR2X2_3050 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5518) );
  OR2X2 OR2X2_3051 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5519) );
  OR2X2 OR2X2_3052 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5521) );
  OR2X2 OR2X2_3053 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5522) );
  OR2X2 OR2X2_3054 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5524) );
  OR2X2 OR2X2_3055 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5525) );
  OR2X2 OR2X2_3056 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5527) );
  OR2X2 OR2X2_3057 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5528) );
  OR2X2 OR2X2_3058 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5530) );
  OR2X2 OR2X2_3059 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5531) );
  OR2X2 OR2X2_306 ( .A(_abc_43815_n1472_1_bF_buf1), .B(_abc_43815_n1563), .Y(_abc_43815_n1564) );
  OR2X2 OR2X2_3060 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5533) );
  OR2X2 OR2X2_3061 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5534) );
  OR2X2 OR2X2_3062 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5441_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .Y(REGFILE_SIM_reg_bank__abc_33898_n5536) );
  OR2X2 OR2X2_3063 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5443_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_33898_n5537) );
  OR2X2 OR2X2_3064 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5546), .B(REGFILE_SIM_reg_bank__abc_33898_n5549), .Y(REGFILE_SIM_reg_bank__abc_33898_n5550) );
  OR2X2 OR2X2_3065 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5555), .B(REGFILE_SIM_reg_bank__abc_33898_n5558), .Y(REGFILE_SIM_reg_bank__abc_33898_n5559) );
  OR2X2 OR2X2_3066 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5559), .B(REGFILE_SIM_reg_bank__abc_33898_n5550), .Y(REGFILE_SIM_reg_bank__abc_33898_n5560) );
  OR2X2 OR2X2_3067 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5566), .B(REGFILE_SIM_reg_bank__abc_33898_n5569), .Y(REGFILE_SIM_reg_bank__abc_33898_n5570) );
  OR2X2 OR2X2_3068 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5574), .B(REGFILE_SIM_reg_bank__abc_33898_n5577), .Y(REGFILE_SIM_reg_bank__abc_33898_n5578) );
  OR2X2 OR2X2_3069 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5570), .B(REGFILE_SIM_reg_bank__abc_33898_n5578), .Y(REGFILE_SIM_reg_bank__abc_33898_n5579) );
  OR2X2 OR2X2_307 ( .A(_abc_43815_n1565), .B(_abc_43815_n1350_bF_buf2), .Y(_abc_43815_n1566_1) );
  OR2X2 OR2X2_3070 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5560), .B(REGFILE_SIM_reg_bank__abc_33898_n5579), .Y(REGFILE_SIM_reg_bank__abc_33898_n5580) );
  OR2X2 OR2X2_3071 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5582), .B(REGFILE_SIM_reg_bank__abc_33898_n5584), .Y(REGFILE_SIM_reg_bank__abc_33898_n5585) );
  OR2X2 OR2X2_3072 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5588), .B(REGFILE_SIM_reg_bank__abc_33898_n5591), .Y(REGFILE_SIM_reg_bank__abc_33898_n5592) );
  OR2X2 OR2X2_3073 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5585), .B(REGFILE_SIM_reg_bank__abc_33898_n5592), .Y(REGFILE_SIM_reg_bank__abc_33898_n5593) );
  OR2X2 OR2X2_3074 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5595), .B(REGFILE_SIM_reg_bank__abc_33898_n5598), .Y(REGFILE_SIM_reg_bank__abc_33898_n5599) );
  OR2X2 OR2X2_3075 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5601), .B(REGFILE_SIM_reg_bank__abc_33898_n5604), .Y(REGFILE_SIM_reg_bank__abc_33898_n5605) );
  OR2X2 OR2X2_3076 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5605), .B(REGFILE_SIM_reg_bank__abc_33898_n5599), .Y(REGFILE_SIM_reg_bank__abc_33898_n5606) );
  OR2X2 OR2X2_3077 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5593), .B(REGFILE_SIM_reg_bank__abc_33898_n5606), .Y(REGFILE_SIM_reg_bank__abc_33898_n5607) );
  OR2X2 OR2X2_3078 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5580), .B(REGFILE_SIM_reg_bank__abc_33898_n5607), .Y(REGFILE_SIM_reg_bank__abc_33898_n5608) );
  OR2X2 OR2X2_3079 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5611), .B(REGFILE_SIM_reg_bank__abc_33898_n5614), .Y(REGFILE_SIM_reg_bank__abc_33898_n5615) );
  OR2X2 OR2X2_308 ( .A(_abc_43815_n1567_1), .B(_abc_43815_n1461_bF_buf1), .Y(_abc_43815_n1568) );
  OR2X2 OR2X2_3080 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5617), .B(REGFILE_SIM_reg_bank__abc_33898_n5619), .Y(REGFILE_SIM_reg_bank__abc_33898_n5620) );
  OR2X2 OR2X2_3081 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5615), .B(REGFILE_SIM_reg_bank__abc_33898_n5620), .Y(REGFILE_SIM_reg_bank__abc_33898_n5621) );
  OR2X2 OR2X2_3082 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5626), .B(REGFILE_SIM_reg_bank__abc_33898_n5628), .Y(REGFILE_SIM_reg_bank__abc_33898_n5629) );
  OR2X2 OR2X2_3083 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5629), .B(REGFILE_SIM_reg_bank__abc_33898_n5624), .Y(REGFILE_SIM_reg_bank__abc_33898_n5630) );
  OR2X2 OR2X2_3084 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5621), .B(REGFILE_SIM_reg_bank__abc_33898_n5630), .Y(REGFILE_SIM_reg_bank__abc_33898_n5631) );
  OR2X2 OR2X2_3085 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5633), .B(REGFILE_SIM_reg_bank__abc_33898_n5635), .Y(REGFILE_SIM_reg_bank__abc_33898_n5636) );
  OR2X2 OR2X2_3086 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5638), .B(REGFILE_SIM_reg_bank__abc_33898_n5640), .Y(REGFILE_SIM_reg_bank__abc_33898_n5641) );
  OR2X2 OR2X2_3087 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5641), .B(REGFILE_SIM_reg_bank__abc_33898_n5636), .Y(REGFILE_SIM_reg_bank__abc_33898_n5642) );
  OR2X2 OR2X2_3088 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5644), .B(REGFILE_SIM_reg_bank__abc_33898_n5646), .Y(REGFILE_SIM_reg_bank__abc_33898_n5647) );
  OR2X2 OR2X2_3089 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5649), .B(REGFILE_SIM_reg_bank__abc_33898_n5651), .Y(REGFILE_SIM_reg_bank__abc_33898_n5652) );
  OR2X2 OR2X2_309 ( .A(_abc_43815_n1351_bF_buf2), .B(_abc_43815_n1563), .Y(_abc_43815_n1569) );
  OR2X2 OR2X2_3090 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5647), .B(REGFILE_SIM_reg_bank__abc_33898_n5652), .Y(REGFILE_SIM_reg_bank__abc_33898_n5653) );
  OR2X2 OR2X2_3091 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5642), .B(REGFILE_SIM_reg_bank__abc_33898_n5653), .Y(REGFILE_SIM_reg_bank__abc_33898_n5654) );
  OR2X2 OR2X2_3092 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5654), .B(REGFILE_SIM_reg_bank__abc_33898_n5631), .Y(REGFILE_SIM_reg_bank__abc_33898_n5655) );
  OR2X2 OR2X2_3093 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5608), .B(REGFILE_SIM_reg_bank__abc_33898_n5655), .Y(REGFILE_SIM_reg_bank_reg_rb_o_0_) );
  OR2X2 OR2X2_3094 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5657), .B(REGFILE_SIM_reg_bank__abc_33898_n5658), .Y(REGFILE_SIM_reg_bank__abc_33898_n5659) );
  OR2X2 OR2X2_3095 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5660), .B(REGFILE_SIM_reg_bank__abc_33898_n5661), .Y(REGFILE_SIM_reg_bank__abc_33898_n5662) );
  OR2X2 OR2X2_3096 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5662), .B(REGFILE_SIM_reg_bank__abc_33898_n5659), .Y(REGFILE_SIM_reg_bank__abc_33898_n5663) );
  OR2X2 OR2X2_3097 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5664), .B(REGFILE_SIM_reg_bank__abc_33898_n5665), .Y(REGFILE_SIM_reg_bank__abc_33898_n5666) );
  OR2X2 OR2X2_3098 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5667), .B(REGFILE_SIM_reg_bank__abc_33898_n5668), .Y(REGFILE_SIM_reg_bank__abc_33898_n5669) );
  OR2X2 OR2X2_3099 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5666), .B(REGFILE_SIM_reg_bank__abc_33898_n5669), .Y(REGFILE_SIM_reg_bank__abc_33898_n5670) );
  OR2X2 OR2X2_31 ( .A(_abc_43815_n747), .B(_abc_43815_n748), .Y(_abc_43815_n749) );
  OR2X2 OR2X2_310 ( .A(_abc_43815_n1570), .B(_abc_43815_n1278_bF_buf5), .Y(_abc_43815_n1571) );
  OR2X2 OR2X2_3100 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5663), .B(REGFILE_SIM_reg_bank__abc_33898_n5670), .Y(REGFILE_SIM_reg_bank__abc_33898_n5671) );
  OR2X2 OR2X2_3101 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5672), .B(REGFILE_SIM_reg_bank__abc_33898_n5673), .Y(REGFILE_SIM_reg_bank__abc_33898_n5674) );
  OR2X2 OR2X2_3102 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5675), .B(REGFILE_SIM_reg_bank__abc_33898_n5676), .Y(REGFILE_SIM_reg_bank__abc_33898_n5677) );
  OR2X2 OR2X2_3103 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5674), .B(REGFILE_SIM_reg_bank__abc_33898_n5677), .Y(REGFILE_SIM_reg_bank__abc_33898_n5678) );
  OR2X2 OR2X2_3104 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5679), .B(REGFILE_SIM_reg_bank__abc_33898_n5680), .Y(REGFILE_SIM_reg_bank__abc_33898_n5681) );
  OR2X2 OR2X2_3105 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5682), .B(REGFILE_SIM_reg_bank__abc_33898_n5683), .Y(REGFILE_SIM_reg_bank__abc_33898_n5684) );
  OR2X2 OR2X2_3106 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5684), .B(REGFILE_SIM_reg_bank__abc_33898_n5681), .Y(REGFILE_SIM_reg_bank__abc_33898_n5685) );
  OR2X2 OR2X2_3107 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5678), .B(REGFILE_SIM_reg_bank__abc_33898_n5685), .Y(REGFILE_SIM_reg_bank__abc_33898_n5686) );
  OR2X2 OR2X2_3108 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5671), .B(REGFILE_SIM_reg_bank__abc_33898_n5686), .Y(REGFILE_SIM_reg_bank__abc_33898_n5687) );
  OR2X2 OR2X2_3109 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5688), .B(REGFILE_SIM_reg_bank__abc_33898_n5689), .Y(REGFILE_SIM_reg_bank__abc_33898_n5690) );
  OR2X2 OR2X2_311 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_4_), .Y(_abc_43815_n1572) );
  OR2X2 OR2X2_3110 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5691), .B(REGFILE_SIM_reg_bank__abc_33898_n5692), .Y(REGFILE_SIM_reg_bank__abc_33898_n5693) );
  OR2X2 OR2X2_3111 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5690), .B(REGFILE_SIM_reg_bank__abc_33898_n5693), .Y(REGFILE_SIM_reg_bank__abc_33898_n5694) );
  OR2X2 OR2X2_3112 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5696), .B(REGFILE_SIM_reg_bank__abc_33898_n5697), .Y(REGFILE_SIM_reg_bank__abc_33898_n5698) );
  OR2X2 OR2X2_3113 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5698), .B(REGFILE_SIM_reg_bank__abc_33898_n5695), .Y(REGFILE_SIM_reg_bank__abc_33898_n5699) );
  OR2X2 OR2X2_3114 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5694), .B(REGFILE_SIM_reg_bank__abc_33898_n5699), .Y(REGFILE_SIM_reg_bank__abc_33898_n5700) );
  OR2X2 OR2X2_3115 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5701), .B(REGFILE_SIM_reg_bank__abc_33898_n5702), .Y(REGFILE_SIM_reg_bank__abc_33898_n5703) );
  OR2X2 OR2X2_3116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5704), .B(REGFILE_SIM_reg_bank__abc_33898_n5705), .Y(REGFILE_SIM_reg_bank__abc_33898_n5706) );
  OR2X2 OR2X2_3117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5706), .B(REGFILE_SIM_reg_bank__abc_33898_n5703), .Y(REGFILE_SIM_reg_bank__abc_33898_n5707) );
  OR2X2 OR2X2_3118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5708), .B(REGFILE_SIM_reg_bank__abc_33898_n5709), .Y(REGFILE_SIM_reg_bank__abc_33898_n5710) );
  OR2X2 OR2X2_3119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5711), .B(REGFILE_SIM_reg_bank__abc_33898_n5712), .Y(REGFILE_SIM_reg_bank__abc_33898_n5713) );
  OR2X2 OR2X2_312 ( .A(_abc_43815_n1418_bF_buf1), .B(epc_q_5_), .Y(_abc_43815_n1575) );
  OR2X2 OR2X2_3120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5710), .B(REGFILE_SIM_reg_bank__abc_33898_n5713), .Y(REGFILE_SIM_reg_bank__abc_33898_n5714) );
  OR2X2 OR2X2_3121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5707), .B(REGFILE_SIM_reg_bank__abc_33898_n5714), .Y(REGFILE_SIM_reg_bank__abc_33898_n5715) );
  OR2X2 OR2X2_3122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5715), .B(REGFILE_SIM_reg_bank__abc_33898_n5700), .Y(REGFILE_SIM_reg_bank__abc_33898_n5716) );
  OR2X2 OR2X2_3123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5687), .B(REGFILE_SIM_reg_bank__abc_33898_n5716), .Y(REGFILE_SIM_reg_bank_reg_rb_o_1_) );
  OR2X2 OR2X2_3124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5718), .B(REGFILE_SIM_reg_bank__abc_33898_n5719), .Y(REGFILE_SIM_reg_bank__abc_33898_n5720) );
  OR2X2 OR2X2_3125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5721), .B(REGFILE_SIM_reg_bank__abc_33898_n5722), .Y(REGFILE_SIM_reg_bank__abc_33898_n5723) );
  OR2X2 OR2X2_3126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5723), .B(REGFILE_SIM_reg_bank__abc_33898_n5720), .Y(REGFILE_SIM_reg_bank__abc_33898_n5724) );
  OR2X2 OR2X2_3127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5725), .B(REGFILE_SIM_reg_bank__abc_33898_n5726), .Y(REGFILE_SIM_reg_bank__abc_33898_n5727) );
  OR2X2 OR2X2_3128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5728), .B(REGFILE_SIM_reg_bank__abc_33898_n5729), .Y(REGFILE_SIM_reg_bank__abc_33898_n5730) );
  OR2X2 OR2X2_3129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5727), .B(REGFILE_SIM_reg_bank__abc_33898_n5730), .Y(REGFILE_SIM_reg_bank__abc_33898_n5731) );
  OR2X2 OR2X2_313 ( .A(_abc_43815_n1413_bF_buf4), .B(_abc_43815_n1579), .Y(_abc_43815_n1580) );
  OR2X2 OR2X2_3130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5724), .B(REGFILE_SIM_reg_bank__abc_33898_n5731), .Y(REGFILE_SIM_reg_bank__abc_33898_n5732) );
  OR2X2 OR2X2_3131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5733), .B(REGFILE_SIM_reg_bank__abc_33898_n5734), .Y(REGFILE_SIM_reg_bank__abc_33898_n5735) );
  OR2X2 OR2X2_3132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5736), .B(REGFILE_SIM_reg_bank__abc_33898_n5737), .Y(REGFILE_SIM_reg_bank__abc_33898_n5738) );
  OR2X2 OR2X2_3133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5735), .B(REGFILE_SIM_reg_bank__abc_33898_n5738), .Y(REGFILE_SIM_reg_bank__abc_33898_n5739) );
  OR2X2 OR2X2_3134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5740), .B(REGFILE_SIM_reg_bank__abc_33898_n5741), .Y(REGFILE_SIM_reg_bank__abc_33898_n5742) );
  OR2X2 OR2X2_3135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5743), .B(REGFILE_SIM_reg_bank__abc_33898_n5744), .Y(REGFILE_SIM_reg_bank__abc_33898_n5745) );
  OR2X2 OR2X2_3136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5745), .B(REGFILE_SIM_reg_bank__abc_33898_n5742), .Y(REGFILE_SIM_reg_bank__abc_33898_n5746) );
  OR2X2 OR2X2_3137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5739), .B(REGFILE_SIM_reg_bank__abc_33898_n5746), .Y(REGFILE_SIM_reg_bank__abc_33898_n5747) );
  OR2X2 OR2X2_3138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5732), .B(REGFILE_SIM_reg_bank__abc_33898_n5747), .Y(REGFILE_SIM_reg_bank__abc_33898_n5748) );
  OR2X2 OR2X2_3139 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5749), .B(REGFILE_SIM_reg_bank__abc_33898_n5750), .Y(REGFILE_SIM_reg_bank__abc_33898_n5751) );
  OR2X2 OR2X2_314 ( .A(alu_op_r_3_), .B(pc_q_5_), .Y(_abc_43815_n1581) );
  OR2X2 OR2X2_3140 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5752), .B(REGFILE_SIM_reg_bank__abc_33898_n5753), .Y(REGFILE_SIM_reg_bank__abc_33898_n5754) );
  OR2X2 OR2X2_3141 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5751), .B(REGFILE_SIM_reg_bank__abc_33898_n5754), .Y(REGFILE_SIM_reg_bank__abc_33898_n5755) );
  OR2X2 OR2X2_3142 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5757), .B(REGFILE_SIM_reg_bank__abc_33898_n5758), .Y(REGFILE_SIM_reg_bank__abc_33898_n5759) );
  OR2X2 OR2X2_3143 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5759), .B(REGFILE_SIM_reg_bank__abc_33898_n5756), .Y(REGFILE_SIM_reg_bank__abc_33898_n5760) );
  OR2X2 OR2X2_3144 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5755), .B(REGFILE_SIM_reg_bank__abc_33898_n5760), .Y(REGFILE_SIM_reg_bank__abc_33898_n5761) );
  OR2X2 OR2X2_3145 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5762), .B(REGFILE_SIM_reg_bank__abc_33898_n5763), .Y(REGFILE_SIM_reg_bank__abc_33898_n5764) );
  OR2X2 OR2X2_3146 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5765), .B(REGFILE_SIM_reg_bank__abc_33898_n5766), .Y(REGFILE_SIM_reg_bank__abc_33898_n5767) );
  OR2X2 OR2X2_3147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5767), .B(REGFILE_SIM_reg_bank__abc_33898_n5764), .Y(REGFILE_SIM_reg_bank__abc_33898_n5768) );
  OR2X2 OR2X2_3148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5769), .B(REGFILE_SIM_reg_bank__abc_33898_n5770), .Y(REGFILE_SIM_reg_bank__abc_33898_n5771) );
  OR2X2 OR2X2_3149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5772), .B(REGFILE_SIM_reg_bank__abc_33898_n5773), .Y(REGFILE_SIM_reg_bank__abc_33898_n5774) );
  OR2X2 OR2X2_315 ( .A(_abc_43815_n1584), .B(_abc_43815_n1547_1), .Y(_abc_43815_n1588) );
  OR2X2 OR2X2_3150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5771), .B(REGFILE_SIM_reg_bank__abc_33898_n5774), .Y(REGFILE_SIM_reg_bank__abc_33898_n5775) );
  OR2X2 OR2X2_3151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5768), .B(REGFILE_SIM_reg_bank__abc_33898_n5775), .Y(REGFILE_SIM_reg_bank__abc_33898_n5776) );
  OR2X2 OR2X2_3152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5776), .B(REGFILE_SIM_reg_bank__abc_33898_n5761), .Y(REGFILE_SIM_reg_bank__abc_33898_n5777) );
  OR2X2 OR2X2_3153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5748), .B(REGFILE_SIM_reg_bank__abc_33898_n5777), .Y(REGFILE_SIM_reg_bank_reg_rb_o_2_) );
  OR2X2 OR2X2_3154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5779), .B(REGFILE_SIM_reg_bank__abc_33898_n5780), .Y(REGFILE_SIM_reg_bank__abc_33898_n5781) );
  OR2X2 OR2X2_3155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5782), .B(REGFILE_SIM_reg_bank__abc_33898_n5783), .Y(REGFILE_SIM_reg_bank__abc_33898_n5784) );
  OR2X2 OR2X2_3156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5784), .B(REGFILE_SIM_reg_bank__abc_33898_n5781), .Y(REGFILE_SIM_reg_bank__abc_33898_n5785) );
  OR2X2 OR2X2_3157 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5786), .B(REGFILE_SIM_reg_bank__abc_33898_n5787), .Y(REGFILE_SIM_reg_bank__abc_33898_n5788) );
  OR2X2 OR2X2_3158 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5789), .B(REGFILE_SIM_reg_bank__abc_33898_n5790), .Y(REGFILE_SIM_reg_bank__abc_33898_n5791) );
  OR2X2 OR2X2_3159 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5788), .B(REGFILE_SIM_reg_bank__abc_33898_n5791), .Y(REGFILE_SIM_reg_bank__abc_33898_n5792) );
  OR2X2 OR2X2_316 ( .A(_abc_43815_n1551), .B(_abc_43815_n1588), .Y(_abc_43815_n1589) );
  OR2X2 OR2X2_3160 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5785), .B(REGFILE_SIM_reg_bank__abc_33898_n5792), .Y(REGFILE_SIM_reg_bank__abc_33898_n5793) );
  OR2X2 OR2X2_3161 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5794), .B(REGFILE_SIM_reg_bank__abc_33898_n5795), .Y(REGFILE_SIM_reg_bank__abc_33898_n5796) );
  OR2X2 OR2X2_3162 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5797), .B(REGFILE_SIM_reg_bank__abc_33898_n5798), .Y(REGFILE_SIM_reg_bank__abc_33898_n5799) );
  OR2X2 OR2X2_3163 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5796), .B(REGFILE_SIM_reg_bank__abc_33898_n5799), .Y(REGFILE_SIM_reg_bank__abc_33898_n5800) );
  OR2X2 OR2X2_3164 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5801), .B(REGFILE_SIM_reg_bank__abc_33898_n5802), .Y(REGFILE_SIM_reg_bank__abc_33898_n5803) );
  OR2X2 OR2X2_3165 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5804), .B(REGFILE_SIM_reg_bank__abc_33898_n5805), .Y(REGFILE_SIM_reg_bank__abc_33898_n5806) );
  OR2X2 OR2X2_3166 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5806), .B(REGFILE_SIM_reg_bank__abc_33898_n5803), .Y(REGFILE_SIM_reg_bank__abc_33898_n5807) );
  OR2X2 OR2X2_3167 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5800), .B(REGFILE_SIM_reg_bank__abc_33898_n5807), .Y(REGFILE_SIM_reg_bank__abc_33898_n5808) );
  OR2X2 OR2X2_3168 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5793), .B(REGFILE_SIM_reg_bank__abc_33898_n5808), .Y(REGFILE_SIM_reg_bank__abc_33898_n5809) );
  OR2X2 OR2X2_3169 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5810), .B(REGFILE_SIM_reg_bank__abc_33898_n5811), .Y(REGFILE_SIM_reg_bank__abc_33898_n5812) );
  OR2X2 OR2X2_317 ( .A(_abc_43815_n1428_bF_buf3), .B(_abc_43815_n1594), .Y(_abc_43815_n1595) );
  OR2X2 OR2X2_3170 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5813), .B(REGFILE_SIM_reg_bank__abc_33898_n5814), .Y(REGFILE_SIM_reg_bank__abc_33898_n5815) );
  OR2X2 OR2X2_3171 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5812), .B(REGFILE_SIM_reg_bank__abc_33898_n5815), .Y(REGFILE_SIM_reg_bank__abc_33898_n5816) );
  OR2X2 OR2X2_3172 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5818), .B(REGFILE_SIM_reg_bank__abc_33898_n5819), .Y(REGFILE_SIM_reg_bank__abc_33898_n5820) );
  OR2X2 OR2X2_3173 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5820), .B(REGFILE_SIM_reg_bank__abc_33898_n5817), .Y(REGFILE_SIM_reg_bank__abc_33898_n5821) );
  OR2X2 OR2X2_3174 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5816), .B(REGFILE_SIM_reg_bank__abc_33898_n5821), .Y(REGFILE_SIM_reg_bank__abc_33898_n5822) );
  OR2X2 OR2X2_3175 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5823), .B(REGFILE_SIM_reg_bank__abc_33898_n5824), .Y(REGFILE_SIM_reg_bank__abc_33898_n5825) );
  OR2X2 OR2X2_3176 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5826), .B(REGFILE_SIM_reg_bank__abc_33898_n5827), .Y(REGFILE_SIM_reg_bank__abc_33898_n5828) );
  OR2X2 OR2X2_3177 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5828), .B(REGFILE_SIM_reg_bank__abc_33898_n5825), .Y(REGFILE_SIM_reg_bank__abc_33898_n5829) );
  OR2X2 OR2X2_3178 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5830), .B(REGFILE_SIM_reg_bank__abc_33898_n5831), .Y(REGFILE_SIM_reg_bank__abc_33898_n5832) );
  OR2X2 OR2X2_3179 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5833), .B(REGFILE_SIM_reg_bank__abc_33898_n5834), .Y(REGFILE_SIM_reg_bank__abc_33898_n5835) );
  OR2X2 OR2X2_318 ( .A(_abc_43815_n1593), .B(_abc_43815_n1595), .Y(_abc_43815_n1596) );
  OR2X2 OR2X2_3180 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5832), .B(REGFILE_SIM_reg_bank__abc_33898_n5835), .Y(REGFILE_SIM_reg_bank__abc_33898_n5836) );
  OR2X2 OR2X2_3181 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5829), .B(REGFILE_SIM_reg_bank__abc_33898_n5836), .Y(REGFILE_SIM_reg_bank__abc_33898_n5837) );
  OR2X2 OR2X2_3182 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5837), .B(REGFILE_SIM_reg_bank__abc_33898_n5822), .Y(REGFILE_SIM_reg_bank__abc_33898_n5838) );
  OR2X2 OR2X2_3183 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5809), .B(REGFILE_SIM_reg_bank__abc_33898_n5838), .Y(REGFILE_SIM_reg_bank_reg_rb_o_3_) );
  OR2X2 OR2X2_3184 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5840), .B(REGFILE_SIM_reg_bank__abc_33898_n5841), .Y(REGFILE_SIM_reg_bank__abc_33898_n5842) );
  OR2X2 OR2X2_3185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5843), .B(REGFILE_SIM_reg_bank__abc_33898_n5844), .Y(REGFILE_SIM_reg_bank__abc_33898_n5845) );
  OR2X2 OR2X2_3186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5845), .B(REGFILE_SIM_reg_bank__abc_33898_n5842), .Y(REGFILE_SIM_reg_bank__abc_33898_n5846) );
  OR2X2 OR2X2_3187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5847), .B(REGFILE_SIM_reg_bank__abc_33898_n5848), .Y(REGFILE_SIM_reg_bank__abc_33898_n5849) );
  OR2X2 OR2X2_3188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5850), .B(REGFILE_SIM_reg_bank__abc_33898_n5851), .Y(REGFILE_SIM_reg_bank__abc_33898_n5852) );
  OR2X2 OR2X2_3189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5849), .B(REGFILE_SIM_reg_bank__abc_33898_n5852), .Y(REGFILE_SIM_reg_bank__abc_33898_n5853) );
  OR2X2 OR2X2_319 ( .A(_abc_43815_n1431_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_43815_n1597) );
  OR2X2 OR2X2_3190 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5846), .B(REGFILE_SIM_reg_bank__abc_33898_n5853), .Y(REGFILE_SIM_reg_bank__abc_33898_n5854) );
  OR2X2 OR2X2_3191 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5855), .B(REGFILE_SIM_reg_bank__abc_33898_n5856), .Y(REGFILE_SIM_reg_bank__abc_33898_n5857) );
  OR2X2 OR2X2_3192 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5858), .B(REGFILE_SIM_reg_bank__abc_33898_n5859), .Y(REGFILE_SIM_reg_bank__abc_33898_n5860) );
  OR2X2 OR2X2_3193 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5857), .B(REGFILE_SIM_reg_bank__abc_33898_n5860), .Y(REGFILE_SIM_reg_bank__abc_33898_n5861) );
  OR2X2 OR2X2_3194 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5862), .B(REGFILE_SIM_reg_bank__abc_33898_n5863), .Y(REGFILE_SIM_reg_bank__abc_33898_n5864) );
  OR2X2 OR2X2_3195 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5865), .B(REGFILE_SIM_reg_bank__abc_33898_n5866), .Y(REGFILE_SIM_reg_bank__abc_33898_n5867) );
  OR2X2 OR2X2_3196 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5867), .B(REGFILE_SIM_reg_bank__abc_33898_n5864), .Y(REGFILE_SIM_reg_bank__abc_33898_n5868) );
  OR2X2 OR2X2_3197 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5861), .B(REGFILE_SIM_reg_bank__abc_33898_n5868), .Y(REGFILE_SIM_reg_bank__abc_33898_n5869) );
  OR2X2 OR2X2_3198 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5854), .B(REGFILE_SIM_reg_bank__abc_33898_n5869), .Y(REGFILE_SIM_reg_bank__abc_33898_n5870) );
  OR2X2 OR2X2_3199 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5871), .B(REGFILE_SIM_reg_bank__abc_33898_n5872), .Y(REGFILE_SIM_reg_bank__abc_33898_n5873) );
  OR2X2 OR2X2_32 ( .A(_abc_43815_n751), .B(_abc_43815_n752), .Y(_abc_43815_n753_1) );
  OR2X2 OR2X2_320 ( .A(_abc_43815_n1473_bF_buf1), .B(_abc_43815_n1598), .Y(_abc_43815_n1599) );
  OR2X2 OR2X2_3200 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5874), .B(REGFILE_SIM_reg_bank__abc_33898_n5875), .Y(REGFILE_SIM_reg_bank__abc_33898_n5876) );
  OR2X2 OR2X2_3201 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5873), .B(REGFILE_SIM_reg_bank__abc_33898_n5876), .Y(REGFILE_SIM_reg_bank__abc_33898_n5877) );
  OR2X2 OR2X2_3202 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5879), .B(REGFILE_SIM_reg_bank__abc_33898_n5880), .Y(REGFILE_SIM_reg_bank__abc_33898_n5881) );
  OR2X2 OR2X2_3203 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5881), .B(REGFILE_SIM_reg_bank__abc_33898_n5878), .Y(REGFILE_SIM_reg_bank__abc_33898_n5882) );
  OR2X2 OR2X2_3204 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5877), .B(REGFILE_SIM_reg_bank__abc_33898_n5882), .Y(REGFILE_SIM_reg_bank__abc_33898_n5883) );
  OR2X2 OR2X2_3205 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5884), .B(REGFILE_SIM_reg_bank__abc_33898_n5885), .Y(REGFILE_SIM_reg_bank__abc_33898_n5886) );
  OR2X2 OR2X2_3206 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5887), .B(REGFILE_SIM_reg_bank__abc_33898_n5888), .Y(REGFILE_SIM_reg_bank__abc_33898_n5889) );
  OR2X2 OR2X2_3207 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5889), .B(REGFILE_SIM_reg_bank__abc_33898_n5886), .Y(REGFILE_SIM_reg_bank__abc_33898_n5890) );
  OR2X2 OR2X2_3208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5891), .B(REGFILE_SIM_reg_bank__abc_33898_n5892), .Y(REGFILE_SIM_reg_bank__abc_33898_n5893) );
  OR2X2 OR2X2_3209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5894), .B(REGFILE_SIM_reg_bank__abc_33898_n5895), .Y(REGFILE_SIM_reg_bank__abc_33898_n5896) );
  OR2X2 OR2X2_321 ( .A(_abc_43815_n1561), .B(pc_q_5_), .Y(_abc_43815_n1600) );
  OR2X2 OR2X2_3210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5893), .B(REGFILE_SIM_reg_bank__abc_33898_n5896), .Y(REGFILE_SIM_reg_bank__abc_33898_n5897) );
  OR2X2 OR2X2_3211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5890), .B(REGFILE_SIM_reg_bank__abc_33898_n5897), .Y(REGFILE_SIM_reg_bank__abc_33898_n5898) );
  OR2X2 OR2X2_3212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5898), .B(REGFILE_SIM_reg_bank__abc_33898_n5883), .Y(REGFILE_SIM_reg_bank__abc_33898_n5899) );
  OR2X2 OR2X2_3213 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5870), .B(REGFILE_SIM_reg_bank__abc_33898_n5899), .Y(REGFILE_SIM_reg_bank_reg_rb_o_4_) );
  OR2X2 OR2X2_3214 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5901), .B(REGFILE_SIM_reg_bank__abc_33898_n5902), .Y(REGFILE_SIM_reg_bank__abc_33898_n5903) );
  OR2X2 OR2X2_3215 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5904), .B(REGFILE_SIM_reg_bank__abc_33898_n5905), .Y(REGFILE_SIM_reg_bank__abc_33898_n5906) );
  OR2X2 OR2X2_3216 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5906), .B(REGFILE_SIM_reg_bank__abc_33898_n5903), .Y(REGFILE_SIM_reg_bank__abc_33898_n5907) );
  OR2X2 OR2X2_3217 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5908), .B(REGFILE_SIM_reg_bank__abc_33898_n5909), .Y(REGFILE_SIM_reg_bank__abc_33898_n5910) );
  OR2X2 OR2X2_3218 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5911), .B(REGFILE_SIM_reg_bank__abc_33898_n5912), .Y(REGFILE_SIM_reg_bank__abc_33898_n5913) );
  OR2X2 OR2X2_3219 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5910), .B(REGFILE_SIM_reg_bank__abc_33898_n5913), .Y(REGFILE_SIM_reg_bank__abc_33898_n5914) );
  OR2X2 OR2X2_322 ( .A(_abc_43815_n1472_1_bF_buf0), .B(_abc_43815_n1603_1), .Y(_abc_43815_n1604) );
  OR2X2 OR2X2_3220 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5907), .B(REGFILE_SIM_reg_bank__abc_33898_n5914), .Y(REGFILE_SIM_reg_bank__abc_33898_n5915) );
  OR2X2 OR2X2_3221 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5916), .B(REGFILE_SIM_reg_bank__abc_33898_n5917), .Y(REGFILE_SIM_reg_bank__abc_33898_n5918) );
  OR2X2 OR2X2_3222 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5919), .B(REGFILE_SIM_reg_bank__abc_33898_n5920), .Y(REGFILE_SIM_reg_bank__abc_33898_n5921) );
  OR2X2 OR2X2_3223 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5918), .B(REGFILE_SIM_reg_bank__abc_33898_n5921), .Y(REGFILE_SIM_reg_bank__abc_33898_n5922) );
  OR2X2 OR2X2_3224 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5923), .B(REGFILE_SIM_reg_bank__abc_33898_n5924), .Y(REGFILE_SIM_reg_bank__abc_33898_n5925) );
  OR2X2 OR2X2_3225 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5926), .B(REGFILE_SIM_reg_bank__abc_33898_n5927), .Y(REGFILE_SIM_reg_bank__abc_33898_n5928) );
  OR2X2 OR2X2_3226 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5928), .B(REGFILE_SIM_reg_bank__abc_33898_n5925), .Y(REGFILE_SIM_reg_bank__abc_33898_n5929) );
  OR2X2 OR2X2_3227 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5922), .B(REGFILE_SIM_reg_bank__abc_33898_n5929), .Y(REGFILE_SIM_reg_bank__abc_33898_n5930) );
  OR2X2 OR2X2_3228 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5915), .B(REGFILE_SIM_reg_bank__abc_33898_n5930), .Y(REGFILE_SIM_reg_bank__abc_33898_n5931) );
  OR2X2 OR2X2_3229 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5932), .B(REGFILE_SIM_reg_bank__abc_33898_n5933), .Y(REGFILE_SIM_reg_bank__abc_33898_n5934) );
  OR2X2 OR2X2_323 ( .A(_abc_43815_n1605), .B(_abc_43815_n1350_bF_buf1), .Y(_abc_43815_n1606) );
  OR2X2 OR2X2_3230 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5935), .B(REGFILE_SIM_reg_bank__abc_33898_n5936), .Y(REGFILE_SIM_reg_bank__abc_33898_n5937) );
  OR2X2 OR2X2_3231 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5934), .B(REGFILE_SIM_reg_bank__abc_33898_n5937), .Y(REGFILE_SIM_reg_bank__abc_33898_n5938) );
  OR2X2 OR2X2_3232 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5940), .B(REGFILE_SIM_reg_bank__abc_33898_n5941), .Y(REGFILE_SIM_reg_bank__abc_33898_n5942) );
  OR2X2 OR2X2_3233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5942), .B(REGFILE_SIM_reg_bank__abc_33898_n5939), .Y(REGFILE_SIM_reg_bank__abc_33898_n5943) );
  OR2X2 OR2X2_3234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5938), .B(REGFILE_SIM_reg_bank__abc_33898_n5943), .Y(REGFILE_SIM_reg_bank__abc_33898_n5944) );
  OR2X2 OR2X2_3235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5945), .B(REGFILE_SIM_reg_bank__abc_33898_n5946), .Y(REGFILE_SIM_reg_bank__abc_33898_n5947) );
  OR2X2 OR2X2_3236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5948), .B(REGFILE_SIM_reg_bank__abc_33898_n5949), .Y(REGFILE_SIM_reg_bank__abc_33898_n5950) );
  OR2X2 OR2X2_3237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5950), .B(REGFILE_SIM_reg_bank__abc_33898_n5947), .Y(REGFILE_SIM_reg_bank__abc_33898_n5951) );
  OR2X2 OR2X2_3238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5952), .B(REGFILE_SIM_reg_bank__abc_33898_n5953), .Y(REGFILE_SIM_reg_bank__abc_33898_n5954) );
  OR2X2 OR2X2_3239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5955), .B(REGFILE_SIM_reg_bank__abc_33898_n5956), .Y(REGFILE_SIM_reg_bank__abc_33898_n5957) );
  OR2X2 OR2X2_324 ( .A(_abc_43815_n1607), .B(_abc_43815_n1461_bF_buf0), .Y(_abc_43815_n1608) );
  OR2X2 OR2X2_3240 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5954), .B(REGFILE_SIM_reg_bank__abc_33898_n5957), .Y(REGFILE_SIM_reg_bank__abc_33898_n5958) );
  OR2X2 OR2X2_3241 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5951), .B(REGFILE_SIM_reg_bank__abc_33898_n5958), .Y(REGFILE_SIM_reg_bank__abc_33898_n5959) );
  OR2X2 OR2X2_3242 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5959), .B(REGFILE_SIM_reg_bank__abc_33898_n5944), .Y(REGFILE_SIM_reg_bank__abc_33898_n5960) );
  OR2X2 OR2X2_3243 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5931), .B(REGFILE_SIM_reg_bank__abc_33898_n5960), .Y(REGFILE_SIM_reg_bank_reg_rb_o_5_) );
  OR2X2 OR2X2_3244 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5962), .B(REGFILE_SIM_reg_bank__abc_33898_n5963), .Y(REGFILE_SIM_reg_bank__abc_33898_n5964) );
  OR2X2 OR2X2_3245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5965), .B(REGFILE_SIM_reg_bank__abc_33898_n5966), .Y(REGFILE_SIM_reg_bank__abc_33898_n5967) );
  OR2X2 OR2X2_3246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5967), .B(REGFILE_SIM_reg_bank__abc_33898_n5964), .Y(REGFILE_SIM_reg_bank__abc_33898_n5968) );
  OR2X2 OR2X2_3247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5969), .B(REGFILE_SIM_reg_bank__abc_33898_n5970), .Y(REGFILE_SIM_reg_bank__abc_33898_n5971) );
  OR2X2 OR2X2_3248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5972), .B(REGFILE_SIM_reg_bank__abc_33898_n5973), .Y(REGFILE_SIM_reg_bank__abc_33898_n5974) );
  OR2X2 OR2X2_3249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5971), .B(REGFILE_SIM_reg_bank__abc_33898_n5974), .Y(REGFILE_SIM_reg_bank__abc_33898_n5975) );
  OR2X2 OR2X2_325 ( .A(_abc_43815_n1351_bF_buf1), .B(_abc_43815_n1603_1), .Y(_abc_43815_n1609) );
  OR2X2 OR2X2_3250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5968), .B(REGFILE_SIM_reg_bank__abc_33898_n5975), .Y(REGFILE_SIM_reg_bank__abc_33898_n5976) );
  OR2X2 OR2X2_3251 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5977), .B(REGFILE_SIM_reg_bank__abc_33898_n5978), .Y(REGFILE_SIM_reg_bank__abc_33898_n5979) );
  OR2X2 OR2X2_3252 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5980), .B(REGFILE_SIM_reg_bank__abc_33898_n5981), .Y(REGFILE_SIM_reg_bank__abc_33898_n5982) );
  OR2X2 OR2X2_3253 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5979), .B(REGFILE_SIM_reg_bank__abc_33898_n5982), .Y(REGFILE_SIM_reg_bank__abc_33898_n5983) );
  OR2X2 OR2X2_3254 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5984), .B(REGFILE_SIM_reg_bank__abc_33898_n5985), .Y(REGFILE_SIM_reg_bank__abc_33898_n5986) );
  OR2X2 OR2X2_3255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5987), .B(REGFILE_SIM_reg_bank__abc_33898_n5988), .Y(REGFILE_SIM_reg_bank__abc_33898_n5989) );
  OR2X2 OR2X2_3256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5989), .B(REGFILE_SIM_reg_bank__abc_33898_n5986), .Y(REGFILE_SIM_reg_bank__abc_33898_n5990) );
  OR2X2 OR2X2_3257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5983), .B(REGFILE_SIM_reg_bank__abc_33898_n5990), .Y(REGFILE_SIM_reg_bank__abc_33898_n5991) );
  OR2X2 OR2X2_3258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5976), .B(REGFILE_SIM_reg_bank__abc_33898_n5991), .Y(REGFILE_SIM_reg_bank__abc_33898_n5992) );
  OR2X2 OR2X2_3259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5993), .B(REGFILE_SIM_reg_bank__abc_33898_n5994), .Y(REGFILE_SIM_reg_bank__abc_33898_n5995) );
  OR2X2 OR2X2_326 ( .A(_abc_43815_n1610), .B(_abc_43815_n1278_bF_buf4), .Y(_abc_43815_n1611) );
  OR2X2 OR2X2_3260 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5996), .B(REGFILE_SIM_reg_bank__abc_33898_n5997), .Y(REGFILE_SIM_reg_bank__abc_33898_n5998) );
  OR2X2 OR2X2_3261 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5995), .B(REGFILE_SIM_reg_bank__abc_33898_n5998), .Y(REGFILE_SIM_reg_bank__abc_33898_n5999) );
  OR2X2 OR2X2_3262 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6001), .B(REGFILE_SIM_reg_bank__abc_33898_n6002), .Y(REGFILE_SIM_reg_bank__abc_33898_n6003) );
  OR2X2 OR2X2_3263 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6003), .B(REGFILE_SIM_reg_bank__abc_33898_n6000), .Y(REGFILE_SIM_reg_bank__abc_33898_n6004) );
  OR2X2 OR2X2_3264 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5999), .B(REGFILE_SIM_reg_bank__abc_33898_n6004), .Y(REGFILE_SIM_reg_bank__abc_33898_n6005) );
  OR2X2 OR2X2_3265 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6006), .B(REGFILE_SIM_reg_bank__abc_33898_n6007), .Y(REGFILE_SIM_reg_bank__abc_33898_n6008) );
  OR2X2 OR2X2_3266 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6009), .B(REGFILE_SIM_reg_bank__abc_33898_n6010), .Y(REGFILE_SIM_reg_bank__abc_33898_n6011) );
  OR2X2 OR2X2_3267 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6011), .B(REGFILE_SIM_reg_bank__abc_33898_n6008), .Y(REGFILE_SIM_reg_bank__abc_33898_n6012) );
  OR2X2 OR2X2_3268 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6013), .B(REGFILE_SIM_reg_bank__abc_33898_n6014), .Y(REGFILE_SIM_reg_bank__abc_33898_n6015) );
  OR2X2 OR2X2_3269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6016), .B(REGFILE_SIM_reg_bank__abc_33898_n6017), .Y(REGFILE_SIM_reg_bank__abc_33898_n6018) );
  OR2X2 OR2X2_327 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_5_), .Y(_abc_43815_n1612) );
  OR2X2 OR2X2_3270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6015), .B(REGFILE_SIM_reg_bank__abc_33898_n6018), .Y(REGFILE_SIM_reg_bank__abc_33898_n6019) );
  OR2X2 OR2X2_3271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6012), .B(REGFILE_SIM_reg_bank__abc_33898_n6019), .Y(REGFILE_SIM_reg_bank__abc_33898_n6020) );
  OR2X2 OR2X2_3272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6020), .B(REGFILE_SIM_reg_bank__abc_33898_n6005), .Y(REGFILE_SIM_reg_bank__abc_33898_n6021) );
  OR2X2 OR2X2_3273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n5992), .B(REGFILE_SIM_reg_bank__abc_33898_n6021), .Y(REGFILE_SIM_reg_bank_reg_rb_o_6_) );
  OR2X2 OR2X2_3274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6023), .B(REGFILE_SIM_reg_bank__abc_33898_n6024), .Y(REGFILE_SIM_reg_bank__abc_33898_n6025) );
  OR2X2 OR2X2_3275 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6026), .B(REGFILE_SIM_reg_bank__abc_33898_n6027), .Y(REGFILE_SIM_reg_bank__abc_33898_n6028) );
  OR2X2 OR2X2_3276 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6028), .B(REGFILE_SIM_reg_bank__abc_33898_n6025), .Y(REGFILE_SIM_reg_bank__abc_33898_n6029) );
  OR2X2 OR2X2_3277 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6030), .B(REGFILE_SIM_reg_bank__abc_33898_n6031), .Y(REGFILE_SIM_reg_bank__abc_33898_n6032) );
  OR2X2 OR2X2_3278 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6033), .B(REGFILE_SIM_reg_bank__abc_33898_n6034), .Y(REGFILE_SIM_reg_bank__abc_33898_n6035) );
  OR2X2 OR2X2_3279 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6032), .B(REGFILE_SIM_reg_bank__abc_33898_n6035), .Y(REGFILE_SIM_reg_bank__abc_33898_n6036) );
  OR2X2 OR2X2_328 ( .A(_abc_43815_n1585), .B(_abc_43815_n1582), .Y(_abc_43815_n1615_1) );
  OR2X2 OR2X2_3280 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6029), .B(REGFILE_SIM_reg_bank__abc_33898_n6036), .Y(REGFILE_SIM_reg_bank__abc_33898_n6037) );
  OR2X2 OR2X2_3281 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6038), .B(REGFILE_SIM_reg_bank__abc_33898_n6039), .Y(REGFILE_SIM_reg_bank__abc_33898_n6040) );
  OR2X2 OR2X2_3282 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6041), .B(REGFILE_SIM_reg_bank__abc_33898_n6042), .Y(REGFILE_SIM_reg_bank__abc_33898_n6043) );
  OR2X2 OR2X2_3283 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6040), .B(REGFILE_SIM_reg_bank__abc_33898_n6043), .Y(REGFILE_SIM_reg_bank__abc_33898_n6044) );
  OR2X2 OR2X2_3284 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6045), .B(REGFILE_SIM_reg_bank__abc_33898_n6046), .Y(REGFILE_SIM_reg_bank__abc_33898_n6047) );
  OR2X2 OR2X2_3285 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6048), .B(REGFILE_SIM_reg_bank__abc_33898_n6049), .Y(REGFILE_SIM_reg_bank__abc_33898_n6050) );
  OR2X2 OR2X2_3286 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6050), .B(REGFILE_SIM_reg_bank__abc_33898_n6047), .Y(REGFILE_SIM_reg_bank__abc_33898_n6051) );
  OR2X2 OR2X2_3287 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6044), .B(REGFILE_SIM_reg_bank__abc_33898_n6051), .Y(REGFILE_SIM_reg_bank__abc_33898_n6052) );
  OR2X2 OR2X2_3288 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6037), .B(REGFILE_SIM_reg_bank__abc_33898_n6052), .Y(REGFILE_SIM_reg_bank__abc_33898_n6053) );
  OR2X2 OR2X2_3289 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6054), .B(REGFILE_SIM_reg_bank__abc_33898_n6055), .Y(REGFILE_SIM_reg_bank__abc_33898_n6056) );
  OR2X2 OR2X2_329 ( .A(_abc_43815_n1590), .B(_abc_43815_n1615_1), .Y(_abc_43815_n1616) );
  OR2X2 OR2X2_3290 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6057), .B(REGFILE_SIM_reg_bank__abc_33898_n6058), .Y(REGFILE_SIM_reg_bank__abc_33898_n6059) );
  OR2X2 OR2X2_3291 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6056), .B(REGFILE_SIM_reg_bank__abc_33898_n6059), .Y(REGFILE_SIM_reg_bank__abc_33898_n6060) );
  OR2X2 OR2X2_3292 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6062), .B(REGFILE_SIM_reg_bank__abc_33898_n6063), .Y(REGFILE_SIM_reg_bank__abc_33898_n6064) );
  OR2X2 OR2X2_3293 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6064), .B(REGFILE_SIM_reg_bank__abc_33898_n6061), .Y(REGFILE_SIM_reg_bank__abc_33898_n6065) );
  OR2X2 OR2X2_3294 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6060), .B(REGFILE_SIM_reg_bank__abc_33898_n6065), .Y(REGFILE_SIM_reg_bank__abc_33898_n6066) );
  OR2X2 OR2X2_3295 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6067), .B(REGFILE_SIM_reg_bank__abc_33898_n6068), .Y(REGFILE_SIM_reg_bank__abc_33898_n6069) );
  OR2X2 OR2X2_3296 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6070), .B(REGFILE_SIM_reg_bank__abc_33898_n6071), .Y(REGFILE_SIM_reg_bank__abc_33898_n6072) );
  OR2X2 OR2X2_3297 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6072), .B(REGFILE_SIM_reg_bank__abc_33898_n6069), .Y(REGFILE_SIM_reg_bank__abc_33898_n6073) );
  OR2X2 OR2X2_3298 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6074), .B(REGFILE_SIM_reg_bank__abc_33898_n6075), .Y(REGFILE_SIM_reg_bank__abc_33898_n6076) );
  OR2X2 OR2X2_3299 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6077), .B(REGFILE_SIM_reg_bank__abc_33898_n6078), .Y(REGFILE_SIM_reg_bank__abc_33898_n6079) );
  OR2X2 OR2X2_33 ( .A(_abc_43815_n754_1), .B(_abc_43815_n755), .Y(_abc_43815_n756) );
  OR2X2 OR2X2_330 ( .A(int32_r_4_), .B(pc_q_6_), .Y(_abc_43815_n1617) );
  OR2X2 OR2X2_3300 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6076), .B(REGFILE_SIM_reg_bank__abc_33898_n6079), .Y(REGFILE_SIM_reg_bank__abc_33898_n6080) );
  OR2X2 OR2X2_3301 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6073), .B(REGFILE_SIM_reg_bank__abc_33898_n6080), .Y(REGFILE_SIM_reg_bank__abc_33898_n6081) );
  OR2X2 OR2X2_3302 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6081), .B(REGFILE_SIM_reg_bank__abc_33898_n6066), .Y(REGFILE_SIM_reg_bank__abc_33898_n6082) );
  OR2X2 OR2X2_3303 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6053), .B(REGFILE_SIM_reg_bank__abc_33898_n6082), .Y(REGFILE_SIM_reg_bank_reg_rb_o_7_) );
  OR2X2 OR2X2_3304 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6084), .B(REGFILE_SIM_reg_bank__abc_33898_n6085), .Y(REGFILE_SIM_reg_bank__abc_33898_n6086) );
  OR2X2 OR2X2_3305 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6087), .B(REGFILE_SIM_reg_bank__abc_33898_n6088), .Y(REGFILE_SIM_reg_bank__abc_33898_n6089) );
  OR2X2 OR2X2_3306 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6089), .B(REGFILE_SIM_reg_bank__abc_33898_n6086), .Y(REGFILE_SIM_reg_bank__abc_33898_n6090) );
  OR2X2 OR2X2_3307 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6091), .B(REGFILE_SIM_reg_bank__abc_33898_n6092), .Y(REGFILE_SIM_reg_bank__abc_33898_n6093) );
  OR2X2 OR2X2_3308 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6094), .B(REGFILE_SIM_reg_bank__abc_33898_n6095), .Y(REGFILE_SIM_reg_bank__abc_33898_n6096) );
  OR2X2 OR2X2_3309 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6093), .B(REGFILE_SIM_reg_bank__abc_33898_n6096), .Y(REGFILE_SIM_reg_bank__abc_33898_n6097) );
  OR2X2 OR2X2_331 ( .A(_abc_43815_n1616), .B(_abc_43815_n1620), .Y(_abc_43815_n1621) );
  OR2X2 OR2X2_3310 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6090), .B(REGFILE_SIM_reg_bank__abc_33898_n6097), .Y(REGFILE_SIM_reg_bank__abc_33898_n6098) );
  OR2X2 OR2X2_3311 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6099), .B(REGFILE_SIM_reg_bank__abc_33898_n6100), .Y(REGFILE_SIM_reg_bank__abc_33898_n6101) );
  OR2X2 OR2X2_3312 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6102), .B(REGFILE_SIM_reg_bank__abc_33898_n6103), .Y(REGFILE_SIM_reg_bank__abc_33898_n6104) );
  OR2X2 OR2X2_3313 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6101), .B(REGFILE_SIM_reg_bank__abc_33898_n6104), .Y(REGFILE_SIM_reg_bank__abc_33898_n6105) );
  OR2X2 OR2X2_3314 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6106), .B(REGFILE_SIM_reg_bank__abc_33898_n6107), .Y(REGFILE_SIM_reg_bank__abc_33898_n6108) );
  OR2X2 OR2X2_3315 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6109), .B(REGFILE_SIM_reg_bank__abc_33898_n6110), .Y(REGFILE_SIM_reg_bank__abc_33898_n6111) );
  OR2X2 OR2X2_3316 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6111), .B(REGFILE_SIM_reg_bank__abc_33898_n6108), .Y(REGFILE_SIM_reg_bank__abc_33898_n6112) );
  OR2X2 OR2X2_3317 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6105), .B(REGFILE_SIM_reg_bank__abc_33898_n6112), .Y(REGFILE_SIM_reg_bank__abc_33898_n6113) );
  OR2X2 OR2X2_3318 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6098), .B(REGFILE_SIM_reg_bank__abc_33898_n6113), .Y(REGFILE_SIM_reg_bank__abc_33898_n6114) );
  OR2X2 OR2X2_3319 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6115), .B(REGFILE_SIM_reg_bank__abc_33898_n6116), .Y(REGFILE_SIM_reg_bank__abc_33898_n6117) );
  OR2X2 OR2X2_332 ( .A(_abc_43815_n1428_bF_buf2), .B(_abc_43815_n1626), .Y(_abc_43815_n1627) );
  OR2X2 OR2X2_3320 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6118), .B(REGFILE_SIM_reg_bank__abc_33898_n6119), .Y(REGFILE_SIM_reg_bank__abc_33898_n6120) );
  OR2X2 OR2X2_3321 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6117), .B(REGFILE_SIM_reg_bank__abc_33898_n6120), .Y(REGFILE_SIM_reg_bank__abc_33898_n6121) );
  OR2X2 OR2X2_3322 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6123), .B(REGFILE_SIM_reg_bank__abc_33898_n6124), .Y(REGFILE_SIM_reg_bank__abc_33898_n6125) );
  OR2X2 OR2X2_3323 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6125), .B(REGFILE_SIM_reg_bank__abc_33898_n6122), .Y(REGFILE_SIM_reg_bank__abc_33898_n6126) );
  OR2X2 OR2X2_3324 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6121), .B(REGFILE_SIM_reg_bank__abc_33898_n6126), .Y(REGFILE_SIM_reg_bank__abc_33898_n6127) );
  OR2X2 OR2X2_3325 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6128), .B(REGFILE_SIM_reg_bank__abc_33898_n6129), .Y(REGFILE_SIM_reg_bank__abc_33898_n6130) );
  OR2X2 OR2X2_3326 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6131), .B(REGFILE_SIM_reg_bank__abc_33898_n6132), .Y(REGFILE_SIM_reg_bank__abc_33898_n6133) );
  OR2X2 OR2X2_3327 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6133), .B(REGFILE_SIM_reg_bank__abc_33898_n6130), .Y(REGFILE_SIM_reg_bank__abc_33898_n6134) );
  OR2X2 OR2X2_3328 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6135), .B(REGFILE_SIM_reg_bank__abc_33898_n6136), .Y(REGFILE_SIM_reg_bank__abc_33898_n6137) );
  OR2X2 OR2X2_3329 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6138), .B(REGFILE_SIM_reg_bank__abc_33898_n6139), .Y(REGFILE_SIM_reg_bank__abc_33898_n6140) );
  OR2X2 OR2X2_333 ( .A(_abc_43815_n1625), .B(_abc_43815_n1627), .Y(_abc_43815_n1628) );
  OR2X2 OR2X2_3330 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6137), .B(REGFILE_SIM_reg_bank__abc_33898_n6140), .Y(REGFILE_SIM_reg_bank__abc_33898_n6141) );
  OR2X2 OR2X2_3331 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6134), .B(REGFILE_SIM_reg_bank__abc_33898_n6141), .Y(REGFILE_SIM_reg_bank__abc_33898_n6142) );
  OR2X2 OR2X2_3332 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6142), .B(REGFILE_SIM_reg_bank__abc_33898_n6127), .Y(REGFILE_SIM_reg_bank__abc_33898_n6143) );
  OR2X2 OR2X2_3333 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6114), .B(REGFILE_SIM_reg_bank__abc_33898_n6143), .Y(REGFILE_SIM_reg_bank_reg_rb_o_8_) );
  OR2X2 OR2X2_3334 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6145), .B(REGFILE_SIM_reg_bank__abc_33898_n6146), .Y(REGFILE_SIM_reg_bank__abc_33898_n6147) );
  OR2X2 OR2X2_3335 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6148), .B(REGFILE_SIM_reg_bank__abc_33898_n6149), .Y(REGFILE_SIM_reg_bank__abc_33898_n6150) );
  OR2X2 OR2X2_3336 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6150), .B(REGFILE_SIM_reg_bank__abc_33898_n6147), .Y(REGFILE_SIM_reg_bank__abc_33898_n6151) );
  OR2X2 OR2X2_3337 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6152), .B(REGFILE_SIM_reg_bank__abc_33898_n6153), .Y(REGFILE_SIM_reg_bank__abc_33898_n6154) );
  OR2X2 OR2X2_3338 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6155), .B(REGFILE_SIM_reg_bank__abc_33898_n6156), .Y(REGFILE_SIM_reg_bank__abc_33898_n6157) );
  OR2X2 OR2X2_3339 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6154), .B(REGFILE_SIM_reg_bank__abc_33898_n6157), .Y(REGFILE_SIM_reg_bank__abc_33898_n6158) );
  OR2X2 OR2X2_334 ( .A(_abc_43815_n1431_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_43815_n1629) );
  OR2X2 OR2X2_3340 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6151), .B(REGFILE_SIM_reg_bank__abc_33898_n6158), .Y(REGFILE_SIM_reg_bank__abc_33898_n6159) );
  OR2X2 OR2X2_3341 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6160), .B(REGFILE_SIM_reg_bank__abc_33898_n6161), .Y(REGFILE_SIM_reg_bank__abc_33898_n6162) );
  OR2X2 OR2X2_3342 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6163), .B(REGFILE_SIM_reg_bank__abc_33898_n6164), .Y(REGFILE_SIM_reg_bank__abc_33898_n6165) );
  OR2X2 OR2X2_3343 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6162), .B(REGFILE_SIM_reg_bank__abc_33898_n6165), .Y(REGFILE_SIM_reg_bank__abc_33898_n6166) );
  OR2X2 OR2X2_3344 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6167), .B(REGFILE_SIM_reg_bank__abc_33898_n6168), .Y(REGFILE_SIM_reg_bank__abc_33898_n6169) );
  OR2X2 OR2X2_3345 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6170), .B(REGFILE_SIM_reg_bank__abc_33898_n6171), .Y(REGFILE_SIM_reg_bank__abc_33898_n6172) );
  OR2X2 OR2X2_3346 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6172), .B(REGFILE_SIM_reg_bank__abc_33898_n6169), .Y(REGFILE_SIM_reg_bank__abc_33898_n6173) );
  OR2X2 OR2X2_3347 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6166), .B(REGFILE_SIM_reg_bank__abc_33898_n6173), .Y(REGFILE_SIM_reg_bank__abc_33898_n6174) );
  OR2X2 OR2X2_3348 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6159), .B(REGFILE_SIM_reg_bank__abc_33898_n6174), .Y(REGFILE_SIM_reg_bank__abc_33898_n6175) );
  OR2X2 OR2X2_3349 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6176), .B(REGFILE_SIM_reg_bank__abc_33898_n6177), .Y(REGFILE_SIM_reg_bank__abc_33898_n6178) );
  OR2X2 OR2X2_335 ( .A(_abc_43815_n1630), .B(_abc_43815_n1473_bF_buf0), .Y(_abc_43815_n1631) );
  OR2X2 OR2X2_3350 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6179), .B(REGFILE_SIM_reg_bank__abc_33898_n6180), .Y(REGFILE_SIM_reg_bank__abc_33898_n6181) );
  OR2X2 OR2X2_3351 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6178), .B(REGFILE_SIM_reg_bank__abc_33898_n6181), .Y(REGFILE_SIM_reg_bank__abc_33898_n6182) );
  OR2X2 OR2X2_3352 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6184), .B(REGFILE_SIM_reg_bank__abc_33898_n6185), .Y(REGFILE_SIM_reg_bank__abc_33898_n6186) );
  OR2X2 OR2X2_3353 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6186), .B(REGFILE_SIM_reg_bank__abc_33898_n6183), .Y(REGFILE_SIM_reg_bank__abc_33898_n6187) );
  OR2X2 OR2X2_3354 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6182), .B(REGFILE_SIM_reg_bank__abc_33898_n6187), .Y(REGFILE_SIM_reg_bank__abc_33898_n6188) );
  OR2X2 OR2X2_3355 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6189), .B(REGFILE_SIM_reg_bank__abc_33898_n6190), .Y(REGFILE_SIM_reg_bank__abc_33898_n6191) );
  OR2X2 OR2X2_3356 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6192), .B(REGFILE_SIM_reg_bank__abc_33898_n6193), .Y(REGFILE_SIM_reg_bank__abc_33898_n6194) );
  OR2X2 OR2X2_3357 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6194), .B(REGFILE_SIM_reg_bank__abc_33898_n6191), .Y(REGFILE_SIM_reg_bank__abc_33898_n6195) );
  OR2X2 OR2X2_3358 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6196), .B(REGFILE_SIM_reg_bank__abc_33898_n6197), .Y(REGFILE_SIM_reg_bank__abc_33898_n6198) );
  OR2X2 OR2X2_3359 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6199), .B(REGFILE_SIM_reg_bank__abc_33898_n6200), .Y(REGFILE_SIM_reg_bank__abc_33898_n6201) );
  OR2X2 OR2X2_336 ( .A(_abc_43815_n1601), .B(pc_q_6_), .Y(_abc_43815_n1632) );
  OR2X2 OR2X2_3360 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6198), .B(REGFILE_SIM_reg_bank__abc_33898_n6201), .Y(REGFILE_SIM_reg_bank__abc_33898_n6202) );
  OR2X2 OR2X2_3361 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6195), .B(REGFILE_SIM_reg_bank__abc_33898_n6202), .Y(REGFILE_SIM_reg_bank__abc_33898_n6203) );
  OR2X2 OR2X2_3362 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6203), .B(REGFILE_SIM_reg_bank__abc_33898_n6188), .Y(REGFILE_SIM_reg_bank__abc_33898_n6204) );
  OR2X2 OR2X2_3363 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6175), .B(REGFILE_SIM_reg_bank__abc_33898_n6204), .Y(REGFILE_SIM_reg_bank_reg_rb_o_9_) );
  OR2X2 OR2X2_3364 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6206), .B(REGFILE_SIM_reg_bank__abc_33898_n6207), .Y(REGFILE_SIM_reg_bank__abc_33898_n6208) );
  OR2X2 OR2X2_3365 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6209), .B(REGFILE_SIM_reg_bank__abc_33898_n6210), .Y(REGFILE_SIM_reg_bank__abc_33898_n6211) );
  OR2X2 OR2X2_3366 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6211), .B(REGFILE_SIM_reg_bank__abc_33898_n6208), .Y(REGFILE_SIM_reg_bank__abc_33898_n6212) );
  OR2X2 OR2X2_3367 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6213), .B(REGFILE_SIM_reg_bank__abc_33898_n6214), .Y(REGFILE_SIM_reg_bank__abc_33898_n6215) );
  OR2X2 OR2X2_3368 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6216), .B(REGFILE_SIM_reg_bank__abc_33898_n6217), .Y(REGFILE_SIM_reg_bank__abc_33898_n6218) );
  OR2X2 OR2X2_3369 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6215), .B(REGFILE_SIM_reg_bank__abc_33898_n6218), .Y(REGFILE_SIM_reg_bank__abc_33898_n6219) );
  OR2X2 OR2X2_337 ( .A(_abc_43815_n1472_1_bF_buf4), .B(_abc_43815_n1635_1), .Y(_abc_43815_n1636) );
  OR2X2 OR2X2_3370 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6212), .B(REGFILE_SIM_reg_bank__abc_33898_n6219), .Y(REGFILE_SIM_reg_bank__abc_33898_n6220) );
  OR2X2 OR2X2_3371 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6221), .B(REGFILE_SIM_reg_bank__abc_33898_n6222), .Y(REGFILE_SIM_reg_bank__abc_33898_n6223) );
  OR2X2 OR2X2_3372 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6224), .B(REGFILE_SIM_reg_bank__abc_33898_n6225), .Y(REGFILE_SIM_reg_bank__abc_33898_n6226) );
  OR2X2 OR2X2_3373 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6223), .B(REGFILE_SIM_reg_bank__abc_33898_n6226), .Y(REGFILE_SIM_reg_bank__abc_33898_n6227) );
  OR2X2 OR2X2_3374 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6228), .B(REGFILE_SIM_reg_bank__abc_33898_n6229), .Y(REGFILE_SIM_reg_bank__abc_33898_n6230) );
  OR2X2 OR2X2_3375 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6231), .B(REGFILE_SIM_reg_bank__abc_33898_n6232), .Y(REGFILE_SIM_reg_bank__abc_33898_n6233) );
  OR2X2 OR2X2_3376 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6233), .B(REGFILE_SIM_reg_bank__abc_33898_n6230), .Y(REGFILE_SIM_reg_bank__abc_33898_n6234) );
  OR2X2 OR2X2_3377 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6227), .B(REGFILE_SIM_reg_bank__abc_33898_n6234), .Y(REGFILE_SIM_reg_bank__abc_33898_n6235) );
  OR2X2 OR2X2_3378 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6220), .B(REGFILE_SIM_reg_bank__abc_33898_n6235), .Y(REGFILE_SIM_reg_bank__abc_33898_n6236) );
  OR2X2 OR2X2_3379 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6237), .B(REGFILE_SIM_reg_bank__abc_33898_n6238), .Y(REGFILE_SIM_reg_bank__abc_33898_n6239) );
  OR2X2 OR2X2_338 ( .A(_abc_43815_n1637), .B(_abc_43815_n1350_bF_buf0), .Y(_abc_43815_n1638) );
  OR2X2 OR2X2_3380 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6240), .B(REGFILE_SIM_reg_bank__abc_33898_n6241), .Y(REGFILE_SIM_reg_bank__abc_33898_n6242) );
  OR2X2 OR2X2_3381 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6239), .B(REGFILE_SIM_reg_bank__abc_33898_n6242), .Y(REGFILE_SIM_reg_bank__abc_33898_n6243) );
  OR2X2 OR2X2_3382 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6245), .B(REGFILE_SIM_reg_bank__abc_33898_n6246), .Y(REGFILE_SIM_reg_bank__abc_33898_n6247) );
  OR2X2 OR2X2_3383 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6247), .B(REGFILE_SIM_reg_bank__abc_33898_n6244), .Y(REGFILE_SIM_reg_bank__abc_33898_n6248) );
  OR2X2 OR2X2_3384 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6243), .B(REGFILE_SIM_reg_bank__abc_33898_n6248), .Y(REGFILE_SIM_reg_bank__abc_33898_n6249) );
  OR2X2 OR2X2_3385 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6250), .B(REGFILE_SIM_reg_bank__abc_33898_n6251), .Y(REGFILE_SIM_reg_bank__abc_33898_n6252) );
  OR2X2 OR2X2_3386 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6253), .B(REGFILE_SIM_reg_bank__abc_33898_n6254), .Y(REGFILE_SIM_reg_bank__abc_33898_n6255) );
  OR2X2 OR2X2_3387 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6255), .B(REGFILE_SIM_reg_bank__abc_33898_n6252), .Y(REGFILE_SIM_reg_bank__abc_33898_n6256) );
  OR2X2 OR2X2_3388 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6257), .B(REGFILE_SIM_reg_bank__abc_33898_n6258), .Y(REGFILE_SIM_reg_bank__abc_33898_n6259) );
  OR2X2 OR2X2_3389 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6260), .B(REGFILE_SIM_reg_bank__abc_33898_n6261), .Y(REGFILE_SIM_reg_bank__abc_33898_n6262) );
  OR2X2 OR2X2_339 ( .A(_abc_43815_n1640), .B(_abc_43815_n1639), .Y(_abc_43815_n1641) );
  OR2X2 OR2X2_3390 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6259), .B(REGFILE_SIM_reg_bank__abc_33898_n6262), .Y(REGFILE_SIM_reg_bank__abc_33898_n6263) );
  OR2X2 OR2X2_3391 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6256), .B(REGFILE_SIM_reg_bank__abc_33898_n6263), .Y(REGFILE_SIM_reg_bank__abc_33898_n6264) );
  OR2X2 OR2X2_3392 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6264), .B(REGFILE_SIM_reg_bank__abc_33898_n6249), .Y(REGFILE_SIM_reg_bank__abc_33898_n6265) );
  OR2X2 OR2X2_3393 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6236), .B(REGFILE_SIM_reg_bank__abc_33898_n6265), .Y(REGFILE_SIM_reg_bank_reg_rb_o_10_) );
  OR2X2 OR2X2_3394 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6267), .B(REGFILE_SIM_reg_bank__abc_33898_n6268), .Y(REGFILE_SIM_reg_bank__abc_33898_n6269) );
  OR2X2 OR2X2_3395 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6270), .B(REGFILE_SIM_reg_bank__abc_33898_n6271), .Y(REGFILE_SIM_reg_bank__abc_33898_n6272) );
  OR2X2 OR2X2_3396 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6272), .B(REGFILE_SIM_reg_bank__abc_33898_n6269), .Y(REGFILE_SIM_reg_bank__abc_33898_n6273) );
  OR2X2 OR2X2_3397 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6274), .B(REGFILE_SIM_reg_bank__abc_33898_n6275), .Y(REGFILE_SIM_reg_bank__abc_33898_n6276) );
  OR2X2 OR2X2_3398 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6277), .B(REGFILE_SIM_reg_bank__abc_33898_n6278), .Y(REGFILE_SIM_reg_bank__abc_33898_n6279) );
  OR2X2 OR2X2_3399 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6276), .B(REGFILE_SIM_reg_bank__abc_33898_n6279), .Y(REGFILE_SIM_reg_bank__abc_33898_n6280) );
  OR2X2 OR2X2_34 ( .A(_abc_43815_n753_1), .B(_abc_43815_n756), .Y(_abc_43815_n757) );
  OR2X2 OR2X2_340 ( .A(_abc_43815_n1413_bF_buf3), .B(_abc_43815_n1641), .Y(_abc_43815_n1642) );
  OR2X2 OR2X2_3400 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6273), .B(REGFILE_SIM_reg_bank__abc_33898_n6280), .Y(REGFILE_SIM_reg_bank__abc_33898_n6281) );
  OR2X2 OR2X2_3401 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6282), .B(REGFILE_SIM_reg_bank__abc_33898_n6283), .Y(REGFILE_SIM_reg_bank__abc_33898_n6284) );
  OR2X2 OR2X2_3402 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6285), .B(REGFILE_SIM_reg_bank__abc_33898_n6286), .Y(REGFILE_SIM_reg_bank__abc_33898_n6287) );
  OR2X2 OR2X2_3403 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6284), .B(REGFILE_SIM_reg_bank__abc_33898_n6287), .Y(REGFILE_SIM_reg_bank__abc_33898_n6288) );
  OR2X2 OR2X2_3404 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6289), .B(REGFILE_SIM_reg_bank__abc_33898_n6290), .Y(REGFILE_SIM_reg_bank__abc_33898_n6291) );
  OR2X2 OR2X2_3405 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6292), .B(REGFILE_SIM_reg_bank__abc_33898_n6293), .Y(REGFILE_SIM_reg_bank__abc_33898_n6294) );
  OR2X2 OR2X2_3406 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6294), .B(REGFILE_SIM_reg_bank__abc_33898_n6291), .Y(REGFILE_SIM_reg_bank__abc_33898_n6295) );
  OR2X2 OR2X2_3407 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6288), .B(REGFILE_SIM_reg_bank__abc_33898_n6295), .Y(REGFILE_SIM_reg_bank__abc_33898_n6296) );
  OR2X2 OR2X2_3408 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6281), .B(REGFILE_SIM_reg_bank__abc_33898_n6296), .Y(REGFILE_SIM_reg_bank__abc_33898_n6297) );
  OR2X2 OR2X2_3409 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6298), .B(REGFILE_SIM_reg_bank__abc_33898_n6299), .Y(REGFILE_SIM_reg_bank__abc_33898_n6300) );
  OR2X2 OR2X2_341 ( .A(_abc_43815_n1643), .B(_abc_43815_n1461_bF_buf3), .Y(_abc_43815_n1644) );
  OR2X2 OR2X2_3410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6301), .B(REGFILE_SIM_reg_bank__abc_33898_n6302), .Y(REGFILE_SIM_reg_bank__abc_33898_n6303) );
  OR2X2 OR2X2_3411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6300), .B(REGFILE_SIM_reg_bank__abc_33898_n6303), .Y(REGFILE_SIM_reg_bank__abc_33898_n6304) );
  OR2X2 OR2X2_3412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6306), .B(REGFILE_SIM_reg_bank__abc_33898_n6307), .Y(REGFILE_SIM_reg_bank__abc_33898_n6308) );
  OR2X2 OR2X2_3413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6308), .B(REGFILE_SIM_reg_bank__abc_33898_n6305), .Y(REGFILE_SIM_reg_bank__abc_33898_n6309) );
  OR2X2 OR2X2_3414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6304), .B(REGFILE_SIM_reg_bank__abc_33898_n6309), .Y(REGFILE_SIM_reg_bank__abc_33898_n6310) );
  OR2X2 OR2X2_3415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6311), .B(REGFILE_SIM_reg_bank__abc_33898_n6312), .Y(REGFILE_SIM_reg_bank__abc_33898_n6313) );
  OR2X2 OR2X2_3416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6314), .B(REGFILE_SIM_reg_bank__abc_33898_n6315), .Y(REGFILE_SIM_reg_bank__abc_33898_n6316) );
  OR2X2 OR2X2_3417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6316), .B(REGFILE_SIM_reg_bank__abc_33898_n6313), .Y(REGFILE_SIM_reg_bank__abc_33898_n6317) );
  OR2X2 OR2X2_3418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6318), .B(REGFILE_SIM_reg_bank__abc_33898_n6319), .Y(REGFILE_SIM_reg_bank__abc_33898_n6320) );
  OR2X2 OR2X2_3419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6321), .B(REGFILE_SIM_reg_bank__abc_33898_n6322), .Y(REGFILE_SIM_reg_bank__abc_33898_n6323) );
  OR2X2 OR2X2_342 ( .A(_abc_43815_n1351_bF_buf0), .B(_abc_43815_n1635_1), .Y(_abc_43815_n1645) );
  OR2X2 OR2X2_3420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6320), .B(REGFILE_SIM_reg_bank__abc_33898_n6323), .Y(REGFILE_SIM_reg_bank__abc_33898_n6324) );
  OR2X2 OR2X2_3421 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6317), .B(REGFILE_SIM_reg_bank__abc_33898_n6324), .Y(REGFILE_SIM_reg_bank__abc_33898_n6325) );
  OR2X2 OR2X2_3422 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6325), .B(REGFILE_SIM_reg_bank__abc_33898_n6310), .Y(REGFILE_SIM_reg_bank__abc_33898_n6326) );
  OR2X2 OR2X2_3423 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6297), .B(REGFILE_SIM_reg_bank__abc_33898_n6326), .Y(REGFILE_SIM_reg_bank_reg_rb_o_11_) );
  OR2X2 OR2X2_3424 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6328), .B(REGFILE_SIM_reg_bank__abc_33898_n6329), .Y(REGFILE_SIM_reg_bank__abc_33898_n6330) );
  OR2X2 OR2X2_3425 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6331), .B(REGFILE_SIM_reg_bank__abc_33898_n6332), .Y(REGFILE_SIM_reg_bank__abc_33898_n6333) );
  OR2X2 OR2X2_3426 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6333), .B(REGFILE_SIM_reg_bank__abc_33898_n6330), .Y(REGFILE_SIM_reg_bank__abc_33898_n6334) );
  OR2X2 OR2X2_3427 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6335), .B(REGFILE_SIM_reg_bank__abc_33898_n6336), .Y(REGFILE_SIM_reg_bank__abc_33898_n6337) );
  OR2X2 OR2X2_3428 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6338), .B(REGFILE_SIM_reg_bank__abc_33898_n6339), .Y(REGFILE_SIM_reg_bank__abc_33898_n6340) );
  OR2X2 OR2X2_3429 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6337), .B(REGFILE_SIM_reg_bank__abc_33898_n6340), .Y(REGFILE_SIM_reg_bank__abc_33898_n6341) );
  OR2X2 OR2X2_343 ( .A(_abc_43815_n1646), .B(_abc_43815_n1278_bF_buf3), .Y(_abc_43815_n1647) );
  OR2X2 OR2X2_3430 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6334), .B(REGFILE_SIM_reg_bank__abc_33898_n6341), .Y(REGFILE_SIM_reg_bank__abc_33898_n6342) );
  OR2X2 OR2X2_3431 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6343), .B(REGFILE_SIM_reg_bank__abc_33898_n6344), .Y(REGFILE_SIM_reg_bank__abc_33898_n6345) );
  OR2X2 OR2X2_3432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6346), .B(REGFILE_SIM_reg_bank__abc_33898_n6347), .Y(REGFILE_SIM_reg_bank__abc_33898_n6348) );
  OR2X2 OR2X2_3433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6345), .B(REGFILE_SIM_reg_bank__abc_33898_n6348), .Y(REGFILE_SIM_reg_bank__abc_33898_n6349) );
  OR2X2 OR2X2_3434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6350), .B(REGFILE_SIM_reg_bank__abc_33898_n6351), .Y(REGFILE_SIM_reg_bank__abc_33898_n6352) );
  OR2X2 OR2X2_3435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6353), .B(REGFILE_SIM_reg_bank__abc_33898_n6354), .Y(REGFILE_SIM_reg_bank__abc_33898_n6355) );
  OR2X2 OR2X2_3436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6355), .B(REGFILE_SIM_reg_bank__abc_33898_n6352), .Y(REGFILE_SIM_reg_bank__abc_33898_n6356) );
  OR2X2 OR2X2_3437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6349), .B(REGFILE_SIM_reg_bank__abc_33898_n6356), .Y(REGFILE_SIM_reg_bank__abc_33898_n6357) );
  OR2X2 OR2X2_3438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6342), .B(REGFILE_SIM_reg_bank__abc_33898_n6357), .Y(REGFILE_SIM_reg_bank__abc_33898_n6358) );
  OR2X2 OR2X2_3439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6359), .B(REGFILE_SIM_reg_bank__abc_33898_n6360), .Y(REGFILE_SIM_reg_bank__abc_33898_n6361) );
  OR2X2 OR2X2_344 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_6_), .Y(_abc_43815_n1648) );
  OR2X2 OR2X2_3440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6362), .B(REGFILE_SIM_reg_bank__abc_33898_n6363), .Y(REGFILE_SIM_reg_bank__abc_33898_n6364) );
  OR2X2 OR2X2_3441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6361), .B(REGFILE_SIM_reg_bank__abc_33898_n6364), .Y(REGFILE_SIM_reg_bank__abc_33898_n6365) );
  OR2X2 OR2X2_3442 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6367), .B(REGFILE_SIM_reg_bank__abc_33898_n6368), .Y(REGFILE_SIM_reg_bank__abc_33898_n6369) );
  OR2X2 OR2X2_3443 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6369), .B(REGFILE_SIM_reg_bank__abc_33898_n6366), .Y(REGFILE_SIM_reg_bank__abc_33898_n6370) );
  OR2X2 OR2X2_3444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6365), .B(REGFILE_SIM_reg_bank__abc_33898_n6370), .Y(REGFILE_SIM_reg_bank__abc_33898_n6371) );
  OR2X2 OR2X2_3445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6372), .B(REGFILE_SIM_reg_bank__abc_33898_n6373), .Y(REGFILE_SIM_reg_bank__abc_33898_n6374) );
  OR2X2 OR2X2_3446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6375), .B(REGFILE_SIM_reg_bank__abc_33898_n6376), .Y(REGFILE_SIM_reg_bank__abc_33898_n6377) );
  OR2X2 OR2X2_3447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6377), .B(REGFILE_SIM_reg_bank__abc_33898_n6374), .Y(REGFILE_SIM_reg_bank__abc_33898_n6378) );
  OR2X2 OR2X2_3448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6379), .B(REGFILE_SIM_reg_bank__abc_33898_n6380), .Y(REGFILE_SIM_reg_bank__abc_33898_n6381) );
  OR2X2 OR2X2_3449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6382), .B(REGFILE_SIM_reg_bank__abc_33898_n6383), .Y(REGFILE_SIM_reg_bank__abc_33898_n6384) );
  OR2X2 OR2X2_345 ( .A(_abc_43815_n1418_bF_buf4), .B(epc_q_7_), .Y(_abc_43815_n1651) );
  OR2X2 OR2X2_3450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6381), .B(REGFILE_SIM_reg_bank__abc_33898_n6384), .Y(REGFILE_SIM_reg_bank__abc_33898_n6385) );
  OR2X2 OR2X2_3451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6378), .B(REGFILE_SIM_reg_bank__abc_33898_n6385), .Y(REGFILE_SIM_reg_bank__abc_33898_n6386) );
  OR2X2 OR2X2_3452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6386), .B(REGFILE_SIM_reg_bank__abc_33898_n6371), .Y(REGFILE_SIM_reg_bank__abc_33898_n6387) );
  OR2X2 OR2X2_3453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6358), .B(REGFILE_SIM_reg_bank__abc_33898_n6387), .Y(REGFILE_SIM_reg_bank_reg_rb_o_12_) );
  OR2X2 OR2X2_3454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6389), .B(REGFILE_SIM_reg_bank__abc_33898_n6390), .Y(REGFILE_SIM_reg_bank__abc_33898_n6391) );
  OR2X2 OR2X2_3455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6392), .B(REGFILE_SIM_reg_bank__abc_33898_n6393), .Y(REGFILE_SIM_reg_bank__abc_33898_n6394) );
  OR2X2 OR2X2_3456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6394), .B(REGFILE_SIM_reg_bank__abc_33898_n6391), .Y(REGFILE_SIM_reg_bank__abc_33898_n6395) );
  OR2X2 OR2X2_3457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6396), .B(REGFILE_SIM_reg_bank__abc_33898_n6397), .Y(REGFILE_SIM_reg_bank__abc_33898_n6398) );
  OR2X2 OR2X2_3458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6399), .B(REGFILE_SIM_reg_bank__abc_33898_n6400), .Y(REGFILE_SIM_reg_bank__abc_33898_n6401) );
  OR2X2 OR2X2_3459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6398), .B(REGFILE_SIM_reg_bank__abc_33898_n6401), .Y(REGFILE_SIM_reg_bank__abc_33898_n6402) );
  OR2X2 OR2X2_346 ( .A(int32_r_5_), .B(pc_q_7_), .Y(_abc_43815_n1657) );
  OR2X2 OR2X2_3460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6395), .B(REGFILE_SIM_reg_bank__abc_33898_n6402), .Y(REGFILE_SIM_reg_bank__abc_33898_n6403) );
  OR2X2 OR2X2_3461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6404), .B(REGFILE_SIM_reg_bank__abc_33898_n6405), .Y(REGFILE_SIM_reg_bank__abc_33898_n6406) );
  OR2X2 OR2X2_3462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6407), .B(REGFILE_SIM_reg_bank__abc_33898_n6408), .Y(REGFILE_SIM_reg_bank__abc_33898_n6409) );
  OR2X2 OR2X2_3463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6406), .B(REGFILE_SIM_reg_bank__abc_33898_n6409), .Y(REGFILE_SIM_reg_bank__abc_33898_n6410) );
  OR2X2 OR2X2_3464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6411), .B(REGFILE_SIM_reg_bank__abc_33898_n6412), .Y(REGFILE_SIM_reg_bank__abc_33898_n6413) );
  OR2X2 OR2X2_3465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6414), .B(REGFILE_SIM_reg_bank__abc_33898_n6415), .Y(REGFILE_SIM_reg_bank__abc_33898_n6416) );
  OR2X2 OR2X2_3466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6416), .B(REGFILE_SIM_reg_bank__abc_33898_n6413), .Y(REGFILE_SIM_reg_bank__abc_33898_n6417) );
  OR2X2 OR2X2_3467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6410), .B(REGFILE_SIM_reg_bank__abc_33898_n6417), .Y(REGFILE_SIM_reg_bank__abc_33898_n6418) );
  OR2X2 OR2X2_3468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6403), .B(REGFILE_SIM_reg_bank__abc_33898_n6418), .Y(REGFILE_SIM_reg_bank__abc_33898_n6419) );
  OR2X2 OR2X2_3469 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6420), .B(REGFILE_SIM_reg_bank__abc_33898_n6421), .Y(REGFILE_SIM_reg_bank__abc_33898_n6422) );
  OR2X2 OR2X2_347 ( .A(_abc_43815_n1660), .B(_abc_43815_n1618_1), .Y(_abc_43815_n1661) );
  OR2X2 OR2X2_3470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6423), .B(REGFILE_SIM_reg_bank__abc_33898_n6424), .Y(REGFILE_SIM_reg_bank__abc_33898_n6425) );
  OR2X2 OR2X2_3471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6422), .B(REGFILE_SIM_reg_bank__abc_33898_n6425), .Y(REGFILE_SIM_reg_bank__abc_33898_n6426) );
  OR2X2 OR2X2_3472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6428), .B(REGFILE_SIM_reg_bank__abc_33898_n6429), .Y(REGFILE_SIM_reg_bank__abc_33898_n6430) );
  OR2X2 OR2X2_3473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6430), .B(REGFILE_SIM_reg_bank__abc_33898_n6427), .Y(REGFILE_SIM_reg_bank__abc_33898_n6431) );
  OR2X2 OR2X2_3474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6426), .B(REGFILE_SIM_reg_bank__abc_33898_n6431), .Y(REGFILE_SIM_reg_bank__abc_33898_n6432) );
  OR2X2 OR2X2_3475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6433), .B(REGFILE_SIM_reg_bank__abc_33898_n6434), .Y(REGFILE_SIM_reg_bank__abc_33898_n6435) );
  OR2X2 OR2X2_3476 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6436), .B(REGFILE_SIM_reg_bank__abc_33898_n6437), .Y(REGFILE_SIM_reg_bank__abc_33898_n6438) );
  OR2X2 OR2X2_3477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6438), .B(REGFILE_SIM_reg_bank__abc_33898_n6435), .Y(REGFILE_SIM_reg_bank__abc_33898_n6439) );
  OR2X2 OR2X2_3478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6440), .B(REGFILE_SIM_reg_bank__abc_33898_n6441), .Y(REGFILE_SIM_reg_bank__abc_33898_n6442) );
  OR2X2 OR2X2_3479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6443), .B(REGFILE_SIM_reg_bank__abc_33898_n6444), .Y(REGFILE_SIM_reg_bank__abc_33898_n6445) );
  OR2X2 OR2X2_348 ( .A(_abc_43815_n1622), .B(_abc_43815_n1661), .Y(_abc_43815_n1662) );
  OR2X2 OR2X2_3480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6442), .B(REGFILE_SIM_reg_bank__abc_33898_n6445), .Y(REGFILE_SIM_reg_bank__abc_33898_n6446) );
  OR2X2 OR2X2_3481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6439), .B(REGFILE_SIM_reg_bank__abc_33898_n6446), .Y(REGFILE_SIM_reg_bank__abc_33898_n6447) );
  OR2X2 OR2X2_3482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6447), .B(REGFILE_SIM_reg_bank__abc_33898_n6432), .Y(REGFILE_SIM_reg_bank__abc_33898_n6448) );
  OR2X2 OR2X2_3483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6419), .B(REGFILE_SIM_reg_bank__abc_33898_n6448), .Y(REGFILE_SIM_reg_bank_reg_rb_o_13_) );
  OR2X2 OR2X2_3484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6450), .B(REGFILE_SIM_reg_bank__abc_33898_n6451), .Y(REGFILE_SIM_reg_bank__abc_33898_n6452) );
  OR2X2 OR2X2_3485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6453), .B(REGFILE_SIM_reg_bank__abc_33898_n6454), .Y(REGFILE_SIM_reg_bank__abc_33898_n6455) );
  OR2X2 OR2X2_3486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6455), .B(REGFILE_SIM_reg_bank__abc_33898_n6452), .Y(REGFILE_SIM_reg_bank__abc_33898_n6456) );
  OR2X2 OR2X2_3487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6457), .B(REGFILE_SIM_reg_bank__abc_33898_n6458), .Y(REGFILE_SIM_reg_bank__abc_33898_n6459) );
  OR2X2 OR2X2_3488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6460), .B(REGFILE_SIM_reg_bank__abc_33898_n6461), .Y(REGFILE_SIM_reg_bank__abc_33898_n6462) );
  OR2X2 OR2X2_3489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6459), .B(REGFILE_SIM_reg_bank__abc_33898_n6462), .Y(REGFILE_SIM_reg_bank__abc_33898_n6463) );
  OR2X2 OR2X2_349 ( .A(_abc_43815_n1428_bF_buf1), .B(_abc_43815_n1671), .Y(_abc_43815_n1672) );
  OR2X2 OR2X2_3490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6456), .B(REGFILE_SIM_reg_bank__abc_33898_n6463), .Y(REGFILE_SIM_reg_bank__abc_33898_n6464) );
  OR2X2 OR2X2_3491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6465), .B(REGFILE_SIM_reg_bank__abc_33898_n6466), .Y(REGFILE_SIM_reg_bank__abc_33898_n6467) );
  OR2X2 OR2X2_3492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6468), .B(REGFILE_SIM_reg_bank__abc_33898_n6469), .Y(REGFILE_SIM_reg_bank__abc_33898_n6470) );
  OR2X2 OR2X2_3493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6467), .B(REGFILE_SIM_reg_bank__abc_33898_n6470), .Y(REGFILE_SIM_reg_bank__abc_33898_n6471) );
  OR2X2 OR2X2_3494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6472), .B(REGFILE_SIM_reg_bank__abc_33898_n6473), .Y(REGFILE_SIM_reg_bank__abc_33898_n6474) );
  OR2X2 OR2X2_3495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6475), .B(REGFILE_SIM_reg_bank__abc_33898_n6476), .Y(REGFILE_SIM_reg_bank__abc_33898_n6477) );
  OR2X2 OR2X2_3496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6477), .B(REGFILE_SIM_reg_bank__abc_33898_n6474), .Y(REGFILE_SIM_reg_bank__abc_33898_n6478) );
  OR2X2 OR2X2_3497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6471), .B(REGFILE_SIM_reg_bank__abc_33898_n6478), .Y(REGFILE_SIM_reg_bank__abc_33898_n6479) );
  OR2X2 OR2X2_3498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6464), .B(REGFILE_SIM_reg_bank__abc_33898_n6479), .Y(REGFILE_SIM_reg_bank__abc_33898_n6480) );
  OR2X2 OR2X2_3499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6481), .B(REGFILE_SIM_reg_bank__abc_33898_n6482), .Y(REGFILE_SIM_reg_bank__abc_33898_n6483) );
  OR2X2 OR2X2_35 ( .A(_abc_43815_n750), .B(_abc_43815_n758), .Y(_abc_43815_n759) );
  OR2X2 OR2X2_350 ( .A(_abc_43815_n1670), .B(_abc_43815_n1672), .Y(_abc_43815_n1673) );
  OR2X2 OR2X2_3500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6484), .B(REGFILE_SIM_reg_bank__abc_33898_n6485), .Y(REGFILE_SIM_reg_bank__abc_33898_n6486) );
  OR2X2 OR2X2_3501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6483), .B(REGFILE_SIM_reg_bank__abc_33898_n6486), .Y(REGFILE_SIM_reg_bank__abc_33898_n6487) );
  OR2X2 OR2X2_3502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6489), .B(REGFILE_SIM_reg_bank__abc_33898_n6490), .Y(REGFILE_SIM_reg_bank__abc_33898_n6491) );
  OR2X2 OR2X2_3503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6491), .B(REGFILE_SIM_reg_bank__abc_33898_n6488), .Y(REGFILE_SIM_reg_bank__abc_33898_n6492) );
  OR2X2 OR2X2_3504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6487), .B(REGFILE_SIM_reg_bank__abc_33898_n6492), .Y(REGFILE_SIM_reg_bank__abc_33898_n6493) );
  OR2X2 OR2X2_3505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6494), .B(REGFILE_SIM_reg_bank__abc_33898_n6495), .Y(REGFILE_SIM_reg_bank__abc_33898_n6496) );
  OR2X2 OR2X2_3506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6497), .B(REGFILE_SIM_reg_bank__abc_33898_n6498), .Y(REGFILE_SIM_reg_bank__abc_33898_n6499) );
  OR2X2 OR2X2_3507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6499), .B(REGFILE_SIM_reg_bank__abc_33898_n6496), .Y(REGFILE_SIM_reg_bank__abc_33898_n6500) );
  OR2X2 OR2X2_3508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6501), .B(REGFILE_SIM_reg_bank__abc_33898_n6502), .Y(REGFILE_SIM_reg_bank__abc_33898_n6503) );
  OR2X2 OR2X2_3509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6504), .B(REGFILE_SIM_reg_bank__abc_33898_n6505), .Y(REGFILE_SIM_reg_bank__abc_33898_n6506) );
  OR2X2 OR2X2_351 ( .A(_abc_43815_n1431_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_43815_n1674_1) );
  OR2X2 OR2X2_3510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6503), .B(REGFILE_SIM_reg_bank__abc_33898_n6506), .Y(REGFILE_SIM_reg_bank__abc_33898_n6507) );
  OR2X2 OR2X2_3511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6500), .B(REGFILE_SIM_reg_bank__abc_33898_n6507), .Y(REGFILE_SIM_reg_bank__abc_33898_n6508) );
  OR2X2 OR2X2_3512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6508), .B(REGFILE_SIM_reg_bank__abc_33898_n6493), .Y(REGFILE_SIM_reg_bank__abc_33898_n6509) );
  OR2X2 OR2X2_3513 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6480), .B(REGFILE_SIM_reg_bank__abc_33898_n6509), .Y(REGFILE_SIM_reg_bank_reg_rb_o_14_) );
  OR2X2 OR2X2_3514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6511), .B(REGFILE_SIM_reg_bank__abc_33898_n6512), .Y(REGFILE_SIM_reg_bank__abc_33898_n6513) );
  OR2X2 OR2X2_3515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6514), .B(REGFILE_SIM_reg_bank__abc_33898_n6515), .Y(REGFILE_SIM_reg_bank__abc_33898_n6516) );
  OR2X2 OR2X2_3516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6516), .B(REGFILE_SIM_reg_bank__abc_33898_n6513), .Y(REGFILE_SIM_reg_bank__abc_33898_n6517) );
  OR2X2 OR2X2_3517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6518), .B(REGFILE_SIM_reg_bank__abc_33898_n6519), .Y(REGFILE_SIM_reg_bank__abc_33898_n6520) );
  OR2X2 OR2X2_3518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6521), .B(REGFILE_SIM_reg_bank__abc_33898_n6522), .Y(REGFILE_SIM_reg_bank__abc_33898_n6523) );
  OR2X2 OR2X2_3519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6520), .B(REGFILE_SIM_reg_bank__abc_33898_n6523), .Y(REGFILE_SIM_reg_bank__abc_33898_n6524) );
  OR2X2 OR2X2_352 ( .A(_abc_43815_n1675_1), .B(_abc_43815_n1473_bF_buf4), .Y(_abc_43815_n1676) );
  OR2X2 OR2X2_3520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6517), .B(REGFILE_SIM_reg_bank__abc_33898_n6524), .Y(REGFILE_SIM_reg_bank__abc_33898_n6525) );
  OR2X2 OR2X2_3521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6526), .B(REGFILE_SIM_reg_bank__abc_33898_n6527), .Y(REGFILE_SIM_reg_bank__abc_33898_n6528) );
  OR2X2 OR2X2_3522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6529), .B(REGFILE_SIM_reg_bank__abc_33898_n6530), .Y(REGFILE_SIM_reg_bank__abc_33898_n6531) );
  OR2X2 OR2X2_3523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6528), .B(REGFILE_SIM_reg_bank__abc_33898_n6531), .Y(REGFILE_SIM_reg_bank__abc_33898_n6532) );
  OR2X2 OR2X2_3524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6533), .B(REGFILE_SIM_reg_bank__abc_33898_n6534), .Y(REGFILE_SIM_reg_bank__abc_33898_n6535) );
  OR2X2 OR2X2_3525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6536), .B(REGFILE_SIM_reg_bank__abc_33898_n6537), .Y(REGFILE_SIM_reg_bank__abc_33898_n6538) );
  OR2X2 OR2X2_3526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6538), .B(REGFILE_SIM_reg_bank__abc_33898_n6535), .Y(REGFILE_SIM_reg_bank__abc_33898_n6539) );
  OR2X2 OR2X2_3527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6532), .B(REGFILE_SIM_reg_bank__abc_33898_n6539), .Y(REGFILE_SIM_reg_bank__abc_33898_n6540) );
  OR2X2 OR2X2_3528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6525), .B(REGFILE_SIM_reg_bank__abc_33898_n6540), .Y(REGFILE_SIM_reg_bank__abc_33898_n6541) );
  OR2X2 OR2X2_3529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6542), .B(REGFILE_SIM_reg_bank__abc_33898_n6543), .Y(REGFILE_SIM_reg_bank__abc_33898_n6544) );
  OR2X2 OR2X2_353 ( .A(_abc_43815_n1633), .B(pc_q_7_), .Y(_abc_43815_n1677) );
  OR2X2 OR2X2_3530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6545), .B(REGFILE_SIM_reg_bank__abc_33898_n6546), .Y(REGFILE_SIM_reg_bank__abc_33898_n6547) );
  OR2X2 OR2X2_3531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6544), .B(REGFILE_SIM_reg_bank__abc_33898_n6547), .Y(REGFILE_SIM_reg_bank__abc_33898_n6548) );
  OR2X2 OR2X2_3532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6550), .B(REGFILE_SIM_reg_bank__abc_33898_n6551), .Y(REGFILE_SIM_reg_bank__abc_33898_n6552) );
  OR2X2 OR2X2_3533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6552), .B(REGFILE_SIM_reg_bank__abc_33898_n6549), .Y(REGFILE_SIM_reg_bank__abc_33898_n6553) );
  OR2X2 OR2X2_3534 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6548), .B(REGFILE_SIM_reg_bank__abc_33898_n6553), .Y(REGFILE_SIM_reg_bank__abc_33898_n6554) );
  OR2X2 OR2X2_3535 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6555), .B(REGFILE_SIM_reg_bank__abc_33898_n6556), .Y(REGFILE_SIM_reg_bank__abc_33898_n6557) );
  OR2X2 OR2X2_3536 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6558), .B(REGFILE_SIM_reg_bank__abc_33898_n6559), .Y(REGFILE_SIM_reg_bank__abc_33898_n6560) );
  OR2X2 OR2X2_3537 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6560), .B(REGFILE_SIM_reg_bank__abc_33898_n6557), .Y(REGFILE_SIM_reg_bank__abc_33898_n6561) );
  OR2X2 OR2X2_3538 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6562), .B(REGFILE_SIM_reg_bank__abc_33898_n6563), .Y(REGFILE_SIM_reg_bank__abc_33898_n6564) );
  OR2X2 OR2X2_3539 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6565), .B(REGFILE_SIM_reg_bank__abc_33898_n6566), .Y(REGFILE_SIM_reg_bank__abc_33898_n6567) );
  OR2X2 OR2X2_354 ( .A(_abc_43815_n1472_1_bF_buf3), .B(_abc_43815_n1680), .Y(_abc_43815_n1681) );
  OR2X2 OR2X2_3540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6564), .B(REGFILE_SIM_reg_bank__abc_33898_n6567), .Y(REGFILE_SIM_reg_bank__abc_33898_n6568) );
  OR2X2 OR2X2_3541 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6561), .B(REGFILE_SIM_reg_bank__abc_33898_n6568), .Y(REGFILE_SIM_reg_bank__abc_33898_n6569) );
  OR2X2 OR2X2_3542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6569), .B(REGFILE_SIM_reg_bank__abc_33898_n6554), .Y(REGFILE_SIM_reg_bank__abc_33898_n6570) );
  OR2X2 OR2X2_3543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6541), .B(REGFILE_SIM_reg_bank__abc_33898_n6570), .Y(REGFILE_SIM_reg_bank_reg_rb_o_15_) );
  OR2X2 OR2X2_3544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6572), .B(REGFILE_SIM_reg_bank__abc_33898_n6573), .Y(REGFILE_SIM_reg_bank__abc_33898_n6574) );
  OR2X2 OR2X2_3545 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6575), .B(REGFILE_SIM_reg_bank__abc_33898_n6576), .Y(REGFILE_SIM_reg_bank__abc_33898_n6577) );
  OR2X2 OR2X2_3546 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6577), .B(REGFILE_SIM_reg_bank__abc_33898_n6574), .Y(REGFILE_SIM_reg_bank__abc_33898_n6578) );
  OR2X2 OR2X2_3547 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6579), .B(REGFILE_SIM_reg_bank__abc_33898_n6580), .Y(REGFILE_SIM_reg_bank__abc_33898_n6581) );
  OR2X2 OR2X2_3548 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6582), .B(REGFILE_SIM_reg_bank__abc_33898_n6583), .Y(REGFILE_SIM_reg_bank__abc_33898_n6584) );
  OR2X2 OR2X2_3549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6581), .B(REGFILE_SIM_reg_bank__abc_33898_n6584), .Y(REGFILE_SIM_reg_bank__abc_33898_n6585) );
  OR2X2 OR2X2_355 ( .A(_abc_43815_n1683), .B(_abc_43815_n1656), .Y(_abc_43815_n1684) );
  OR2X2 OR2X2_3550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6578), .B(REGFILE_SIM_reg_bank__abc_33898_n6585), .Y(REGFILE_SIM_reg_bank__abc_33898_n6586) );
  OR2X2 OR2X2_3551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6587), .B(REGFILE_SIM_reg_bank__abc_33898_n6588), .Y(REGFILE_SIM_reg_bank__abc_33898_n6589) );
  OR2X2 OR2X2_3552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6590), .B(REGFILE_SIM_reg_bank__abc_33898_n6591), .Y(REGFILE_SIM_reg_bank__abc_33898_n6592) );
  OR2X2 OR2X2_3553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6589), .B(REGFILE_SIM_reg_bank__abc_33898_n6592), .Y(REGFILE_SIM_reg_bank__abc_33898_n6593) );
  OR2X2 OR2X2_3554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6594), .B(REGFILE_SIM_reg_bank__abc_33898_n6595), .Y(REGFILE_SIM_reg_bank__abc_33898_n6596) );
  OR2X2 OR2X2_3555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6597), .B(REGFILE_SIM_reg_bank__abc_33898_n6598), .Y(REGFILE_SIM_reg_bank__abc_33898_n6599) );
  OR2X2 OR2X2_3556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6599), .B(REGFILE_SIM_reg_bank__abc_33898_n6596), .Y(REGFILE_SIM_reg_bank__abc_33898_n6600) );
  OR2X2 OR2X2_3557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6593), .B(REGFILE_SIM_reg_bank__abc_33898_n6600), .Y(REGFILE_SIM_reg_bank__abc_33898_n6601) );
  OR2X2 OR2X2_3558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6586), .B(REGFILE_SIM_reg_bank__abc_33898_n6601), .Y(REGFILE_SIM_reg_bank__abc_33898_n6602) );
  OR2X2 OR2X2_3559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6603), .B(REGFILE_SIM_reg_bank__abc_33898_n6604), .Y(REGFILE_SIM_reg_bank__abc_33898_n6605) );
  OR2X2 OR2X2_356 ( .A(_abc_43815_n1686_1), .B(_abc_43815_n1278_bF_buf2), .Y(_abc_43815_n1687) );
  OR2X2 OR2X2_3560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6606), .B(REGFILE_SIM_reg_bank__abc_33898_n6607), .Y(REGFILE_SIM_reg_bank__abc_33898_n6608) );
  OR2X2 OR2X2_3561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6605), .B(REGFILE_SIM_reg_bank__abc_33898_n6608), .Y(REGFILE_SIM_reg_bank__abc_33898_n6609) );
  OR2X2 OR2X2_3562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6611), .B(REGFILE_SIM_reg_bank__abc_33898_n6612), .Y(REGFILE_SIM_reg_bank__abc_33898_n6613) );
  OR2X2 OR2X2_3563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6613), .B(REGFILE_SIM_reg_bank__abc_33898_n6610), .Y(REGFILE_SIM_reg_bank__abc_33898_n6614) );
  OR2X2 OR2X2_3564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6609), .B(REGFILE_SIM_reg_bank__abc_33898_n6614), .Y(REGFILE_SIM_reg_bank__abc_33898_n6615) );
  OR2X2 OR2X2_3565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6616), .B(REGFILE_SIM_reg_bank__abc_33898_n6617), .Y(REGFILE_SIM_reg_bank__abc_33898_n6618) );
  OR2X2 OR2X2_3566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6619), .B(REGFILE_SIM_reg_bank__abc_33898_n6620), .Y(REGFILE_SIM_reg_bank__abc_33898_n6621) );
  OR2X2 OR2X2_3567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6621), .B(REGFILE_SIM_reg_bank__abc_33898_n6618), .Y(REGFILE_SIM_reg_bank__abc_33898_n6622) );
  OR2X2 OR2X2_3568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6623), .B(REGFILE_SIM_reg_bank__abc_33898_n6624), .Y(REGFILE_SIM_reg_bank__abc_33898_n6625) );
  OR2X2 OR2X2_3569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6626), .B(REGFILE_SIM_reg_bank__abc_33898_n6627), .Y(REGFILE_SIM_reg_bank__abc_33898_n6628) );
  OR2X2 OR2X2_357 ( .A(_abc_43815_n1685), .B(_abc_43815_n1687), .Y(_abc_43815_n1688) );
  OR2X2 OR2X2_3570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6625), .B(REGFILE_SIM_reg_bank__abc_33898_n6628), .Y(REGFILE_SIM_reg_bank__abc_33898_n6629) );
  OR2X2 OR2X2_3571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6622), .B(REGFILE_SIM_reg_bank__abc_33898_n6629), .Y(REGFILE_SIM_reg_bank__abc_33898_n6630) );
  OR2X2 OR2X2_3572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6630), .B(REGFILE_SIM_reg_bank__abc_33898_n6615), .Y(REGFILE_SIM_reg_bank__abc_33898_n6631) );
  OR2X2 OR2X2_3573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6602), .B(REGFILE_SIM_reg_bank__abc_33898_n6631), .Y(REGFILE_SIM_reg_bank_reg_rb_o_16_) );
  OR2X2 OR2X2_3574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6633), .B(REGFILE_SIM_reg_bank__abc_33898_n6634), .Y(REGFILE_SIM_reg_bank__abc_33898_n6635) );
  OR2X2 OR2X2_3575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6636), .B(REGFILE_SIM_reg_bank__abc_33898_n6637), .Y(REGFILE_SIM_reg_bank__abc_33898_n6638) );
  OR2X2 OR2X2_3576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6638), .B(REGFILE_SIM_reg_bank__abc_33898_n6635), .Y(REGFILE_SIM_reg_bank__abc_33898_n6639) );
  OR2X2 OR2X2_3577 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6640), .B(REGFILE_SIM_reg_bank__abc_33898_n6641), .Y(REGFILE_SIM_reg_bank__abc_33898_n6642) );
  OR2X2 OR2X2_3578 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6643), .B(REGFILE_SIM_reg_bank__abc_33898_n6644), .Y(REGFILE_SIM_reg_bank__abc_33898_n6645) );
  OR2X2 OR2X2_3579 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6642), .B(REGFILE_SIM_reg_bank__abc_33898_n6645), .Y(REGFILE_SIM_reg_bank__abc_33898_n6646) );
  OR2X2 OR2X2_358 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_7_), .Y(_abc_43815_n1689_1) );
  OR2X2 OR2X2_3580 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6639), .B(REGFILE_SIM_reg_bank__abc_33898_n6646), .Y(REGFILE_SIM_reg_bank__abc_33898_n6647) );
  OR2X2 OR2X2_3581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6648), .B(REGFILE_SIM_reg_bank__abc_33898_n6649), .Y(REGFILE_SIM_reg_bank__abc_33898_n6650) );
  OR2X2 OR2X2_3582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6651), .B(REGFILE_SIM_reg_bank__abc_33898_n6652), .Y(REGFILE_SIM_reg_bank__abc_33898_n6653) );
  OR2X2 OR2X2_3583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6650), .B(REGFILE_SIM_reg_bank__abc_33898_n6653), .Y(REGFILE_SIM_reg_bank__abc_33898_n6654) );
  OR2X2 OR2X2_3584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6655), .B(REGFILE_SIM_reg_bank__abc_33898_n6656), .Y(REGFILE_SIM_reg_bank__abc_33898_n6657) );
  OR2X2 OR2X2_3585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6658), .B(REGFILE_SIM_reg_bank__abc_33898_n6659), .Y(REGFILE_SIM_reg_bank__abc_33898_n6660) );
  OR2X2 OR2X2_3586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6660), .B(REGFILE_SIM_reg_bank__abc_33898_n6657), .Y(REGFILE_SIM_reg_bank__abc_33898_n6661) );
  OR2X2 OR2X2_3587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6654), .B(REGFILE_SIM_reg_bank__abc_33898_n6661), .Y(REGFILE_SIM_reg_bank__abc_33898_n6662) );
  OR2X2 OR2X2_3588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6647), .B(REGFILE_SIM_reg_bank__abc_33898_n6662), .Y(REGFILE_SIM_reg_bank__abc_33898_n6663) );
  OR2X2 OR2X2_3589 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6664), .B(REGFILE_SIM_reg_bank__abc_33898_n6665), .Y(REGFILE_SIM_reg_bank__abc_33898_n6666) );
  OR2X2 OR2X2_359 ( .A(_abc_43815_n1678), .B(pc_q_8_), .Y(_abc_43815_n1693) );
  OR2X2 OR2X2_3590 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6667), .B(REGFILE_SIM_reg_bank__abc_33898_n6668), .Y(REGFILE_SIM_reg_bank__abc_33898_n6669) );
  OR2X2 OR2X2_3591 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6666), .B(REGFILE_SIM_reg_bank__abc_33898_n6669), .Y(REGFILE_SIM_reg_bank__abc_33898_n6670) );
  OR2X2 OR2X2_3592 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6672), .B(REGFILE_SIM_reg_bank__abc_33898_n6673), .Y(REGFILE_SIM_reg_bank__abc_33898_n6674) );
  OR2X2 OR2X2_3593 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6674), .B(REGFILE_SIM_reg_bank__abc_33898_n6671), .Y(REGFILE_SIM_reg_bank__abc_33898_n6675) );
  OR2X2 OR2X2_3594 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6670), .B(REGFILE_SIM_reg_bank__abc_33898_n6675), .Y(REGFILE_SIM_reg_bank__abc_33898_n6676) );
  OR2X2 OR2X2_3595 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6677), .B(REGFILE_SIM_reg_bank__abc_33898_n6678), .Y(REGFILE_SIM_reg_bank__abc_33898_n6679) );
  OR2X2 OR2X2_3596 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6680), .B(REGFILE_SIM_reg_bank__abc_33898_n6681), .Y(REGFILE_SIM_reg_bank__abc_33898_n6682) );
  OR2X2 OR2X2_3597 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6682), .B(REGFILE_SIM_reg_bank__abc_33898_n6679), .Y(REGFILE_SIM_reg_bank__abc_33898_n6683) );
  OR2X2 OR2X2_3598 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6684), .B(REGFILE_SIM_reg_bank__abc_33898_n6685), .Y(REGFILE_SIM_reg_bank__abc_33898_n6686) );
  OR2X2 OR2X2_3599 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6687), .B(REGFILE_SIM_reg_bank__abc_33898_n6688), .Y(REGFILE_SIM_reg_bank__abc_33898_n6689) );
  OR2X2 OR2X2_36 ( .A(_abc_43815_n760_1), .B(_abc_43815_n746), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_) );
  OR2X2 OR2X2_360 ( .A(_abc_43815_n1696), .B(_abc_43815_n1278_bF_buf1), .Y(_abc_43815_n1697) );
  OR2X2 OR2X2_3600 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6686), .B(REGFILE_SIM_reg_bank__abc_33898_n6689), .Y(REGFILE_SIM_reg_bank__abc_33898_n6690) );
  OR2X2 OR2X2_3601 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6683), .B(REGFILE_SIM_reg_bank__abc_33898_n6690), .Y(REGFILE_SIM_reg_bank__abc_33898_n6691) );
  OR2X2 OR2X2_3602 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6691), .B(REGFILE_SIM_reg_bank__abc_33898_n6676), .Y(REGFILE_SIM_reg_bank__abc_33898_n6692) );
  OR2X2 OR2X2_3603 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6663), .B(REGFILE_SIM_reg_bank__abc_33898_n6692), .Y(REGFILE_SIM_reg_bank_reg_rb_o_17_) );
  OR2X2 OR2X2_3604 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6694), .B(REGFILE_SIM_reg_bank__abc_33898_n6695), .Y(REGFILE_SIM_reg_bank__abc_33898_n6696) );
  OR2X2 OR2X2_3605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6697), .B(REGFILE_SIM_reg_bank__abc_33898_n6698), .Y(REGFILE_SIM_reg_bank__abc_33898_n6699) );
  OR2X2 OR2X2_3606 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6699), .B(REGFILE_SIM_reg_bank__abc_33898_n6696), .Y(REGFILE_SIM_reg_bank__abc_33898_n6700) );
  OR2X2 OR2X2_3607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6701), .B(REGFILE_SIM_reg_bank__abc_33898_n6702), .Y(REGFILE_SIM_reg_bank__abc_33898_n6703) );
  OR2X2 OR2X2_3608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6704), .B(REGFILE_SIM_reg_bank__abc_33898_n6705), .Y(REGFILE_SIM_reg_bank__abc_33898_n6706) );
  OR2X2 OR2X2_3609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6703), .B(REGFILE_SIM_reg_bank__abc_33898_n6706), .Y(REGFILE_SIM_reg_bank__abc_33898_n6707) );
  OR2X2 OR2X2_361 ( .A(_abc_43815_n1472_1_bF_buf2), .B(_abc_43815_n1696), .Y(_abc_43815_n1699) );
  OR2X2 OR2X2_3610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6700), .B(REGFILE_SIM_reg_bank__abc_33898_n6707), .Y(REGFILE_SIM_reg_bank__abc_33898_n6708) );
  OR2X2 OR2X2_3611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6709), .B(REGFILE_SIM_reg_bank__abc_33898_n6710), .Y(REGFILE_SIM_reg_bank__abc_33898_n6711) );
  OR2X2 OR2X2_3612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6712), .B(REGFILE_SIM_reg_bank__abc_33898_n6713), .Y(REGFILE_SIM_reg_bank__abc_33898_n6714) );
  OR2X2 OR2X2_3613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6711), .B(REGFILE_SIM_reg_bank__abc_33898_n6714), .Y(REGFILE_SIM_reg_bank__abc_33898_n6715) );
  OR2X2 OR2X2_3614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6716), .B(REGFILE_SIM_reg_bank__abc_33898_n6717), .Y(REGFILE_SIM_reg_bank__abc_33898_n6718) );
  OR2X2 OR2X2_3615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6719), .B(REGFILE_SIM_reg_bank__abc_33898_n6720), .Y(REGFILE_SIM_reg_bank__abc_33898_n6721) );
  OR2X2 OR2X2_3616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6721), .B(REGFILE_SIM_reg_bank__abc_33898_n6718), .Y(REGFILE_SIM_reg_bank__abc_33898_n6722) );
  OR2X2 OR2X2_3617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6715), .B(REGFILE_SIM_reg_bank__abc_33898_n6722), .Y(REGFILE_SIM_reg_bank__abc_33898_n6723) );
  OR2X2 OR2X2_3618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6708), .B(REGFILE_SIM_reg_bank__abc_33898_n6723), .Y(REGFILE_SIM_reg_bank__abc_33898_n6724) );
  OR2X2 OR2X2_3619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6725), .B(REGFILE_SIM_reg_bank__abc_33898_n6726), .Y(REGFILE_SIM_reg_bank__abc_33898_n6727) );
  OR2X2 OR2X2_362 ( .A(_abc_43815_n1664), .B(_abc_43815_n1702), .Y(_abc_43815_n1703) );
  OR2X2 OR2X2_3620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6728), .B(REGFILE_SIM_reg_bank__abc_33898_n6729), .Y(REGFILE_SIM_reg_bank__abc_33898_n6730) );
  OR2X2 OR2X2_3621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6727), .B(REGFILE_SIM_reg_bank__abc_33898_n6730), .Y(REGFILE_SIM_reg_bank__abc_33898_n6731) );
  OR2X2 OR2X2_3622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6733), .B(REGFILE_SIM_reg_bank__abc_33898_n6734), .Y(REGFILE_SIM_reg_bank__abc_33898_n6735) );
  OR2X2 OR2X2_3623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6735), .B(REGFILE_SIM_reg_bank__abc_33898_n6732), .Y(REGFILE_SIM_reg_bank__abc_33898_n6736) );
  OR2X2 OR2X2_3624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6731), .B(REGFILE_SIM_reg_bank__abc_33898_n6736), .Y(REGFILE_SIM_reg_bank__abc_33898_n6737) );
  OR2X2 OR2X2_3625 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6738), .B(REGFILE_SIM_reg_bank__abc_33898_n6739), .Y(REGFILE_SIM_reg_bank__abc_33898_n6740) );
  OR2X2 OR2X2_3626 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6741), .B(REGFILE_SIM_reg_bank__abc_33898_n6742), .Y(REGFILE_SIM_reg_bank__abc_33898_n6743) );
  OR2X2 OR2X2_3627 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6743), .B(REGFILE_SIM_reg_bank__abc_33898_n6740), .Y(REGFILE_SIM_reg_bank__abc_33898_n6744) );
  OR2X2 OR2X2_3628 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6745), .B(REGFILE_SIM_reg_bank__abc_33898_n6746), .Y(REGFILE_SIM_reg_bank__abc_33898_n6747) );
  OR2X2 OR2X2_3629 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6748), .B(REGFILE_SIM_reg_bank__abc_33898_n6749), .Y(REGFILE_SIM_reg_bank__abc_33898_n6750) );
  OR2X2 OR2X2_363 ( .A(alu_op_r_4_), .B(pc_q_8_), .Y(_abc_43815_n1704) );
  OR2X2 OR2X2_3630 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6747), .B(REGFILE_SIM_reg_bank__abc_33898_n6750), .Y(REGFILE_SIM_reg_bank__abc_33898_n6751) );
  OR2X2 OR2X2_3631 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6744), .B(REGFILE_SIM_reg_bank__abc_33898_n6751), .Y(REGFILE_SIM_reg_bank__abc_33898_n6752) );
  OR2X2 OR2X2_3632 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6752), .B(REGFILE_SIM_reg_bank__abc_33898_n6737), .Y(REGFILE_SIM_reg_bank__abc_33898_n6753) );
  OR2X2 OR2X2_3633 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6724), .B(REGFILE_SIM_reg_bank__abc_33898_n6753), .Y(REGFILE_SIM_reg_bank_reg_rb_o_18_) );
  OR2X2 OR2X2_3634 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6755), .B(REGFILE_SIM_reg_bank__abc_33898_n6756), .Y(REGFILE_SIM_reg_bank__abc_33898_n6757) );
  OR2X2 OR2X2_3635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6758), .B(REGFILE_SIM_reg_bank__abc_33898_n6759), .Y(REGFILE_SIM_reg_bank__abc_33898_n6760) );
  OR2X2 OR2X2_3636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6760), .B(REGFILE_SIM_reg_bank__abc_33898_n6757), .Y(REGFILE_SIM_reg_bank__abc_33898_n6761) );
  OR2X2 OR2X2_3637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6762), .B(REGFILE_SIM_reg_bank__abc_33898_n6763), .Y(REGFILE_SIM_reg_bank__abc_33898_n6764) );
  OR2X2 OR2X2_3638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6765), .B(REGFILE_SIM_reg_bank__abc_33898_n6766), .Y(REGFILE_SIM_reg_bank__abc_33898_n6767) );
  OR2X2 OR2X2_3639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6764), .B(REGFILE_SIM_reg_bank__abc_33898_n6767), .Y(REGFILE_SIM_reg_bank__abc_33898_n6768) );
  OR2X2 OR2X2_364 ( .A(_abc_43815_n1703), .B(_abc_43815_n1707), .Y(_abc_43815_n1708) );
  OR2X2 OR2X2_3640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6761), .B(REGFILE_SIM_reg_bank__abc_33898_n6768), .Y(REGFILE_SIM_reg_bank__abc_33898_n6769) );
  OR2X2 OR2X2_3641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6770), .B(REGFILE_SIM_reg_bank__abc_33898_n6771), .Y(REGFILE_SIM_reg_bank__abc_33898_n6772) );
  OR2X2 OR2X2_3642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6773), .B(REGFILE_SIM_reg_bank__abc_33898_n6774), .Y(REGFILE_SIM_reg_bank__abc_33898_n6775) );
  OR2X2 OR2X2_3643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6772), .B(REGFILE_SIM_reg_bank__abc_33898_n6775), .Y(REGFILE_SIM_reg_bank__abc_33898_n6776) );
  OR2X2 OR2X2_3644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6777), .B(REGFILE_SIM_reg_bank__abc_33898_n6778), .Y(REGFILE_SIM_reg_bank__abc_33898_n6779) );
  OR2X2 OR2X2_3645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6780), .B(REGFILE_SIM_reg_bank__abc_33898_n6781), .Y(REGFILE_SIM_reg_bank__abc_33898_n6782) );
  OR2X2 OR2X2_3646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6782), .B(REGFILE_SIM_reg_bank__abc_33898_n6779), .Y(REGFILE_SIM_reg_bank__abc_33898_n6783) );
  OR2X2 OR2X2_3647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6776), .B(REGFILE_SIM_reg_bank__abc_33898_n6783), .Y(REGFILE_SIM_reg_bank__abc_33898_n6784) );
  OR2X2 OR2X2_3648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6769), .B(REGFILE_SIM_reg_bank__abc_33898_n6784), .Y(REGFILE_SIM_reg_bank__abc_33898_n6785) );
  OR2X2 OR2X2_3649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6786), .B(REGFILE_SIM_reg_bank__abc_33898_n6787), .Y(REGFILE_SIM_reg_bank__abc_33898_n6788) );
  OR2X2 OR2X2_365 ( .A(_abc_43815_n1712), .B(_abc_43815_n1700), .Y(_abc_43815_n1713) );
  OR2X2 OR2X2_3650 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6789), .B(REGFILE_SIM_reg_bank__abc_33898_n6790), .Y(REGFILE_SIM_reg_bank__abc_33898_n6791) );
  OR2X2 OR2X2_3651 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6788), .B(REGFILE_SIM_reg_bank__abc_33898_n6791), .Y(REGFILE_SIM_reg_bank__abc_33898_n6792) );
  OR2X2 OR2X2_3652 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6794), .B(REGFILE_SIM_reg_bank__abc_33898_n6795), .Y(REGFILE_SIM_reg_bank__abc_33898_n6796) );
  OR2X2 OR2X2_3653 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6796), .B(REGFILE_SIM_reg_bank__abc_33898_n6793), .Y(REGFILE_SIM_reg_bank__abc_33898_n6797) );
  OR2X2 OR2X2_3654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6792), .B(REGFILE_SIM_reg_bank__abc_33898_n6797), .Y(REGFILE_SIM_reg_bank__abc_33898_n6798) );
  OR2X2 OR2X2_3655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6799), .B(REGFILE_SIM_reg_bank__abc_33898_n6800), .Y(REGFILE_SIM_reg_bank__abc_33898_n6801) );
  OR2X2 OR2X2_3656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6802), .B(REGFILE_SIM_reg_bank__abc_33898_n6803), .Y(REGFILE_SIM_reg_bank__abc_33898_n6804) );
  OR2X2 OR2X2_3657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6804), .B(REGFILE_SIM_reg_bank__abc_33898_n6801), .Y(REGFILE_SIM_reg_bank__abc_33898_n6805) );
  OR2X2 OR2X2_3658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6806), .B(REGFILE_SIM_reg_bank__abc_33898_n6807), .Y(REGFILE_SIM_reg_bank__abc_33898_n6808) );
  OR2X2 OR2X2_3659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6809), .B(REGFILE_SIM_reg_bank__abc_33898_n6810), .Y(REGFILE_SIM_reg_bank__abc_33898_n6811) );
  OR2X2 OR2X2_366 ( .A(_abc_43815_n1473_bF_buf3), .B(_abc_43815_n1715), .Y(_abc_43815_n1716) );
  OR2X2 OR2X2_3660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6808), .B(REGFILE_SIM_reg_bank__abc_33898_n6811), .Y(REGFILE_SIM_reg_bank__abc_33898_n6812) );
  OR2X2 OR2X2_3661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6805), .B(REGFILE_SIM_reg_bank__abc_33898_n6812), .Y(REGFILE_SIM_reg_bank__abc_33898_n6813) );
  OR2X2 OR2X2_3662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6813), .B(REGFILE_SIM_reg_bank__abc_33898_n6798), .Y(REGFILE_SIM_reg_bank__abc_33898_n6814) );
  OR2X2 OR2X2_3663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6785), .B(REGFILE_SIM_reg_bank__abc_33898_n6814), .Y(REGFILE_SIM_reg_bank_reg_rb_o_19_) );
  OR2X2 OR2X2_3664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6816), .B(REGFILE_SIM_reg_bank__abc_33898_n6817), .Y(REGFILE_SIM_reg_bank__abc_33898_n6818) );
  OR2X2 OR2X2_3665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6819), .B(REGFILE_SIM_reg_bank__abc_33898_n6820), .Y(REGFILE_SIM_reg_bank__abc_33898_n6821) );
  OR2X2 OR2X2_3666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6821), .B(REGFILE_SIM_reg_bank__abc_33898_n6818), .Y(REGFILE_SIM_reg_bank__abc_33898_n6822) );
  OR2X2 OR2X2_3667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6823), .B(REGFILE_SIM_reg_bank__abc_33898_n6824), .Y(REGFILE_SIM_reg_bank__abc_33898_n6825) );
  OR2X2 OR2X2_3668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6826), .B(REGFILE_SIM_reg_bank__abc_33898_n6827), .Y(REGFILE_SIM_reg_bank__abc_33898_n6828) );
  OR2X2 OR2X2_3669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6825), .B(REGFILE_SIM_reg_bank__abc_33898_n6828), .Y(REGFILE_SIM_reg_bank__abc_33898_n6829) );
  OR2X2 OR2X2_367 ( .A(_abc_43815_n1714), .B(_abc_43815_n1716), .Y(_abc_43815_n1717) );
  OR2X2 OR2X2_3670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6822), .B(REGFILE_SIM_reg_bank__abc_33898_n6829), .Y(REGFILE_SIM_reg_bank__abc_33898_n6830) );
  OR2X2 OR2X2_3671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6831), .B(REGFILE_SIM_reg_bank__abc_33898_n6832), .Y(REGFILE_SIM_reg_bank__abc_33898_n6833) );
  OR2X2 OR2X2_3672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6834), .B(REGFILE_SIM_reg_bank__abc_33898_n6835), .Y(REGFILE_SIM_reg_bank__abc_33898_n6836) );
  OR2X2 OR2X2_3673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6833), .B(REGFILE_SIM_reg_bank__abc_33898_n6836), .Y(REGFILE_SIM_reg_bank__abc_33898_n6837) );
  OR2X2 OR2X2_3674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6838), .B(REGFILE_SIM_reg_bank__abc_33898_n6839), .Y(REGFILE_SIM_reg_bank__abc_33898_n6840) );
  OR2X2 OR2X2_3675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6841), .B(REGFILE_SIM_reg_bank__abc_33898_n6842), .Y(REGFILE_SIM_reg_bank__abc_33898_n6843) );
  OR2X2 OR2X2_3676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6843), .B(REGFILE_SIM_reg_bank__abc_33898_n6840), .Y(REGFILE_SIM_reg_bank__abc_33898_n6844) );
  OR2X2 OR2X2_3677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6837), .B(REGFILE_SIM_reg_bank__abc_33898_n6844), .Y(REGFILE_SIM_reg_bank__abc_33898_n6845) );
  OR2X2 OR2X2_3678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6830), .B(REGFILE_SIM_reg_bank__abc_33898_n6845), .Y(REGFILE_SIM_reg_bank__abc_33898_n6846) );
  OR2X2 OR2X2_3679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6847), .B(REGFILE_SIM_reg_bank__abc_33898_n6848), .Y(REGFILE_SIM_reg_bank__abc_33898_n6849) );
  OR2X2 OR2X2_368 ( .A(_abc_43815_n1718), .B(_abc_43815_n1350_bF_buf3), .Y(_abc_43815_n1719_1) );
  OR2X2 OR2X2_3680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6850), .B(REGFILE_SIM_reg_bank__abc_33898_n6851), .Y(REGFILE_SIM_reg_bank__abc_33898_n6852) );
  OR2X2 OR2X2_3681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6849), .B(REGFILE_SIM_reg_bank__abc_33898_n6852), .Y(REGFILE_SIM_reg_bank__abc_33898_n6853) );
  OR2X2 OR2X2_3682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6855), .B(REGFILE_SIM_reg_bank__abc_33898_n6856), .Y(REGFILE_SIM_reg_bank__abc_33898_n6857) );
  OR2X2 OR2X2_3683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6857), .B(REGFILE_SIM_reg_bank__abc_33898_n6854), .Y(REGFILE_SIM_reg_bank__abc_33898_n6858) );
  OR2X2 OR2X2_3684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6853), .B(REGFILE_SIM_reg_bank__abc_33898_n6858), .Y(REGFILE_SIM_reg_bank__abc_33898_n6859) );
  OR2X2 OR2X2_3685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6860), .B(REGFILE_SIM_reg_bank__abc_33898_n6861), .Y(REGFILE_SIM_reg_bank__abc_33898_n6862) );
  OR2X2 OR2X2_3686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6863), .B(REGFILE_SIM_reg_bank__abc_33898_n6864), .Y(REGFILE_SIM_reg_bank__abc_33898_n6865) );
  OR2X2 OR2X2_3687 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6865), .B(REGFILE_SIM_reg_bank__abc_33898_n6862), .Y(REGFILE_SIM_reg_bank__abc_33898_n6866) );
  OR2X2 OR2X2_3688 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6867), .B(REGFILE_SIM_reg_bank__abc_33898_n6868), .Y(REGFILE_SIM_reg_bank__abc_33898_n6869) );
  OR2X2 OR2X2_3689 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6870), .B(REGFILE_SIM_reg_bank__abc_33898_n6871), .Y(REGFILE_SIM_reg_bank__abc_33898_n6872) );
  OR2X2 OR2X2_369 ( .A(_abc_43815_n1720), .B(_abc_43815_n1721), .Y(_abc_43815_n1722_1) );
  OR2X2 OR2X2_3690 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6869), .B(REGFILE_SIM_reg_bank__abc_33898_n6872), .Y(REGFILE_SIM_reg_bank__abc_33898_n6873) );
  OR2X2 OR2X2_3691 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6866), .B(REGFILE_SIM_reg_bank__abc_33898_n6873), .Y(REGFILE_SIM_reg_bank__abc_33898_n6874) );
  OR2X2 OR2X2_3692 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6874), .B(REGFILE_SIM_reg_bank__abc_33898_n6859), .Y(REGFILE_SIM_reg_bank__abc_33898_n6875) );
  OR2X2 OR2X2_3693 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6846), .B(REGFILE_SIM_reg_bank__abc_33898_n6875), .Y(REGFILE_SIM_reg_bank_reg_rb_o_20_) );
  OR2X2 OR2X2_3694 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6877), .B(REGFILE_SIM_reg_bank__abc_33898_n6878), .Y(REGFILE_SIM_reg_bank__abc_33898_n6879) );
  OR2X2 OR2X2_3695 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6880), .B(REGFILE_SIM_reg_bank__abc_33898_n6881), .Y(REGFILE_SIM_reg_bank__abc_33898_n6882) );
  OR2X2 OR2X2_3696 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6882), .B(REGFILE_SIM_reg_bank__abc_33898_n6879), .Y(REGFILE_SIM_reg_bank__abc_33898_n6883) );
  OR2X2 OR2X2_3697 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6884), .B(REGFILE_SIM_reg_bank__abc_33898_n6885), .Y(REGFILE_SIM_reg_bank__abc_33898_n6886) );
  OR2X2 OR2X2_3698 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6887), .B(REGFILE_SIM_reg_bank__abc_33898_n6888), .Y(REGFILE_SIM_reg_bank__abc_33898_n6889) );
  OR2X2 OR2X2_3699 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6886), .B(REGFILE_SIM_reg_bank__abc_33898_n6889), .Y(REGFILE_SIM_reg_bank__abc_33898_n6890) );
  OR2X2 OR2X2_37 ( .A(_abc_43815_n763), .B(_abc_43815_n764), .Y(_abc_43815_n765_1) );
  OR2X2 OR2X2_370 ( .A(_abc_43815_n1413_bF_buf1), .B(_abc_43815_n1722_1), .Y(_abc_43815_n1723) );
  OR2X2 OR2X2_3700 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6883), .B(REGFILE_SIM_reg_bank__abc_33898_n6890), .Y(REGFILE_SIM_reg_bank__abc_33898_n6891) );
  OR2X2 OR2X2_3701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6892), .B(REGFILE_SIM_reg_bank__abc_33898_n6893), .Y(REGFILE_SIM_reg_bank__abc_33898_n6894) );
  OR2X2 OR2X2_3702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6895), .B(REGFILE_SIM_reg_bank__abc_33898_n6896), .Y(REGFILE_SIM_reg_bank__abc_33898_n6897) );
  OR2X2 OR2X2_3703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6894), .B(REGFILE_SIM_reg_bank__abc_33898_n6897), .Y(REGFILE_SIM_reg_bank__abc_33898_n6898) );
  OR2X2 OR2X2_3704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6899), .B(REGFILE_SIM_reg_bank__abc_33898_n6900), .Y(REGFILE_SIM_reg_bank__abc_33898_n6901) );
  OR2X2 OR2X2_3705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6902), .B(REGFILE_SIM_reg_bank__abc_33898_n6903), .Y(REGFILE_SIM_reg_bank__abc_33898_n6904) );
  OR2X2 OR2X2_3706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6904), .B(REGFILE_SIM_reg_bank__abc_33898_n6901), .Y(REGFILE_SIM_reg_bank__abc_33898_n6905) );
  OR2X2 OR2X2_3707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6898), .B(REGFILE_SIM_reg_bank__abc_33898_n6905), .Y(REGFILE_SIM_reg_bank__abc_33898_n6906) );
  OR2X2 OR2X2_3708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6891), .B(REGFILE_SIM_reg_bank__abc_33898_n6906), .Y(REGFILE_SIM_reg_bank__abc_33898_n6907) );
  OR2X2 OR2X2_3709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6908), .B(REGFILE_SIM_reg_bank__abc_33898_n6909), .Y(REGFILE_SIM_reg_bank__abc_33898_n6910) );
  OR2X2 OR2X2_371 ( .A(_abc_43815_n1725), .B(_abc_43815_n1698), .Y(_abc_43815_n1726) );
  OR2X2 OR2X2_3710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6911), .B(REGFILE_SIM_reg_bank__abc_33898_n6912), .Y(REGFILE_SIM_reg_bank__abc_33898_n6913) );
  OR2X2 OR2X2_3711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6910), .B(REGFILE_SIM_reg_bank__abc_33898_n6913), .Y(REGFILE_SIM_reg_bank__abc_33898_n6914) );
  OR2X2 OR2X2_3712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6916), .B(REGFILE_SIM_reg_bank__abc_33898_n6917), .Y(REGFILE_SIM_reg_bank__abc_33898_n6918) );
  OR2X2 OR2X2_3713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6918), .B(REGFILE_SIM_reg_bank__abc_33898_n6915), .Y(REGFILE_SIM_reg_bank__abc_33898_n6919) );
  OR2X2 OR2X2_3714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6914), .B(REGFILE_SIM_reg_bank__abc_33898_n6919), .Y(REGFILE_SIM_reg_bank__abc_33898_n6920) );
  OR2X2 OR2X2_3715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6921), .B(REGFILE_SIM_reg_bank__abc_33898_n6922), .Y(REGFILE_SIM_reg_bank__abc_33898_n6923) );
  OR2X2 OR2X2_3716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6924), .B(REGFILE_SIM_reg_bank__abc_33898_n6925), .Y(REGFILE_SIM_reg_bank__abc_33898_n6926) );
  OR2X2 OR2X2_3717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6926), .B(REGFILE_SIM_reg_bank__abc_33898_n6923), .Y(REGFILE_SIM_reg_bank__abc_33898_n6927) );
  OR2X2 OR2X2_3718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6928), .B(REGFILE_SIM_reg_bank__abc_33898_n6929), .Y(REGFILE_SIM_reg_bank__abc_33898_n6930) );
  OR2X2 OR2X2_3719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6931), .B(REGFILE_SIM_reg_bank__abc_33898_n6932), .Y(REGFILE_SIM_reg_bank__abc_33898_n6933) );
  OR2X2 OR2X2_372 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_8_), .Y(_abc_43815_n1727) );
  OR2X2 OR2X2_3720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6930), .B(REGFILE_SIM_reg_bank__abc_33898_n6933), .Y(REGFILE_SIM_reg_bank__abc_33898_n6934) );
  OR2X2 OR2X2_3721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6927), .B(REGFILE_SIM_reg_bank__abc_33898_n6934), .Y(REGFILE_SIM_reg_bank__abc_33898_n6935) );
  OR2X2 OR2X2_3722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6935), .B(REGFILE_SIM_reg_bank__abc_33898_n6920), .Y(REGFILE_SIM_reg_bank__abc_33898_n6936) );
  OR2X2 OR2X2_3723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6907), .B(REGFILE_SIM_reg_bank__abc_33898_n6936), .Y(REGFILE_SIM_reg_bank_reg_rb_o_21_) );
  OR2X2 OR2X2_3724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6938), .B(REGFILE_SIM_reg_bank__abc_33898_n6939), .Y(REGFILE_SIM_reg_bank__abc_33898_n6940) );
  OR2X2 OR2X2_3725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6941), .B(REGFILE_SIM_reg_bank__abc_33898_n6942), .Y(REGFILE_SIM_reg_bank__abc_33898_n6943) );
  OR2X2 OR2X2_3726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6943), .B(REGFILE_SIM_reg_bank__abc_33898_n6940), .Y(REGFILE_SIM_reg_bank__abc_33898_n6944) );
  OR2X2 OR2X2_3727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6945), .B(REGFILE_SIM_reg_bank__abc_33898_n6946), .Y(REGFILE_SIM_reg_bank__abc_33898_n6947) );
  OR2X2 OR2X2_3728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6948), .B(REGFILE_SIM_reg_bank__abc_33898_n6949), .Y(REGFILE_SIM_reg_bank__abc_33898_n6950) );
  OR2X2 OR2X2_3729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6947), .B(REGFILE_SIM_reg_bank__abc_33898_n6950), .Y(REGFILE_SIM_reg_bank__abc_33898_n6951) );
  OR2X2 OR2X2_373 ( .A(_abc_43815_n1694), .B(pc_q_9_), .Y(_abc_43815_n1730) );
  OR2X2 OR2X2_3730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6944), .B(REGFILE_SIM_reg_bank__abc_33898_n6951), .Y(REGFILE_SIM_reg_bank__abc_33898_n6952) );
  OR2X2 OR2X2_3731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6953), .B(REGFILE_SIM_reg_bank__abc_33898_n6954), .Y(REGFILE_SIM_reg_bank__abc_33898_n6955) );
  OR2X2 OR2X2_3732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6956), .B(REGFILE_SIM_reg_bank__abc_33898_n6957), .Y(REGFILE_SIM_reg_bank__abc_33898_n6958) );
  OR2X2 OR2X2_3733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6955), .B(REGFILE_SIM_reg_bank__abc_33898_n6958), .Y(REGFILE_SIM_reg_bank__abc_33898_n6959) );
  OR2X2 OR2X2_3734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6960), .B(REGFILE_SIM_reg_bank__abc_33898_n6961), .Y(REGFILE_SIM_reg_bank__abc_33898_n6962) );
  OR2X2 OR2X2_3735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6963), .B(REGFILE_SIM_reg_bank__abc_33898_n6964), .Y(REGFILE_SIM_reg_bank__abc_33898_n6965) );
  OR2X2 OR2X2_3736 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6965), .B(REGFILE_SIM_reg_bank__abc_33898_n6962), .Y(REGFILE_SIM_reg_bank__abc_33898_n6966) );
  OR2X2 OR2X2_3737 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6959), .B(REGFILE_SIM_reg_bank__abc_33898_n6966), .Y(REGFILE_SIM_reg_bank__abc_33898_n6967) );
  OR2X2 OR2X2_3738 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6952), .B(REGFILE_SIM_reg_bank__abc_33898_n6967), .Y(REGFILE_SIM_reg_bank__abc_33898_n6968) );
  OR2X2 OR2X2_3739 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6969), .B(REGFILE_SIM_reg_bank__abc_33898_n6970), .Y(REGFILE_SIM_reg_bank__abc_33898_n6971) );
  OR2X2 OR2X2_374 ( .A(_abc_43815_n1733), .B(_abc_43815_n1278_bF_buf0), .Y(_abc_43815_n1734) );
  OR2X2 OR2X2_3740 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6972), .B(REGFILE_SIM_reg_bank__abc_33898_n6973), .Y(REGFILE_SIM_reg_bank__abc_33898_n6974) );
  OR2X2 OR2X2_3741 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6971), .B(REGFILE_SIM_reg_bank__abc_33898_n6974), .Y(REGFILE_SIM_reg_bank__abc_33898_n6975) );
  OR2X2 OR2X2_3742 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6977), .B(REGFILE_SIM_reg_bank__abc_33898_n6978), .Y(REGFILE_SIM_reg_bank__abc_33898_n6979) );
  OR2X2 OR2X2_3743 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6979), .B(REGFILE_SIM_reg_bank__abc_33898_n6976), .Y(REGFILE_SIM_reg_bank__abc_33898_n6980) );
  OR2X2 OR2X2_3744 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6975), .B(REGFILE_SIM_reg_bank__abc_33898_n6980), .Y(REGFILE_SIM_reg_bank__abc_33898_n6981) );
  OR2X2 OR2X2_3745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6982), .B(REGFILE_SIM_reg_bank__abc_33898_n6983), .Y(REGFILE_SIM_reg_bank__abc_33898_n6984) );
  OR2X2 OR2X2_3746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6985), .B(REGFILE_SIM_reg_bank__abc_33898_n6986), .Y(REGFILE_SIM_reg_bank__abc_33898_n6987) );
  OR2X2 OR2X2_3747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6987), .B(REGFILE_SIM_reg_bank__abc_33898_n6984), .Y(REGFILE_SIM_reg_bank__abc_33898_n6988) );
  OR2X2 OR2X2_3748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6989), .B(REGFILE_SIM_reg_bank__abc_33898_n6990), .Y(REGFILE_SIM_reg_bank__abc_33898_n6991) );
  OR2X2 OR2X2_3749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6992), .B(REGFILE_SIM_reg_bank__abc_33898_n6993), .Y(REGFILE_SIM_reg_bank__abc_33898_n6994) );
  OR2X2 OR2X2_375 ( .A(_abc_43815_n1737), .B(_abc_43815_n1736), .Y(_abc_43815_n1738_1) );
  OR2X2 OR2X2_3750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6991), .B(REGFILE_SIM_reg_bank__abc_33898_n6994), .Y(REGFILE_SIM_reg_bank__abc_33898_n6995) );
  OR2X2 OR2X2_3751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6988), .B(REGFILE_SIM_reg_bank__abc_33898_n6995), .Y(REGFILE_SIM_reg_bank__abc_33898_n6996) );
  OR2X2 OR2X2_3752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6996), .B(REGFILE_SIM_reg_bank__abc_33898_n6981), .Y(REGFILE_SIM_reg_bank__abc_33898_n6997) );
  OR2X2 OR2X2_3753 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6968), .B(REGFILE_SIM_reg_bank__abc_33898_n6997), .Y(REGFILE_SIM_reg_bank_reg_rb_o_22_) );
  OR2X2 OR2X2_3754 ( .A(REGFILE_SIM_reg_bank__abc_33898_n6999), .B(REGFILE_SIM_reg_bank__abc_33898_n7000), .Y(REGFILE_SIM_reg_bank__abc_33898_n7001) );
  OR2X2 OR2X2_3755 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7002), .B(REGFILE_SIM_reg_bank__abc_33898_n7003), .Y(REGFILE_SIM_reg_bank__abc_33898_n7004) );
  OR2X2 OR2X2_3756 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7004), .B(REGFILE_SIM_reg_bank__abc_33898_n7001), .Y(REGFILE_SIM_reg_bank__abc_33898_n7005) );
  OR2X2 OR2X2_3757 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7006), .B(REGFILE_SIM_reg_bank__abc_33898_n7007), .Y(REGFILE_SIM_reg_bank__abc_33898_n7008) );
  OR2X2 OR2X2_3758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7009), .B(REGFILE_SIM_reg_bank__abc_33898_n7010), .Y(REGFILE_SIM_reg_bank__abc_33898_n7011) );
  OR2X2 OR2X2_3759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7008), .B(REGFILE_SIM_reg_bank__abc_33898_n7011), .Y(REGFILE_SIM_reg_bank__abc_33898_n7012) );
  OR2X2 OR2X2_376 ( .A(alu_op_r_5_), .B(pc_q_9_), .Y(_abc_43815_n1744) );
  OR2X2 OR2X2_3760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7005), .B(REGFILE_SIM_reg_bank__abc_33898_n7012), .Y(REGFILE_SIM_reg_bank__abc_33898_n7013) );
  OR2X2 OR2X2_3761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7014), .B(REGFILE_SIM_reg_bank__abc_33898_n7015), .Y(REGFILE_SIM_reg_bank__abc_33898_n7016) );
  OR2X2 OR2X2_3762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7017), .B(REGFILE_SIM_reg_bank__abc_33898_n7018), .Y(REGFILE_SIM_reg_bank__abc_33898_n7019) );
  OR2X2 OR2X2_3763 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7016), .B(REGFILE_SIM_reg_bank__abc_33898_n7019), .Y(REGFILE_SIM_reg_bank__abc_33898_n7020) );
  OR2X2 OR2X2_3764 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7021), .B(REGFILE_SIM_reg_bank__abc_33898_n7022), .Y(REGFILE_SIM_reg_bank__abc_33898_n7023) );
  OR2X2 OR2X2_3765 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7024), .B(REGFILE_SIM_reg_bank__abc_33898_n7025), .Y(REGFILE_SIM_reg_bank__abc_33898_n7026) );
  OR2X2 OR2X2_3766 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7026), .B(REGFILE_SIM_reg_bank__abc_33898_n7023), .Y(REGFILE_SIM_reg_bank__abc_33898_n7027) );
  OR2X2 OR2X2_3767 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7020), .B(REGFILE_SIM_reg_bank__abc_33898_n7027), .Y(REGFILE_SIM_reg_bank__abc_33898_n7028) );
  OR2X2 OR2X2_3768 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7013), .B(REGFILE_SIM_reg_bank__abc_33898_n7028), .Y(REGFILE_SIM_reg_bank__abc_33898_n7029) );
  OR2X2 OR2X2_3769 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7030), .B(REGFILE_SIM_reg_bank__abc_33898_n7031), .Y(REGFILE_SIM_reg_bank__abc_33898_n7032) );
  OR2X2 OR2X2_377 ( .A(_abc_43815_n1750_1), .B(inst_trap_w), .Y(_abc_43815_n1751) );
  OR2X2 OR2X2_3770 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7033), .B(REGFILE_SIM_reg_bank__abc_33898_n7034), .Y(REGFILE_SIM_reg_bank__abc_33898_n7035) );
  OR2X2 OR2X2_3771 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7032), .B(REGFILE_SIM_reg_bank__abc_33898_n7035), .Y(REGFILE_SIM_reg_bank__abc_33898_n7036) );
  OR2X2 OR2X2_3772 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7038), .B(REGFILE_SIM_reg_bank__abc_33898_n7039), .Y(REGFILE_SIM_reg_bank__abc_33898_n7040) );
  OR2X2 OR2X2_3773 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7040), .B(REGFILE_SIM_reg_bank__abc_33898_n7037), .Y(REGFILE_SIM_reg_bank__abc_33898_n7041) );
  OR2X2 OR2X2_3774 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7036), .B(REGFILE_SIM_reg_bank__abc_33898_n7041), .Y(REGFILE_SIM_reg_bank__abc_33898_n7042) );
  OR2X2 OR2X2_3775 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7043), .B(REGFILE_SIM_reg_bank__abc_33898_n7044), .Y(REGFILE_SIM_reg_bank__abc_33898_n7045) );
  OR2X2 OR2X2_3776 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7046), .B(REGFILE_SIM_reg_bank__abc_33898_n7047), .Y(REGFILE_SIM_reg_bank__abc_33898_n7048) );
  OR2X2 OR2X2_3777 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7048), .B(REGFILE_SIM_reg_bank__abc_33898_n7045), .Y(REGFILE_SIM_reg_bank__abc_33898_n7049) );
  OR2X2 OR2X2_3778 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7050), .B(REGFILE_SIM_reg_bank__abc_33898_n7051), .Y(REGFILE_SIM_reg_bank__abc_33898_n7052) );
  OR2X2 OR2X2_3779 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7053), .B(REGFILE_SIM_reg_bank__abc_33898_n7054), .Y(REGFILE_SIM_reg_bank__abc_33898_n7055) );
  OR2X2 OR2X2_378 ( .A(_abc_43815_n1751), .B(_abc_43815_n1749), .Y(_abc_43815_n1752) );
  OR2X2 OR2X2_3780 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7052), .B(REGFILE_SIM_reg_bank__abc_33898_n7055), .Y(REGFILE_SIM_reg_bank__abc_33898_n7056) );
  OR2X2 OR2X2_3781 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7049), .B(REGFILE_SIM_reg_bank__abc_33898_n7056), .Y(REGFILE_SIM_reg_bank__abc_33898_n7057) );
  OR2X2 OR2X2_3782 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7057), .B(REGFILE_SIM_reg_bank__abc_33898_n7042), .Y(REGFILE_SIM_reg_bank__abc_33898_n7058) );
  OR2X2 OR2X2_3783 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7029), .B(REGFILE_SIM_reg_bank__abc_33898_n7058), .Y(REGFILE_SIM_reg_bank_reg_rb_o_23_) );
  OR2X2 OR2X2_3784 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7060), .B(REGFILE_SIM_reg_bank__abc_33898_n7061), .Y(REGFILE_SIM_reg_bank__abc_33898_n7062) );
  OR2X2 OR2X2_3785 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7063), .B(REGFILE_SIM_reg_bank__abc_33898_n7064), .Y(REGFILE_SIM_reg_bank__abc_33898_n7065) );
  OR2X2 OR2X2_3786 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7065), .B(REGFILE_SIM_reg_bank__abc_33898_n7062), .Y(REGFILE_SIM_reg_bank__abc_33898_n7066) );
  OR2X2 OR2X2_3787 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7067), .B(REGFILE_SIM_reg_bank__abc_33898_n7068), .Y(REGFILE_SIM_reg_bank__abc_33898_n7069) );
  OR2X2 OR2X2_3788 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7070), .B(REGFILE_SIM_reg_bank__abc_33898_n7071), .Y(REGFILE_SIM_reg_bank__abc_33898_n7072) );
  OR2X2 OR2X2_3789 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7069), .B(REGFILE_SIM_reg_bank__abc_33898_n7072), .Y(REGFILE_SIM_reg_bank__abc_33898_n7073) );
  OR2X2 OR2X2_379 ( .A(_abc_43815_n1428_bF_buf4), .B(_abc_43815_n1754), .Y(_abc_43815_n1755) );
  OR2X2 OR2X2_3790 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7066), .B(REGFILE_SIM_reg_bank__abc_33898_n7073), .Y(REGFILE_SIM_reg_bank__abc_33898_n7074) );
  OR2X2 OR2X2_3791 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7075), .B(REGFILE_SIM_reg_bank__abc_33898_n7076), .Y(REGFILE_SIM_reg_bank__abc_33898_n7077) );
  OR2X2 OR2X2_3792 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7078), .B(REGFILE_SIM_reg_bank__abc_33898_n7079), .Y(REGFILE_SIM_reg_bank__abc_33898_n7080) );
  OR2X2 OR2X2_3793 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7077), .B(REGFILE_SIM_reg_bank__abc_33898_n7080), .Y(REGFILE_SIM_reg_bank__abc_33898_n7081) );
  OR2X2 OR2X2_3794 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7082), .B(REGFILE_SIM_reg_bank__abc_33898_n7083), .Y(REGFILE_SIM_reg_bank__abc_33898_n7084) );
  OR2X2 OR2X2_3795 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7085), .B(REGFILE_SIM_reg_bank__abc_33898_n7086), .Y(REGFILE_SIM_reg_bank__abc_33898_n7087) );
  OR2X2 OR2X2_3796 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7087), .B(REGFILE_SIM_reg_bank__abc_33898_n7084), .Y(REGFILE_SIM_reg_bank__abc_33898_n7088) );
  OR2X2 OR2X2_3797 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7081), .B(REGFILE_SIM_reg_bank__abc_33898_n7088), .Y(REGFILE_SIM_reg_bank__abc_33898_n7089) );
  OR2X2 OR2X2_3798 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7074), .B(REGFILE_SIM_reg_bank__abc_33898_n7089), .Y(REGFILE_SIM_reg_bank__abc_33898_n7090) );
  OR2X2 OR2X2_3799 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7091), .B(REGFILE_SIM_reg_bank__abc_33898_n7092), .Y(REGFILE_SIM_reg_bank__abc_33898_n7093) );
  OR2X2 OR2X2_38 ( .A(_abc_43815_n767), .B(_abc_43815_n768), .Y(_abc_43815_n769) );
  OR2X2 OR2X2_380 ( .A(_abc_43815_n1753_1), .B(_abc_43815_n1755), .Y(_abc_43815_n1756) );
  OR2X2 OR2X2_3800 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7094), .B(REGFILE_SIM_reg_bank__abc_33898_n7095), .Y(REGFILE_SIM_reg_bank__abc_33898_n7096) );
  OR2X2 OR2X2_3801 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7093), .B(REGFILE_SIM_reg_bank__abc_33898_n7096), .Y(REGFILE_SIM_reg_bank__abc_33898_n7097) );
  OR2X2 OR2X2_3802 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7099), .B(REGFILE_SIM_reg_bank__abc_33898_n7100), .Y(REGFILE_SIM_reg_bank__abc_33898_n7101) );
  OR2X2 OR2X2_3803 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7101), .B(REGFILE_SIM_reg_bank__abc_33898_n7098), .Y(REGFILE_SIM_reg_bank__abc_33898_n7102) );
  OR2X2 OR2X2_3804 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7097), .B(REGFILE_SIM_reg_bank__abc_33898_n7102), .Y(REGFILE_SIM_reg_bank__abc_33898_n7103) );
  OR2X2 OR2X2_3805 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7104), .B(REGFILE_SIM_reg_bank__abc_33898_n7105), .Y(REGFILE_SIM_reg_bank__abc_33898_n7106) );
  OR2X2 OR2X2_3806 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7107), .B(REGFILE_SIM_reg_bank__abc_33898_n7108), .Y(REGFILE_SIM_reg_bank__abc_33898_n7109) );
  OR2X2 OR2X2_3807 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7109), .B(REGFILE_SIM_reg_bank__abc_33898_n7106), .Y(REGFILE_SIM_reg_bank__abc_33898_n7110) );
  OR2X2 OR2X2_3808 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7111), .B(REGFILE_SIM_reg_bank__abc_33898_n7112), .Y(REGFILE_SIM_reg_bank__abc_33898_n7113) );
  OR2X2 OR2X2_3809 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7114), .B(REGFILE_SIM_reg_bank__abc_33898_n7115), .Y(REGFILE_SIM_reg_bank__abc_33898_n7116) );
  OR2X2 OR2X2_381 ( .A(_abc_43815_n1431_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_43815_n1757) );
  OR2X2 OR2X2_3810 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7113), .B(REGFILE_SIM_reg_bank__abc_33898_n7116), .Y(REGFILE_SIM_reg_bank__abc_33898_n7117) );
  OR2X2 OR2X2_3811 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7110), .B(REGFILE_SIM_reg_bank__abc_33898_n7117), .Y(REGFILE_SIM_reg_bank__abc_33898_n7118) );
  OR2X2 OR2X2_3812 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7118), .B(REGFILE_SIM_reg_bank__abc_33898_n7103), .Y(REGFILE_SIM_reg_bank__abc_33898_n7119) );
  OR2X2 OR2X2_3813 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7090), .B(REGFILE_SIM_reg_bank__abc_33898_n7119), .Y(REGFILE_SIM_reg_bank_reg_rb_o_24_) );
  OR2X2 OR2X2_3814 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7121), .B(REGFILE_SIM_reg_bank__abc_33898_n7122), .Y(REGFILE_SIM_reg_bank__abc_33898_n7123) );
  OR2X2 OR2X2_3815 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7124), .B(REGFILE_SIM_reg_bank__abc_33898_n7125), .Y(REGFILE_SIM_reg_bank__abc_33898_n7126) );
  OR2X2 OR2X2_3816 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7126), .B(REGFILE_SIM_reg_bank__abc_33898_n7123), .Y(REGFILE_SIM_reg_bank__abc_33898_n7127) );
  OR2X2 OR2X2_3817 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7128), .B(REGFILE_SIM_reg_bank__abc_33898_n7129), .Y(REGFILE_SIM_reg_bank__abc_33898_n7130) );
  OR2X2 OR2X2_3818 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7131), .B(REGFILE_SIM_reg_bank__abc_33898_n7132), .Y(REGFILE_SIM_reg_bank__abc_33898_n7133) );
  OR2X2 OR2X2_3819 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7130), .B(REGFILE_SIM_reg_bank__abc_33898_n7133), .Y(REGFILE_SIM_reg_bank__abc_33898_n7134) );
  OR2X2 OR2X2_382 ( .A(_abc_43815_n1759), .B(_abc_43815_n1760), .Y(_abc_43815_n1761) );
  OR2X2 OR2X2_3820 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7127), .B(REGFILE_SIM_reg_bank__abc_33898_n7134), .Y(REGFILE_SIM_reg_bank__abc_33898_n7135) );
  OR2X2 OR2X2_3821 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7136), .B(REGFILE_SIM_reg_bank__abc_33898_n7137), .Y(REGFILE_SIM_reg_bank__abc_33898_n7138) );
  OR2X2 OR2X2_3822 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7139), .B(REGFILE_SIM_reg_bank__abc_33898_n7140), .Y(REGFILE_SIM_reg_bank__abc_33898_n7141) );
  OR2X2 OR2X2_3823 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7138), .B(REGFILE_SIM_reg_bank__abc_33898_n7141), .Y(REGFILE_SIM_reg_bank__abc_33898_n7142) );
  OR2X2 OR2X2_3824 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7143), .B(REGFILE_SIM_reg_bank__abc_33898_n7144), .Y(REGFILE_SIM_reg_bank__abc_33898_n7145) );
  OR2X2 OR2X2_3825 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7146), .B(REGFILE_SIM_reg_bank__abc_33898_n7147), .Y(REGFILE_SIM_reg_bank__abc_33898_n7148) );
  OR2X2 OR2X2_3826 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7148), .B(REGFILE_SIM_reg_bank__abc_33898_n7145), .Y(REGFILE_SIM_reg_bank__abc_33898_n7149) );
  OR2X2 OR2X2_3827 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7142), .B(REGFILE_SIM_reg_bank__abc_33898_n7149), .Y(REGFILE_SIM_reg_bank__abc_33898_n7150) );
  OR2X2 OR2X2_3828 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7135), .B(REGFILE_SIM_reg_bank__abc_33898_n7150), .Y(REGFILE_SIM_reg_bank__abc_33898_n7151) );
  OR2X2 OR2X2_3829 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7152), .B(REGFILE_SIM_reg_bank__abc_33898_n7153), .Y(REGFILE_SIM_reg_bank__abc_33898_n7154) );
  OR2X2 OR2X2_383 ( .A(_abc_43815_n1762), .B(_abc_43815_n1739_1), .Y(_abc_43815_n1763) );
  OR2X2 OR2X2_3830 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7155), .B(REGFILE_SIM_reg_bank__abc_33898_n7156), .Y(REGFILE_SIM_reg_bank__abc_33898_n7157) );
  OR2X2 OR2X2_3831 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7154), .B(REGFILE_SIM_reg_bank__abc_33898_n7157), .Y(REGFILE_SIM_reg_bank__abc_33898_n7158) );
  OR2X2 OR2X2_3832 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7160), .B(REGFILE_SIM_reg_bank__abc_33898_n7161), .Y(REGFILE_SIM_reg_bank__abc_33898_n7162) );
  OR2X2 OR2X2_3833 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7162), .B(REGFILE_SIM_reg_bank__abc_33898_n7159), .Y(REGFILE_SIM_reg_bank__abc_33898_n7163) );
  OR2X2 OR2X2_3834 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7158), .B(REGFILE_SIM_reg_bank__abc_33898_n7163), .Y(REGFILE_SIM_reg_bank__abc_33898_n7164) );
  OR2X2 OR2X2_3835 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7165), .B(REGFILE_SIM_reg_bank__abc_33898_n7166), .Y(REGFILE_SIM_reg_bank__abc_33898_n7167) );
  OR2X2 OR2X2_3836 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7168), .B(REGFILE_SIM_reg_bank__abc_33898_n7169), .Y(REGFILE_SIM_reg_bank__abc_33898_n7170) );
  OR2X2 OR2X2_3837 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7170), .B(REGFILE_SIM_reg_bank__abc_33898_n7167), .Y(REGFILE_SIM_reg_bank__abc_33898_n7171) );
  OR2X2 OR2X2_3838 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7172), .B(REGFILE_SIM_reg_bank__abc_33898_n7173), .Y(REGFILE_SIM_reg_bank__abc_33898_n7174) );
  OR2X2 OR2X2_3839 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7175), .B(REGFILE_SIM_reg_bank__abc_33898_n7176), .Y(REGFILE_SIM_reg_bank__abc_33898_n7177) );
  OR2X2 OR2X2_384 ( .A(_abc_43815_n1764), .B(_abc_43815_n1735), .Y(_abc_43815_n1765) );
  OR2X2 OR2X2_3840 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7174), .B(REGFILE_SIM_reg_bank__abc_33898_n7177), .Y(REGFILE_SIM_reg_bank__abc_33898_n7178) );
  OR2X2 OR2X2_3841 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7171), .B(REGFILE_SIM_reg_bank__abc_33898_n7178), .Y(REGFILE_SIM_reg_bank__abc_33898_n7179) );
  OR2X2 OR2X2_3842 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7179), .B(REGFILE_SIM_reg_bank__abc_33898_n7164), .Y(REGFILE_SIM_reg_bank__abc_33898_n7180) );
  OR2X2 OR2X2_3843 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7151), .B(REGFILE_SIM_reg_bank__abc_33898_n7180), .Y(REGFILE_SIM_reg_bank_reg_rb_o_25_) );
  OR2X2 OR2X2_3844 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7182), .B(REGFILE_SIM_reg_bank__abc_33898_n7183), .Y(REGFILE_SIM_reg_bank__abc_33898_n7184) );
  OR2X2 OR2X2_3845 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7185), .B(REGFILE_SIM_reg_bank__abc_33898_n7186), .Y(REGFILE_SIM_reg_bank__abc_33898_n7187) );
  OR2X2 OR2X2_3846 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7187), .B(REGFILE_SIM_reg_bank__abc_33898_n7184), .Y(REGFILE_SIM_reg_bank__abc_33898_n7188) );
  OR2X2 OR2X2_3847 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7189), .B(REGFILE_SIM_reg_bank__abc_33898_n7190), .Y(REGFILE_SIM_reg_bank__abc_33898_n7191) );
  OR2X2 OR2X2_3848 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7192), .B(REGFILE_SIM_reg_bank__abc_33898_n7193), .Y(REGFILE_SIM_reg_bank__abc_33898_n7194) );
  OR2X2 OR2X2_3849 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7191), .B(REGFILE_SIM_reg_bank__abc_33898_n7194), .Y(REGFILE_SIM_reg_bank__abc_33898_n7195) );
  OR2X2 OR2X2_385 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_9_), .Y(_abc_43815_n1766) );
  OR2X2 OR2X2_3850 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7188), .B(REGFILE_SIM_reg_bank__abc_33898_n7195), .Y(REGFILE_SIM_reg_bank__abc_33898_n7196) );
  OR2X2 OR2X2_3851 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7197), .B(REGFILE_SIM_reg_bank__abc_33898_n7198), .Y(REGFILE_SIM_reg_bank__abc_33898_n7199) );
  OR2X2 OR2X2_3852 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7200), .B(REGFILE_SIM_reg_bank__abc_33898_n7201), .Y(REGFILE_SIM_reg_bank__abc_33898_n7202) );
  OR2X2 OR2X2_3853 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7199), .B(REGFILE_SIM_reg_bank__abc_33898_n7202), .Y(REGFILE_SIM_reg_bank__abc_33898_n7203) );
  OR2X2 OR2X2_3854 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7204), .B(REGFILE_SIM_reg_bank__abc_33898_n7205), .Y(REGFILE_SIM_reg_bank__abc_33898_n7206) );
  OR2X2 OR2X2_3855 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7207), .B(REGFILE_SIM_reg_bank__abc_33898_n7208), .Y(REGFILE_SIM_reg_bank__abc_33898_n7209) );
  OR2X2 OR2X2_3856 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7209), .B(REGFILE_SIM_reg_bank__abc_33898_n7206), .Y(REGFILE_SIM_reg_bank__abc_33898_n7210) );
  OR2X2 OR2X2_3857 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7203), .B(REGFILE_SIM_reg_bank__abc_33898_n7210), .Y(REGFILE_SIM_reg_bank__abc_33898_n7211) );
  OR2X2 OR2X2_3858 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7196), .B(REGFILE_SIM_reg_bank__abc_33898_n7211), .Y(REGFILE_SIM_reg_bank__abc_33898_n7212) );
  OR2X2 OR2X2_3859 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7213), .B(REGFILE_SIM_reg_bank__abc_33898_n7214), .Y(REGFILE_SIM_reg_bank__abc_33898_n7215) );
  OR2X2 OR2X2_386 ( .A(_abc_43815_n1731), .B(pc_q_10_), .Y(_abc_43815_n1769_1) );
  OR2X2 OR2X2_3860 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7216), .B(REGFILE_SIM_reg_bank__abc_33898_n7217), .Y(REGFILE_SIM_reg_bank__abc_33898_n7218) );
  OR2X2 OR2X2_3861 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7215), .B(REGFILE_SIM_reg_bank__abc_33898_n7218), .Y(REGFILE_SIM_reg_bank__abc_33898_n7219) );
  OR2X2 OR2X2_3862 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7221), .B(REGFILE_SIM_reg_bank__abc_33898_n7222), .Y(REGFILE_SIM_reg_bank__abc_33898_n7223) );
  OR2X2 OR2X2_3863 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7223), .B(REGFILE_SIM_reg_bank__abc_33898_n7220), .Y(REGFILE_SIM_reg_bank__abc_33898_n7224) );
  OR2X2 OR2X2_3864 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7219), .B(REGFILE_SIM_reg_bank__abc_33898_n7224), .Y(REGFILE_SIM_reg_bank__abc_33898_n7225) );
  OR2X2 OR2X2_3865 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7226), .B(REGFILE_SIM_reg_bank__abc_33898_n7227), .Y(REGFILE_SIM_reg_bank__abc_33898_n7228) );
  OR2X2 OR2X2_3866 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7229), .B(REGFILE_SIM_reg_bank__abc_33898_n7230), .Y(REGFILE_SIM_reg_bank__abc_33898_n7231) );
  OR2X2 OR2X2_3867 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7231), .B(REGFILE_SIM_reg_bank__abc_33898_n7228), .Y(REGFILE_SIM_reg_bank__abc_33898_n7232) );
  OR2X2 OR2X2_3868 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7233), .B(REGFILE_SIM_reg_bank__abc_33898_n7234), .Y(REGFILE_SIM_reg_bank__abc_33898_n7235) );
  OR2X2 OR2X2_3869 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7236), .B(REGFILE_SIM_reg_bank__abc_33898_n7237), .Y(REGFILE_SIM_reg_bank__abc_33898_n7238) );
  OR2X2 OR2X2_387 ( .A(_abc_43815_n1772), .B(_abc_43815_n1278_bF_buf7), .Y(_abc_43815_n1773) );
  OR2X2 OR2X2_3870 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7235), .B(REGFILE_SIM_reg_bank__abc_33898_n7238), .Y(REGFILE_SIM_reg_bank__abc_33898_n7239) );
  OR2X2 OR2X2_3871 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7232), .B(REGFILE_SIM_reg_bank__abc_33898_n7239), .Y(REGFILE_SIM_reg_bank__abc_33898_n7240) );
  OR2X2 OR2X2_3872 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7240), .B(REGFILE_SIM_reg_bank__abc_33898_n7225), .Y(REGFILE_SIM_reg_bank__abc_33898_n7241) );
  OR2X2 OR2X2_3873 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7212), .B(REGFILE_SIM_reg_bank__abc_33898_n7241), .Y(REGFILE_SIM_reg_bank_reg_rb_o_26_) );
  OR2X2 OR2X2_3874 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7243), .B(REGFILE_SIM_reg_bank__abc_33898_n7244), .Y(REGFILE_SIM_reg_bank__abc_33898_n7245) );
  OR2X2 OR2X2_3875 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7246), .B(REGFILE_SIM_reg_bank__abc_33898_n7247), .Y(REGFILE_SIM_reg_bank__abc_33898_n7248) );
  OR2X2 OR2X2_3876 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7248), .B(REGFILE_SIM_reg_bank__abc_33898_n7245), .Y(REGFILE_SIM_reg_bank__abc_33898_n7249) );
  OR2X2 OR2X2_3877 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7250), .B(REGFILE_SIM_reg_bank__abc_33898_n7251), .Y(REGFILE_SIM_reg_bank__abc_33898_n7252) );
  OR2X2 OR2X2_3878 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7253), .B(REGFILE_SIM_reg_bank__abc_33898_n7254), .Y(REGFILE_SIM_reg_bank__abc_33898_n7255) );
  OR2X2 OR2X2_3879 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7252), .B(REGFILE_SIM_reg_bank__abc_33898_n7255), .Y(REGFILE_SIM_reg_bank__abc_33898_n7256) );
  OR2X2 OR2X2_388 ( .A(_abc_43815_n1776), .B(_abc_43815_n1775_1), .Y(_abc_43815_n1777) );
  OR2X2 OR2X2_3880 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7249), .B(REGFILE_SIM_reg_bank__abc_33898_n7256), .Y(REGFILE_SIM_reg_bank__abc_33898_n7257) );
  OR2X2 OR2X2_3881 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7258), .B(REGFILE_SIM_reg_bank__abc_33898_n7259), .Y(REGFILE_SIM_reg_bank__abc_33898_n7260) );
  OR2X2 OR2X2_3882 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7261), .B(REGFILE_SIM_reg_bank__abc_33898_n7262), .Y(REGFILE_SIM_reg_bank__abc_33898_n7263) );
  OR2X2 OR2X2_3883 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7260), .B(REGFILE_SIM_reg_bank__abc_33898_n7263), .Y(REGFILE_SIM_reg_bank__abc_33898_n7264) );
  OR2X2 OR2X2_3884 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7265), .B(REGFILE_SIM_reg_bank__abc_33898_n7266), .Y(REGFILE_SIM_reg_bank__abc_33898_n7267) );
  OR2X2 OR2X2_3885 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7268), .B(REGFILE_SIM_reg_bank__abc_33898_n7269), .Y(REGFILE_SIM_reg_bank__abc_33898_n7270) );
  OR2X2 OR2X2_3886 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7270), .B(REGFILE_SIM_reg_bank__abc_33898_n7267), .Y(REGFILE_SIM_reg_bank__abc_33898_n7271) );
  OR2X2 OR2X2_3887 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7264), .B(REGFILE_SIM_reg_bank__abc_33898_n7271), .Y(REGFILE_SIM_reg_bank__abc_33898_n7272) );
  OR2X2 OR2X2_3888 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7257), .B(REGFILE_SIM_reg_bank__abc_33898_n7272), .Y(REGFILE_SIM_reg_bank__abc_33898_n7273) );
  OR2X2 OR2X2_3889 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7274), .B(REGFILE_SIM_reg_bank__abc_33898_n7275), .Y(REGFILE_SIM_reg_bank__abc_33898_n7276) );
  OR2X2 OR2X2_389 ( .A(alu_op_r_6_), .B(pc_q_10_), .Y(_abc_43815_n1780) );
  OR2X2 OR2X2_3890 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7277), .B(REGFILE_SIM_reg_bank__abc_33898_n7278), .Y(REGFILE_SIM_reg_bank__abc_33898_n7279) );
  OR2X2 OR2X2_3891 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7276), .B(REGFILE_SIM_reg_bank__abc_33898_n7279), .Y(REGFILE_SIM_reg_bank__abc_33898_n7280) );
  OR2X2 OR2X2_3892 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7282), .B(REGFILE_SIM_reg_bank__abc_33898_n7283), .Y(REGFILE_SIM_reg_bank__abc_33898_n7284) );
  OR2X2 OR2X2_3893 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7284), .B(REGFILE_SIM_reg_bank__abc_33898_n7281), .Y(REGFILE_SIM_reg_bank__abc_33898_n7285) );
  OR2X2 OR2X2_3894 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7280), .B(REGFILE_SIM_reg_bank__abc_33898_n7285), .Y(REGFILE_SIM_reg_bank__abc_33898_n7286) );
  OR2X2 OR2X2_3895 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7287), .B(REGFILE_SIM_reg_bank__abc_33898_n7288), .Y(REGFILE_SIM_reg_bank__abc_33898_n7289) );
  OR2X2 OR2X2_3896 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7290), .B(REGFILE_SIM_reg_bank__abc_33898_n7291), .Y(REGFILE_SIM_reg_bank__abc_33898_n7292) );
  OR2X2 OR2X2_3897 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7292), .B(REGFILE_SIM_reg_bank__abc_33898_n7289), .Y(REGFILE_SIM_reg_bank__abc_33898_n7293) );
  OR2X2 OR2X2_3898 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7294), .B(REGFILE_SIM_reg_bank__abc_33898_n7295), .Y(REGFILE_SIM_reg_bank__abc_33898_n7296) );
  OR2X2 OR2X2_3899 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7297), .B(REGFILE_SIM_reg_bank__abc_33898_n7298), .Y(REGFILE_SIM_reg_bank__abc_33898_n7299) );
  OR2X2 OR2X2_39 ( .A(_abc_43815_n770), .B(_abc_43815_n771), .Y(_abc_43815_n772) );
  OR2X2 OR2X2_390 ( .A(_abc_43815_n1748), .B(_abc_43815_n1706_1), .Y(_abc_43815_n1784) );
  OR2X2 OR2X2_3900 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7296), .B(REGFILE_SIM_reg_bank__abc_33898_n7299), .Y(REGFILE_SIM_reg_bank__abc_33898_n7300) );
  OR2X2 OR2X2_3901 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7293), .B(REGFILE_SIM_reg_bank__abc_33898_n7300), .Y(REGFILE_SIM_reg_bank__abc_33898_n7301) );
  OR2X2 OR2X2_3902 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7301), .B(REGFILE_SIM_reg_bank__abc_33898_n7286), .Y(REGFILE_SIM_reg_bank__abc_33898_n7302) );
  OR2X2 OR2X2_3903 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7273), .B(REGFILE_SIM_reg_bank__abc_33898_n7302), .Y(REGFILE_SIM_reg_bank_reg_rb_o_27_) );
  OR2X2 OR2X2_3904 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7304), .B(REGFILE_SIM_reg_bank__abc_33898_n7305), .Y(REGFILE_SIM_reg_bank__abc_33898_n7306) );
  OR2X2 OR2X2_3905 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7307), .B(REGFILE_SIM_reg_bank__abc_33898_n7308), .Y(REGFILE_SIM_reg_bank__abc_33898_n7309) );
  OR2X2 OR2X2_3906 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7309), .B(REGFILE_SIM_reg_bank__abc_33898_n7306), .Y(REGFILE_SIM_reg_bank__abc_33898_n7310) );
  OR2X2 OR2X2_3907 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7311), .B(REGFILE_SIM_reg_bank__abc_33898_n7312), .Y(REGFILE_SIM_reg_bank__abc_33898_n7313) );
  OR2X2 OR2X2_3908 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7314), .B(REGFILE_SIM_reg_bank__abc_33898_n7315), .Y(REGFILE_SIM_reg_bank__abc_33898_n7316) );
  OR2X2 OR2X2_3909 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7313), .B(REGFILE_SIM_reg_bank__abc_33898_n7316), .Y(REGFILE_SIM_reg_bank__abc_33898_n7317) );
  OR2X2 OR2X2_391 ( .A(_abc_43815_n1788_1), .B(_abc_43815_n1786), .Y(_abc_43815_n1789) );
  OR2X2 OR2X2_3910 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7310), .B(REGFILE_SIM_reg_bank__abc_33898_n7317), .Y(REGFILE_SIM_reg_bank__abc_33898_n7318) );
  OR2X2 OR2X2_3911 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7319), .B(REGFILE_SIM_reg_bank__abc_33898_n7320), .Y(REGFILE_SIM_reg_bank__abc_33898_n7321) );
  OR2X2 OR2X2_3912 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7322), .B(REGFILE_SIM_reg_bank__abc_33898_n7323), .Y(REGFILE_SIM_reg_bank__abc_33898_n7324) );
  OR2X2 OR2X2_3913 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7321), .B(REGFILE_SIM_reg_bank__abc_33898_n7324), .Y(REGFILE_SIM_reg_bank__abc_33898_n7325) );
  OR2X2 OR2X2_3914 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7326), .B(REGFILE_SIM_reg_bank__abc_33898_n7327), .Y(REGFILE_SIM_reg_bank__abc_33898_n7328) );
  OR2X2 OR2X2_3915 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7329), .B(REGFILE_SIM_reg_bank__abc_33898_n7330), .Y(REGFILE_SIM_reg_bank__abc_33898_n7331) );
  OR2X2 OR2X2_3916 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7331), .B(REGFILE_SIM_reg_bank__abc_33898_n7328), .Y(REGFILE_SIM_reg_bank__abc_33898_n7332) );
  OR2X2 OR2X2_3917 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7325), .B(REGFILE_SIM_reg_bank__abc_33898_n7332), .Y(REGFILE_SIM_reg_bank__abc_33898_n7333) );
  OR2X2 OR2X2_3918 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7318), .B(REGFILE_SIM_reg_bank__abc_33898_n7333), .Y(REGFILE_SIM_reg_bank__abc_33898_n7334) );
  OR2X2 OR2X2_3919 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7335), .B(REGFILE_SIM_reg_bank__abc_33898_n7336), .Y(REGFILE_SIM_reg_bank__abc_33898_n7337) );
  OR2X2 OR2X2_392 ( .A(_abc_43815_n1789), .B(_abc_43815_n1783), .Y(_abc_43815_n1792) );
  OR2X2 OR2X2_3920 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7338), .B(REGFILE_SIM_reg_bank__abc_33898_n7339), .Y(REGFILE_SIM_reg_bank__abc_33898_n7340) );
  OR2X2 OR2X2_3921 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7337), .B(REGFILE_SIM_reg_bank__abc_33898_n7340), .Y(REGFILE_SIM_reg_bank__abc_33898_n7341) );
  OR2X2 OR2X2_3922 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7343), .B(REGFILE_SIM_reg_bank__abc_33898_n7344), .Y(REGFILE_SIM_reg_bank__abc_33898_n7345) );
  OR2X2 OR2X2_3923 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7345), .B(REGFILE_SIM_reg_bank__abc_33898_n7342), .Y(REGFILE_SIM_reg_bank__abc_33898_n7346) );
  OR2X2 OR2X2_3924 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7341), .B(REGFILE_SIM_reg_bank__abc_33898_n7346), .Y(REGFILE_SIM_reg_bank__abc_33898_n7347) );
  OR2X2 OR2X2_3925 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7348), .B(REGFILE_SIM_reg_bank__abc_33898_n7349), .Y(REGFILE_SIM_reg_bank__abc_33898_n7350) );
  OR2X2 OR2X2_3926 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7351), .B(REGFILE_SIM_reg_bank__abc_33898_n7352), .Y(REGFILE_SIM_reg_bank__abc_33898_n7353) );
  OR2X2 OR2X2_3927 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7353), .B(REGFILE_SIM_reg_bank__abc_33898_n7350), .Y(REGFILE_SIM_reg_bank__abc_33898_n7354) );
  OR2X2 OR2X2_3928 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7355), .B(REGFILE_SIM_reg_bank__abc_33898_n7356), .Y(REGFILE_SIM_reg_bank__abc_33898_n7357) );
  OR2X2 OR2X2_3929 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7358), .B(REGFILE_SIM_reg_bank__abc_33898_n7359), .Y(REGFILE_SIM_reg_bank__abc_33898_n7360) );
  OR2X2 OR2X2_393 ( .A(_abc_43815_n1793), .B(_abc_43815_n1779), .Y(_abc_43815_n1794_1) );
  OR2X2 OR2X2_3930 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7357), .B(REGFILE_SIM_reg_bank__abc_33898_n7360), .Y(REGFILE_SIM_reg_bank__abc_33898_n7361) );
  OR2X2 OR2X2_3931 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7354), .B(REGFILE_SIM_reg_bank__abc_33898_n7361), .Y(REGFILE_SIM_reg_bank__abc_33898_n7362) );
  OR2X2 OR2X2_3932 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7362), .B(REGFILE_SIM_reg_bank__abc_33898_n7347), .Y(REGFILE_SIM_reg_bank__abc_33898_n7363) );
  OR2X2 OR2X2_3933 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7334), .B(REGFILE_SIM_reg_bank__abc_33898_n7363), .Y(REGFILE_SIM_reg_bank_reg_rb_o_28_) );
  OR2X2 OR2X2_3934 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7365), .B(REGFILE_SIM_reg_bank__abc_33898_n7366), .Y(REGFILE_SIM_reg_bank__abc_33898_n7367) );
  OR2X2 OR2X2_3935 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7368), .B(REGFILE_SIM_reg_bank__abc_33898_n7369), .Y(REGFILE_SIM_reg_bank__abc_33898_n7370) );
  OR2X2 OR2X2_3936 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7370), .B(REGFILE_SIM_reg_bank__abc_33898_n7367), .Y(REGFILE_SIM_reg_bank__abc_33898_n7371) );
  OR2X2 OR2X2_3937 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7372), .B(REGFILE_SIM_reg_bank__abc_33898_n7373), .Y(REGFILE_SIM_reg_bank__abc_33898_n7374) );
  OR2X2 OR2X2_3938 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7375), .B(REGFILE_SIM_reg_bank__abc_33898_n7376), .Y(REGFILE_SIM_reg_bank__abc_33898_n7377) );
  OR2X2 OR2X2_3939 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7374), .B(REGFILE_SIM_reg_bank__abc_33898_n7377), .Y(REGFILE_SIM_reg_bank__abc_33898_n7378) );
  OR2X2 OR2X2_394 ( .A(_abc_43815_n1066), .B(epc_q_10_), .Y(_abc_43815_n1795) );
  OR2X2 OR2X2_3940 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7371), .B(REGFILE_SIM_reg_bank__abc_33898_n7378), .Y(REGFILE_SIM_reg_bank__abc_33898_n7379) );
  OR2X2 OR2X2_3941 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7380), .B(REGFILE_SIM_reg_bank__abc_33898_n7381), .Y(REGFILE_SIM_reg_bank__abc_33898_n7382) );
  OR2X2 OR2X2_3942 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7383), .B(REGFILE_SIM_reg_bank__abc_33898_n7384), .Y(REGFILE_SIM_reg_bank__abc_33898_n7385) );
  OR2X2 OR2X2_3943 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7382), .B(REGFILE_SIM_reg_bank__abc_33898_n7385), .Y(REGFILE_SIM_reg_bank__abc_33898_n7386) );
  OR2X2 OR2X2_3944 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7387), .B(REGFILE_SIM_reg_bank__abc_33898_n7388), .Y(REGFILE_SIM_reg_bank__abc_33898_n7389) );
  OR2X2 OR2X2_3945 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7390), .B(REGFILE_SIM_reg_bank__abc_33898_n7391), .Y(REGFILE_SIM_reg_bank__abc_33898_n7392) );
  OR2X2 OR2X2_3946 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7392), .B(REGFILE_SIM_reg_bank__abc_33898_n7389), .Y(REGFILE_SIM_reg_bank__abc_33898_n7393) );
  OR2X2 OR2X2_3947 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7386), .B(REGFILE_SIM_reg_bank__abc_33898_n7393), .Y(REGFILE_SIM_reg_bank__abc_33898_n7394) );
  OR2X2 OR2X2_3948 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7379), .B(REGFILE_SIM_reg_bank__abc_33898_n7394), .Y(REGFILE_SIM_reg_bank__abc_33898_n7395) );
  OR2X2 OR2X2_3949 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7396), .B(REGFILE_SIM_reg_bank__abc_33898_n7397), .Y(REGFILE_SIM_reg_bank__abc_33898_n7398) );
  OR2X2 OR2X2_395 ( .A(_abc_43815_n1473_bF_buf1), .B(_abc_43815_n1798), .Y(_abc_43815_n1799) );
  OR2X2 OR2X2_3950 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7399), .B(REGFILE_SIM_reg_bank__abc_33898_n7400), .Y(REGFILE_SIM_reg_bank__abc_33898_n7401) );
  OR2X2 OR2X2_3951 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7398), .B(REGFILE_SIM_reg_bank__abc_33898_n7401), .Y(REGFILE_SIM_reg_bank__abc_33898_n7402) );
  OR2X2 OR2X2_3952 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7404), .B(REGFILE_SIM_reg_bank__abc_33898_n7405), .Y(REGFILE_SIM_reg_bank__abc_33898_n7406) );
  OR2X2 OR2X2_3953 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7406), .B(REGFILE_SIM_reg_bank__abc_33898_n7403), .Y(REGFILE_SIM_reg_bank__abc_33898_n7407) );
  OR2X2 OR2X2_3954 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7402), .B(REGFILE_SIM_reg_bank__abc_33898_n7407), .Y(REGFILE_SIM_reg_bank__abc_33898_n7408) );
  OR2X2 OR2X2_3955 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7409), .B(REGFILE_SIM_reg_bank__abc_33898_n7410), .Y(REGFILE_SIM_reg_bank__abc_33898_n7411) );
  OR2X2 OR2X2_3956 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7412), .B(REGFILE_SIM_reg_bank__abc_33898_n7413), .Y(REGFILE_SIM_reg_bank__abc_33898_n7414) );
  OR2X2 OR2X2_3957 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7414), .B(REGFILE_SIM_reg_bank__abc_33898_n7411), .Y(REGFILE_SIM_reg_bank__abc_33898_n7415) );
  OR2X2 OR2X2_3958 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7416), .B(REGFILE_SIM_reg_bank__abc_33898_n7417), .Y(REGFILE_SIM_reg_bank__abc_33898_n7418) );
  OR2X2 OR2X2_3959 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7419), .B(REGFILE_SIM_reg_bank__abc_33898_n7420), .Y(REGFILE_SIM_reg_bank__abc_33898_n7421) );
  OR2X2 OR2X2_396 ( .A(_abc_43815_n1797_1), .B(_abc_43815_n1799), .Y(_abc_43815_n1800) );
  OR2X2 OR2X2_3960 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7418), .B(REGFILE_SIM_reg_bank__abc_33898_n7421), .Y(REGFILE_SIM_reg_bank__abc_33898_n7422) );
  OR2X2 OR2X2_3961 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7415), .B(REGFILE_SIM_reg_bank__abc_33898_n7422), .Y(REGFILE_SIM_reg_bank__abc_33898_n7423) );
  OR2X2 OR2X2_3962 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7423), .B(REGFILE_SIM_reg_bank__abc_33898_n7408), .Y(REGFILE_SIM_reg_bank__abc_33898_n7424) );
  OR2X2 OR2X2_3963 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7395), .B(REGFILE_SIM_reg_bank__abc_33898_n7424), .Y(REGFILE_SIM_reg_bank_reg_rb_o_29_) );
  OR2X2 OR2X2_3964 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7426), .B(REGFILE_SIM_reg_bank__abc_33898_n7427), .Y(REGFILE_SIM_reg_bank__abc_33898_n7428) );
  OR2X2 OR2X2_3965 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7429), .B(REGFILE_SIM_reg_bank__abc_33898_n7430), .Y(REGFILE_SIM_reg_bank__abc_33898_n7431) );
  OR2X2 OR2X2_3966 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7431), .B(REGFILE_SIM_reg_bank__abc_33898_n7428), .Y(REGFILE_SIM_reg_bank__abc_33898_n7432) );
  OR2X2 OR2X2_3967 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7433), .B(REGFILE_SIM_reg_bank__abc_33898_n7434), .Y(REGFILE_SIM_reg_bank__abc_33898_n7435) );
  OR2X2 OR2X2_3968 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7436), .B(REGFILE_SIM_reg_bank__abc_33898_n7437), .Y(REGFILE_SIM_reg_bank__abc_33898_n7438) );
  OR2X2 OR2X2_3969 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7435), .B(REGFILE_SIM_reg_bank__abc_33898_n7438), .Y(REGFILE_SIM_reg_bank__abc_33898_n7439) );
  OR2X2 OR2X2_397 ( .A(_abc_43815_n1472_1_bF_buf0), .B(_abc_43815_n1772), .Y(_abc_43815_n1801) );
  OR2X2 OR2X2_3970 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7432), .B(REGFILE_SIM_reg_bank__abc_33898_n7439), .Y(REGFILE_SIM_reg_bank__abc_33898_n7440) );
  OR2X2 OR2X2_3971 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7441), .B(REGFILE_SIM_reg_bank__abc_33898_n7442), .Y(REGFILE_SIM_reg_bank__abc_33898_n7443) );
  OR2X2 OR2X2_3972 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7444), .B(REGFILE_SIM_reg_bank__abc_33898_n7445), .Y(REGFILE_SIM_reg_bank__abc_33898_n7446) );
  OR2X2 OR2X2_3973 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7443), .B(REGFILE_SIM_reg_bank__abc_33898_n7446), .Y(REGFILE_SIM_reg_bank__abc_33898_n7447) );
  OR2X2 OR2X2_3974 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7448), .B(REGFILE_SIM_reg_bank__abc_33898_n7449), .Y(REGFILE_SIM_reg_bank__abc_33898_n7450) );
  OR2X2 OR2X2_3975 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7451), .B(REGFILE_SIM_reg_bank__abc_33898_n7452), .Y(REGFILE_SIM_reg_bank__abc_33898_n7453) );
  OR2X2 OR2X2_3976 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7453), .B(REGFILE_SIM_reg_bank__abc_33898_n7450), .Y(REGFILE_SIM_reg_bank__abc_33898_n7454) );
  OR2X2 OR2X2_3977 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7447), .B(REGFILE_SIM_reg_bank__abc_33898_n7454), .Y(REGFILE_SIM_reg_bank__abc_33898_n7455) );
  OR2X2 OR2X2_3978 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7440), .B(REGFILE_SIM_reg_bank__abc_33898_n7455), .Y(REGFILE_SIM_reg_bank__abc_33898_n7456) );
  OR2X2 OR2X2_3979 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7457), .B(REGFILE_SIM_reg_bank__abc_33898_n7458), .Y(REGFILE_SIM_reg_bank__abc_33898_n7459) );
  OR2X2 OR2X2_398 ( .A(_abc_43815_n1803), .B(_abc_43815_n1778_1), .Y(_abc_43815_n1804) );
  OR2X2 OR2X2_3980 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7460), .B(REGFILE_SIM_reg_bank__abc_33898_n7461), .Y(REGFILE_SIM_reg_bank__abc_33898_n7462) );
  OR2X2 OR2X2_3981 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7459), .B(REGFILE_SIM_reg_bank__abc_33898_n7462), .Y(REGFILE_SIM_reg_bank__abc_33898_n7463) );
  OR2X2 OR2X2_3982 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7465), .B(REGFILE_SIM_reg_bank__abc_33898_n7466), .Y(REGFILE_SIM_reg_bank__abc_33898_n7467) );
  OR2X2 OR2X2_3983 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7467), .B(REGFILE_SIM_reg_bank__abc_33898_n7464), .Y(REGFILE_SIM_reg_bank__abc_33898_n7468) );
  OR2X2 OR2X2_3984 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7463), .B(REGFILE_SIM_reg_bank__abc_33898_n7468), .Y(REGFILE_SIM_reg_bank__abc_33898_n7469) );
  OR2X2 OR2X2_3985 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7470), .B(REGFILE_SIM_reg_bank__abc_33898_n7471), .Y(REGFILE_SIM_reg_bank__abc_33898_n7472) );
  OR2X2 OR2X2_3986 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7473), .B(REGFILE_SIM_reg_bank__abc_33898_n7474), .Y(REGFILE_SIM_reg_bank__abc_33898_n7475) );
  OR2X2 OR2X2_3987 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7475), .B(REGFILE_SIM_reg_bank__abc_33898_n7472), .Y(REGFILE_SIM_reg_bank__abc_33898_n7476) );
  OR2X2 OR2X2_3988 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7477), .B(REGFILE_SIM_reg_bank__abc_33898_n7478), .Y(REGFILE_SIM_reg_bank__abc_33898_n7479) );
  OR2X2 OR2X2_3989 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7480), .B(REGFILE_SIM_reg_bank__abc_33898_n7481), .Y(REGFILE_SIM_reg_bank__abc_33898_n7482) );
  OR2X2 OR2X2_399 ( .A(_abc_43815_n1805), .B(_abc_43815_n1774), .Y(_abc_43815_n1806) );
  OR2X2 OR2X2_3990 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7479), .B(REGFILE_SIM_reg_bank__abc_33898_n7482), .Y(REGFILE_SIM_reg_bank__abc_33898_n7483) );
  OR2X2 OR2X2_3991 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7476), .B(REGFILE_SIM_reg_bank__abc_33898_n7483), .Y(REGFILE_SIM_reg_bank__abc_33898_n7484) );
  OR2X2 OR2X2_3992 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7484), .B(REGFILE_SIM_reg_bank__abc_33898_n7469), .Y(REGFILE_SIM_reg_bank__abc_33898_n7485) );
  OR2X2 OR2X2_3993 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7456), .B(REGFILE_SIM_reg_bank__abc_33898_n7485), .Y(REGFILE_SIM_reg_bank_reg_rb_o_30_) );
  OR2X2 OR2X2_3994 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7487), .B(REGFILE_SIM_reg_bank__abc_33898_n7488), .Y(REGFILE_SIM_reg_bank__abc_33898_n7489) );
  OR2X2 OR2X2_3995 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7490), .B(REGFILE_SIM_reg_bank__abc_33898_n7491), .Y(REGFILE_SIM_reg_bank__abc_33898_n7492) );
  OR2X2 OR2X2_3996 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7492), .B(REGFILE_SIM_reg_bank__abc_33898_n7489), .Y(REGFILE_SIM_reg_bank__abc_33898_n7493) );
  OR2X2 OR2X2_3997 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7494), .B(REGFILE_SIM_reg_bank__abc_33898_n7495), .Y(REGFILE_SIM_reg_bank__abc_33898_n7496) );
  OR2X2 OR2X2_3998 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7497), .B(REGFILE_SIM_reg_bank__abc_33898_n7498), .Y(REGFILE_SIM_reg_bank__abc_33898_n7499) );
  OR2X2 OR2X2_3999 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7496), .B(REGFILE_SIM_reg_bank__abc_33898_n7499), .Y(REGFILE_SIM_reg_bank__abc_33898_n7500) );
  OR2X2 OR2X2_4 ( .A(_abc_43815_n661), .B(_abc_43815_n655), .Y(_abc_43815_n662) );
  OR2X2 OR2X2_40 ( .A(_abc_43815_n769), .B(_abc_43815_n772), .Y(_abc_43815_n773) );
  OR2X2 OR2X2_400 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_10_), .Y(_abc_43815_n1807) );
  OR2X2 OR2X2_4000 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7493), .B(REGFILE_SIM_reg_bank__abc_33898_n7500), .Y(REGFILE_SIM_reg_bank__abc_33898_n7501) );
  OR2X2 OR2X2_4001 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7502), .B(REGFILE_SIM_reg_bank__abc_33898_n7503), .Y(REGFILE_SIM_reg_bank__abc_33898_n7504) );
  OR2X2 OR2X2_4002 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7505), .B(REGFILE_SIM_reg_bank__abc_33898_n7506), .Y(REGFILE_SIM_reg_bank__abc_33898_n7507) );
  OR2X2 OR2X2_4003 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7504), .B(REGFILE_SIM_reg_bank__abc_33898_n7507), .Y(REGFILE_SIM_reg_bank__abc_33898_n7508) );
  OR2X2 OR2X2_4004 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7509), .B(REGFILE_SIM_reg_bank__abc_33898_n7510), .Y(REGFILE_SIM_reg_bank__abc_33898_n7511) );
  OR2X2 OR2X2_4005 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7512), .B(REGFILE_SIM_reg_bank__abc_33898_n7513), .Y(REGFILE_SIM_reg_bank__abc_33898_n7514) );
  OR2X2 OR2X2_4006 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7514), .B(REGFILE_SIM_reg_bank__abc_33898_n7511), .Y(REGFILE_SIM_reg_bank__abc_33898_n7515) );
  OR2X2 OR2X2_4007 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7508), .B(REGFILE_SIM_reg_bank__abc_33898_n7515), .Y(REGFILE_SIM_reg_bank__abc_33898_n7516) );
  OR2X2 OR2X2_4008 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7501), .B(REGFILE_SIM_reg_bank__abc_33898_n7516), .Y(REGFILE_SIM_reg_bank__abc_33898_n7517) );
  OR2X2 OR2X2_4009 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7518), .B(REGFILE_SIM_reg_bank__abc_33898_n7519), .Y(REGFILE_SIM_reg_bank__abc_33898_n7520) );
  OR2X2 OR2X2_401 ( .A(_abc_43815_n1770), .B(pc_q_11_), .Y(_abc_43815_n1810_1) );
  OR2X2 OR2X2_4010 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7521), .B(REGFILE_SIM_reg_bank__abc_33898_n7522), .Y(REGFILE_SIM_reg_bank__abc_33898_n7523) );
  OR2X2 OR2X2_4011 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7520), .B(REGFILE_SIM_reg_bank__abc_33898_n7523), .Y(REGFILE_SIM_reg_bank__abc_33898_n7524) );
  OR2X2 OR2X2_4012 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7526), .B(REGFILE_SIM_reg_bank__abc_33898_n7527), .Y(REGFILE_SIM_reg_bank__abc_33898_n7528) );
  OR2X2 OR2X2_4013 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7528), .B(REGFILE_SIM_reg_bank__abc_33898_n7525), .Y(REGFILE_SIM_reg_bank__abc_33898_n7529) );
  OR2X2 OR2X2_4014 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7524), .B(REGFILE_SIM_reg_bank__abc_33898_n7529), .Y(REGFILE_SIM_reg_bank__abc_33898_n7530) );
  OR2X2 OR2X2_4015 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7531), .B(REGFILE_SIM_reg_bank__abc_33898_n7532), .Y(REGFILE_SIM_reg_bank__abc_33898_n7533) );
  OR2X2 OR2X2_4016 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7534), .B(REGFILE_SIM_reg_bank__abc_33898_n7535), .Y(REGFILE_SIM_reg_bank__abc_33898_n7536) );
  OR2X2 OR2X2_4017 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7536), .B(REGFILE_SIM_reg_bank__abc_33898_n7533), .Y(REGFILE_SIM_reg_bank__abc_33898_n7537) );
  OR2X2 OR2X2_4018 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7538), .B(REGFILE_SIM_reg_bank__abc_33898_n7539), .Y(REGFILE_SIM_reg_bank__abc_33898_n7540) );
  OR2X2 OR2X2_4019 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7541), .B(REGFILE_SIM_reg_bank__abc_33898_n7542), .Y(REGFILE_SIM_reg_bank__abc_33898_n7543) );
  OR2X2 OR2X2_402 ( .A(_abc_43815_n1813), .B(_abc_43815_n1278_bF_buf6), .Y(_abc_43815_n1814) );
  OR2X2 OR2X2_4020 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7540), .B(REGFILE_SIM_reg_bank__abc_33898_n7543), .Y(REGFILE_SIM_reg_bank__abc_33898_n7544) );
  OR2X2 OR2X2_4021 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7537), .B(REGFILE_SIM_reg_bank__abc_33898_n7544), .Y(REGFILE_SIM_reg_bank__abc_33898_n7545) );
  OR2X2 OR2X2_4022 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7545), .B(REGFILE_SIM_reg_bank__abc_33898_n7530), .Y(REGFILE_SIM_reg_bank__abc_33898_n7546) );
  OR2X2 OR2X2_4023 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7517), .B(REGFILE_SIM_reg_bank__abc_33898_n7546), .Y(REGFILE_SIM_reg_bank_reg_rb_o_31_) );
  OR2X2 OR2X2_4024 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7555), .B(REGFILE_SIM_reg_bank__abc_33898_n7558), .Y(REGFILE_SIM_reg_bank__abc_33898_n7559) );
  OR2X2 OR2X2_4025 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7564), .B(REGFILE_SIM_reg_bank__abc_33898_n7567), .Y(REGFILE_SIM_reg_bank__abc_33898_n7568) );
  OR2X2 OR2X2_4026 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7568), .B(REGFILE_SIM_reg_bank__abc_33898_n7559), .Y(REGFILE_SIM_reg_bank__abc_33898_n7569) );
  OR2X2 OR2X2_4027 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7575), .B(REGFILE_SIM_reg_bank__abc_33898_n7578), .Y(REGFILE_SIM_reg_bank__abc_33898_n7579) );
  OR2X2 OR2X2_4028 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7583), .B(REGFILE_SIM_reg_bank__abc_33898_n7586), .Y(REGFILE_SIM_reg_bank__abc_33898_n7587) );
  OR2X2 OR2X2_4029 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7579), .B(REGFILE_SIM_reg_bank__abc_33898_n7587), .Y(REGFILE_SIM_reg_bank__abc_33898_n7588) );
  OR2X2 OR2X2_403 ( .A(_abc_43815_n1472_1_bF_buf4), .B(_abc_43815_n1813), .Y(_abc_43815_n1816) );
  OR2X2 OR2X2_4030 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7569), .B(REGFILE_SIM_reg_bank__abc_33898_n7588), .Y(REGFILE_SIM_reg_bank__abc_33898_n7589) );
  OR2X2 OR2X2_4031 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7591), .B(REGFILE_SIM_reg_bank__abc_33898_n7593), .Y(REGFILE_SIM_reg_bank__abc_33898_n7594) );
  OR2X2 OR2X2_4032 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7597), .B(REGFILE_SIM_reg_bank__abc_33898_n7600), .Y(REGFILE_SIM_reg_bank__abc_33898_n7601) );
  OR2X2 OR2X2_4033 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7594), .B(REGFILE_SIM_reg_bank__abc_33898_n7601), .Y(REGFILE_SIM_reg_bank__abc_33898_n7602) );
  OR2X2 OR2X2_4034 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7604), .B(REGFILE_SIM_reg_bank__abc_33898_n7607), .Y(REGFILE_SIM_reg_bank__abc_33898_n7608) );
  OR2X2 OR2X2_4035 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7610), .B(REGFILE_SIM_reg_bank__abc_33898_n7613), .Y(REGFILE_SIM_reg_bank__abc_33898_n7614) );
  OR2X2 OR2X2_4036 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7614), .B(REGFILE_SIM_reg_bank__abc_33898_n7608), .Y(REGFILE_SIM_reg_bank__abc_33898_n7615) );
  OR2X2 OR2X2_4037 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7602), .B(REGFILE_SIM_reg_bank__abc_33898_n7615), .Y(REGFILE_SIM_reg_bank__abc_33898_n7616) );
  OR2X2 OR2X2_4038 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7589), .B(REGFILE_SIM_reg_bank__abc_33898_n7616), .Y(REGFILE_SIM_reg_bank__abc_33898_n7617) );
  OR2X2 OR2X2_4039 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7620), .B(REGFILE_SIM_reg_bank__abc_33898_n7623), .Y(REGFILE_SIM_reg_bank__abc_33898_n7624) );
  OR2X2 OR2X2_404 ( .A(alu_op_r_7_), .B(pc_q_11_), .Y(_abc_43815_n1820_1) );
  OR2X2 OR2X2_4040 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7626), .B(REGFILE_SIM_reg_bank__abc_33898_n7628), .Y(REGFILE_SIM_reg_bank__abc_33898_n7629) );
  OR2X2 OR2X2_4041 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7624), .B(REGFILE_SIM_reg_bank__abc_33898_n7629), .Y(REGFILE_SIM_reg_bank__abc_33898_n7630) );
  OR2X2 OR2X2_4042 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7635), .B(REGFILE_SIM_reg_bank__abc_33898_n7637), .Y(REGFILE_SIM_reg_bank__abc_33898_n7638) );
  OR2X2 OR2X2_4043 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7638), .B(REGFILE_SIM_reg_bank__abc_33898_n7633), .Y(REGFILE_SIM_reg_bank__abc_33898_n7639) );
  OR2X2 OR2X2_4044 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7630), .B(REGFILE_SIM_reg_bank__abc_33898_n7639), .Y(REGFILE_SIM_reg_bank__abc_33898_n7640) );
  OR2X2 OR2X2_4045 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7642), .B(REGFILE_SIM_reg_bank__abc_33898_n7644), .Y(REGFILE_SIM_reg_bank__abc_33898_n7645) );
  OR2X2 OR2X2_4046 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7647), .B(REGFILE_SIM_reg_bank__abc_33898_n7649), .Y(REGFILE_SIM_reg_bank__abc_33898_n7650) );
  OR2X2 OR2X2_4047 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7650), .B(REGFILE_SIM_reg_bank__abc_33898_n7645), .Y(REGFILE_SIM_reg_bank__abc_33898_n7651) );
  OR2X2 OR2X2_4048 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7653), .B(REGFILE_SIM_reg_bank__abc_33898_n7655), .Y(REGFILE_SIM_reg_bank__abc_33898_n7656) );
  OR2X2 OR2X2_4049 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7658), .B(REGFILE_SIM_reg_bank__abc_33898_n7660), .Y(REGFILE_SIM_reg_bank__abc_33898_n7661) );
  OR2X2 OR2X2_405 ( .A(_abc_43815_n1819), .B(_abc_43815_n1823_1), .Y(_abc_43815_n1824) );
  OR2X2 OR2X2_4050 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7656), .B(REGFILE_SIM_reg_bank__abc_33898_n7661), .Y(REGFILE_SIM_reg_bank__abc_33898_n7662) );
  OR2X2 OR2X2_4051 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7651), .B(REGFILE_SIM_reg_bank__abc_33898_n7662), .Y(REGFILE_SIM_reg_bank__abc_33898_n7663) );
  OR2X2 OR2X2_4052 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7663), .B(REGFILE_SIM_reg_bank__abc_33898_n7640), .Y(REGFILE_SIM_reg_bank__abc_33898_n7664) );
  OR2X2 OR2X2_4053 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7617), .B(REGFILE_SIM_reg_bank__abc_33898_n7664), .Y(REGFILE_SIM_reg_bank_reg_ra_o_0_) );
  OR2X2 OR2X2_4054 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7666), .B(REGFILE_SIM_reg_bank__abc_33898_n7667), .Y(REGFILE_SIM_reg_bank__abc_33898_n7668) );
  OR2X2 OR2X2_4055 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7669), .B(REGFILE_SIM_reg_bank__abc_33898_n7670), .Y(REGFILE_SIM_reg_bank__abc_33898_n7671) );
  OR2X2 OR2X2_4056 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7671), .B(REGFILE_SIM_reg_bank__abc_33898_n7668), .Y(REGFILE_SIM_reg_bank__abc_33898_n7672) );
  OR2X2 OR2X2_4057 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7673), .B(REGFILE_SIM_reg_bank__abc_33898_n7674), .Y(REGFILE_SIM_reg_bank__abc_33898_n7675) );
  OR2X2 OR2X2_4058 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7676), .B(REGFILE_SIM_reg_bank__abc_33898_n7677), .Y(REGFILE_SIM_reg_bank__abc_33898_n7678) );
  OR2X2 OR2X2_4059 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7675), .B(REGFILE_SIM_reg_bank__abc_33898_n7678), .Y(REGFILE_SIM_reg_bank__abc_33898_n7679) );
  OR2X2 OR2X2_406 ( .A(_abc_43815_n1818), .B(_abc_43815_n1825), .Y(_abc_43815_n1826_1) );
  OR2X2 OR2X2_4060 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7672), .B(REGFILE_SIM_reg_bank__abc_33898_n7679), .Y(REGFILE_SIM_reg_bank__abc_33898_n7680) );
  OR2X2 OR2X2_4061 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7681), .B(REGFILE_SIM_reg_bank__abc_33898_n7682), .Y(REGFILE_SIM_reg_bank__abc_33898_n7683) );
  OR2X2 OR2X2_4062 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7684), .B(REGFILE_SIM_reg_bank__abc_33898_n7685), .Y(REGFILE_SIM_reg_bank__abc_33898_n7686) );
  OR2X2 OR2X2_4063 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7683), .B(REGFILE_SIM_reg_bank__abc_33898_n7686), .Y(REGFILE_SIM_reg_bank__abc_33898_n7687) );
  OR2X2 OR2X2_4064 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7688), .B(REGFILE_SIM_reg_bank__abc_33898_n7689), .Y(REGFILE_SIM_reg_bank__abc_33898_n7690) );
  OR2X2 OR2X2_4065 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7691), .B(REGFILE_SIM_reg_bank__abc_33898_n7692), .Y(REGFILE_SIM_reg_bank__abc_33898_n7693) );
  OR2X2 OR2X2_4066 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7693), .B(REGFILE_SIM_reg_bank__abc_33898_n7690), .Y(REGFILE_SIM_reg_bank__abc_33898_n7694) );
  OR2X2 OR2X2_4067 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7687), .B(REGFILE_SIM_reg_bank__abc_33898_n7694), .Y(REGFILE_SIM_reg_bank__abc_33898_n7695) );
  OR2X2 OR2X2_4068 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7680), .B(REGFILE_SIM_reg_bank__abc_33898_n7695), .Y(REGFILE_SIM_reg_bank__abc_33898_n7696) );
  OR2X2 OR2X2_4069 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7697), .B(REGFILE_SIM_reg_bank__abc_33898_n7698), .Y(REGFILE_SIM_reg_bank__abc_33898_n7699) );
  OR2X2 OR2X2_407 ( .A(_abc_43815_n1828), .B(_abc_43815_n1817), .Y(_abc_43815_n1829_1) );
  OR2X2 OR2X2_4070 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7700), .B(REGFILE_SIM_reg_bank__abc_33898_n7701), .Y(REGFILE_SIM_reg_bank__abc_33898_n7702) );
  OR2X2 OR2X2_4071 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7699), .B(REGFILE_SIM_reg_bank__abc_33898_n7702), .Y(REGFILE_SIM_reg_bank__abc_33898_n7703) );
  OR2X2 OR2X2_4072 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7705), .B(REGFILE_SIM_reg_bank__abc_33898_n7706), .Y(REGFILE_SIM_reg_bank__abc_33898_n7707) );
  OR2X2 OR2X2_4073 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7707), .B(REGFILE_SIM_reg_bank__abc_33898_n7704), .Y(REGFILE_SIM_reg_bank__abc_33898_n7708) );
  OR2X2 OR2X2_4074 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7703), .B(REGFILE_SIM_reg_bank__abc_33898_n7708), .Y(REGFILE_SIM_reg_bank__abc_33898_n7709) );
  OR2X2 OR2X2_4075 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7710), .B(REGFILE_SIM_reg_bank__abc_33898_n7711), .Y(REGFILE_SIM_reg_bank__abc_33898_n7712) );
  OR2X2 OR2X2_4076 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7713), .B(REGFILE_SIM_reg_bank__abc_33898_n7714), .Y(REGFILE_SIM_reg_bank__abc_33898_n7715) );
  OR2X2 OR2X2_4077 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7715), .B(REGFILE_SIM_reg_bank__abc_33898_n7712), .Y(REGFILE_SIM_reg_bank__abc_33898_n7716) );
  OR2X2 OR2X2_4078 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7717), .B(REGFILE_SIM_reg_bank__abc_33898_n7718), .Y(REGFILE_SIM_reg_bank__abc_33898_n7719) );
  OR2X2 OR2X2_4079 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7720), .B(REGFILE_SIM_reg_bank__abc_33898_n7721), .Y(REGFILE_SIM_reg_bank__abc_33898_n7722) );
  OR2X2 OR2X2_408 ( .A(_abc_43815_n1473_bF_buf0), .B(_abc_43815_n1831), .Y(_abc_43815_n1832_1) );
  OR2X2 OR2X2_4080 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7719), .B(REGFILE_SIM_reg_bank__abc_33898_n7722), .Y(REGFILE_SIM_reg_bank__abc_33898_n7723) );
  OR2X2 OR2X2_4081 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7716), .B(REGFILE_SIM_reg_bank__abc_33898_n7723), .Y(REGFILE_SIM_reg_bank__abc_33898_n7724) );
  OR2X2 OR2X2_4082 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7724), .B(REGFILE_SIM_reg_bank__abc_33898_n7709), .Y(REGFILE_SIM_reg_bank__abc_33898_n7725) );
  OR2X2 OR2X2_4083 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7696), .B(REGFILE_SIM_reg_bank__abc_33898_n7725), .Y(REGFILE_SIM_reg_bank_reg_ra_o_1_) );
  OR2X2 OR2X2_4084 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7727), .B(REGFILE_SIM_reg_bank__abc_33898_n7728), .Y(REGFILE_SIM_reg_bank__abc_33898_n7729) );
  OR2X2 OR2X2_4085 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7730), .B(REGFILE_SIM_reg_bank__abc_33898_n7731), .Y(REGFILE_SIM_reg_bank__abc_33898_n7732) );
  OR2X2 OR2X2_4086 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7732), .B(REGFILE_SIM_reg_bank__abc_33898_n7729), .Y(REGFILE_SIM_reg_bank__abc_33898_n7733) );
  OR2X2 OR2X2_4087 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7734), .B(REGFILE_SIM_reg_bank__abc_33898_n7735), .Y(REGFILE_SIM_reg_bank__abc_33898_n7736) );
  OR2X2 OR2X2_4088 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7737), .B(REGFILE_SIM_reg_bank__abc_33898_n7738), .Y(REGFILE_SIM_reg_bank__abc_33898_n7739) );
  OR2X2 OR2X2_4089 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7736), .B(REGFILE_SIM_reg_bank__abc_33898_n7739), .Y(REGFILE_SIM_reg_bank__abc_33898_n7740) );
  OR2X2 OR2X2_409 ( .A(_abc_43815_n1830), .B(_abc_43815_n1832_1), .Y(_abc_43815_n1833) );
  OR2X2 OR2X2_4090 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7733), .B(REGFILE_SIM_reg_bank__abc_33898_n7740), .Y(REGFILE_SIM_reg_bank__abc_33898_n7741) );
  OR2X2 OR2X2_4091 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7742), .B(REGFILE_SIM_reg_bank__abc_33898_n7743), .Y(REGFILE_SIM_reg_bank__abc_33898_n7744) );
  OR2X2 OR2X2_4092 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7745), .B(REGFILE_SIM_reg_bank__abc_33898_n7746), .Y(REGFILE_SIM_reg_bank__abc_33898_n7747) );
  OR2X2 OR2X2_4093 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7744), .B(REGFILE_SIM_reg_bank__abc_33898_n7747), .Y(REGFILE_SIM_reg_bank__abc_33898_n7748) );
  OR2X2 OR2X2_4094 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7749), .B(REGFILE_SIM_reg_bank__abc_33898_n7750), .Y(REGFILE_SIM_reg_bank__abc_33898_n7751) );
  OR2X2 OR2X2_4095 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7752), .B(REGFILE_SIM_reg_bank__abc_33898_n7753), .Y(REGFILE_SIM_reg_bank__abc_33898_n7754) );
  OR2X2 OR2X2_4096 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7754), .B(REGFILE_SIM_reg_bank__abc_33898_n7751), .Y(REGFILE_SIM_reg_bank__abc_33898_n7755) );
  OR2X2 OR2X2_4097 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7748), .B(REGFILE_SIM_reg_bank__abc_33898_n7755), .Y(REGFILE_SIM_reg_bank__abc_33898_n7756) );
  OR2X2 OR2X2_4098 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7741), .B(REGFILE_SIM_reg_bank__abc_33898_n7756), .Y(REGFILE_SIM_reg_bank__abc_33898_n7757) );
  OR2X2 OR2X2_4099 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7758), .B(REGFILE_SIM_reg_bank__abc_33898_n7759), .Y(REGFILE_SIM_reg_bank__abc_33898_n7760) );
  OR2X2 OR2X2_41 ( .A(_abc_43815_n766), .B(_abc_43815_n774), .Y(_abc_43815_n775) );
  OR2X2 OR2X2_410 ( .A(_abc_43815_n1834), .B(_abc_43815_n1350_bF_buf0), .Y(_abc_43815_n1835_1) );
  OR2X2 OR2X2_4100 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7761), .B(REGFILE_SIM_reg_bank__abc_33898_n7762), .Y(REGFILE_SIM_reg_bank__abc_33898_n7763) );
  OR2X2 OR2X2_4101 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7760), .B(REGFILE_SIM_reg_bank__abc_33898_n7763), .Y(REGFILE_SIM_reg_bank__abc_33898_n7764) );
  OR2X2 OR2X2_4102 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7766), .B(REGFILE_SIM_reg_bank__abc_33898_n7767), .Y(REGFILE_SIM_reg_bank__abc_33898_n7768) );
  OR2X2 OR2X2_4103 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7768), .B(REGFILE_SIM_reg_bank__abc_33898_n7765), .Y(REGFILE_SIM_reg_bank__abc_33898_n7769) );
  OR2X2 OR2X2_4104 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7764), .B(REGFILE_SIM_reg_bank__abc_33898_n7769), .Y(REGFILE_SIM_reg_bank__abc_33898_n7770) );
  OR2X2 OR2X2_4105 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7771), .B(REGFILE_SIM_reg_bank__abc_33898_n7772), .Y(REGFILE_SIM_reg_bank__abc_33898_n7773) );
  OR2X2 OR2X2_4106 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7774), .B(REGFILE_SIM_reg_bank__abc_33898_n7775), .Y(REGFILE_SIM_reg_bank__abc_33898_n7776) );
  OR2X2 OR2X2_4107 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7776), .B(REGFILE_SIM_reg_bank__abc_33898_n7773), .Y(REGFILE_SIM_reg_bank__abc_33898_n7777) );
  OR2X2 OR2X2_4108 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7778), .B(REGFILE_SIM_reg_bank__abc_33898_n7779), .Y(REGFILE_SIM_reg_bank__abc_33898_n7780) );
  OR2X2 OR2X2_4109 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7781), .B(REGFILE_SIM_reg_bank__abc_33898_n7782), .Y(REGFILE_SIM_reg_bank__abc_33898_n7783) );
  OR2X2 OR2X2_411 ( .A(_abc_43815_n1836), .B(_abc_43815_n1837), .Y(_abc_43815_n1838_1) );
  OR2X2 OR2X2_4110 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7780), .B(REGFILE_SIM_reg_bank__abc_33898_n7783), .Y(REGFILE_SIM_reg_bank__abc_33898_n7784) );
  OR2X2 OR2X2_4111 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7777), .B(REGFILE_SIM_reg_bank__abc_33898_n7784), .Y(REGFILE_SIM_reg_bank__abc_33898_n7785) );
  OR2X2 OR2X2_4112 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7785), .B(REGFILE_SIM_reg_bank__abc_33898_n7770), .Y(REGFILE_SIM_reg_bank__abc_33898_n7786) );
  OR2X2 OR2X2_4113 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7757), .B(REGFILE_SIM_reg_bank__abc_33898_n7786), .Y(REGFILE_SIM_reg_bank_reg_ra_o_2_) );
  OR2X2 OR2X2_4114 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7788), .B(REGFILE_SIM_reg_bank__abc_33898_n7789), .Y(REGFILE_SIM_reg_bank__abc_33898_n7790) );
  OR2X2 OR2X2_4115 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7791), .B(REGFILE_SIM_reg_bank__abc_33898_n7792), .Y(REGFILE_SIM_reg_bank__abc_33898_n7793) );
  OR2X2 OR2X2_4116 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7793), .B(REGFILE_SIM_reg_bank__abc_33898_n7790), .Y(REGFILE_SIM_reg_bank__abc_33898_n7794) );
  OR2X2 OR2X2_4117 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7795), .B(REGFILE_SIM_reg_bank__abc_33898_n7796), .Y(REGFILE_SIM_reg_bank__abc_33898_n7797) );
  OR2X2 OR2X2_4118 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7798), .B(REGFILE_SIM_reg_bank__abc_33898_n7799), .Y(REGFILE_SIM_reg_bank__abc_33898_n7800) );
  OR2X2 OR2X2_4119 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7797), .B(REGFILE_SIM_reg_bank__abc_33898_n7800), .Y(REGFILE_SIM_reg_bank__abc_33898_n7801) );
  OR2X2 OR2X2_412 ( .A(_abc_43815_n1413_bF_buf3), .B(_abc_43815_n1838_1), .Y(_abc_43815_n1839) );
  OR2X2 OR2X2_4120 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7794), .B(REGFILE_SIM_reg_bank__abc_33898_n7801), .Y(REGFILE_SIM_reg_bank__abc_33898_n7802) );
  OR2X2 OR2X2_4121 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7803), .B(REGFILE_SIM_reg_bank__abc_33898_n7804), .Y(REGFILE_SIM_reg_bank__abc_33898_n7805) );
  OR2X2 OR2X2_4122 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7806), .B(REGFILE_SIM_reg_bank__abc_33898_n7807), .Y(REGFILE_SIM_reg_bank__abc_33898_n7808) );
  OR2X2 OR2X2_4123 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7805), .B(REGFILE_SIM_reg_bank__abc_33898_n7808), .Y(REGFILE_SIM_reg_bank__abc_33898_n7809) );
  OR2X2 OR2X2_4124 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7810), .B(REGFILE_SIM_reg_bank__abc_33898_n7811), .Y(REGFILE_SIM_reg_bank__abc_33898_n7812) );
  OR2X2 OR2X2_4125 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7813), .B(REGFILE_SIM_reg_bank__abc_33898_n7814), .Y(REGFILE_SIM_reg_bank__abc_33898_n7815) );
  OR2X2 OR2X2_4126 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7815), .B(REGFILE_SIM_reg_bank__abc_33898_n7812), .Y(REGFILE_SIM_reg_bank__abc_33898_n7816) );
  OR2X2 OR2X2_4127 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7809), .B(REGFILE_SIM_reg_bank__abc_33898_n7816), .Y(REGFILE_SIM_reg_bank__abc_33898_n7817) );
  OR2X2 OR2X2_4128 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7802), .B(REGFILE_SIM_reg_bank__abc_33898_n7817), .Y(REGFILE_SIM_reg_bank__abc_33898_n7818) );
  OR2X2 OR2X2_4129 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7819), .B(REGFILE_SIM_reg_bank__abc_33898_n7820), .Y(REGFILE_SIM_reg_bank__abc_33898_n7821) );
  OR2X2 OR2X2_413 ( .A(_abc_43815_n1841_1), .B(_abc_43815_n1815_1), .Y(_abc_43815_n1842) );
  OR2X2 OR2X2_4130 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7822), .B(REGFILE_SIM_reg_bank__abc_33898_n7823), .Y(REGFILE_SIM_reg_bank__abc_33898_n7824) );
  OR2X2 OR2X2_4131 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7821), .B(REGFILE_SIM_reg_bank__abc_33898_n7824), .Y(REGFILE_SIM_reg_bank__abc_33898_n7825) );
  OR2X2 OR2X2_4132 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7827), .B(REGFILE_SIM_reg_bank__abc_33898_n7828), .Y(REGFILE_SIM_reg_bank__abc_33898_n7829) );
  OR2X2 OR2X2_4133 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7829), .B(REGFILE_SIM_reg_bank__abc_33898_n7826), .Y(REGFILE_SIM_reg_bank__abc_33898_n7830) );
  OR2X2 OR2X2_4134 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7825), .B(REGFILE_SIM_reg_bank__abc_33898_n7830), .Y(REGFILE_SIM_reg_bank__abc_33898_n7831) );
  OR2X2 OR2X2_4135 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7832), .B(REGFILE_SIM_reg_bank__abc_33898_n7833), .Y(REGFILE_SIM_reg_bank__abc_33898_n7834) );
  OR2X2 OR2X2_4136 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7835), .B(REGFILE_SIM_reg_bank__abc_33898_n7836), .Y(REGFILE_SIM_reg_bank__abc_33898_n7837) );
  OR2X2 OR2X2_4137 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7837), .B(REGFILE_SIM_reg_bank__abc_33898_n7834), .Y(REGFILE_SIM_reg_bank__abc_33898_n7838) );
  OR2X2 OR2X2_4138 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7839), .B(REGFILE_SIM_reg_bank__abc_33898_n7840), .Y(REGFILE_SIM_reg_bank__abc_33898_n7841) );
  OR2X2 OR2X2_4139 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7842), .B(REGFILE_SIM_reg_bank__abc_33898_n7843), .Y(REGFILE_SIM_reg_bank__abc_33898_n7844) );
  OR2X2 OR2X2_414 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_11_), .Y(_abc_43815_n1843) );
  OR2X2 OR2X2_4140 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7841), .B(REGFILE_SIM_reg_bank__abc_33898_n7844), .Y(REGFILE_SIM_reg_bank__abc_33898_n7845) );
  OR2X2 OR2X2_4141 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7838), .B(REGFILE_SIM_reg_bank__abc_33898_n7845), .Y(REGFILE_SIM_reg_bank__abc_33898_n7846) );
  OR2X2 OR2X2_4142 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7846), .B(REGFILE_SIM_reg_bank__abc_33898_n7831), .Y(REGFILE_SIM_reg_bank__abc_33898_n7847) );
  OR2X2 OR2X2_4143 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7818), .B(REGFILE_SIM_reg_bank__abc_33898_n7847), .Y(REGFILE_SIM_reg_bank_reg_ra_o_3_) );
  OR2X2 OR2X2_4144 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7849), .B(REGFILE_SIM_reg_bank__abc_33898_n7850), .Y(REGFILE_SIM_reg_bank__abc_33898_n7851) );
  OR2X2 OR2X2_4145 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7852), .B(REGFILE_SIM_reg_bank__abc_33898_n7853), .Y(REGFILE_SIM_reg_bank__abc_33898_n7854) );
  OR2X2 OR2X2_4146 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7854), .B(REGFILE_SIM_reg_bank__abc_33898_n7851), .Y(REGFILE_SIM_reg_bank__abc_33898_n7855) );
  OR2X2 OR2X2_4147 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7856), .B(REGFILE_SIM_reg_bank__abc_33898_n7857), .Y(REGFILE_SIM_reg_bank__abc_33898_n7858) );
  OR2X2 OR2X2_4148 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7859), .B(REGFILE_SIM_reg_bank__abc_33898_n7860), .Y(REGFILE_SIM_reg_bank__abc_33898_n7861) );
  OR2X2 OR2X2_4149 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7858), .B(REGFILE_SIM_reg_bank__abc_33898_n7861), .Y(REGFILE_SIM_reg_bank__abc_33898_n7862) );
  OR2X2 OR2X2_415 ( .A(_abc_43815_n1811), .B(pc_q_12_), .Y(_abc_43815_n1846) );
  OR2X2 OR2X2_4150 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7855), .B(REGFILE_SIM_reg_bank__abc_33898_n7862), .Y(REGFILE_SIM_reg_bank__abc_33898_n7863) );
  OR2X2 OR2X2_4151 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7864), .B(REGFILE_SIM_reg_bank__abc_33898_n7865), .Y(REGFILE_SIM_reg_bank__abc_33898_n7866) );
  OR2X2 OR2X2_4152 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7867), .B(REGFILE_SIM_reg_bank__abc_33898_n7868), .Y(REGFILE_SIM_reg_bank__abc_33898_n7869) );
  OR2X2 OR2X2_4153 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7866), .B(REGFILE_SIM_reg_bank__abc_33898_n7869), .Y(REGFILE_SIM_reg_bank__abc_33898_n7870) );
  OR2X2 OR2X2_4154 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7871), .B(REGFILE_SIM_reg_bank__abc_33898_n7872), .Y(REGFILE_SIM_reg_bank__abc_33898_n7873) );
  OR2X2 OR2X2_4155 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7874), .B(REGFILE_SIM_reg_bank__abc_33898_n7875), .Y(REGFILE_SIM_reg_bank__abc_33898_n7876) );
  OR2X2 OR2X2_4156 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7876), .B(REGFILE_SIM_reg_bank__abc_33898_n7873), .Y(REGFILE_SIM_reg_bank__abc_33898_n7877) );
  OR2X2 OR2X2_4157 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7870), .B(REGFILE_SIM_reg_bank__abc_33898_n7877), .Y(REGFILE_SIM_reg_bank__abc_33898_n7878) );
  OR2X2 OR2X2_4158 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7863), .B(REGFILE_SIM_reg_bank__abc_33898_n7878), .Y(REGFILE_SIM_reg_bank__abc_33898_n7879) );
  OR2X2 OR2X2_4159 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7880), .B(REGFILE_SIM_reg_bank__abc_33898_n7881), .Y(REGFILE_SIM_reg_bank__abc_33898_n7882) );
  OR2X2 OR2X2_416 ( .A(_abc_43815_n1849), .B(_abc_43815_n1278_bF_buf5), .Y(_abc_43815_n1850_1) );
  OR2X2 OR2X2_4160 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7883), .B(REGFILE_SIM_reg_bank__abc_33898_n7884), .Y(REGFILE_SIM_reg_bank__abc_33898_n7885) );
  OR2X2 OR2X2_4161 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7882), .B(REGFILE_SIM_reg_bank__abc_33898_n7885), .Y(REGFILE_SIM_reg_bank__abc_33898_n7886) );
  OR2X2 OR2X2_4162 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7888), .B(REGFILE_SIM_reg_bank__abc_33898_n7889), .Y(REGFILE_SIM_reg_bank__abc_33898_n7890) );
  OR2X2 OR2X2_4163 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7890), .B(REGFILE_SIM_reg_bank__abc_33898_n7887), .Y(REGFILE_SIM_reg_bank__abc_33898_n7891) );
  OR2X2 OR2X2_4164 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7886), .B(REGFILE_SIM_reg_bank__abc_33898_n7891), .Y(REGFILE_SIM_reg_bank__abc_33898_n7892) );
  OR2X2 OR2X2_4165 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7893), .B(REGFILE_SIM_reg_bank__abc_33898_n7894), .Y(REGFILE_SIM_reg_bank__abc_33898_n7895) );
  OR2X2 OR2X2_4166 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7896), .B(REGFILE_SIM_reg_bank__abc_33898_n7897), .Y(REGFILE_SIM_reg_bank__abc_33898_n7898) );
  OR2X2 OR2X2_4167 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7898), .B(REGFILE_SIM_reg_bank__abc_33898_n7895), .Y(REGFILE_SIM_reg_bank__abc_33898_n7899) );
  OR2X2 OR2X2_4168 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7900), .B(REGFILE_SIM_reg_bank__abc_33898_n7901), .Y(REGFILE_SIM_reg_bank__abc_33898_n7902) );
  OR2X2 OR2X2_4169 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7903), .B(REGFILE_SIM_reg_bank__abc_33898_n7904), .Y(REGFILE_SIM_reg_bank__abc_33898_n7905) );
  OR2X2 OR2X2_417 ( .A(_abc_43815_n1853_1), .B(_abc_43815_n1852), .Y(_abc_43815_n1854) );
  OR2X2 OR2X2_4170 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7902), .B(REGFILE_SIM_reg_bank__abc_33898_n7905), .Y(REGFILE_SIM_reg_bank__abc_33898_n7906) );
  OR2X2 OR2X2_4171 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7899), .B(REGFILE_SIM_reg_bank__abc_33898_n7906), .Y(REGFILE_SIM_reg_bank__abc_33898_n7907) );
  OR2X2 OR2X2_4172 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7907), .B(REGFILE_SIM_reg_bank__abc_33898_n7892), .Y(REGFILE_SIM_reg_bank__abc_33898_n7908) );
  OR2X2 OR2X2_4173 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7879), .B(REGFILE_SIM_reg_bank__abc_33898_n7908), .Y(REGFILE_SIM_reg_bank_reg_ra_o_4_) );
  OR2X2 OR2X2_4174 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7910), .B(REGFILE_SIM_reg_bank__abc_33898_n7911), .Y(REGFILE_SIM_reg_bank__abc_33898_n7912) );
  OR2X2 OR2X2_4175 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7913), .B(REGFILE_SIM_reg_bank__abc_33898_n7914), .Y(REGFILE_SIM_reg_bank__abc_33898_n7915) );
  OR2X2 OR2X2_4176 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7915), .B(REGFILE_SIM_reg_bank__abc_33898_n7912), .Y(REGFILE_SIM_reg_bank__abc_33898_n7916) );
  OR2X2 OR2X2_4177 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7917), .B(REGFILE_SIM_reg_bank__abc_33898_n7918), .Y(REGFILE_SIM_reg_bank__abc_33898_n7919) );
  OR2X2 OR2X2_4178 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7920), .B(REGFILE_SIM_reg_bank__abc_33898_n7921), .Y(REGFILE_SIM_reg_bank__abc_33898_n7922) );
  OR2X2 OR2X2_4179 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7919), .B(REGFILE_SIM_reg_bank__abc_33898_n7922), .Y(REGFILE_SIM_reg_bank__abc_33898_n7923) );
  OR2X2 OR2X2_418 ( .A(_abc_43815_n1431_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_43815_n1856_1) );
  OR2X2 OR2X2_4180 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7916), .B(REGFILE_SIM_reg_bank__abc_33898_n7923), .Y(REGFILE_SIM_reg_bank__abc_33898_n7924) );
  OR2X2 OR2X2_4181 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7925), .B(REGFILE_SIM_reg_bank__abc_33898_n7926), .Y(REGFILE_SIM_reg_bank__abc_33898_n7927) );
  OR2X2 OR2X2_4182 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7928), .B(REGFILE_SIM_reg_bank__abc_33898_n7929), .Y(REGFILE_SIM_reg_bank__abc_33898_n7930) );
  OR2X2 OR2X2_4183 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7927), .B(REGFILE_SIM_reg_bank__abc_33898_n7930), .Y(REGFILE_SIM_reg_bank__abc_33898_n7931) );
  OR2X2 OR2X2_4184 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7932), .B(REGFILE_SIM_reg_bank__abc_33898_n7933), .Y(REGFILE_SIM_reg_bank__abc_33898_n7934) );
  OR2X2 OR2X2_4185 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7935), .B(REGFILE_SIM_reg_bank__abc_33898_n7936), .Y(REGFILE_SIM_reg_bank__abc_33898_n7937) );
  OR2X2 OR2X2_4186 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7937), .B(REGFILE_SIM_reg_bank__abc_33898_n7934), .Y(REGFILE_SIM_reg_bank__abc_33898_n7938) );
  OR2X2 OR2X2_4187 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7931), .B(REGFILE_SIM_reg_bank__abc_33898_n7938), .Y(REGFILE_SIM_reg_bank__abc_33898_n7939) );
  OR2X2 OR2X2_4188 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7924), .B(REGFILE_SIM_reg_bank__abc_33898_n7939), .Y(REGFILE_SIM_reg_bank__abc_33898_n7940) );
  OR2X2 OR2X2_4189 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7941), .B(REGFILE_SIM_reg_bank__abc_33898_n7942), .Y(REGFILE_SIM_reg_bank__abc_33898_n7943) );
  OR2X2 OR2X2_419 ( .A(_abc_43815_n1825), .B(_abc_43815_n1782), .Y(_abc_43815_n1862_1) );
  OR2X2 OR2X2_4190 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7944), .B(REGFILE_SIM_reg_bank__abc_33898_n7945), .Y(REGFILE_SIM_reg_bank__abc_33898_n7946) );
  OR2X2 OR2X2_4191 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7943), .B(REGFILE_SIM_reg_bank__abc_33898_n7946), .Y(REGFILE_SIM_reg_bank__abc_33898_n7947) );
  OR2X2 OR2X2_4192 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7949), .B(REGFILE_SIM_reg_bank__abc_33898_n7950), .Y(REGFILE_SIM_reg_bank__abc_33898_n7951) );
  OR2X2 OR2X2_4193 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7951), .B(REGFILE_SIM_reg_bank__abc_33898_n7948), .Y(REGFILE_SIM_reg_bank__abc_33898_n7952) );
  OR2X2 OR2X2_4194 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7947), .B(REGFILE_SIM_reg_bank__abc_33898_n7952), .Y(REGFILE_SIM_reg_bank__abc_33898_n7953) );
  OR2X2 OR2X2_4195 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7954), .B(REGFILE_SIM_reg_bank__abc_33898_n7955), .Y(REGFILE_SIM_reg_bank__abc_33898_n7956) );
  OR2X2 OR2X2_4196 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7957), .B(REGFILE_SIM_reg_bank__abc_33898_n7958), .Y(REGFILE_SIM_reg_bank__abc_33898_n7959) );
  OR2X2 OR2X2_4197 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7959), .B(REGFILE_SIM_reg_bank__abc_33898_n7956), .Y(REGFILE_SIM_reg_bank__abc_33898_n7960) );
  OR2X2 OR2X2_4198 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7961), .B(REGFILE_SIM_reg_bank__abc_33898_n7962), .Y(REGFILE_SIM_reg_bank__abc_33898_n7963) );
  OR2X2 OR2X2_4199 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7964), .B(REGFILE_SIM_reg_bank__abc_33898_n7965), .Y(REGFILE_SIM_reg_bank__abc_33898_n7966) );
  OR2X2 OR2X2_42 ( .A(_abc_43815_n776), .B(_abc_43815_n762), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_) );
  OR2X2 OR2X2_420 ( .A(_abc_43815_n1859_1), .B(_abc_43815_n1865_1), .Y(_abc_43815_n1866) );
  OR2X2 OR2X2_4200 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7963), .B(REGFILE_SIM_reg_bank__abc_33898_n7966), .Y(REGFILE_SIM_reg_bank__abc_33898_n7967) );
  OR2X2 OR2X2_4201 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7960), .B(REGFILE_SIM_reg_bank__abc_33898_n7967), .Y(REGFILE_SIM_reg_bank__abc_33898_n7968) );
  OR2X2 OR2X2_4202 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7968), .B(REGFILE_SIM_reg_bank__abc_33898_n7953), .Y(REGFILE_SIM_reg_bank__abc_33898_n7969) );
  OR2X2 OR2X2_4203 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7940), .B(REGFILE_SIM_reg_bank__abc_33898_n7969), .Y(REGFILE_SIM_reg_bank_reg_ra_o_5_) );
  OR2X2 OR2X2_4204 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7971), .B(REGFILE_SIM_reg_bank__abc_33898_n7972), .Y(REGFILE_SIM_reg_bank__abc_33898_n7973) );
  OR2X2 OR2X2_4205 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7974), .B(REGFILE_SIM_reg_bank__abc_33898_n7975), .Y(REGFILE_SIM_reg_bank__abc_33898_n7976) );
  OR2X2 OR2X2_4206 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7976), .B(REGFILE_SIM_reg_bank__abc_33898_n7973), .Y(REGFILE_SIM_reg_bank__abc_33898_n7977) );
  OR2X2 OR2X2_4207 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7978), .B(REGFILE_SIM_reg_bank__abc_33898_n7979), .Y(REGFILE_SIM_reg_bank__abc_33898_n7980) );
  OR2X2 OR2X2_4208 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7981), .B(REGFILE_SIM_reg_bank__abc_33898_n7982), .Y(REGFILE_SIM_reg_bank__abc_33898_n7983) );
  OR2X2 OR2X2_4209 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7980), .B(REGFILE_SIM_reg_bank__abc_33898_n7983), .Y(REGFILE_SIM_reg_bank__abc_33898_n7984) );
  OR2X2 OR2X2_421 ( .A(int32_r_10_), .B(pc_q_12_), .Y(_abc_43815_n1867) );
  OR2X2 OR2X2_4210 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7977), .B(REGFILE_SIM_reg_bank__abc_33898_n7984), .Y(REGFILE_SIM_reg_bank__abc_33898_n7985) );
  OR2X2 OR2X2_4211 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7986), .B(REGFILE_SIM_reg_bank__abc_33898_n7987), .Y(REGFILE_SIM_reg_bank__abc_33898_n7988) );
  OR2X2 OR2X2_4212 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7989), .B(REGFILE_SIM_reg_bank__abc_33898_n7990), .Y(REGFILE_SIM_reg_bank__abc_33898_n7991) );
  OR2X2 OR2X2_4213 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7988), .B(REGFILE_SIM_reg_bank__abc_33898_n7991), .Y(REGFILE_SIM_reg_bank__abc_33898_n7992) );
  OR2X2 OR2X2_4214 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7993), .B(REGFILE_SIM_reg_bank__abc_33898_n7994), .Y(REGFILE_SIM_reg_bank__abc_33898_n7995) );
  OR2X2 OR2X2_4215 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7996), .B(REGFILE_SIM_reg_bank__abc_33898_n7997), .Y(REGFILE_SIM_reg_bank__abc_33898_n7998) );
  OR2X2 OR2X2_4216 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7998), .B(REGFILE_SIM_reg_bank__abc_33898_n7995), .Y(REGFILE_SIM_reg_bank__abc_33898_n7999) );
  OR2X2 OR2X2_4217 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7992), .B(REGFILE_SIM_reg_bank__abc_33898_n7999), .Y(REGFILE_SIM_reg_bank__abc_33898_n8000) );
  OR2X2 OR2X2_4218 ( .A(REGFILE_SIM_reg_bank__abc_33898_n7985), .B(REGFILE_SIM_reg_bank__abc_33898_n8000), .Y(REGFILE_SIM_reg_bank__abc_33898_n8001) );
  OR2X2 OR2X2_4219 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8002), .B(REGFILE_SIM_reg_bank__abc_33898_n8003), .Y(REGFILE_SIM_reg_bank__abc_33898_n8004) );
  OR2X2 OR2X2_422 ( .A(_abc_43815_n1866), .B(_abc_43815_n1870), .Y(_abc_43815_n1873) );
  OR2X2 OR2X2_4220 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8005), .B(REGFILE_SIM_reg_bank__abc_33898_n8006), .Y(REGFILE_SIM_reg_bank__abc_33898_n8007) );
  OR2X2 OR2X2_4221 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8004), .B(REGFILE_SIM_reg_bank__abc_33898_n8007), .Y(REGFILE_SIM_reg_bank__abc_33898_n8008) );
  OR2X2 OR2X2_4222 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8010), .B(REGFILE_SIM_reg_bank__abc_33898_n8011), .Y(REGFILE_SIM_reg_bank__abc_33898_n8012) );
  OR2X2 OR2X2_4223 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8012), .B(REGFILE_SIM_reg_bank__abc_33898_n8009), .Y(REGFILE_SIM_reg_bank__abc_33898_n8013) );
  OR2X2 OR2X2_4224 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8008), .B(REGFILE_SIM_reg_bank__abc_33898_n8013), .Y(REGFILE_SIM_reg_bank__abc_33898_n8014) );
  OR2X2 OR2X2_4225 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8015), .B(REGFILE_SIM_reg_bank__abc_33898_n8016), .Y(REGFILE_SIM_reg_bank__abc_33898_n8017) );
  OR2X2 OR2X2_4226 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8018), .B(REGFILE_SIM_reg_bank__abc_33898_n8019), .Y(REGFILE_SIM_reg_bank__abc_33898_n8020) );
  OR2X2 OR2X2_4227 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8020), .B(REGFILE_SIM_reg_bank__abc_33898_n8017), .Y(REGFILE_SIM_reg_bank__abc_33898_n8021) );
  OR2X2 OR2X2_4228 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8022), .B(REGFILE_SIM_reg_bank__abc_33898_n8023), .Y(REGFILE_SIM_reg_bank__abc_33898_n8024) );
  OR2X2 OR2X2_4229 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8025), .B(REGFILE_SIM_reg_bank__abc_33898_n8026), .Y(REGFILE_SIM_reg_bank__abc_33898_n8027) );
  OR2X2 OR2X2_423 ( .A(_abc_43815_n1428_bF_buf1), .B(_abc_43815_n1876), .Y(_abc_43815_n1877_1) );
  OR2X2 OR2X2_4230 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8024), .B(REGFILE_SIM_reg_bank__abc_33898_n8027), .Y(REGFILE_SIM_reg_bank__abc_33898_n8028) );
  OR2X2 OR2X2_4231 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8021), .B(REGFILE_SIM_reg_bank__abc_33898_n8028), .Y(REGFILE_SIM_reg_bank__abc_33898_n8029) );
  OR2X2 OR2X2_4232 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8029), .B(REGFILE_SIM_reg_bank__abc_33898_n8014), .Y(REGFILE_SIM_reg_bank__abc_33898_n8030) );
  OR2X2 OR2X2_4233 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8001), .B(REGFILE_SIM_reg_bank__abc_33898_n8030), .Y(REGFILE_SIM_reg_bank_reg_ra_o_6_) );
  OR2X2 OR2X2_4234 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8032), .B(REGFILE_SIM_reg_bank__abc_33898_n8033), .Y(REGFILE_SIM_reg_bank__abc_33898_n8034) );
  OR2X2 OR2X2_4235 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8035), .B(REGFILE_SIM_reg_bank__abc_33898_n8036), .Y(REGFILE_SIM_reg_bank__abc_33898_n8037) );
  OR2X2 OR2X2_4236 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8037), .B(REGFILE_SIM_reg_bank__abc_33898_n8034), .Y(REGFILE_SIM_reg_bank__abc_33898_n8038) );
  OR2X2 OR2X2_4237 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8039), .B(REGFILE_SIM_reg_bank__abc_33898_n8040), .Y(REGFILE_SIM_reg_bank__abc_33898_n8041) );
  OR2X2 OR2X2_4238 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8042), .B(REGFILE_SIM_reg_bank__abc_33898_n8043), .Y(REGFILE_SIM_reg_bank__abc_33898_n8044) );
  OR2X2 OR2X2_4239 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8041), .B(REGFILE_SIM_reg_bank__abc_33898_n8044), .Y(REGFILE_SIM_reg_bank__abc_33898_n8045) );
  OR2X2 OR2X2_424 ( .A(_abc_43815_n1875), .B(_abc_43815_n1877_1), .Y(_abc_43815_n1878) );
  OR2X2 OR2X2_4240 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8038), .B(REGFILE_SIM_reg_bank__abc_33898_n8045), .Y(REGFILE_SIM_reg_bank__abc_33898_n8046) );
  OR2X2 OR2X2_4241 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8047), .B(REGFILE_SIM_reg_bank__abc_33898_n8048), .Y(REGFILE_SIM_reg_bank__abc_33898_n8049) );
  OR2X2 OR2X2_4242 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8050), .B(REGFILE_SIM_reg_bank__abc_33898_n8051), .Y(REGFILE_SIM_reg_bank__abc_33898_n8052) );
  OR2X2 OR2X2_4243 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8049), .B(REGFILE_SIM_reg_bank__abc_33898_n8052), .Y(REGFILE_SIM_reg_bank__abc_33898_n8053) );
  OR2X2 OR2X2_4244 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8054), .B(REGFILE_SIM_reg_bank__abc_33898_n8055), .Y(REGFILE_SIM_reg_bank__abc_33898_n8056) );
  OR2X2 OR2X2_4245 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8057), .B(REGFILE_SIM_reg_bank__abc_33898_n8058), .Y(REGFILE_SIM_reg_bank__abc_33898_n8059) );
  OR2X2 OR2X2_4246 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8059), .B(REGFILE_SIM_reg_bank__abc_33898_n8056), .Y(REGFILE_SIM_reg_bank__abc_33898_n8060) );
  OR2X2 OR2X2_4247 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8053), .B(REGFILE_SIM_reg_bank__abc_33898_n8060), .Y(REGFILE_SIM_reg_bank__abc_33898_n8061) );
  OR2X2 OR2X2_4248 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8046), .B(REGFILE_SIM_reg_bank__abc_33898_n8061), .Y(REGFILE_SIM_reg_bank__abc_33898_n8062) );
  OR2X2 OR2X2_4249 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8063), .B(REGFILE_SIM_reg_bank__abc_33898_n8064), .Y(REGFILE_SIM_reg_bank__abc_33898_n8065) );
  OR2X2 OR2X2_425 ( .A(_abc_43815_n1879), .B(_abc_43815_n1473_bF_buf4), .Y(_abc_43815_n1880_1) );
  OR2X2 OR2X2_4250 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8066), .B(REGFILE_SIM_reg_bank__abc_33898_n8067), .Y(REGFILE_SIM_reg_bank__abc_33898_n8068) );
  OR2X2 OR2X2_4251 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8065), .B(REGFILE_SIM_reg_bank__abc_33898_n8068), .Y(REGFILE_SIM_reg_bank__abc_33898_n8069) );
  OR2X2 OR2X2_4252 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8071), .B(REGFILE_SIM_reg_bank__abc_33898_n8072), .Y(REGFILE_SIM_reg_bank__abc_33898_n8073) );
  OR2X2 OR2X2_4253 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8073), .B(REGFILE_SIM_reg_bank__abc_33898_n8070), .Y(REGFILE_SIM_reg_bank__abc_33898_n8074) );
  OR2X2 OR2X2_4254 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8069), .B(REGFILE_SIM_reg_bank__abc_33898_n8074), .Y(REGFILE_SIM_reg_bank__abc_33898_n8075) );
  OR2X2 OR2X2_4255 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8076), .B(REGFILE_SIM_reg_bank__abc_33898_n8077), .Y(REGFILE_SIM_reg_bank__abc_33898_n8078) );
  OR2X2 OR2X2_4256 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8079), .B(REGFILE_SIM_reg_bank__abc_33898_n8080), .Y(REGFILE_SIM_reg_bank__abc_33898_n8081) );
  OR2X2 OR2X2_4257 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8081), .B(REGFILE_SIM_reg_bank__abc_33898_n8078), .Y(REGFILE_SIM_reg_bank__abc_33898_n8082) );
  OR2X2 OR2X2_4258 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8083), .B(REGFILE_SIM_reg_bank__abc_33898_n8084), .Y(REGFILE_SIM_reg_bank__abc_33898_n8085) );
  OR2X2 OR2X2_4259 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8086), .B(REGFILE_SIM_reg_bank__abc_33898_n8087), .Y(REGFILE_SIM_reg_bank__abc_33898_n8088) );
  OR2X2 OR2X2_426 ( .A(_abc_43815_n1472_1_bF_buf3), .B(_abc_43815_n1849), .Y(_abc_43815_n1881) );
  OR2X2 OR2X2_4260 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8085), .B(REGFILE_SIM_reg_bank__abc_33898_n8088), .Y(REGFILE_SIM_reg_bank__abc_33898_n8089) );
  OR2X2 OR2X2_4261 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8082), .B(REGFILE_SIM_reg_bank__abc_33898_n8089), .Y(REGFILE_SIM_reg_bank__abc_33898_n8090) );
  OR2X2 OR2X2_4262 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8090), .B(REGFILE_SIM_reg_bank__abc_33898_n8075), .Y(REGFILE_SIM_reg_bank__abc_33898_n8091) );
  OR2X2 OR2X2_4263 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8062), .B(REGFILE_SIM_reg_bank__abc_33898_n8091), .Y(REGFILE_SIM_reg_bank_reg_ra_o_7_) );
  OR2X2 OR2X2_4264 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8093), .B(REGFILE_SIM_reg_bank__abc_33898_n8094), .Y(REGFILE_SIM_reg_bank__abc_33898_n8095) );
  OR2X2 OR2X2_4265 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8096), .B(REGFILE_SIM_reg_bank__abc_33898_n8097), .Y(REGFILE_SIM_reg_bank__abc_33898_n8098) );
  OR2X2 OR2X2_4266 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8098), .B(REGFILE_SIM_reg_bank__abc_33898_n8095), .Y(REGFILE_SIM_reg_bank__abc_33898_n8099) );
  OR2X2 OR2X2_4267 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8100), .B(REGFILE_SIM_reg_bank__abc_33898_n8101), .Y(REGFILE_SIM_reg_bank__abc_33898_n8102) );
  OR2X2 OR2X2_4268 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8103), .B(REGFILE_SIM_reg_bank__abc_33898_n8104), .Y(REGFILE_SIM_reg_bank__abc_33898_n8105) );
  OR2X2 OR2X2_4269 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8102), .B(REGFILE_SIM_reg_bank__abc_33898_n8105), .Y(REGFILE_SIM_reg_bank__abc_33898_n8106) );
  OR2X2 OR2X2_427 ( .A(_abc_43815_n1883), .B(_abc_43815_n1855), .Y(_abc_43815_n1884) );
  OR2X2 OR2X2_4270 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8099), .B(REGFILE_SIM_reg_bank__abc_33898_n8106), .Y(REGFILE_SIM_reg_bank__abc_33898_n8107) );
  OR2X2 OR2X2_4271 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8108), .B(REGFILE_SIM_reg_bank__abc_33898_n8109), .Y(REGFILE_SIM_reg_bank__abc_33898_n8110) );
  OR2X2 OR2X2_4272 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8111), .B(REGFILE_SIM_reg_bank__abc_33898_n8112), .Y(REGFILE_SIM_reg_bank__abc_33898_n8113) );
  OR2X2 OR2X2_4273 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8110), .B(REGFILE_SIM_reg_bank__abc_33898_n8113), .Y(REGFILE_SIM_reg_bank__abc_33898_n8114) );
  OR2X2 OR2X2_4274 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8115), .B(REGFILE_SIM_reg_bank__abc_33898_n8116), .Y(REGFILE_SIM_reg_bank__abc_33898_n8117) );
  OR2X2 OR2X2_4275 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8118), .B(REGFILE_SIM_reg_bank__abc_33898_n8119), .Y(REGFILE_SIM_reg_bank__abc_33898_n8120) );
  OR2X2 OR2X2_4276 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8120), .B(REGFILE_SIM_reg_bank__abc_33898_n8117), .Y(REGFILE_SIM_reg_bank__abc_33898_n8121) );
  OR2X2 OR2X2_4277 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8114), .B(REGFILE_SIM_reg_bank__abc_33898_n8121), .Y(REGFILE_SIM_reg_bank__abc_33898_n8122) );
  OR2X2 OR2X2_4278 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8107), .B(REGFILE_SIM_reg_bank__abc_33898_n8122), .Y(REGFILE_SIM_reg_bank__abc_33898_n8123) );
  OR2X2 OR2X2_4279 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8124), .B(REGFILE_SIM_reg_bank__abc_33898_n8125), .Y(REGFILE_SIM_reg_bank__abc_33898_n8126) );
  OR2X2 OR2X2_428 ( .A(_abc_43815_n1885), .B(_abc_43815_n1851), .Y(_abc_43815_n1886) );
  OR2X2 OR2X2_4280 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8127), .B(REGFILE_SIM_reg_bank__abc_33898_n8128), .Y(REGFILE_SIM_reg_bank__abc_33898_n8129) );
  OR2X2 OR2X2_4281 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8126), .B(REGFILE_SIM_reg_bank__abc_33898_n8129), .Y(REGFILE_SIM_reg_bank__abc_33898_n8130) );
  OR2X2 OR2X2_4282 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8132), .B(REGFILE_SIM_reg_bank__abc_33898_n8133), .Y(REGFILE_SIM_reg_bank__abc_33898_n8134) );
  OR2X2 OR2X2_4283 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8134), .B(REGFILE_SIM_reg_bank__abc_33898_n8131), .Y(REGFILE_SIM_reg_bank__abc_33898_n8135) );
  OR2X2 OR2X2_4284 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8130), .B(REGFILE_SIM_reg_bank__abc_33898_n8135), .Y(REGFILE_SIM_reg_bank__abc_33898_n8136) );
  OR2X2 OR2X2_4285 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8137), .B(REGFILE_SIM_reg_bank__abc_33898_n8138), .Y(REGFILE_SIM_reg_bank__abc_33898_n8139) );
  OR2X2 OR2X2_4286 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8140), .B(REGFILE_SIM_reg_bank__abc_33898_n8141), .Y(REGFILE_SIM_reg_bank__abc_33898_n8142) );
  OR2X2 OR2X2_4287 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8142), .B(REGFILE_SIM_reg_bank__abc_33898_n8139), .Y(REGFILE_SIM_reg_bank__abc_33898_n8143) );
  OR2X2 OR2X2_4288 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8144), .B(REGFILE_SIM_reg_bank__abc_33898_n8145), .Y(REGFILE_SIM_reg_bank__abc_33898_n8146) );
  OR2X2 OR2X2_4289 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8147), .B(REGFILE_SIM_reg_bank__abc_33898_n8148), .Y(REGFILE_SIM_reg_bank__abc_33898_n8149) );
  OR2X2 OR2X2_429 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_12_), .Y(_abc_43815_n1887) );
  OR2X2 OR2X2_4290 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8146), .B(REGFILE_SIM_reg_bank__abc_33898_n8149), .Y(REGFILE_SIM_reg_bank__abc_33898_n8150) );
  OR2X2 OR2X2_4291 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8143), .B(REGFILE_SIM_reg_bank__abc_33898_n8150), .Y(REGFILE_SIM_reg_bank__abc_33898_n8151) );
  OR2X2 OR2X2_4292 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8151), .B(REGFILE_SIM_reg_bank__abc_33898_n8136), .Y(REGFILE_SIM_reg_bank__abc_33898_n8152) );
  OR2X2 OR2X2_4293 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8123), .B(REGFILE_SIM_reg_bank__abc_33898_n8152), .Y(REGFILE_SIM_reg_bank_reg_ra_o_8_) );
  OR2X2 OR2X2_4294 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8154), .B(REGFILE_SIM_reg_bank__abc_33898_n8155), .Y(REGFILE_SIM_reg_bank__abc_33898_n8156) );
  OR2X2 OR2X2_4295 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8157), .B(REGFILE_SIM_reg_bank__abc_33898_n8158), .Y(REGFILE_SIM_reg_bank__abc_33898_n8159) );
  OR2X2 OR2X2_4296 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8159), .B(REGFILE_SIM_reg_bank__abc_33898_n8156), .Y(REGFILE_SIM_reg_bank__abc_33898_n8160) );
  OR2X2 OR2X2_4297 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8161), .B(REGFILE_SIM_reg_bank__abc_33898_n8162), .Y(REGFILE_SIM_reg_bank__abc_33898_n8163) );
  OR2X2 OR2X2_4298 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8164), .B(REGFILE_SIM_reg_bank__abc_33898_n8165), .Y(REGFILE_SIM_reg_bank__abc_33898_n8166) );
  OR2X2 OR2X2_4299 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8163), .B(REGFILE_SIM_reg_bank__abc_33898_n8166), .Y(REGFILE_SIM_reg_bank__abc_33898_n8167) );
  OR2X2 OR2X2_43 ( .A(_abc_43815_n779), .B(_abc_43815_n780), .Y(_abc_43815_n781_1) );
  OR2X2 OR2X2_430 ( .A(_abc_43815_n1847_1), .B(pc_q_13_), .Y(_abc_43815_n1890) );
  OR2X2 OR2X2_4300 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8160), .B(REGFILE_SIM_reg_bank__abc_33898_n8167), .Y(REGFILE_SIM_reg_bank__abc_33898_n8168) );
  OR2X2 OR2X2_4301 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8169), .B(REGFILE_SIM_reg_bank__abc_33898_n8170), .Y(REGFILE_SIM_reg_bank__abc_33898_n8171) );
  OR2X2 OR2X2_4302 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8172), .B(REGFILE_SIM_reg_bank__abc_33898_n8173), .Y(REGFILE_SIM_reg_bank__abc_33898_n8174) );
  OR2X2 OR2X2_4303 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8171), .B(REGFILE_SIM_reg_bank__abc_33898_n8174), .Y(REGFILE_SIM_reg_bank__abc_33898_n8175) );
  OR2X2 OR2X2_4304 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8176), .B(REGFILE_SIM_reg_bank__abc_33898_n8177), .Y(REGFILE_SIM_reg_bank__abc_33898_n8178) );
  OR2X2 OR2X2_4305 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8179), .B(REGFILE_SIM_reg_bank__abc_33898_n8180), .Y(REGFILE_SIM_reg_bank__abc_33898_n8181) );
  OR2X2 OR2X2_4306 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8181), .B(REGFILE_SIM_reg_bank__abc_33898_n8178), .Y(REGFILE_SIM_reg_bank__abc_33898_n8182) );
  OR2X2 OR2X2_4307 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8175), .B(REGFILE_SIM_reg_bank__abc_33898_n8182), .Y(REGFILE_SIM_reg_bank__abc_33898_n8183) );
  OR2X2 OR2X2_4308 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8168), .B(REGFILE_SIM_reg_bank__abc_33898_n8183), .Y(REGFILE_SIM_reg_bank__abc_33898_n8184) );
  OR2X2 OR2X2_4309 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8185), .B(REGFILE_SIM_reg_bank__abc_33898_n8186), .Y(REGFILE_SIM_reg_bank__abc_33898_n8187) );
  OR2X2 OR2X2_431 ( .A(_abc_43815_n1893), .B(_abc_43815_n1278_bF_buf4), .Y(_abc_43815_n1894) );
  OR2X2 OR2X2_4310 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8188), .B(REGFILE_SIM_reg_bank__abc_33898_n8189), .Y(REGFILE_SIM_reg_bank__abc_33898_n8190) );
  OR2X2 OR2X2_4311 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8187), .B(REGFILE_SIM_reg_bank__abc_33898_n8190), .Y(REGFILE_SIM_reg_bank__abc_33898_n8191) );
  OR2X2 OR2X2_4312 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8193), .B(REGFILE_SIM_reg_bank__abc_33898_n8194), .Y(REGFILE_SIM_reg_bank__abc_33898_n8195) );
  OR2X2 OR2X2_4313 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8195), .B(REGFILE_SIM_reg_bank__abc_33898_n8192), .Y(REGFILE_SIM_reg_bank__abc_33898_n8196) );
  OR2X2 OR2X2_4314 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8191), .B(REGFILE_SIM_reg_bank__abc_33898_n8196), .Y(REGFILE_SIM_reg_bank__abc_33898_n8197) );
  OR2X2 OR2X2_4315 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8198), .B(REGFILE_SIM_reg_bank__abc_33898_n8199), .Y(REGFILE_SIM_reg_bank__abc_33898_n8200) );
  OR2X2 OR2X2_4316 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8201), .B(REGFILE_SIM_reg_bank__abc_33898_n8202), .Y(REGFILE_SIM_reg_bank__abc_33898_n8203) );
  OR2X2 OR2X2_4317 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8203), .B(REGFILE_SIM_reg_bank__abc_33898_n8200), .Y(REGFILE_SIM_reg_bank__abc_33898_n8204) );
  OR2X2 OR2X2_4318 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8205), .B(REGFILE_SIM_reg_bank__abc_33898_n8206), .Y(REGFILE_SIM_reg_bank__abc_33898_n8207) );
  OR2X2 OR2X2_4319 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8208), .B(REGFILE_SIM_reg_bank__abc_33898_n8209), .Y(REGFILE_SIM_reg_bank__abc_33898_n8210) );
  OR2X2 OR2X2_432 ( .A(_abc_43815_n1897), .B(_abc_43815_n1896), .Y(_abc_43815_n1898) );
  OR2X2 OR2X2_4320 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8207), .B(REGFILE_SIM_reg_bank__abc_33898_n8210), .Y(REGFILE_SIM_reg_bank__abc_33898_n8211) );
  OR2X2 OR2X2_4321 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8204), .B(REGFILE_SIM_reg_bank__abc_33898_n8211), .Y(REGFILE_SIM_reg_bank__abc_33898_n8212) );
  OR2X2 OR2X2_4322 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8212), .B(REGFILE_SIM_reg_bank__abc_33898_n8197), .Y(REGFILE_SIM_reg_bank__abc_33898_n8213) );
  OR2X2 OR2X2_4323 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8184), .B(REGFILE_SIM_reg_bank__abc_33898_n8213), .Y(REGFILE_SIM_reg_bank_reg_ra_o_9_) );
  OR2X2 OR2X2_4324 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8215), .B(REGFILE_SIM_reg_bank__abc_33898_n8216), .Y(REGFILE_SIM_reg_bank__abc_33898_n8217) );
  OR2X2 OR2X2_4325 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8218), .B(REGFILE_SIM_reg_bank__abc_33898_n8219), .Y(REGFILE_SIM_reg_bank__abc_33898_n8220) );
  OR2X2 OR2X2_4326 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8220), .B(REGFILE_SIM_reg_bank__abc_33898_n8217), .Y(REGFILE_SIM_reg_bank__abc_33898_n8221) );
  OR2X2 OR2X2_4327 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8222), .B(REGFILE_SIM_reg_bank__abc_33898_n8223), .Y(REGFILE_SIM_reg_bank__abc_33898_n8224) );
  OR2X2 OR2X2_4328 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8225), .B(REGFILE_SIM_reg_bank__abc_33898_n8226), .Y(REGFILE_SIM_reg_bank__abc_33898_n8227) );
  OR2X2 OR2X2_4329 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8224), .B(REGFILE_SIM_reg_bank__abc_33898_n8227), .Y(REGFILE_SIM_reg_bank__abc_33898_n8228) );
  OR2X2 OR2X2_433 ( .A(_abc_43815_n1431_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_43815_n1900) );
  OR2X2 OR2X2_4330 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8221), .B(REGFILE_SIM_reg_bank__abc_33898_n8228), .Y(REGFILE_SIM_reg_bank__abc_33898_n8229) );
  OR2X2 OR2X2_4331 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8230), .B(REGFILE_SIM_reg_bank__abc_33898_n8231), .Y(REGFILE_SIM_reg_bank__abc_33898_n8232) );
  OR2X2 OR2X2_4332 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8233), .B(REGFILE_SIM_reg_bank__abc_33898_n8234), .Y(REGFILE_SIM_reg_bank__abc_33898_n8235) );
  OR2X2 OR2X2_4333 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8232), .B(REGFILE_SIM_reg_bank__abc_33898_n8235), .Y(REGFILE_SIM_reg_bank__abc_33898_n8236) );
  OR2X2 OR2X2_4334 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8237), .B(REGFILE_SIM_reg_bank__abc_33898_n8238), .Y(REGFILE_SIM_reg_bank__abc_33898_n8239) );
  OR2X2 OR2X2_4335 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8240), .B(REGFILE_SIM_reg_bank__abc_33898_n8241), .Y(REGFILE_SIM_reg_bank__abc_33898_n8242) );
  OR2X2 OR2X2_4336 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8242), .B(REGFILE_SIM_reg_bank__abc_33898_n8239), .Y(REGFILE_SIM_reg_bank__abc_33898_n8243) );
  OR2X2 OR2X2_4337 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8236), .B(REGFILE_SIM_reg_bank__abc_33898_n8243), .Y(REGFILE_SIM_reg_bank__abc_33898_n8244) );
  OR2X2 OR2X2_4338 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8229), .B(REGFILE_SIM_reg_bank__abc_33898_n8244), .Y(REGFILE_SIM_reg_bank__abc_33898_n8245) );
  OR2X2 OR2X2_4339 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8246), .B(REGFILE_SIM_reg_bank__abc_33898_n8247), .Y(REGFILE_SIM_reg_bank__abc_33898_n8248) );
  OR2X2 OR2X2_434 ( .A(pc_q_13_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_43815_n1901) );
  OR2X2 OR2X2_4340 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8249), .B(REGFILE_SIM_reg_bank__abc_33898_n8250), .Y(REGFILE_SIM_reg_bank__abc_33898_n8251) );
  OR2X2 OR2X2_4341 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8248), .B(REGFILE_SIM_reg_bank__abc_33898_n8251), .Y(REGFILE_SIM_reg_bank__abc_33898_n8252) );
  OR2X2 OR2X2_4342 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8254), .B(REGFILE_SIM_reg_bank__abc_33898_n8255), .Y(REGFILE_SIM_reg_bank__abc_33898_n8256) );
  OR2X2 OR2X2_4343 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8256), .B(REGFILE_SIM_reg_bank__abc_33898_n8253), .Y(REGFILE_SIM_reg_bank__abc_33898_n8257) );
  OR2X2 OR2X2_4344 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8252), .B(REGFILE_SIM_reg_bank__abc_33898_n8257), .Y(REGFILE_SIM_reg_bank__abc_33898_n8258) );
  OR2X2 OR2X2_4345 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8259), .B(REGFILE_SIM_reg_bank__abc_33898_n8260), .Y(REGFILE_SIM_reg_bank__abc_33898_n8261) );
  OR2X2 OR2X2_4346 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8262), .B(REGFILE_SIM_reg_bank__abc_33898_n8263), .Y(REGFILE_SIM_reg_bank__abc_33898_n8264) );
  OR2X2 OR2X2_4347 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8264), .B(REGFILE_SIM_reg_bank__abc_33898_n8261), .Y(REGFILE_SIM_reg_bank__abc_33898_n8265) );
  OR2X2 OR2X2_4348 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8266), .B(REGFILE_SIM_reg_bank__abc_33898_n8267), .Y(REGFILE_SIM_reg_bank__abc_33898_n8268) );
  OR2X2 OR2X2_4349 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8269), .B(REGFILE_SIM_reg_bank__abc_33898_n8270), .Y(REGFILE_SIM_reg_bank__abc_33898_n8271) );
  OR2X2 OR2X2_435 ( .A(_abc_43815_n1904), .B(_abc_43815_n1868_1), .Y(_abc_43815_n1905) );
  OR2X2 OR2X2_4350 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8268), .B(REGFILE_SIM_reg_bank__abc_33898_n8271), .Y(REGFILE_SIM_reg_bank__abc_33898_n8272) );
  OR2X2 OR2X2_4351 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8265), .B(REGFILE_SIM_reg_bank__abc_33898_n8272), .Y(REGFILE_SIM_reg_bank__abc_33898_n8273) );
  OR2X2 OR2X2_4352 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8273), .B(REGFILE_SIM_reg_bank__abc_33898_n8258), .Y(REGFILE_SIM_reg_bank__abc_33898_n8274) );
  OR2X2 OR2X2_4353 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8245), .B(REGFILE_SIM_reg_bank__abc_33898_n8274), .Y(REGFILE_SIM_reg_bank_reg_ra_o_10_) );
  OR2X2 OR2X2_4354 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8276), .B(REGFILE_SIM_reg_bank__abc_33898_n8277), .Y(REGFILE_SIM_reg_bank__abc_33898_n8278) );
  OR2X2 OR2X2_4355 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8279), .B(REGFILE_SIM_reg_bank__abc_33898_n8280), .Y(REGFILE_SIM_reg_bank__abc_33898_n8281) );
  OR2X2 OR2X2_4356 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8281), .B(REGFILE_SIM_reg_bank__abc_33898_n8278), .Y(REGFILE_SIM_reg_bank__abc_33898_n8282) );
  OR2X2 OR2X2_4357 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8283), .B(REGFILE_SIM_reg_bank__abc_33898_n8284), .Y(REGFILE_SIM_reg_bank__abc_33898_n8285) );
  OR2X2 OR2X2_4358 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8286), .B(REGFILE_SIM_reg_bank__abc_33898_n8287), .Y(REGFILE_SIM_reg_bank__abc_33898_n8288) );
  OR2X2 OR2X2_4359 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8285), .B(REGFILE_SIM_reg_bank__abc_33898_n8288), .Y(REGFILE_SIM_reg_bank__abc_33898_n8289) );
  OR2X2 OR2X2_436 ( .A(_abc_43815_n1871_1), .B(_abc_43815_n1905), .Y(_abc_43815_n1906) );
  OR2X2 OR2X2_4360 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8282), .B(REGFILE_SIM_reg_bank__abc_33898_n8289), .Y(REGFILE_SIM_reg_bank__abc_33898_n8290) );
  OR2X2 OR2X2_4361 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8291), .B(REGFILE_SIM_reg_bank__abc_33898_n8292), .Y(REGFILE_SIM_reg_bank__abc_33898_n8293) );
  OR2X2 OR2X2_4362 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8294), .B(REGFILE_SIM_reg_bank__abc_33898_n8295), .Y(REGFILE_SIM_reg_bank__abc_33898_n8296) );
  OR2X2 OR2X2_4363 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8293), .B(REGFILE_SIM_reg_bank__abc_33898_n8296), .Y(REGFILE_SIM_reg_bank__abc_33898_n8297) );
  OR2X2 OR2X2_4364 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8298), .B(REGFILE_SIM_reg_bank__abc_33898_n8299), .Y(REGFILE_SIM_reg_bank__abc_33898_n8300) );
  OR2X2 OR2X2_4365 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8301), .B(REGFILE_SIM_reg_bank__abc_33898_n8302), .Y(REGFILE_SIM_reg_bank__abc_33898_n8303) );
  OR2X2 OR2X2_4366 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8303), .B(REGFILE_SIM_reg_bank__abc_33898_n8300), .Y(REGFILE_SIM_reg_bank__abc_33898_n8304) );
  OR2X2 OR2X2_4367 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8297), .B(REGFILE_SIM_reg_bank__abc_33898_n8304), .Y(REGFILE_SIM_reg_bank__abc_33898_n8305) );
  OR2X2 OR2X2_4368 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8290), .B(REGFILE_SIM_reg_bank__abc_33898_n8305), .Y(REGFILE_SIM_reg_bank__abc_33898_n8306) );
  OR2X2 OR2X2_4369 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8307), .B(REGFILE_SIM_reg_bank__abc_33898_n8308), .Y(REGFILE_SIM_reg_bank__abc_33898_n8309) );
  OR2X2 OR2X2_437 ( .A(_abc_43815_n1428_bF_buf0), .B(_abc_43815_n1915), .Y(_abc_43815_n1916) );
  OR2X2 OR2X2_4370 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8310), .B(REGFILE_SIM_reg_bank__abc_33898_n8311), .Y(REGFILE_SIM_reg_bank__abc_33898_n8312) );
  OR2X2 OR2X2_4371 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8309), .B(REGFILE_SIM_reg_bank__abc_33898_n8312), .Y(REGFILE_SIM_reg_bank__abc_33898_n8313) );
  OR2X2 OR2X2_4372 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8315), .B(REGFILE_SIM_reg_bank__abc_33898_n8316), .Y(REGFILE_SIM_reg_bank__abc_33898_n8317) );
  OR2X2 OR2X2_4373 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8317), .B(REGFILE_SIM_reg_bank__abc_33898_n8314), .Y(REGFILE_SIM_reg_bank__abc_33898_n8318) );
  OR2X2 OR2X2_4374 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8313), .B(REGFILE_SIM_reg_bank__abc_33898_n8318), .Y(REGFILE_SIM_reg_bank__abc_33898_n8319) );
  OR2X2 OR2X2_4375 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8320), .B(REGFILE_SIM_reg_bank__abc_33898_n8321), .Y(REGFILE_SIM_reg_bank__abc_33898_n8322) );
  OR2X2 OR2X2_4376 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8323), .B(REGFILE_SIM_reg_bank__abc_33898_n8324), .Y(REGFILE_SIM_reg_bank__abc_33898_n8325) );
  OR2X2 OR2X2_4377 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8325), .B(REGFILE_SIM_reg_bank__abc_33898_n8322), .Y(REGFILE_SIM_reg_bank__abc_33898_n8326) );
  OR2X2 OR2X2_4378 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8327), .B(REGFILE_SIM_reg_bank__abc_33898_n8328), .Y(REGFILE_SIM_reg_bank__abc_33898_n8329) );
  OR2X2 OR2X2_4379 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8330), .B(REGFILE_SIM_reg_bank__abc_33898_n8331), .Y(REGFILE_SIM_reg_bank__abc_33898_n8332) );
  OR2X2 OR2X2_438 ( .A(_abc_43815_n1914), .B(_abc_43815_n1916), .Y(_abc_43815_n1917) );
  OR2X2 OR2X2_4380 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8329), .B(REGFILE_SIM_reg_bank__abc_33898_n8332), .Y(REGFILE_SIM_reg_bank__abc_33898_n8333) );
  OR2X2 OR2X2_4381 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8326), .B(REGFILE_SIM_reg_bank__abc_33898_n8333), .Y(REGFILE_SIM_reg_bank__abc_33898_n8334) );
  OR2X2 OR2X2_4382 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8334), .B(REGFILE_SIM_reg_bank__abc_33898_n8319), .Y(REGFILE_SIM_reg_bank__abc_33898_n8335) );
  OR2X2 OR2X2_4383 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8306), .B(REGFILE_SIM_reg_bank__abc_33898_n8335), .Y(REGFILE_SIM_reg_bank_reg_ra_o_11_) );
  OR2X2 OR2X2_4384 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8337), .B(REGFILE_SIM_reg_bank__abc_33898_n8338), .Y(REGFILE_SIM_reg_bank__abc_33898_n8339) );
  OR2X2 OR2X2_4385 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8340), .B(REGFILE_SIM_reg_bank__abc_33898_n8341), .Y(REGFILE_SIM_reg_bank__abc_33898_n8342) );
  OR2X2 OR2X2_4386 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8342), .B(REGFILE_SIM_reg_bank__abc_33898_n8339), .Y(REGFILE_SIM_reg_bank__abc_33898_n8343) );
  OR2X2 OR2X2_4387 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8344), .B(REGFILE_SIM_reg_bank__abc_33898_n8345), .Y(REGFILE_SIM_reg_bank__abc_33898_n8346) );
  OR2X2 OR2X2_4388 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8347), .B(REGFILE_SIM_reg_bank__abc_33898_n8348), .Y(REGFILE_SIM_reg_bank__abc_33898_n8349) );
  OR2X2 OR2X2_4389 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8346), .B(REGFILE_SIM_reg_bank__abc_33898_n8349), .Y(REGFILE_SIM_reg_bank__abc_33898_n8350) );
  OR2X2 OR2X2_439 ( .A(_abc_43815_n1918_1), .B(_abc_43815_n1473_bF_buf3), .Y(_abc_43815_n1919) );
  OR2X2 OR2X2_4390 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8343), .B(REGFILE_SIM_reg_bank__abc_33898_n8350), .Y(REGFILE_SIM_reg_bank__abc_33898_n8351) );
  OR2X2 OR2X2_4391 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8352), .B(REGFILE_SIM_reg_bank__abc_33898_n8353), .Y(REGFILE_SIM_reg_bank__abc_33898_n8354) );
  OR2X2 OR2X2_4392 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8355), .B(REGFILE_SIM_reg_bank__abc_33898_n8356), .Y(REGFILE_SIM_reg_bank__abc_33898_n8357) );
  OR2X2 OR2X2_4393 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8354), .B(REGFILE_SIM_reg_bank__abc_33898_n8357), .Y(REGFILE_SIM_reg_bank__abc_33898_n8358) );
  OR2X2 OR2X2_4394 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8359), .B(REGFILE_SIM_reg_bank__abc_33898_n8360), .Y(REGFILE_SIM_reg_bank__abc_33898_n8361) );
  OR2X2 OR2X2_4395 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8362), .B(REGFILE_SIM_reg_bank__abc_33898_n8363), .Y(REGFILE_SIM_reg_bank__abc_33898_n8364) );
  OR2X2 OR2X2_4396 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8364), .B(REGFILE_SIM_reg_bank__abc_33898_n8361), .Y(REGFILE_SIM_reg_bank__abc_33898_n8365) );
  OR2X2 OR2X2_4397 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8358), .B(REGFILE_SIM_reg_bank__abc_33898_n8365), .Y(REGFILE_SIM_reg_bank__abc_33898_n8366) );
  OR2X2 OR2X2_4398 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8351), .B(REGFILE_SIM_reg_bank__abc_33898_n8366), .Y(REGFILE_SIM_reg_bank__abc_33898_n8367) );
  OR2X2 OR2X2_4399 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8368), .B(REGFILE_SIM_reg_bank__abc_33898_n8369), .Y(REGFILE_SIM_reg_bank__abc_33898_n8370) );
  OR2X2 OR2X2_44 ( .A(_abc_43815_n783), .B(_abc_43815_n784), .Y(_abc_43815_n785) );
  OR2X2 OR2X2_440 ( .A(_abc_43815_n1893), .B(_abc_43815_n1472_1_bF_buf2), .Y(_abc_43815_n1920_1) );
  OR2X2 OR2X2_4400 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8371), .B(REGFILE_SIM_reg_bank__abc_33898_n8372), .Y(REGFILE_SIM_reg_bank__abc_33898_n8373) );
  OR2X2 OR2X2_4401 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8370), .B(REGFILE_SIM_reg_bank__abc_33898_n8373), .Y(REGFILE_SIM_reg_bank__abc_33898_n8374) );
  OR2X2 OR2X2_4402 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8376), .B(REGFILE_SIM_reg_bank__abc_33898_n8377), .Y(REGFILE_SIM_reg_bank__abc_33898_n8378) );
  OR2X2 OR2X2_4403 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8378), .B(REGFILE_SIM_reg_bank__abc_33898_n8375), .Y(REGFILE_SIM_reg_bank__abc_33898_n8379) );
  OR2X2 OR2X2_4404 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8374), .B(REGFILE_SIM_reg_bank__abc_33898_n8379), .Y(REGFILE_SIM_reg_bank__abc_33898_n8380) );
  OR2X2 OR2X2_4405 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8381), .B(REGFILE_SIM_reg_bank__abc_33898_n8382), .Y(REGFILE_SIM_reg_bank__abc_33898_n8383) );
  OR2X2 OR2X2_4406 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8384), .B(REGFILE_SIM_reg_bank__abc_33898_n8385), .Y(REGFILE_SIM_reg_bank__abc_33898_n8386) );
  OR2X2 OR2X2_4407 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8386), .B(REGFILE_SIM_reg_bank__abc_33898_n8383), .Y(REGFILE_SIM_reg_bank__abc_33898_n8387) );
  OR2X2 OR2X2_4408 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8388), .B(REGFILE_SIM_reg_bank__abc_33898_n8389), .Y(REGFILE_SIM_reg_bank__abc_33898_n8390) );
  OR2X2 OR2X2_4409 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8391), .B(REGFILE_SIM_reg_bank__abc_33898_n8392), .Y(REGFILE_SIM_reg_bank__abc_33898_n8393) );
  OR2X2 OR2X2_441 ( .A(_abc_43815_n1922_1), .B(_abc_43815_n1899), .Y(_abc_43815_n1923_1) );
  OR2X2 OR2X2_4410 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8390), .B(REGFILE_SIM_reg_bank__abc_33898_n8393), .Y(REGFILE_SIM_reg_bank__abc_33898_n8394) );
  OR2X2 OR2X2_4411 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8387), .B(REGFILE_SIM_reg_bank__abc_33898_n8394), .Y(REGFILE_SIM_reg_bank__abc_33898_n8395) );
  OR2X2 OR2X2_4412 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8395), .B(REGFILE_SIM_reg_bank__abc_33898_n8380), .Y(REGFILE_SIM_reg_bank__abc_33898_n8396) );
  OR2X2 OR2X2_4413 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8367), .B(REGFILE_SIM_reg_bank__abc_33898_n8396), .Y(REGFILE_SIM_reg_bank_reg_ra_o_12_) );
  OR2X2 OR2X2_4414 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8398), .B(REGFILE_SIM_reg_bank__abc_33898_n8399), .Y(REGFILE_SIM_reg_bank__abc_33898_n8400) );
  OR2X2 OR2X2_4415 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8401), .B(REGFILE_SIM_reg_bank__abc_33898_n8402), .Y(REGFILE_SIM_reg_bank__abc_33898_n8403) );
  OR2X2 OR2X2_4416 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8403), .B(REGFILE_SIM_reg_bank__abc_33898_n8400), .Y(REGFILE_SIM_reg_bank__abc_33898_n8404) );
  OR2X2 OR2X2_4417 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8405), .B(REGFILE_SIM_reg_bank__abc_33898_n8406), .Y(REGFILE_SIM_reg_bank__abc_33898_n8407) );
  OR2X2 OR2X2_4418 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8408), .B(REGFILE_SIM_reg_bank__abc_33898_n8409), .Y(REGFILE_SIM_reg_bank__abc_33898_n8410) );
  OR2X2 OR2X2_4419 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8407), .B(REGFILE_SIM_reg_bank__abc_33898_n8410), .Y(REGFILE_SIM_reg_bank__abc_33898_n8411) );
  OR2X2 OR2X2_442 ( .A(_abc_43815_n1924), .B(_abc_43815_n1895), .Y(_abc_43815_n1925_1) );
  OR2X2 OR2X2_4420 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8404), .B(REGFILE_SIM_reg_bank__abc_33898_n8411), .Y(REGFILE_SIM_reg_bank__abc_33898_n8412) );
  OR2X2 OR2X2_4421 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8413), .B(REGFILE_SIM_reg_bank__abc_33898_n8414), .Y(REGFILE_SIM_reg_bank__abc_33898_n8415) );
  OR2X2 OR2X2_4422 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8416), .B(REGFILE_SIM_reg_bank__abc_33898_n8417), .Y(REGFILE_SIM_reg_bank__abc_33898_n8418) );
  OR2X2 OR2X2_4423 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8415), .B(REGFILE_SIM_reg_bank__abc_33898_n8418), .Y(REGFILE_SIM_reg_bank__abc_33898_n8419) );
  OR2X2 OR2X2_4424 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8420), .B(REGFILE_SIM_reg_bank__abc_33898_n8421), .Y(REGFILE_SIM_reg_bank__abc_33898_n8422) );
  OR2X2 OR2X2_4425 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8423), .B(REGFILE_SIM_reg_bank__abc_33898_n8424), .Y(REGFILE_SIM_reg_bank__abc_33898_n8425) );
  OR2X2 OR2X2_4426 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8425), .B(REGFILE_SIM_reg_bank__abc_33898_n8422), .Y(REGFILE_SIM_reg_bank__abc_33898_n8426) );
  OR2X2 OR2X2_4427 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8419), .B(REGFILE_SIM_reg_bank__abc_33898_n8426), .Y(REGFILE_SIM_reg_bank__abc_33898_n8427) );
  OR2X2 OR2X2_4428 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8412), .B(REGFILE_SIM_reg_bank__abc_33898_n8427), .Y(REGFILE_SIM_reg_bank__abc_33898_n8428) );
  OR2X2 OR2X2_4429 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8429), .B(REGFILE_SIM_reg_bank__abc_33898_n8430), .Y(REGFILE_SIM_reg_bank__abc_33898_n8431) );
  OR2X2 OR2X2_443 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_13_), .Y(_abc_43815_n1926) );
  OR2X2 OR2X2_4430 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8432), .B(REGFILE_SIM_reg_bank__abc_33898_n8433), .Y(REGFILE_SIM_reg_bank__abc_33898_n8434) );
  OR2X2 OR2X2_4431 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8431), .B(REGFILE_SIM_reg_bank__abc_33898_n8434), .Y(REGFILE_SIM_reg_bank__abc_33898_n8435) );
  OR2X2 OR2X2_4432 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8437), .B(REGFILE_SIM_reg_bank__abc_33898_n8438), .Y(REGFILE_SIM_reg_bank__abc_33898_n8439) );
  OR2X2 OR2X2_4433 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8439), .B(REGFILE_SIM_reg_bank__abc_33898_n8436), .Y(REGFILE_SIM_reg_bank__abc_33898_n8440) );
  OR2X2 OR2X2_4434 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8435), .B(REGFILE_SIM_reg_bank__abc_33898_n8440), .Y(REGFILE_SIM_reg_bank__abc_33898_n8441) );
  OR2X2 OR2X2_4435 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8442), .B(REGFILE_SIM_reg_bank__abc_33898_n8443), .Y(REGFILE_SIM_reg_bank__abc_33898_n8444) );
  OR2X2 OR2X2_4436 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8445), .B(REGFILE_SIM_reg_bank__abc_33898_n8446), .Y(REGFILE_SIM_reg_bank__abc_33898_n8447) );
  OR2X2 OR2X2_4437 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8447), .B(REGFILE_SIM_reg_bank__abc_33898_n8444), .Y(REGFILE_SIM_reg_bank__abc_33898_n8448) );
  OR2X2 OR2X2_4438 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8449), .B(REGFILE_SIM_reg_bank__abc_33898_n8450), .Y(REGFILE_SIM_reg_bank__abc_33898_n8451) );
  OR2X2 OR2X2_4439 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8452), .B(REGFILE_SIM_reg_bank__abc_33898_n8453), .Y(REGFILE_SIM_reg_bank__abc_33898_n8454) );
  OR2X2 OR2X2_444 ( .A(_abc_43815_n1891), .B(pc_q_14_), .Y(_abc_43815_n1929) );
  OR2X2 OR2X2_4440 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8451), .B(REGFILE_SIM_reg_bank__abc_33898_n8454), .Y(REGFILE_SIM_reg_bank__abc_33898_n8455) );
  OR2X2 OR2X2_4441 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8448), .B(REGFILE_SIM_reg_bank__abc_33898_n8455), .Y(REGFILE_SIM_reg_bank__abc_33898_n8456) );
  OR2X2 OR2X2_4442 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8456), .B(REGFILE_SIM_reg_bank__abc_33898_n8441), .Y(REGFILE_SIM_reg_bank__abc_33898_n8457) );
  OR2X2 OR2X2_4443 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8428), .B(REGFILE_SIM_reg_bank__abc_33898_n8457), .Y(REGFILE_SIM_reg_bank_reg_ra_o_13_) );
  OR2X2 OR2X2_4444 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8459), .B(REGFILE_SIM_reg_bank__abc_33898_n8460), .Y(REGFILE_SIM_reg_bank__abc_33898_n8461) );
  OR2X2 OR2X2_4445 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8462), .B(REGFILE_SIM_reg_bank__abc_33898_n8463), .Y(REGFILE_SIM_reg_bank__abc_33898_n8464) );
  OR2X2 OR2X2_4446 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8464), .B(REGFILE_SIM_reg_bank__abc_33898_n8461), .Y(REGFILE_SIM_reg_bank__abc_33898_n8465) );
  OR2X2 OR2X2_4447 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8466), .B(REGFILE_SIM_reg_bank__abc_33898_n8467), .Y(REGFILE_SIM_reg_bank__abc_33898_n8468) );
  OR2X2 OR2X2_4448 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8469), .B(REGFILE_SIM_reg_bank__abc_33898_n8470), .Y(REGFILE_SIM_reg_bank__abc_33898_n8471) );
  OR2X2 OR2X2_4449 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8468), .B(REGFILE_SIM_reg_bank__abc_33898_n8471), .Y(REGFILE_SIM_reg_bank__abc_33898_n8472) );
  OR2X2 OR2X2_445 ( .A(_abc_43815_n1932), .B(_abc_43815_n1278_bF_buf3), .Y(_abc_43815_n1933) );
  OR2X2 OR2X2_4450 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8465), .B(REGFILE_SIM_reg_bank__abc_33898_n8472), .Y(REGFILE_SIM_reg_bank__abc_33898_n8473) );
  OR2X2 OR2X2_4451 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8474), .B(REGFILE_SIM_reg_bank__abc_33898_n8475), .Y(REGFILE_SIM_reg_bank__abc_33898_n8476) );
  OR2X2 OR2X2_4452 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8477), .B(REGFILE_SIM_reg_bank__abc_33898_n8478), .Y(REGFILE_SIM_reg_bank__abc_33898_n8479) );
  OR2X2 OR2X2_4453 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8476), .B(REGFILE_SIM_reg_bank__abc_33898_n8479), .Y(REGFILE_SIM_reg_bank__abc_33898_n8480) );
  OR2X2 OR2X2_4454 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8481), .B(REGFILE_SIM_reg_bank__abc_33898_n8482), .Y(REGFILE_SIM_reg_bank__abc_33898_n8483) );
  OR2X2 OR2X2_4455 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8484), .B(REGFILE_SIM_reg_bank__abc_33898_n8485), .Y(REGFILE_SIM_reg_bank__abc_33898_n8486) );
  OR2X2 OR2X2_4456 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8486), .B(REGFILE_SIM_reg_bank__abc_33898_n8483), .Y(REGFILE_SIM_reg_bank__abc_33898_n8487) );
  OR2X2 OR2X2_4457 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8480), .B(REGFILE_SIM_reg_bank__abc_33898_n8487), .Y(REGFILE_SIM_reg_bank__abc_33898_n8488) );
  OR2X2 OR2X2_4458 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8473), .B(REGFILE_SIM_reg_bank__abc_33898_n8488), .Y(REGFILE_SIM_reg_bank__abc_33898_n8489) );
  OR2X2 OR2X2_4459 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8490), .B(REGFILE_SIM_reg_bank__abc_33898_n8491), .Y(REGFILE_SIM_reg_bank__abc_33898_n8492) );
  OR2X2 OR2X2_446 ( .A(_abc_43815_n1936), .B(_abc_43815_n1935), .Y(_abc_43815_n1937) );
  OR2X2 OR2X2_4460 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8493), .B(REGFILE_SIM_reg_bank__abc_33898_n8494), .Y(REGFILE_SIM_reg_bank__abc_33898_n8495) );
  OR2X2 OR2X2_4461 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8492), .B(REGFILE_SIM_reg_bank__abc_33898_n8495), .Y(REGFILE_SIM_reg_bank__abc_33898_n8496) );
  OR2X2 OR2X2_4462 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8498), .B(REGFILE_SIM_reg_bank__abc_33898_n8499), .Y(REGFILE_SIM_reg_bank__abc_33898_n8500) );
  OR2X2 OR2X2_4463 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8500), .B(REGFILE_SIM_reg_bank__abc_33898_n8497), .Y(REGFILE_SIM_reg_bank__abc_33898_n8501) );
  OR2X2 OR2X2_4464 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8496), .B(REGFILE_SIM_reg_bank__abc_33898_n8501), .Y(REGFILE_SIM_reg_bank__abc_33898_n8502) );
  OR2X2 OR2X2_4465 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8503), .B(REGFILE_SIM_reg_bank__abc_33898_n8504), .Y(REGFILE_SIM_reg_bank__abc_33898_n8505) );
  OR2X2 OR2X2_4466 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8506), .B(REGFILE_SIM_reg_bank__abc_33898_n8507), .Y(REGFILE_SIM_reg_bank__abc_33898_n8508) );
  OR2X2 OR2X2_4467 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8508), .B(REGFILE_SIM_reg_bank__abc_33898_n8505), .Y(REGFILE_SIM_reg_bank__abc_33898_n8509) );
  OR2X2 OR2X2_4468 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8510), .B(REGFILE_SIM_reg_bank__abc_33898_n8511), .Y(REGFILE_SIM_reg_bank__abc_33898_n8512) );
  OR2X2 OR2X2_4469 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8513), .B(REGFILE_SIM_reg_bank__abc_33898_n8514), .Y(REGFILE_SIM_reg_bank__abc_33898_n8515) );
  OR2X2 OR2X2_447 ( .A(_abc_43815_n1431_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_43815_n1939) );
  OR2X2 OR2X2_4470 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8512), .B(REGFILE_SIM_reg_bank__abc_33898_n8515), .Y(REGFILE_SIM_reg_bank__abc_33898_n8516) );
  OR2X2 OR2X2_4471 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8509), .B(REGFILE_SIM_reg_bank__abc_33898_n8516), .Y(REGFILE_SIM_reg_bank__abc_33898_n8517) );
  OR2X2 OR2X2_4472 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8517), .B(REGFILE_SIM_reg_bank__abc_33898_n8502), .Y(REGFILE_SIM_reg_bank__abc_33898_n8518) );
  OR2X2 OR2X2_4473 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8489), .B(REGFILE_SIM_reg_bank__abc_33898_n8518), .Y(REGFILE_SIM_reg_bank_reg_ra_o_14_) );
  OR2X2 OR2X2_4474 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8520), .B(REGFILE_SIM_reg_bank__abc_33898_n8521), .Y(REGFILE_SIM_reg_bank__abc_33898_n8522) );
  OR2X2 OR2X2_4475 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8523), .B(REGFILE_SIM_reg_bank__abc_33898_n8524), .Y(REGFILE_SIM_reg_bank__abc_33898_n8525) );
  OR2X2 OR2X2_4476 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8525), .B(REGFILE_SIM_reg_bank__abc_33898_n8522), .Y(REGFILE_SIM_reg_bank__abc_33898_n8526) );
  OR2X2 OR2X2_4477 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8527), .B(REGFILE_SIM_reg_bank__abc_33898_n8528), .Y(REGFILE_SIM_reg_bank__abc_33898_n8529) );
  OR2X2 OR2X2_4478 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8530), .B(REGFILE_SIM_reg_bank__abc_33898_n8531), .Y(REGFILE_SIM_reg_bank__abc_33898_n8532) );
  OR2X2 OR2X2_4479 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8529), .B(REGFILE_SIM_reg_bank__abc_33898_n8532), .Y(REGFILE_SIM_reg_bank__abc_33898_n8533) );
  OR2X2 OR2X2_448 ( .A(pc_q_14_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_43815_n1943) );
  OR2X2 OR2X2_4480 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8526), .B(REGFILE_SIM_reg_bank__abc_33898_n8533), .Y(REGFILE_SIM_reg_bank__abc_33898_n8534) );
  OR2X2 OR2X2_4481 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8535), .B(REGFILE_SIM_reg_bank__abc_33898_n8536), .Y(REGFILE_SIM_reg_bank__abc_33898_n8537) );
  OR2X2 OR2X2_4482 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8538), .B(REGFILE_SIM_reg_bank__abc_33898_n8539), .Y(REGFILE_SIM_reg_bank__abc_33898_n8540) );
  OR2X2 OR2X2_4483 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8537), .B(REGFILE_SIM_reg_bank__abc_33898_n8540), .Y(REGFILE_SIM_reg_bank__abc_33898_n8541) );
  OR2X2 OR2X2_4484 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8542), .B(REGFILE_SIM_reg_bank__abc_33898_n8543), .Y(REGFILE_SIM_reg_bank__abc_33898_n8544) );
  OR2X2 OR2X2_4485 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8545), .B(REGFILE_SIM_reg_bank__abc_33898_n8546), .Y(REGFILE_SIM_reg_bank__abc_33898_n8547) );
  OR2X2 OR2X2_4486 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8547), .B(REGFILE_SIM_reg_bank__abc_33898_n8544), .Y(REGFILE_SIM_reg_bank__abc_33898_n8548) );
  OR2X2 OR2X2_4487 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8541), .B(REGFILE_SIM_reg_bank__abc_33898_n8548), .Y(REGFILE_SIM_reg_bank__abc_33898_n8549) );
  OR2X2 OR2X2_4488 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8534), .B(REGFILE_SIM_reg_bank__abc_33898_n8549), .Y(REGFILE_SIM_reg_bank__abc_33898_n8550) );
  OR2X2 OR2X2_4489 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8551), .B(REGFILE_SIM_reg_bank__abc_33898_n8552), .Y(REGFILE_SIM_reg_bank__abc_33898_n8553) );
  OR2X2 OR2X2_449 ( .A(_abc_43815_n1942), .B(_abc_43815_n1946), .Y(_abc_43815_n1949) );
  OR2X2 OR2X2_4490 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8554), .B(REGFILE_SIM_reg_bank__abc_33898_n8555), .Y(REGFILE_SIM_reg_bank__abc_33898_n8556) );
  OR2X2 OR2X2_4491 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8553), .B(REGFILE_SIM_reg_bank__abc_33898_n8556), .Y(REGFILE_SIM_reg_bank__abc_33898_n8557) );
  OR2X2 OR2X2_4492 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8559), .B(REGFILE_SIM_reg_bank__abc_33898_n8560), .Y(REGFILE_SIM_reg_bank__abc_33898_n8561) );
  OR2X2 OR2X2_4493 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8561), .B(REGFILE_SIM_reg_bank__abc_33898_n8558), .Y(REGFILE_SIM_reg_bank__abc_33898_n8562) );
  OR2X2 OR2X2_4494 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8557), .B(REGFILE_SIM_reg_bank__abc_33898_n8562), .Y(REGFILE_SIM_reg_bank__abc_33898_n8563) );
  OR2X2 OR2X2_4495 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8564), .B(REGFILE_SIM_reg_bank__abc_33898_n8565), .Y(REGFILE_SIM_reg_bank__abc_33898_n8566) );
  OR2X2 OR2X2_4496 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8567), .B(REGFILE_SIM_reg_bank__abc_33898_n8568), .Y(REGFILE_SIM_reg_bank__abc_33898_n8569) );
  OR2X2 OR2X2_4497 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8569), .B(REGFILE_SIM_reg_bank__abc_33898_n8566), .Y(REGFILE_SIM_reg_bank__abc_33898_n8570) );
  OR2X2 OR2X2_4498 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8571), .B(REGFILE_SIM_reg_bank__abc_33898_n8572), .Y(REGFILE_SIM_reg_bank__abc_33898_n8573) );
  OR2X2 OR2X2_4499 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8574), .B(REGFILE_SIM_reg_bank__abc_33898_n8575), .Y(REGFILE_SIM_reg_bank__abc_33898_n8576) );
  OR2X2 OR2X2_45 ( .A(_abc_43815_n786), .B(_abc_43815_n787), .Y(_abc_43815_n788) );
  OR2X2 OR2X2_450 ( .A(_abc_43815_n1428_bF_buf4), .B(_abc_43815_n1952), .Y(_abc_43815_n1953) );
  OR2X2 OR2X2_4500 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8573), .B(REGFILE_SIM_reg_bank__abc_33898_n8576), .Y(REGFILE_SIM_reg_bank__abc_33898_n8577) );
  OR2X2 OR2X2_4501 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8570), .B(REGFILE_SIM_reg_bank__abc_33898_n8577), .Y(REGFILE_SIM_reg_bank__abc_33898_n8578) );
  OR2X2 OR2X2_4502 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8578), .B(REGFILE_SIM_reg_bank__abc_33898_n8563), .Y(REGFILE_SIM_reg_bank__abc_33898_n8579) );
  OR2X2 OR2X2_4503 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8550), .B(REGFILE_SIM_reg_bank__abc_33898_n8579), .Y(REGFILE_SIM_reg_bank_reg_ra_o_15_) );
  OR2X2 OR2X2_4504 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8581), .B(REGFILE_SIM_reg_bank__abc_33898_n8582), .Y(REGFILE_SIM_reg_bank__abc_33898_n8583) );
  OR2X2 OR2X2_4505 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8584), .B(REGFILE_SIM_reg_bank__abc_33898_n8585), .Y(REGFILE_SIM_reg_bank__abc_33898_n8586) );
  OR2X2 OR2X2_4506 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8586), .B(REGFILE_SIM_reg_bank__abc_33898_n8583), .Y(REGFILE_SIM_reg_bank__abc_33898_n8587) );
  OR2X2 OR2X2_4507 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8588), .B(REGFILE_SIM_reg_bank__abc_33898_n8589), .Y(REGFILE_SIM_reg_bank__abc_33898_n8590) );
  OR2X2 OR2X2_4508 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8591), .B(REGFILE_SIM_reg_bank__abc_33898_n8592), .Y(REGFILE_SIM_reg_bank__abc_33898_n8593) );
  OR2X2 OR2X2_4509 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8590), .B(REGFILE_SIM_reg_bank__abc_33898_n8593), .Y(REGFILE_SIM_reg_bank__abc_33898_n8594) );
  OR2X2 OR2X2_451 ( .A(_abc_43815_n1951), .B(_abc_43815_n1953), .Y(_abc_43815_n1954_1) );
  OR2X2 OR2X2_4510 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8587), .B(REGFILE_SIM_reg_bank__abc_33898_n8594), .Y(REGFILE_SIM_reg_bank__abc_33898_n8595) );
  OR2X2 OR2X2_4511 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8596), .B(REGFILE_SIM_reg_bank__abc_33898_n8597), .Y(REGFILE_SIM_reg_bank__abc_33898_n8598) );
  OR2X2 OR2X2_4512 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8599), .B(REGFILE_SIM_reg_bank__abc_33898_n8600), .Y(REGFILE_SIM_reg_bank__abc_33898_n8601) );
  OR2X2 OR2X2_4513 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8598), .B(REGFILE_SIM_reg_bank__abc_33898_n8601), .Y(REGFILE_SIM_reg_bank__abc_33898_n8602) );
  OR2X2 OR2X2_4514 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8603), .B(REGFILE_SIM_reg_bank__abc_33898_n8604), .Y(REGFILE_SIM_reg_bank__abc_33898_n8605) );
  OR2X2 OR2X2_4515 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8606), .B(REGFILE_SIM_reg_bank__abc_33898_n8607), .Y(REGFILE_SIM_reg_bank__abc_33898_n8608) );
  OR2X2 OR2X2_4516 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8608), .B(REGFILE_SIM_reg_bank__abc_33898_n8605), .Y(REGFILE_SIM_reg_bank__abc_33898_n8609) );
  OR2X2 OR2X2_4517 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8602), .B(REGFILE_SIM_reg_bank__abc_33898_n8609), .Y(REGFILE_SIM_reg_bank__abc_33898_n8610) );
  OR2X2 OR2X2_4518 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8595), .B(REGFILE_SIM_reg_bank__abc_33898_n8610), .Y(REGFILE_SIM_reg_bank__abc_33898_n8611) );
  OR2X2 OR2X2_4519 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8612), .B(REGFILE_SIM_reg_bank__abc_33898_n8613), .Y(REGFILE_SIM_reg_bank__abc_33898_n8614) );
  OR2X2 OR2X2_452 ( .A(_abc_43815_n1955), .B(_abc_43815_n1473_bF_buf2), .Y(_abc_43815_n1956) );
  OR2X2 OR2X2_4520 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8615), .B(REGFILE_SIM_reg_bank__abc_33898_n8616), .Y(REGFILE_SIM_reg_bank__abc_33898_n8617) );
  OR2X2 OR2X2_4521 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8614), .B(REGFILE_SIM_reg_bank__abc_33898_n8617), .Y(REGFILE_SIM_reg_bank__abc_33898_n8618) );
  OR2X2 OR2X2_4522 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8620), .B(REGFILE_SIM_reg_bank__abc_33898_n8621), .Y(REGFILE_SIM_reg_bank__abc_33898_n8622) );
  OR2X2 OR2X2_4523 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8622), .B(REGFILE_SIM_reg_bank__abc_33898_n8619), .Y(REGFILE_SIM_reg_bank__abc_33898_n8623) );
  OR2X2 OR2X2_4524 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8618), .B(REGFILE_SIM_reg_bank__abc_33898_n8623), .Y(REGFILE_SIM_reg_bank__abc_33898_n8624) );
  OR2X2 OR2X2_4525 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8625), .B(REGFILE_SIM_reg_bank__abc_33898_n8626), .Y(REGFILE_SIM_reg_bank__abc_33898_n8627) );
  OR2X2 OR2X2_4526 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8628), .B(REGFILE_SIM_reg_bank__abc_33898_n8629), .Y(REGFILE_SIM_reg_bank__abc_33898_n8630) );
  OR2X2 OR2X2_4527 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8630), .B(REGFILE_SIM_reg_bank__abc_33898_n8627), .Y(REGFILE_SIM_reg_bank__abc_33898_n8631) );
  OR2X2 OR2X2_4528 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8632), .B(REGFILE_SIM_reg_bank__abc_33898_n8633), .Y(REGFILE_SIM_reg_bank__abc_33898_n8634) );
  OR2X2 OR2X2_4529 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8635), .B(REGFILE_SIM_reg_bank__abc_33898_n8636), .Y(REGFILE_SIM_reg_bank__abc_33898_n8637) );
  OR2X2 OR2X2_453 ( .A(_abc_43815_n1932), .B(_abc_43815_n1472_1_bF_buf1), .Y(_abc_43815_n1957) );
  OR2X2 OR2X2_4530 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8634), .B(REGFILE_SIM_reg_bank__abc_33898_n8637), .Y(REGFILE_SIM_reg_bank__abc_33898_n8638) );
  OR2X2 OR2X2_4531 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8631), .B(REGFILE_SIM_reg_bank__abc_33898_n8638), .Y(REGFILE_SIM_reg_bank__abc_33898_n8639) );
  OR2X2 OR2X2_4532 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8639), .B(REGFILE_SIM_reg_bank__abc_33898_n8624), .Y(REGFILE_SIM_reg_bank__abc_33898_n8640) );
  OR2X2 OR2X2_4533 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8611), .B(REGFILE_SIM_reg_bank__abc_33898_n8640), .Y(REGFILE_SIM_reg_bank_reg_ra_o_16_) );
  OR2X2 OR2X2_4534 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8642), .B(REGFILE_SIM_reg_bank__abc_33898_n8643), .Y(REGFILE_SIM_reg_bank__abc_33898_n8644) );
  OR2X2 OR2X2_4535 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8645), .B(REGFILE_SIM_reg_bank__abc_33898_n8646), .Y(REGFILE_SIM_reg_bank__abc_33898_n8647) );
  OR2X2 OR2X2_4536 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8647), .B(REGFILE_SIM_reg_bank__abc_33898_n8644), .Y(REGFILE_SIM_reg_bank__abc_33898_n8648) );
  OR2X2 OR2X2_4537 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8649), .B(REGFILE_SIM_reg_bank__abc_33898_n8650), .Y(REGFILE_SIM_reg_bank__abc_33898_n8651) );
  OR2X2 OR2X2_4538 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8652), .B(REGFILE_SIM_reg_bank__abc_33898_n8653), .Y(REGFILE_SIM_reg_bank__abc_33898_n8654) );
  OR2X2 OR2X2_4539 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8651), .B(REGFILE_SIM_reg_bank__abc_33898_n8654), .Y(REGFILE_SIM_reg_bank__abc_33898_n8655) );
  OR2X2 OR2X2_454 ( .A(_abc_43815_n1959), .B(_abc_43815_n1938), .Y(_abc_43815_n1960) );
  OR2X2 OR2X2_4540 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8648), .B(REGFILE_SIM_reg_bank__abc_33898_n8655), .Y(REGFILE_SIM_reg_bank__abc_33898_n8656) );
  OR2X2 OR2X2_4541 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8657), .B(REGFILE_SIM_reg_bank__abc_33898_n8658), .Y(REGFILE_SIM_reg_bank__abc_33898_n8659) );
  OR2X2 OR2X2_4542 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8660), .B(REGFILE_SIM_reg_bank__abc_33898_n8661), .Y(REGFILE_SIM_reg_bank__abc_33898_n8662) );
  OR2X2 OR2X2_4543 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8659), .B(REGFILE_SIM_reg_bank__abc_33898_n8662), .Y(REGFILE_SIM_reg_bank__abc_33898_n8663) );
  OR2X2 OR2X2_4544 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8664), .B(REGFILE_SIM_reg_bank__abc_33898_n8665), .Y(REGFILE_SIM_reg_bank__abc_33898_n8666) );
  OR2X2 OR2X2_4545 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8667), .B(REGFILE_SIM_reg_bank__abc_33898_n8668), .Y(REGFILE_SIM_reg_bank__abc_33898_n8669) );
  OR2X2 OR2X2_4546 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8669), .B(REGFILE_SIM_reg_bank__abc_33898_n8666), .Y(REGFILE_SIM_reg_bank__abc_33898_n8670) );
  OR2X2 OR2X2_4547 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8663), .B(REGFILE_SIM_reg_bank__abc_33898_n8670), .Y(REGFILE_SIM_reg_bank__abc_33898_n8671) );
  OR2X2 OR2X2_4548 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8656), .B(REGFILE_SIM_reg_bank__abc_33898_n8671), .Y(REGFILE_SIM_reg_bank__abc_33898_n8672) );
  OR2X2 OR2X2_4549 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8673), .B(REGFILE_SIM_reg_bank__abc_33898_n8674), .Y(REGFILE_SIM_reg_bank__abc_33898_n8675) );
  OR2X2 OR2X2_455 ( .A(_abc_43815_n1961), .B(_abc_43815_n1934), .Y(_abc_43815_n1962) );
  OR2X2 OR2X2_4550 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8676), .B(REGFILE_SIM_reg_bank__abc_33898_n8677), .Y(REGFILE_SIM_reg_bank__abc_33898_n8678) );
  OR2X2 OR2X2_4551 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8675), .B(REGFILE_SIM_reg_bank__abc_33898_n8678), .Y(REGFILE_SIM_reg_bank__abc_33898_n8679) );
  OR2X2 OR2X2_4552 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8681), .B(REGFILE_SIM_reg_bank__abc_33898_n8682), .Y(REGFILE_SIM_reg_bank__abc_33898_n8683) );
  OR2X2 OR2X2_4553 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8683), .B(REGFILE_SIM_reg_bank__abc_33898_n8680), .Y(REGFILE_SIM_reg_bank__abc_33898_n8684) );
  OR2X2 OR2X2_4554 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8679), .B(REGFILE_SIM_reg_bank__abc_33898_n8684), .Y(REGFILE_SIM_reg_bank__abc_33898_n8685) );
  OR2X2 OR2X2_4555 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8686), .B(REGFILE_SIM_reg_bank__abc_33898_n8687), .Y(REGFILE_SIM_reg_bank__abc_33898_n8688) );
  OR2X2 OR2X2_4556 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8689), .B(REGFILE_SIM_reg_bank__abc_33898_n8690), .Y(REGFILE_SIM_reg_bank__abc_33898_n8691) );
  OR2X2 OR2X2_4557 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8691), .B(REGFILE_SIM_reg_bank__abc_33898_n8688), .Y(REGFILE_SIM_reg_bank__abc_33898_n8692) );
  OR2X2 OR2X2_4558 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8693), .B(REGFILE_SIM_reg_bank__abc_33898_n8694), .Y(REGFILE_SIM_reg_bank__abc_33898_n8695) );
  OR2X2 OR2X2_4559 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8696), .B(REGFILE_SIM_reg_bank__abc_33898_n8697), .Y(REGFILE_SIM_reg_bank__abc_33898_n8698) );
  OR2X2 OR2X2_456 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_14_), .Y(_abc_43815_n1963) );
  OR2X2 OR2X2_4560 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8695), .B(REGFILE_SIM_reg_bank__abc_33898_n8698), .Y(REGFILE_SIM_reg_bank__abc_33898_n8699) );
  OR2X2 OR2X2_4561 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8692), .B(REGFILE_SIM_reg_bank__abc_33898_n8699), .Y(REGFILE_SIM_reg_bank__abc_33898_n8700) );
  OR2X2 OR2X2_4562 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8700), .B(REGFILE_SIM_reg_bank__abc_33898_n8685), .Y(REGFILE_SIM_reg_bank__abc_33898_n8701) );
  OR2X2 OR2X2_4563 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8672), .B(REGFILE_SIM_reg_bank__abc_33898_n8701), .Y(REGFILE_SIM_reg_bank_reg_ra_o_17_) );
  OR2X2 OR2X2_4564 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8703), .B(REGFILE_SIM_reg_bank__abc_33898_n8704), .Y(REGFILE_SIM_reg_bank__abc_33898_n8705) );
  OR2X2 OR2X2_4565 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8706), .B(REGFILE_SIM_reg_bank__abc_33898_n8707), .Y(REGFILE_SIM_reg_bank__abc_33898_n8708) );
  OR2X2 OR2X2_4566 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8708), .B(REGFILE_SIM_reg_bank__abc_33898_n8705), .Y(REGFILE_SIM_reg_bank__abc_33898_n8709) );
  OR2X2 OR2X2_4567 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8710), .B(REGFILE_SIM_reg_bank__abc_33898_n8711), .Y(REGFILE_SIM_reg_bank__abc_33898_n8712) );
  OR2X2 OR2X2_4568 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8713), .B(REGFILE_SIM_reg_bank__abc_33898_n8714), .Y(REGFILE_SIM_reg_bank__abc_33898_n8715) );
  OR2X2 OR2X2_4569 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8712), .B(REGFILE_SIM_reg_bank__abc_33898_n8715), .Y(REGFILE_SIM_reg_bank__abc_33898_n8716) );
  OR2X2 OR2X2_457 ( .A(_abc_43815_n1930), .B(pc_q_15_), .Y(_abc_43815_n1966) );
  OR2X2 OR2X2_4570 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8709), .B(REGFILE_SIM_reg_bank__abc_33898_n8716), .Y(REGFILE_SIM_reg_bank__abc_33898_n8717) );
  OR2X2 OR2X2_4571 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8718), .B(REGFILE_SIM_reg_bank__abc_33898_n8719), .Y(REGFILE_SIM_reg_bank__abc_33898_n8720) );
  OR2X2 OR2X2_4572 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8721), .B(REGFILE_SIM_reg_bank__abc_33898_n8722), .Y(REGFILE_SIM_reg_bank__abc_33898_n8723) );
  OR2X2 OR2X2_4573 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8720), .B(REGFILE_SIM_reg_bank__abc_33898_n8723), .Y(REGFILE_SIM_reg_bank__abc_33898_n8724) );
  OR2X2 OR2X2_4574 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8725), .B(REGFILE_SIM_reg_bank__abc_33898_n8726), .Y(REGFILE_SIM_reg_bank__abc_33898_n8727) );
  OR2X2 OR2X2_4575 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8728), .B(REGFILE_SIM_reg_bank__abc_33898_n8729), .Y(REGFILE_SIM_reg_bank__abc_33898_n8730) );
  OR2X2 OR2X2_4576 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8730), .B(REGFILE_SIM_reg_bank__abc_33898_n8727), .Y(REGFILE_SIM_reg_bank__abc_33898_n8731) );
  OR2X2 OR2X2_4577 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8724), .B(REGFILE_SIM_reg_bank__abc_33898_n8731), .Y(REGFILE_SIM_reg_bank__abc_33898_n8732) );
  OR2X2 OR2X2_4578 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8717), .B(REGFILE_SIM_reg_bank__abc_33898_n8732), .Y(REGFILE_SIM_reg_bank__abc_33898_n8733) );
  OR2X2 OR2X2_4579 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8734), .B(REGFILE_SIM_reg_bank__abc_33898_n8735), .Y(REGFILE_SIM_reg_bank__abc_33898_n8736) );
  OR2X2 OR2X2_458 ( .A(_abc_43815_n1969), .B(_abc_43815_n1278_bF_buf2), .Y(_abc_43815_n1970) );
  OR2X2 OR2X2_4580 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8737), .B(REGFILE_SIM_reg_bank__abc_33898_n8738), .Y(REGFILE_SIM_reg_bank__abc_33898_n8739) );
  OR2X2 OR2X2_4581 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8736), .B(REGFILE_SIM_reg_bank__abc_33898_n8739), .Y(REGFILE_SIM_reg_bank__abc_33898_n8740) );
  OR2X2 OR2X2_4582 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8742), .B(REGFILE_SIM_reg_bank__abc_33898_n8743), .Y(REGFILE_SIM_reg_bank__abc_33898_n8744) );
  OR2X2 OR2X2_4583 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8744), .B(REGFILE_SIM_reg_bank__abc_33898_n8741), .Y(REGFILE_SIM_reg_bank__abc_33898_n8745) );
  OR2X2 OR2X2_4584 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8740), .B(REGFILE_SIM_reg_bank__abc_33898_n8745), .Y(REGFILE_SIM_reg_bank__abc_33898_n8746) );
  OR2X2 OR2X2_4585 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8747), .B(REGFILE_SIM_reg_bank__abc_33898_n8748), .Y(REGFILE_SIM_reg_bank__abc_33898_n8749) );
  OR2X2 OR2X2_4586 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8750), .B(REGFILE_SIM_reg_bank__abc_33898_n8751), .Y(REGFILE_SIM_reg_bank__abc_33898_n8752) );
  OR2X2 OR2X2_4587 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8752), .B(REGFILE_SIM_reg_bank__abc_33898_n8749), .Y(REGFILE_SIM_reg_bank__abc_33898_n8753) );
  OR2X2 OR2X2_4588 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8754), .B(REGFILE_SIM_reg_bank__abc_33898_n8755), .Y(REGFILE_SIM_reg_bank__abc_33898_n8756) );
  OR2X2 OR2X2_4589 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8757), .B(REGFILE_SIM_reg_bank__abc_33898_n8758), .Y(REGFILE_SIM_reg_bank__abc_33898_n8759) );
  OR2X2 OR2X2_459 ( .A(pc_q_15_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_43815_n1974_1) );
  OR2X2 OR2X2_4590 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8756), .B(REGFILE_SIM_reg_bank__abc_33898_n8759), .Y(REGFILE_SIM_reg_bank__abc_33898_n8760) );
  OR2X2 OR2X2_4591 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8753), .B(REGFILE_SIM_reg_bank__abc_33898_n8760), .Y(REGFILE_SIM_reg_bank__abc_33898_n8761) );
  OR2X2 OR2X2_4592 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8761), .B(REGFILE_SIM_reg_bank__abc_33898_n8746), .Y(REGFILE_SIM_reg_bank__abc_33898_n8762) );
  OR2X2 OR2X2_4593 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8733), .B(REGFILE_SIM_reg_bank__abc_33898_n8762), .Y(REGFILE_SIM_reg_bank_reg_ra_o_18_) );
  OR2X2 OR2X2_4594 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8764), .B(REGFILE_SIM_reg_bank__abc_33898_n8765), .Y(REGFILE_SIM_reg_bank__abc_33898_n8766) );
  OR2X2 OR2X2_4595 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8767), .B(REGFILE_SIM_reg_bank__abc_33898_n8768), .Y(REGFILE_SIM_reg_bank__abc_33898_n8769) );
  OR2X2 OR2X2_4596 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8769), .B(REGFILE_SIM_reg_bank__abc_33898_n8766), .Y(REGFILE_SIM_reg_bank__abc_33898_n8770) );
  OR2X2 OR2X2_4597 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8771), .B(REGFILE_SIM_reg_bank__abc_33898_n8772), .Y(REGFILE_SIM_reg_bank__abc_33898_n8773) );
  OR2X2 OR2X2_4598 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8774), .B(REGFILE_SIM_reg_bank__abc_33898_n8775), .Y(REGFILE_SIM_reg_bank__abc_33898_n8776) );
  OR2X2 OR2X2_4599 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8773), .B(REGFILE_SIM_reg_bank__abc_33898_n8776), .Y(REGFILE_SIM_reg_bank__abc_33898_n8777) );
  OR2X2 OR2X2_46 ( .A(_abc_43815_n785), .B(_abc_43815_n788), .Y(_abc_43815_n789) );
  OR2X2 OR2X2_460 ( .A(_abc_43815_n1973), .B(_abc_43815_n1977), .Y(_abc_43815_n1978) );
  OR2X2 OR2X2_4600 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8770), .B(REGFILE_SIM_reg_bank__abc_33898_n8777), .Y(REGFILE_SIM_reg_bank__abc_33898_n8778) );
  OR2X2 OR2X2_4601 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8779), .B(REGFILE_SIM_reg_bank__abc_33898_n8780), .Y(REGFILE_SIM_reg_bank__abc_33898_n8781) );
  OR2X2 OR2X2_4602 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8782), .B(REGFILE_SIM_reg_bank__abc_33898_n8783), .Y(REGFILE_SIM_reg_bank__abc_33898_n8784) );
  OR2X2 OR2X2_4603 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8781), .B(REGFILE_SIM_reg_bank__abc_33898_n8784), .Y(REGFILE_SIM_reg_bank__abc_33898_n8785) );
  OR2X2 OR2X2_4604 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8786), .B(REGFILE_SIM_reg_bank__abc_33898_n8787), .Y(REGFILE_SIM_reg_bank__abc_33898_n8788) );
  OR2X2 OR2X2_4605 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8789), .B(REGFILE_SIM_reg_bank__abc_33898_n8790), .Y(REGFILE_SIM_reg_bank__abc_33898_n8791) );
  OR2X2 OR2X2_4606 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8791), .B(REGFILE_SIM_reg_bank__abc_33898_n8788), .Y(REGFILE_SIM_reg_bank__abc_33898_n8792) );
  OR2X2 OR2X2_4607 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8785), .B(REGFILE_SIM_reg_bank__abc_33898_n8792), .Y(REGFILE_SIM_reg_bank__abc_33898_n8793) );
  OR2X2 OR2X2_4608 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8778), .B(REGFILE_SIM_reg_bank__abc_33898_n8793), .Y(REGFILE_SIM_reg_bank__abc_33898_n8794) );
  OR2X2 OR2X2_4609 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8795), .B(REGFILE_SIM_reg_bank__abc_33898_n8796), .Y(REGFILE_SIM_reg_bank__abc_33898_n8797) );
  OR2X2 OR2X2_461 ( .A(_abc_43815_n1972), .B(_abc_43815_n1979), .Y(_abc_43815_n1980) );
  OR2X2 OR2X2_4610 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8798), .B(REGFILE_SIM_reg_bank__abc_33898_n8799), .Y(REGFILE_SIM_reg_bank__abc_33898_n8800) );
  OR2X2 OR2X2_4611 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8797), .B(REGFILE_SIM_reg_bank__abc_33898_n8800), .Y(REGFILE_SIM_reg_bank__abc_33898_n8801) );
  OR2X2 OR2X2_4612 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8803), .B(REGFILE_SIM_reg_bank__abc_33898_n8804), .Y(REGFILE_SIM_reg_bank__abc_33898_n8805) );
  OR2X2 OR2X2_4613 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8805), .B(REGFILE_SIM_reg_bank__abc_33898_n8802), .Y(REGFILE_SIM_reg_bank__abc_33898_n8806) );
  OR2X2 OR2X2_4614 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8801), .B(REGFILE_SIM_reg_bank__abc_33898_n8806), .Y(REGFILE_SIM_reg_bank__abc_33898_n8807) );
  OR2X2 OR2X2_4615 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8808), .B(REGFILE_SIM_reg_bank__abc_33898_n8809), .Y(REGFILE_SIM_reg_bank__abc_33898_n8810) );
  OR2X2 OR2X2_4616 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8811), .B(REGFILE_SIM_reg_bank__abc_33898_n8812), .Y(REGFILE_SIM_reg_bank__abc_33898_n8813) );
  OR2X2 OR2X2_4617 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8813), .B(REGFILE_SIM_reg_bank__abc_33898_n8810), .Y(REGFILE_SIM_reg_bank__abc_33898_n8814) );
  OR2X2 OR2X2_4618 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8815), .B(REGFILE_SIM_reg_bank__abc_33898_n8816), .Y(REGFILE_SIM_reg_bank__abc_33898_n8817) );
  OR2X2 OR2X2_4619 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8818), .B(REGFILE_SIM_reg_bank__abc_33898_n8819), .Y(REGFILE_SIM_reg_bank__abc_33898_n8820) );
  OR2X2 OR2X2_462 ( .A(_abc_43815_n1428_bF_buf3), .B(_abc_43815_n1983), .Y(_abc_43815_n1984) );
  OR2X2 OR2X2_4620 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8817), .B(REGFILE_SIM_reg_bank__abc_33898_n8820), .Y(REGFILE_SIM_reg_bank__abc_33898_n8821) );
  OR2X2 OR2X2_4621 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8814), .B(REGFILE_SIM_reg_bank__abc_33898_n8821), .Y(REGFILE_SIM_reg_bank__abc_33898_n8822) );
  OR2X2 OR2X2_4622 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8822), .B(REGFILE_SIM_reg_bank__abc_33898_n8807), .Y(REGFILE_SIM_reg_bank__abc_33898_n8823) );
  OR2X2 OR2X2_4623 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8794), .B(REGFILE_SIM_reg_bank__abc_33898_n8823), .Y(REGFILE_SIM_reg_bank_reg_ra_o_19_) );
  OR2X2 OR2X2_4624 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8825), .B(REGFILE_SIM_reg_bank__abc_33898_n8826), .Y(REGFILE_SIM_reg_bank__abc_33898_n8827) );
  OR2X2 OR2X2_4625 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8828), .B(REGFILE_SIM_reg_bank__abc_33898_n8829), .Y(REGFILE_SIM_reg_bank__abc_33898_n8830) );
  OR2X2 OR2X2_4626 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8830), .B(REGFILE_SIM_reg_bank__abc_33898_n8827), .Y(REGFILE_SIM_reg_bank__abc_33898_n8831) );
  OR2X2 OR2X2_4627 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8832), .B(REGFILE_SIM_reg_bank__abc_33898_n8833), .Y(REGFILE_SIM_reg_bank__abc_33898_n8834) );
  OR2X2 OR2X2_4628 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8835), .B(REGFILE_SIM_reg_bank__abc_33898_n8836), .Y(REGFILE_SIM_reg_bank__abc_33898_n8837) );
  OR2X2 OR2X2_4629 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8834), .B(REGFILE_SIM_reg_bank__abc_33898_n8837), .Y(REGFILE_SIM_reg_bank__abc_33898_n8838) );
  OR2X2 OR2X2_463 ( .A(_abc_43815_n1982), .B(_abc_43815_n1984), .Y(_abc_43815_n1985) );
  OR2X2 OR2X2_4630 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8831), .B(REGFILE_SIM_reg_bank__abc_33898_n8838), .Y(REGFILE_SIM_reg_bank__abc_33898_n8839) );
  OR2X2 OR2X2_4631 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8840), .B(REGFILE_SIM_reg_bank__abc_33898_n8841), .Y(REGFILE_SIM_reg_bank__abc_33898_n8842) );
  OR2X2 OR2X2_4632 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8843), .B(REGFILE_SIM_reg_bank__abc_33898_n8844), .Y(REGFILE_SIM_reg_bank__abc_33898_n8845) );
  OR2X2 OR2X2_4633 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8842), .B(REGFILE_SIM_reg_bank__abc_33898_n8845), .Y(REGFILE_SIM_reg_bank__abc_33898_n8846) );
  OR2X2 OR2X2_4634 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8847), .B(REGFILE_SIM_reg_bank__abc_33898_n8848), .Y(REGFILE_SIM_reg_bank__abc_33898_n8849) );
  OR2X2 OR2X2_4635 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8850), .B(REGFILE_SIM_reg_bank__abc_33898_n8851), .Y(REGFILE_SIM_reg_bank__abc_33898_n8852) );
  OR2X2 OR2X2_4636 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8852), .B(REGFILE_SIM_reg_bank__abc_33898_n8849), .Y(REGFILE_SIM_reg_bank__abc_33898_n8853) );
  OR2X2 OR2X2_4637 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8846), .B(REGFILE_SIM_reg_bank__abc_33898_n8853), .Y(REGFILE_SIM_reg_bank__abc_33898_n8854) );
  OR2X2 OR2X2_4638 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8839), .B(REGFILE_SIM_reg_bank__abc_33898_n8854), .Y(REGFILE_SIM_reg_bank__abc_33898_n8855) );
  OR2X2 OR2X2_4639 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8856), .B(REGFILE_SIM_reg_bank__abc_33898_n8857), .Y(REGFILE_SIM_reg_bank__abc_33898_n8858) );
  OR2X2 OR2X2_464 ( .A(_abc_43815_n1431_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_43815_n1986) );
  OR2X2 OR2X2_4640 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8859), .B(REGFILE_SIM_reg_bank__abc_33898_n8860), .Y(REGFILE_SIM_reg_bank__abc_33898_n8861) );
  OR2X2 OR2X2_4641 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8858), .B(REGFILE_SIM_reg_bank__abc_33898_n8861), .Y(REGFILE_SIM_reg_bank__abc_33898_n8862) );
  OR2X2 OR2X2_4642 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8864), .B(REGFILE_SIM_reg_bank__abc_33898_n8865), .Y(REGFILE_SIM_reg_bank__abc_33898_n8866) );
  OR2X2 OR2X2_4643 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8866), .B(REGFILE_SIM_reg_bank__abc_33898_n8863), .Y(REGFILE_SIM_reg_bank__abc_33898_n8867) );
  OR2X2 OR2X2_4644 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8862), .B(REGFILE_SIM_reg_bank__abc_33898_n8867), .Y(REGFILE_SIM_reg_bank__abc_33898_n8868) );
  OR2X2 OR2X2_4645 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8869), .B(REGFILE_SIM_reg_bank__abc_33898_n8870), .Y(REGFILE_SIM_reg_bank__abc_33898_n8871) );
  OR2X2 OR2X2_4646 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8872), .B(REGFILE_SIM_reg_bank__abc_33898_n8873), .Y(REGFILE_SIM_reg_bank__abc_33898_n8874) );
  OR2X2 OR2X2_4647 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8874), .B(REGFILE_SIM_reg_bank__abc_33898_n8871), .Y(REGFILE_SIM_reg_bank__abc_33898_n8875) );
  OR2X2 OR2X2_4648 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8876), .B(REGFILE_SIM_reg_bank__abc_33898_n8877), .Y(REGFILE_SIM_reg_bank__abc_33898_n8878) );
  OR2X2 OR2X2_4649 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8879), .B(REGFILE_SIM_reg_bank__abc_33898_n8880), .Y(REGFILE_SIM_reg_bank__abc_33898_n8881) );
  OR2X2 OR2X2_465 ( .A(_abc_43815_n1987), .B(_abc_43815_n1473_bF_buf1), .Y(_abc_43815_n1988) );
  OR2X2 OR2X2_4650 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8878), .B(REGFILE_SIM_reg_bank__abc_33898_n8881), .Y(REGFILE_SIM_reg_bank__abc_33898_n8882) );
  OR2X2 OR2X2_4651 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8875), .B(REGFILE_SIM_reg_bank__abc_33898_n8882), .Y(REGFILE_SIM_reg_bank__abc_33898_n8883) );
  OR2X2 OR2X2_4652 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8883), .B(REGFILE_SIM_reg_bank__abc_33898_n8868), .Y(REGFILE_SIM_reg_bank__abc_33898_n8884) );
  OR2X2 OR2X2_4653 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8855), .B(REGFILE_SIM_reg_bank__abc_33898_n8884), .Y(REGFILE_SIM_reg_bank_reg_ra_o_20_) );
  OR2X2 OR2X2_4654 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8886), .B(REGFILE_SIM_reg_bank__abc_33898_n8887), .Y(REGFILE_SIM_reg_bank__abc_33898_n8888) );
  OR2X2 OR2X2_4655 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8889), .B(REGFILE_SIM_reg_bank__abc_33898_n8890), .Y(REGFILE_SIM_reg_bank__abc_33898_n8891) );
  OR2X2 OR2X2_4656 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8891), .B(REGFILE_SIM_reg_bank__abc_33898_n8888), .Y(REGFILE_SIM_reg_bank__abc_33898_n8892) );
  OR2X2 OR2X2_4657 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8893), .B(REGFILE_SIM_reg_bank__abc_33898_n8894), .Y(REGFILE_SIM_reg_bank__abc_33898_n8895) );
  OR2X2 OR2X2_4658 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8896), .B(REGFILE_SIM_reg_bank__abc_33898_n8897), .Y(REGFILE_SIM_reg_bank__abc_33898_n8898) );
  OR2X2 OR2X2_4659 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8895), .B(REGFILE_SIM_reg_bank__abc_33898_n8898), .Y(REGFILE_SIM_reg_bank__abc_33898_n8899) );
  OR2X2 OR2X2_466 ( .A(_abc_43815_n1969), .B(_abc_43815_n1472_1_bF_buf0), .Y(_abc_43815_n1989) );
  OR2X2 OR2X2_4660 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8892), .B(REGFILE_SIM_reg_bank__abc_33898_n8899), .Y(REGFILE_SIM_reg_bank__abc_33898_n8900) );
  OR2X2 OR2X2_4661 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8901), .B(REGFILE_SIM_reg_bank__abc_33898_n8902), .Y(REGFILE_SIM_reg_bank__abc_33898_n8903) );
  OR2X2 OR2X2_4662 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8904), .B(REGFILE_SIM_reg_bank__abc_33898_n8905), .Y(REGFILE_SIM_reg_bank__abc_33898_n8906) );
  OR2X2 OR2X2_4663 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8903), .B(REGFILE_SIM_reg_bank__abc_33898_n8906), .Y(REGFILE_SIM_reg_bank__abc_33898_n8907) );
  OR2X2 OR2X2_4664 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8908), .B(REGFILE_SIM_reg_bank__abc_33898_n8909), .Y(REGFILE_SIM_reg_bank__abc_33898_n8910) );
  OR2X2 OR2X2_4665 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8911), .B(REGFILE_SIM_reg_bank__abc_33898_n8912), .Y(REGFILE_SIM_reg_bank__abc_33898_n8913) );
  OR2X2 OR2X2_4666 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8913), .B(REGFILE_SIM_reg_bank__abc_33898_n8910), .Y(REGFILE_SIM_reg_bank__abc_33898_n8914) );
  OR2X2 OR2X2_4667 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8907), .B(REGFILE_SIM_reg_bank__abc_33898_n8914), .Y(REGFILE_SIM_reg_bank__abc_33898_n8915) );
  OR2X2 OR2X2_4668 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8900), .B(REGFILE_SIM_reg_bank__abc_33898_n8915), .Y(REGFILE_SIM_reg_bank__abc_33898_n8916) );
  OR2X2 OR2X2_4669 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8917), .B(REGFILE_SIM_reg_bank__abc_33898_n8918), .Y(REGFILE_SIM_reg_bank__abc_33898_n8919) );
  OR2X2 OR2X2_467 ( .A(_abc_43815_n1990), .B(_abc_43815_n1350_bF_buf1), .Y(_abc_43815_n1991) );
  OR2X2 OR2X2_4670 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8920), .B(REGFILE_SIM_reg_bank__abc_33898_n8921), .Y(REGFILE_SIM_reg_bank__abc_33898_n8922) );
  OR2X2 OR2X2_4671 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8919), .B(REGFILE_SIM_reg_bank__abc_33898_n8922), .Y(REGFILE_SIM_reg_bank__abc_33898_n8923) );
  OR2X2 OR2X2_4672 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8925), .B(REGFILE_SIM_reg_bank__abc_33898_n8926), .Y(REGFILE_SIM_reg_bank__abc_33898_n8927) );
  OR2X2 OR2X2_4673 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8927), .B(REGFILE_SIM_reg_bank__abc_33898_n8924), .Y(REGFILE_SIM_reg_bank__abc_33898_n8928) );
  OR2X2 OR2X2_4674 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8923), .B(REGFILE_SIM_reg_bank__abc_33898_n8928), .Y(REGFILE_SIM_reg_bank__abc_33898_n8929) );
  OR2X2 OR2X2_4675 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8930), .B(REGFILE_SIM_reg_bank__abc_33898_n8931), .Y(REGFILE_SIM_reg_bank__abc_33898_n8932) );
  OR2X2 OR2X2_4676 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8933), .B(REGFILE_SIM_reg_bank__abc_33898_n8934), .Y(REGFILE_SIM_reg_bank__abc_33898_n8935) );
  OR2X2 OR2X2_4677 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8935), .B(REGFILE_SIM_reg_bank__abc_33898_n8932), .Y(REGFILE_SIM_reg_bank__abc_33898_n8936) );
  OR2X2 OR2X2_4678 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8937), .B(REGFILE_SIM_reg_bank__abc_33898_n8938), .Y(REGFILE_SIM_reg_bank__abc_33898_n8939) );
  OR2X2 OR2X2_4679 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8940), .B(REGFILE_SIM_reg_bank__abc_33898_n8941), .Y(REGFILE_SIM_reg_bank__abc_33898_n8942) );
  OR2X2 OR2X2_468 ( .A(_abc_43815_n1993_1), .B(_abc_43815_n1992), .Y(_abc_43815_n1994) );
  OR2X2 OR2X2_4680 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8939), .B(REGFILE_SIM_reg_bank__abc_33898_n8942), .Y(REGFILE_SIM_reg_bank__abc_33898_n8943) );
  OR2X2 OR2X2_4681 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8936), .B(REGFILE_SIM_reg_bank__abc_33898_n8943), .Y(REGFILE_SIM_reg_bank__abc_33898_n8944) );
  OR2X2 OR2X2_4682 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8944), .B(REGFILE_SIM_reg_bank__abc_33898_n8929), .Y(REGFILE_SIM_reg_bank__abc_33898_n8945) );
  OR2X2 OR2X2_4683 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8916), .B(REGFILE_SIM_reg_bank__abc_33898_n8945), .Y(REGFILE_SIM_reg_bank_reg_ra_o_21_) );
  OR2X2 OR2X2_4684 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8947), .B(REGFILE_SIM_reg_bank__abc_33898_n8948), .Y(REGFILE_SIM_reg_bank__abc_33898_n8949) );
  OR2X2 OR2X2_4685 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8950), .B(REGFILE_SIM_reg_bank__abc_33898_n8951), .Y(REGFILE_SIM_reg_bank__abc_33898_n8952) );
  OR2X2 OR2X2_4686 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8952), .B(REGFILE_SIM_reg_bank__abc_33898_n8949), .Y(REGFILE_SIM_reg_bank__abc_33898_n8953) );
  OR2X2 OR2X2_4687 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8954), .B(REGFILE_SIM_reg_bank__abc_33898_n8955), .Y(REGFILE_SIM_reg_bank__abc_33898_n8956) );
  OR2X2 OR2X2_4688 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8957), .B(REGFILE_SIM_reg_bank__abc_33898_n8958), .Y(REGFILE_SIM_reg_bank__abc_33898_n8959) );
  OR2X2 OR2X2_4689 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8956), .B(REGFILE_SIM_reg_bank__abc_33898_n8959), .Y(REGFILE_SIM_reg_bank__abc_33898_n8960) );
  OR2X2 OR2X2_469 ( .A(_abc_43815_n1413_bF_buf4), .B(_abc_43815_n1994), .Y(_abc_43815_n1995) );
  OR2X2 OR2X2_4690 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8953), .B(REGFILE_SIM_reg_bank__abc_33898_n8960), .Y(REGFILE_SIM_reg_bank__abc_33898_n8961) );
  OR2X2 OR2X2_4691 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8962), .B(REGFILE_SIM_reg_bank__abc_33898_n8963), .Y(REGFILE_SIM_reg_bank__abc_33898_n8964) );
  OR2X2 OR2X2_4692 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8965), .B(REGFILE_SIM_reg_bank__abc_33898_n8966), .Y(REGFILE_SIM_reg_bank__abc_33898_n8967) );
  OR2X2 OR2X2_4693 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8964), .B(REGFILE_SIM_reg_bank__abc_33898_n8967), .Y(REGFILE_SIM_reg_bank__abc_33898_n8968) );
  OR2X2 OR2X2_4694 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8969), .B(REGFILE_SIM_reg_bank__abc_33898_n8970), .Y(REGFILE_SIM_reg_bank__abc_33898_n8971) );
  OR2X2 OR2X2_4695 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8972), .B(REGFILE_SIM_reg_bank__abc_33898_n8973), .Y(REGFILE_SIM_reg_bank__abc_33898_n8974) );
  OR2X2 OR2X2_4696 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8974), .B(REGFILE_SIM_reg_bank__abc_33898_n8971), .Y(REGFILE_SIM_reg_bank__abc_33898_n8975) );
  OR2X2 OR2X2_4697 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8968), .B(REGFILE_SIM_reg_bank__abc_33898_n8975), .Y(REGFILE_SIM_reg_bank__abc_33898_n8976) );
  OR2X2 OR2X2_4698 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8961), .B(REGFILE_SIM_reg_bank__abc_33898_n8976), .Y(REGFILE_SIM_reg_bank__abc_33898_n8977) );
  OR2X2 OR2X2_4699 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8978), .B(REGFILE_SIM_reg_bank__abc_33898_n8979), .Y(REGFILE_SIM_reg_bank__abc_33898_n8980) );
  OR2X2 OR2X2_47 ( .A(_abc_43815_n782_1), .B(_abc_43815_n790), .Y(_abc_43815_n791) );
  OR2X2 OR2X2_470 ( .A(_abc_43815_n1997), .B(_abc_43815_n1971), .Y(_abc_43815_n1998) );
  OR2X2 OR2X2_4700 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8981), .B(REGFILE_SIM_reg_bank__abc_33898_n8982), .Y(REGFILE_SIM_reg_bank__abc_33898_n8983) );
  OR2X2 OR2X2_4701 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8980), .B(REGFILE_SIM_reg_bank__abc_33898_n8983), .Y(REGFILE_SIM_reg_bank__abc_33898_n8984) );
  OR2X2 OR2X2_4702 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8986), .B(REGFILE_SIM_reg_bank__abc_33898_n8987), .Y(REGFILE_SIM_reg_bank__abc_33898_n8988) );
  OR2X2 OR2X2_4703 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8988), .B(REGFILE_SIM_reg_bank__abc_33898_n8985), .Y(REGFILE_SIM_reg_bank__abc_33898_n8989) );
  OR2X2 OR2X2_4704 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8984), .B(REGFILE_SIM_reg_bank__abc_33898_n8989), .Y(REGFILE_SIM_reg_bank__abc_33898_n8990) );
  OR2X2 OR2X2_4705 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8991), .B(REGFILE_SIM_reg_bank__abc_33898_n8992), .Y(REGFILE_SIM_reg_bank__abc_33898_n8993) );
  OR2X2 OR2X2_4706 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8994), .B(REGFILE_SIM_reg_bank__abc_33898_n8995), .Y(REGFILE_SIM_reg_bank__abc_33898_n8996) );
  OR2X2 OR2X2_4707 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8996), .B(REGFILE_SIM_reg_bank__abc_33898_n8993), .Y(REGFILE_SIM_reg_bank__abc_33898_n8997) );
  OR2X2 OR2X2_4708 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8998), .B(REGFILE_SIM_reg_bank__abc_33898_n8999), .Y(REGFILE_SIM_reg_bank__abc_33898_n9000) );
  OR2X2 OR2X2_4709 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9001), .B(REGFILE_SIM_reg_bank__abc_33898_n9002), .Y(REGFILE_SIM_reg_bank__abc_33898_n9003) );
  OR2X2 OR2X2_471 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_15_), .Y(_abc_43815_n1999) );
  OR2X2 OR2X2_4710 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9000), .B(REGFILE_SIM_reg_bank__abc_33898_n9003), .Y(REGFILE_SIM_reg_bank__abc_33898_n9004) );
  OR2X2 OR2X2_4711 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8997), .B(REGFILE_SIM_reg_bank__abc_33898_n9004), .Y(REGFILE_SIM_reg_bank__abc_33898_n9005) );
  OR2X2 OR2X2_4712 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9005), .B(REGFILE_SIM_reg_bank__abc_33898_n8990), .Y(REGFILE_SIM_reg_bank__abc_33898_n9006) );
  OR2X2 OR2X2_4713 ( .A(REGFILE_SIM_reg_bank__abc_33898_n8977), .B(REGFILE_SIM_reg_bank__abc_33898_n9006), .Y(REGFILE_SIM_reg_bank_reg_ra_o_22_) );
  OR2X2 OR2X2_4714 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9008), .B(REGFILE_SIM_reg_bank__abc_33898_n9009), .Y(REGFILE_SIM_reg_bank__abc_33898_n9010) );
  OR2X2 OR2X2_4715 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9011), .B(REGFILE_SIM_reg_bank__abc_33898_n9012), .Y(REGFILE_SIM_reg_bank__abc_33898_n9013) );
  OR2X2 OR2X2_4716 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9013), .B(REGFILE_SIM_reg_bank__abc_33898_n9010), .Y(REGFILE_SIM_reg_bank__abc_33898_n9014) );
  OR2X2 OR2X2_4717 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9015), .B(REGFILE_SIM_reg_bank__abc_33898_n9016), .Y(REGFILE_SIM_reg_bank__abc_33898_n9017) );
  OR2X2 OR2X2_4718 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9018), .B(REGFILE_SIM_reg_bank__abc_33898_n9019), .Y(REGFILE_SIM_reg_bank__abc_33898_n9020) );
  OR2X2 OR2X2_4719 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9017), .B(REGFILE_SIM_reg_bank__abc_33898_n9020), .Y(REGFILE_SIM_reg_bank__abc_33898_n9021) );
  OR2X2 OR2X2_472 ( .A(_abc_43815_n1967), .B(pc_q_16_), .Y(_abc_43815_n2002) );
  OR2X2 OR2X2_4720 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9014), .B(REGFILE_SIM_reg_bank__abc_33898_n9021), .Y(REGFILE_SIM_reg_bank__abc_33898_n9022) );
  OR2X2 OR2X2_4721 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9023), .B(REGFILE_SIM_reg_bank__abc_33898_n9024), .Y(REGFILE_SIM_reg_bank__abc_33898_n9025) );
  OR2X2 OR2X2_4722 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9026), .B(REGFILE_SIM_reg_bank__abc_33898_n9027), .Y(REGFILE_SIM_reg_bank__abc_33898_n9028) );
  OR2X2 OR2X2_4723 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9025), .B(REGFILE_SIM_reg_bank__abc_33898_n9028), .Y(REGFILE_SIM_reg_bank__abc_33898_n9029) );
  OR2X2 OR2X2_4724 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9030), .B(REGFILE_SIM_reg_bank__abc_33898_n9031), .Y(REGFILE_SIM_reg_bank__abc_33898_n9032) );
  OR2X2 OR2X2_4725 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9033), .B(REGFILE_SIM_reg_bank__abc_33898_n9034), .Y(REGFILE_SIM_reg_bank__abc_33898_n9035) );
  OR2X2 OR2X2_4726 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9035), .B(REGFILE_SIM_reg_bank__abc_33898_n9032), .Y(REGFILE_SIM_reg_bank__abc_33898_n9036) );
  OR2X2 OR2X2_4727 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9029), .B(REGFILE_SIM_reg_bank__abc_33898_n9036), .Y(REGFILE_SIM_reg_bank__abc_33898_n9037) );
  OR2X2 OR2X2_4728 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9022), .B(REGFILE_SIM_reg_bank__abc_33898_n9037), .Y(REGFILE_SIM_reg_bank__abc_33898_n9038) );
  OR2X2 OR2X2_4729 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9039), .B(REGFILE_SIM_reg_bank__abc_33898_n9040), .Y(REGFILE_SIM_reg_bank__abc_33898_n9041) );
  OR2X2 OR2X2_473 ( .A(_abc_43815_n2005), .B(_abc_43815_n1278_bF_buf1), .Y(_abc_43815_n2006) );
  OR2X2 OR2X2_4730 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9042), .B(REGFILE_SIM_reg_bank__abc_33898_n9043), .Y(REGFILE_SIM_reg_bank__abc_33898_n9044) );
  OR2X2 OR2X2_4731 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9041), .B(REGFILE_SIM_reg_bank__abc_33898_n9044), .Y(REGFILE_SIM_reg_bank__abc_33898_n9045) );
  OR2X2 OR2X2_4732 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9047), .B(REGFILE_SIM_reg_bank__abc_33898_n9048), .Y(REGFILE_SIM_reg_bank__abc_33898_n9049) );
  OR2X2 OR2X2_4733 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9049), .B(REGFILE_SIM_reg_bank__abc_33898_n9046), .Y(REGFILE_SIM_reg_bank__abc_33898_n9050) );
  OR2X2 OR2X2_4734 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9045), .B(REGFILE_SIM_reg_bank__abc_33898_n9050), .Y(REGFILE_SIM_reg_bank__abc_33898_n9051) );
  OR2X2 OR2X2_4735 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9052), .B(REGFILE_SIM_reg_bank__abc_33898_n9053), .Y(REGFILE_SIM_reg_bank__abc_33898_n9054) );
  OR2X2 OR2X2_4736 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9055), .B(REGFILE_SIM_reg_bank__abc_33898_n9056), .Y(REGFILE_SIM_reg_bank__abc_33898_n9057) );
  OR2X2 OR2X2_4737 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9057), .B(REGFILE_SIM_reg_bank__abc_33898_n9054), .Y(REGFILE_SIM_reg_bank__abc_33898_n9058) );
  OR2X2 OR2X2_4738 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9059), .B(REGFILE_SIM_reg_bank__abc_33898_n9060), .Y(REGFILE_SIM_reg_bank__abc_33898_n9061) );
  OR2X2 OR2X2_4739 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9062), .B(REGFILE_SIM_reg_bank__abc_33898_n9063), .Y(REGFILE_SIM_reg_bank__abc_33898_n9064) );
  OR2X2 OR2X2_474 ( .A(_abc_43815_n2009), .B(_abc_43815_n2008), .Y(_abc_43815_n2010) );
  OR2X2 OR2X2_4740 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9061), .B(REGFILE_SIM_reg_bank__abc_33898_n9064), .Y(REGFILE_SIM_reg_bank__abc_33898_n9065) );
  OR2X2 OR2X2_4741 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9058), .B(REGFILE_SIM_reg_bank__abc_33898_n9065), .Y(REGFILE_SIM_reg_bank__abc_33898_n9066) );
  OR2X2 OR2X2_4742 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9066), .B(REGFILE_SIM_reg_bank__abc_33898_n9051), .Y(REGFILE_SIM_reg_bank__abc_33898_n9067) );
  OR2X2 OR2X2_4743 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9038), .B(REGFILE_SIM_reg_bank__abc_33898_n9067), .Y(REGFILE_SIM_reg_bank_reg_ra_o_23_) );
  OR2X2 OR2X2_4744 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9069), .B(REGFILE_SIM_reg_bank__abc_33898_n9070), .Y(REGFILE_SIM_reg_bank__abc_33898_n9071) );
  OR2X2 OR2X2_4745 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9072), .B(REGFILE_SIM_reg_bank__abc_33898_n9073), .Y(REGFILE_SIM_reg_bank__abc_33898_n9074) );
  OR2X2 OR2X2_4746 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9074), .B(REGFILE_SIM_reg_bank__abc_33898_n9071), .Y(REGFILE_SIM_reg_bank__abc_33898_n9075) );
  OR2X2 OR2X2_4747 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9076), .B(REGFILE_SIM_reg_bank__abc_33898_n9077), .Y(REGFILE_SIM_reg_bank__abc_33898_n9078) );
  OR2X2 OR2X2_4748 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9079), .B(REGFILE_SIM_reg_bank__abc_33898_n9080), .Y(REGFILE_SIM_reg_bank__abc_33898_n9081) );
  OR2X2 OR2X2_4749 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9078), .B(REGFILE_SIM_reg_bank__abc_33898_n9081), .Y(REGFILE_SIM_reg_bank__abc_33898_n9082) );
  OR2X2 OR2X2_475 ( .A(_abc_43815_n1940), .B(_abc_43815_n2013_1), .Y(_abc_43815_n2014) );
  OR2X2 OR2X2_4750 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9075), .B(REGFILE_SIM_reg_bank__abc_33898_n9082), .Y(REGFILE_SIM_reg_bank__abc_33898_n9083) );
  OR2X2 OR2X2_4751 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9084), .B(REGFILE_SIM_reg_bank__abc_33898_n9085), .Y(REGFILE_SIM_reg_bank__abc_33898_n9086) );
  OR2X2 OR2X2_4752 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9087), .B(REGFILE_SIM_reg_bank__abc_33898_n9088), .Y(REGFILE_SIM_reg_bank__abc_33898_n9089) );
  OR2X2 OR2X2_4753 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9086), .B(REGFILE_SIM_reg_bank__abc_33898_n9089), .Y(REGFILE_SIM_reg_bank__abc_33898_n9090) );
  OR2X2 OR2X2_4754 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9091), .B(REGFILE_SIM_reg_bank__abc_33898_n9092), .Y(REGFILE_SIM_reg_bank__abc_33898_n9093) );
  OR2X2 OR2X2_4755 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9094), .B(REGFILE_SIM_reg_bank__abc_33898_n9095), .Y(REGFILE_SIM_reg_bank__abc_33898_n9096) );
  OR2X2 OR2X2_4756 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9096), .B(REGFILE_SIM_reg_bank__abc_33898_n9093), .Y(REGFILE_SIM_reg_bank__abc_33898_n9097) );
  OR2X2 OR2X2_4757 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9090), .B(REGFILE_SIM_reg_bank__abc_33898_n9097), .Y(REGFILE_SIM_reg_bank__abc_33898_n9098) );
  OR2X2 OR2X2_4758 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9083), .B(REGFILE_SIM_reg_bank__abc_33898_n9098), .Y(REGFILE_SIM_reg_bank__abc_33898_n9099) );
  OR2X2 OR2X2_4759 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9100), .B(REGFILE_SIM_reg_bank__abc_33898_n9101), .Y(REGFILE_SIM_reg_bank__abc_33898_n9102) );
  OR2X2 OR2X2_476 ( .A(_abc_43815_n2015), .B(_abc_43815_n1975), .Y(_abc_43815_n2016) );
  OR2X2 OR2X2_4760 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9103), .B(REGFILE_SIM_reg_bank__abc_33898_n9104), .Y(REGFILE_SIM_reg_bank__abc_33898_n9105) );
  OR2X2 OR2X2_4761 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9102), .B(REGFILE_SIM_reg_bank__abc_33898_n9105), .Y(REGFILE_SIM_reg_bank__abc_33898_n9106) );
  OR2X2 OR2X2_4762 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9108), .B(REGFILE_SIM_reg_bank__abc_33898_n9109), .Y(REGFILE_SIM_reg_bank__abc_33898_n9110) );
  OR2X2 OR2X2_4763 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9110), .B(REGFILE_SIM_reg_bank__abc_33898_n9107), .Y(REGFILE_SIM_reg_bank__abc_33898_n9111) );
  OR2X2 OR2X2_4764 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9106), .B(REGFILE_SIM_reg_bank__abc_33898_n9111), .Y(REGFILE_SIM_reg_bank__abc_33898_n9112) );
  OR2X2 OR2X2_4765 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9113), .B(REGFILE_SIM_reg_bank__abc_33898_n9114), .Y(REGFILE_SIM_reg_bank__abc_33898_n9115) );
  OR2X2 OR2X2_4766 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9116), .B(REGFILE_SIM_reg_bank__abc_33898_n9117), .Y(REGFILE_SIM_reg_bank__abc_33898_n9118) );
  OR2X2 OR2X2_4767 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9118), .B(REGFILE_SIM_reg_bank__abc_33898_n9115), .Y(REGFILE_SIM_reg_bank__abc_33898_n9119) );
  OR2X2 OR2X2_4768 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9120), .B(REGFILE_SIM_reg_bank__abc_33898_n9121), .Y(REGFILE_SIM_reg_bank__abc_33898_n9122) );
  OR2X2 OR2X2_4769 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9123), .B(REGFILE_SIM_reg_bank__abc_33898_n9124), .Y(REGFILE_SIM_reg_bank__abc_33898_n9125) );
  OR2X2 OR2X2_477 ( .A(_abc_43815_n2021), .B(_abc_43815_n2019), .Y(_abc_43815_n2022) );
  OR2X2 OR2X2_4770 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9122), .B(REGFILE_SIM_reg_bank__abc_33898_n9125), .Y(REGFILE_SIM_reg_bank__abc_33898_n9126) );
  OR2X2 OR2X2_4771 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9119), .B(REGFILE_SIM_reg_bank__abc_33898_n9126), .Y(REGFILE_SIM_reg_bank__abc_33898_n9127) );
  OR2X2 OR2X2_4772 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9127), .B(REGFILE_SIM_reg_bank__abc_33898_n9112), .Y(REGFILE_SIM_reg_bank__abc_33898_n9128) );
  OR2X2 OR2X2_4773 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9099), .B(REGFILE_SIM_reg_bank__abc_33898_n9128), .Y(REGFILE_SIM_reg_bank_reg_ra_o_24_) );
  OR2X2 OR2X2_4774 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9130), .B(REGFILE_SIM_reg_bank__abc_33898_n9131), .Y(REGFILE_SIM_reg_bank__abc_33898_n9132) );
  OR2X2 OR2X2_4775 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9133), .B(REGFILE_SIM_reg_bank__abc_33898_n9134), .Y(REGFILE_SIM_reg_bank__abc_33898_n9135) );
  OR2X2 OR2X2_4776 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9135), .B(REGFILE_SIM_reg_bank__abc_33898_n9132), .Y(REGFILE_SIM_reg_bank__abc_33898_n9136) );
  OR2X2 OR2X2_4777 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9137), .B(REGFILE_SIM_reg_bank__abc_33898_n9138), .Y(REGFILE_SIM_reg_bank__abc_33898_n9139) );
  OR2X2 OR2X2_4778 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9140), .B(REGFILE_SIM_reg_bank__abc_33898_n9141), .Y(REGFILE_SIM_reg_bank__abc_33898_n9142) );
  OR2X2 OR2X2_4779 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9139), .B(REGFILE_SIM_reg_bank__abc_33898_n9142), .Y(REGFILE_SIM_reg_bank__abc_33898_n9143) );
  OR2X2 OR2X2_478 ( .A(pc_q_16_), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_43815_n2023) );
  OR2X2 OR2X2_4780 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9136), .B(REGFILE_SIM_reg_bank__abc_33898_n9143), .Y(REGFILE_SIM_reg_bank__abc_33898_n9144) );
  OR2X2 OR2X2_4781 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9145), .B(REGFILE_SIM_reg_bank__abc_33898_n9146), .Y(REGFILE_SIM_reg_bank__abc_33898_n9147) );
  OR2X2 OR2X2_4782 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9148), .B(REGFILE_SIM_reg_bank__abc_33898_n9149), .Y(REGFILE_SIM_reg_bank__abc_33898_n9150) );
  OR2X2 OR2X2_4783 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9147), .B(REGFILE_SIM_reg_bank__abc_33898_n9150), .Y(REGFILE_SIM_reg_bank__abc_33898_n9151) );
  OR2X2 OR2X2_4784 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9152), .B(REGFILE_SIM_reg_bank__abc_33898_n9153), .Y(REGFILE_SIM_reg_bank__abc_33898_n9154) );
  OR2X2 OR2X2_4785 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9155), .B(REGFILE_SIM_reg_bank__abc_33898_n9156), .Y(REGFILE_SIM_reg_bank__abc_33898_n9157) );
  OR2X2 OR2X2_4786 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9157), .B(REGFILE_SIM_reg_bank__abc_33898_n9154), .Y(REGFILE_SIM_reg_bank__abc_33898_n9158) );
  OR2X2 OR2X2_4787 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9151), .B(REGFILE_SIM_reg_bank__abc_33898_n9158), .Y(REGFILE_SIM_reg_bank__abc_33898_n9159) );
  OR2X2 OR2X2_4788 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9144), .B(REGFILE_SIM_reg_bank__abc_33898_n9159), .Y(REGFILE_SIM_reg_bank__abc_33898_n9160) );
  OR2X2 OR2X2_4789 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9161), .B(REGFILE_SIM_reg_bank__abc_33898_n9162), .Y(REGFILE_SIM_reg_bank__abc_33898_n9163) );
  OR2X2 OR2X2_479 ( .A(_abc_43815_n2022), .B(_abc_43815_n2026), .Y(_abc_43815_n2027) );
  OR2X2 OR2X2_4790 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9164), .B(REGFILE_SIM_reg_bank__abc_33898_n9165), .Y(REGFILE_SIM_reg_bank__abc_33898_n9166) );
  OR2X2 OR2X2_4791 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9163), .B(REGFILE_SIM_reg_bank__abc_33898_n9166), .Y(REGFILE_SIM_reg_bank__abc_33898_n9167) );
  OR2X2 OR2X2_4792 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9169), .B(REGFILE_SIM_reg_bank__abc_33898_n9170), .Y(REGFILE_SIM_reg_bank__abc_33898_n9171) );
  OR2X2 OR2X2_4793 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9171), .B(REGFILE_SIM_reg_bank__abc_33898_n9168), .Y(REGFILE_SIM_reg_bank__abc_33898_n9172) );
  OR2X2 OR2X2_4794 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9167), .B(REGFILE_SIM_reg_bank__abc_33898_n9172), .Y(REGFILE_SIM_reg_bank__abc_33898_n9173) );
  OR2X2 OR2X2_4795 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9174), .B(REGFILE_SIM_reg_bank__abc_33898_n9175), .Y(REGFILE_SIM_reg_bank__abc_33898_n9176) );
  OR2X2 OR2X2_4796 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9177), .B(REGFILE_SIM_reg_bank__abc_33898_n9178), .Y(REGFILE_SIM_reg_bank__abc_33898_n9179) );
  OR2X2 OR2X2_4797 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9179), .B(REGFILE_SIM_reg_bank__abc_33898_n9176), .Y(REGFILE_SIM_reg_bank__abc_33898_n9180) );
  OR2X2 OR2X2_4798 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9181), .B(REGFILE_SIM_reg_bank__abc_33898_n9182), .Y(REGFILE_SIM_reg_bank__abc_33898_n9183) );
  OR2X2 OR2X2_4799 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9184), .B(REGFILE_SIM_reg_bank__abc_33898_n9185), .Y(REGFILE_SIM_reg_bank__abc_33898_n9186) );
  OR2X2 OR2X2_48 ( .A(_abc_43815_n792), .B(_abc_43815_n778), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_) );
  OR2X2 OR2X2_480 ( .A(_abc_43815_n1428_bF_buf2), .B(_abc_43815_n2032), .Y(_abc_43815_n2033) );
  OR2X2 OR2X2_4800 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9183), .B(REGFILE_SIM_reg_bank__abc_33898_n9186), .Y(REGFILE_SIM_reg_bank__abc_33898_n9187) );
  OR2X2 OR2X2_4801 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9180), .B(REGFILE_SIM_reg_bank__abc_33898_n9187), .Y(REGFILE_SIM_reg_bank__abc_33898_n9188) );
  OR2X2 OR2X2_4802 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9188), .B(REGFILE_SIM_reg_bank__abc_33898_n9173), .Y(REGFILE_SIM_reg_bank__abc_33898_n9189) );
  OR2X2 OR2X2_4803 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9160), .B(REGFILE_SIM_reg_bank__abc_33898_n9189), .Y(REGFILE_SIM_reg_bank_reg_ra_o_25_) );
  OR2X2 OR2X2_4804 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9191), .B(REGFILE_SIM_reg_bank__abc_33898_n9192), .Y(REGFILE_SIM_reg_bank__abc_33898_n9193) );
  OR2X2 OR2X2_4805 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9194), .B(REGFILE_SIM_reg_bank__abc_33898_n9195), .Y(REGFILE_SIM_reg_bank__abc_33898_n9196) );
  OR2X2 OR2X2_4806 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9196), .B(REGFILE_SIM_reg_bank__abc_33898_n9193), .Y(REGFILE_SIM_reg_bank__abc_33898_n9197) );
  OR2X2 OR2X2_4807 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9198), .B(REGFILE_SIM_reg_bank__abc_33898_n9199), .Y(REGFILE_SIM_reg_bank__abc_33898_n9200) );
  OR2X2 OR2X2_4808 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9201), .B(REGFILE_SIM_reg_bank__abc_33898_n9202), .Y(REGFILE_SIM_reg_bank__abc_33898_n9203) );
  OR2X2 OR2X2_4809 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9200), .B(REGFILE_SIM_reg_bank__abc_33898_n9203), .Y(REGFILE_SIM_reg_bank__abc_33898_n9204) );
  OR2X2 OR2X2_481 ( .A(_abc_43815_n2031), .B(_abc_43815_n2033), .Y(_abc_43815_n2034_1) );
  OR2X2 OR2X2_4810 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9197), .B(REGFILE_SIM_reg_bank__abc_33898_n9204), .Y(REGFILE_SIM_reg_bank__abc_33898_n9205) );
  OR2X2 OR2X2_4811 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9206), .B(REGFILE_SIM_reg_bank__abc_33898_n9207), .Y(REGFILE_SIM_reg_bank__abc_33898_n9208) );
  OR2X2 OR2X2_4812 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9209), .B(REGFILE_SIM_reg_bank__abc_33898_n9210), .Y(REGFILE_SIM_reg_bank__abc_33898_n9211) );
  OR2X2 OR2X2_4813 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9208), .B(REGFILE_SIM_reg_bank__abc_33898_n9211), .Y(REGFILE_SIM_reg_bank__abc_33898_n9212) );
  OR2X2 OR2X2_4814 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9213), .B(REGFILE_SIM_reg_bank__abc_33898_n9214), .Y(REGFILE_SIM_reg_bank__abc_33898_n9215) );
  OR2X2 OR2X2_4815 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9216), .B(REGFILE_SIM_reg_bank__abc_33898_n9217), .Y(REGFILE_SIM_reg_bank__abc_33898_n9218) );
  OR2X2 OR2X2_4816 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9218), .B(REGFILE_SIM_reg_bank__abc_33898_n9215), .Y(REGFILE_SIM_reg_bank__abc_33898_n9219) );
  OR2X2 OR2X2_4817 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9212), .B(REGFILE_SIM_reg_bank__abc_33898_n9219), .Y(REGFILE_SIM_reg_bank__abc_33898_n9220) );
  OR2X2 OR2X2_4818 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9205), .B(REGFILE_SIM_reg_bank__abc_33898_n9220), .Y(REGFILE_SIM_reg_bank__abc_33898_n9221) );
  OR2X2 OR2X2_4819 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9222), .B(REGFILE_SIM_reg_bank__abc_33898_n9223), .Y(REGFILE_SIM_reg_bank__abc_33898_n9224) );
  OR2X2 OR2X2_482 ( .A(_abc_43815_n1431_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_43815_n2035) );
  OR2X2 OR2X2_4820 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9225), .B(REGFILE_SIM_reg_bank__abc_33898_n9226), .Y(REGFILE_SIM_reg_bank__abc_33898_n9227) );
  OR2X2 OR2X2_4821 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9224), .B(REGFILE_SIM_reg_bank__abc_33898_n9227), .Y(REGFILE_SIM_reg_bank__abc_33898_n9228) );
  OR2X2 OR2X2_4822 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9230), .B(REGFILE_SIM_reg_bank__abc_33898_n9231), .Y(REGFILE_SIM_reg_bank__abc_33898_n9232) );
  OR2X2 OR2X2_4823 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9232), .B(REGFILE_SIM_reg_bank__abc_33898_n9229), .Y(REGFILE_SIM_reg_bank__abc_33898_n9233) );
  OR2X2 OR2X2_4824 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9228), .B(REGFILE_SIM_reg_bank__abc_33898_n9233), .Y(REGFILE_SIM_reg_bank__abc_33898_n9234) );
  OR2X2 OR2X2_4825 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9235), .B(REGFILE_SIM_reg_bank__abc_33898_n9236), .Y(REGFILE_SIM_reg_bank__abc_33898_n9237) );
  OR2X2 OR2X2_4826 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9238), .B(REGFILE_SIM_reg_bank__abc_33898_n9239), .Y(REGFILE_SIM_reg_bank__abc_33898_n9240) );
  OR2X2 OR2X2_4827 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9240), .B(REGFILE_SIM_reg_bank__abc_33898_n9237), .Y(REGFILE_SIM_reg_bank__abc_33898_n9241) );
  OR2X2 OR2X2_4828 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9242), .B(REGFILE_SIM_reg_bank__abc_33898_n9243), .Y(REGFILE_SIM_reg_bank__abc_33898_n9244) );
  OR2X2 OR2X2_4829 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9245), .B(REGFILE_SIM_reg_bank__abc_33898_n9246), .Y(REGFILE_SIM_reg_bank__abc_33898_n9247) );
  OR2X2 OR2X2_483 ( .A(_abc_43815_n2037), .B(_abc_43815_n2038), .Y(_abc_43815_n2039) );
  OR2X2 OR2X2_4830 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9244), .B(REGFILE_SIM_reg_bank__abc_33898_n9247), .Y(REGFILE_SIM_reg_bank__abc_33898_n9248) );
  OR2X2 OR2X2_4831 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9241), .B(REGFILE_SIM_reg_bank__abc_33898_n9248), .Y(REGFILE_SIM_reg_bank__abc_33898_n9249) );
  OR2X2 OR2X2_4832 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9249), .B(REGFILE_SIM_reg_bank__abc_33898_n9234), .Y(REGFILE_SIM_reg_bank__abc_33898_n9250) );
  OR2X2 OR2X2_4833 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9221), .B(REGFILE_SIM_reg_bank__abc_33898_n9250), .Y(REGFILE_SIM_reg_bank_reg_ra_o_26_) );
  OR2X2 OR2X2_4834 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9252), .B(REGFILE_SIM_reg_bank__abc_33898_n9253), .Y(REGFILE_SIM_reg_bank__abc_33898_n9254) );
  OR2X2 OR2X2_4835 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9255), .B(REGFILE_SIM_reg_bank__abc_33898_n9256), .Y(REGFILE_SIM_reg_bank__abc_33898_n9257) );
  OR2X2 OR2X2_4836 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9257), .B(REGFILE_SIM_reg_bank__abc_33898_n9254), .Y(REGFILE_SIM_reg_bank__abc_33898_n9258) );
  OR2X2 OR2X2_4837 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9259), .B(REGFILE_SIM_reg_bank__abc_33898_n9260), .Y(REGFILE_SIM_reg_bank__abc_33898_n9261) );
  OR2X2 OR2X2_4838 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9262), .B(REGFILE_SIM_reg_bank__abc_33898_n9263), .Y(REGFILE_SIM_reg_bank__abc_33898_n9264) );
  OR2X2 OR2X2_4839 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9261), .B(REGFILE_SIM_reg_bank__abc_33898_n9264), .Y(REGFILE_SIM_reg_bank__abc_33898_n9265) );
  OR2X2 OR2X2_484 ( .A(_abc_43815_n2040), .B(_abc_43815_n2011), .Y(_abc_43815_n2041) );
  OR2X2 OR2X2_4840 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9258), .B(REGFILE_SIM_reg_bank__abc_33898_n9265), .Y(REGFILE_SIM_reg_bank__abc_33898_n9266) );
  OR2X2 OR2X2_4841 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9267), .B(REGFILE_SIM_reg_bank__abc_33898_n9268), .Y(REGFILE_SIM_reg_bank__abc_33898_n9269) );
  OR2X2 OR2X2_4842 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9270), .B(REGFILE_SIM_reg_bank__abc_33898_n9271), .Y(REGFILE_SIM_reg_bank__abc_33898_n9272) );
  OR2X2 OR2X2_4843 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9269), .B(REGFILE_SIM_reg_bank__abc_33898_n9272), .Y(REGFILE_SIM_reg_bank__abc_33898_n9273) );
  OR2X2 OR2X2_4844 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9274), .B(REGFILE_SIM_reg_bank__abc_33898_n9275), .Y(REGFILE_SIM_reg_bank__abc_33898_n9276) );
  OR2X2 OR2X2_4845 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9277), .B(REGFILE_SIM_reg_bank__abc_33898_n9278), .Y(REGFILE_SIM_reg_bank__abc_33898_n9279) );
  OR2X2 OR2X2_4846 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9279), .B(REGFILE_SIM_reg_bank__abc_33898_n9276), .Y(REGFILE_SIM_reg_bank__abc_33898_n9280) );
  OR2X2 OR2X2_4847 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9273), .B(REGFILE_SIM_reg_bank__abc_33898_n9280), .Y(REGFILE_SIM_reg_bank__abc_33898_n9281) );
  OR2X2 OR2X2_4848 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9266), .B(REGFILE_SIM_reg_bank__abc_33898_n9281), .Y(REGFILE_SIM_reg_bank__abc_33898_n9282) );
  OR2X2 OR2X2_4849 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9283), .B(REGFILE_SIM_reg_bank__abc_33898_n9284), .Y(REGFILE_SIM_reg_bank__abc_33898_n9285) );
  OR2X2 OR2X2_485 ( .A(_abc_43815_n2042), .B(_abc_43815_n2007), .Y(_abc_43815_n2043) );
  OR2X2 OR2X2_4850 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9286), .B(REGFILE_SIM_reg_bank__abc_33898_n9287), .Y(REGFILE_SIM_reg_bank__abc_33898_n9288) );
  OR2X2 OR2X2_4851 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9285), .B(REGFILE_SIM_reg_bank__abc_33898_n9288), .Y(REGFILE_SIM_reg_bank__abc_33898_n9289) );
  OR2X2 OR2X2_4852 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9291), .B(REGFILE_SIM_reg_bank__abc_33898_n9292), .Y(REGFILE_SIM_reg_bank__abc_33898_n9293) );
  OR2X2 OR2X2_4853 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9293), .B(REGFILE_SIM_reg_bank__abc_33898_n9290), .Y(REGFILE_SIM_reg_bank__abc_33898_n9294) );
  OR2X2 OR2X2_4854 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9289), .B(REGFILE_SIM_reg_bank__abc_33898_n9294), .Y(REGFILE_SIM_reg_bank__abc_33898_n9295) );
  OR2X2 OR2X2_4855 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9296), .B(REGFILE_SIM_reg_bank__abc_33898_n9297), .Y(REGFILE_SIM_reg_bank__abc_33898_n9298) );
  OR2X2 OR2X2_4856 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9299), .B(REGFILE_SIM_reg_bank__abc_33898_n9300), .Y(REGFILE_SIM_reg_bank__abc_33898_n9301) );
  OR2X2 OR2X2_4857 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9301), .B(REGFILE_SIM_reg_bank__abc_33898_n9298), .Y(REGFILE_SIM_reg_bank__abc_33898_n9302) );
  OR2X2 OR2X2_4858 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9303), .B(REGFILE_SIM_reg_bank__abc_33898_n9304), .Y(REGFILE_SIM_reg_bank__abc_33898_n9305) );
  OR2X2 OR2X2_4859 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9306), .B(REGFILE_SIM_reg_bank__abc_33898_n9307), .Y(REGFILE_SIM_reg_bank__abc_33898_n9308) );
  OR2X2 OR2X2_486 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_16_), .Y(_abc_43815_n2044) );
  OR2X2 OR2X2_4860 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9305), .B(REGFILE_SIM_reg_bank__abc_33898_n9308), .Y(REGFILE_SIM_reg_bank__abc_33898_n9309) );
  OR2X2 OR2X2_4861 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9302), .B(REGFILE_SIM_reg_bank__abc_33898_n9309), .Y(REGFILE_SIM_reg_bank__abc_33898_n9310) );
  OR2X2 OR2X2_4862 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9310), .B(REGFILE_SIM_reg_bank__abc_33898_n9295), .Y(REGFILE_SIM_reg_bank__abc_33898_n9311) );
  OR2X2 OR2X2_4863 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9282), .B(REGFILE_SIM_reg_bank__abc_33898_n9311), .Y(REGFILE_SIM_reg_bank_reg_ra_o_27_) );
  OR2X2 OR2X2_4864 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9313), .B(REGFILE_SIM_reg_bank__abc_33898_n9314), .Y(REGFILE_SIM_reg_bank__abc_33898_n9315) );
  OR2X2 OR2X2_4865 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9316), .B(REGFILE_SIM_reg_bank__abc_33898_n9317), .Y(REGFILE_SIM_reg_bank__abc_33898_n9318) );
  OR2X2 OR2X2_4866 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9318), .B(REGFILE_SIM_reg_bank__abc_33898_n9315), .Y(REGFILE_SIM_reg_bank__abc_33898_n9319) );
  OR2X2 OR2X2_4867 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9320), .B(REGFILE_SIM_reg_bank__abc_33898_n9321), .Y(REGFILE_SIM_reg_bank__abc_33898_n9322) );
  OR2X2 OR2X2_4868 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9323), .B(REGFILE_SIM_reg_bank__abc_33898_n9324), .Y(REGFILE_SIM_reg_bank__abc_33898_n9325) );
  OR2X2 OR2X2_4869 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9322), .B(REGFILE_SIM_reg_bank__abc_33898_n9325), .Y(REGFILE_SIM_reg_bank__abc_33898_n9326) );
  OR2X2 OR2X2_487 ( .A(_abc_43815_n2003), .B(pc_q_17_), .Y(_abc_43815_n2047) );
  OR2X2 OR2X2_4870 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9319), .B(REGFILE_SIM_reg_bank__abc_33898_n9326), .Y(REGFILE_SIM_reg_bank__abc_33898_n9327) );
  OR2X2 OR2X2_4871 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9328), .B(REGFILE_SIM_reg_bank__abc_33898_n9329), .Y(REGFILE_SIM_reg_bank__abc_33898_n9330) );
  OR2X2 OR2X2_4872 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9331), .B(REGFILE_SIM_reg_bank__abc_33898_n9332), .Y(REGFILE_SIM_reg_bank__abc_33898_n9333) );
  OR2X2 OR2X2_4873 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9330), .B(REGFILE_SIM_reg_bank__abc_33898_n9333), .Y(REGFILE_SIM_reg_bank__abc_33898_n9334) );
  OR2X2 OR2X2_4874 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9335), .B(REGFILE_SIM_reg_bank__abc_33898_n9336), .Y(REGFILE_SIM_reg_bank__abc_33898_n9337) );
  OR2X2 OR2X2_4875 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9338), .B(REGFILE_SIM_reg_bank__abc_33898_n9339), .Y(REGFILE_SIM_reg_bank__abc_33898_n9340) );
  OR2X2 OR2X2_4876 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9340), .B(REGFILE_SIM_reg_bank__abc_33898_n9337), .Y(REGFILE_SIM_reg_bank__abc_33898_n9341) );
  OR2X2 OR2X2_4877 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9334), .B(REGFILE_SIM_reg_bank__abc_33898_n9341), .Y(REGFILE_SIM_reg_bank__abc_33898_n9342) );
  OR2X2 OR2X2_4878 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9327), .B(REGFILE_SIM_reg_bank__abc_33898_n9342), .Y(REGFILE_SIM_reg_bank__abc_33898_n9343) );
  OR2X2 OR2X2_4879 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9344), .B(REGFILE_SIM_reg_bank__abc_33898_n9345), .Y(REGFILE_SIM_reg_bank__abc_33898_n9346) );
  OR2X2 OR2X2_488 ( .A(_abc_43815_n2051), .B(_abc_43815_n1278_bF_buf0), .Y(_abc_43815_n2052) );
  OR2X2 OR2X2_4880 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9347), .B(REGFILE_SIM_reg_bank__abc_33898_n9348), .Y(REGFILE_SIM_reg_bank__abc_33898_n9349) );
  OR2X2 OR2X2_4881 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9346), .B(REGFILE_SIM_reg_bank__abc_33898_n9349), .Y(REGFILE_SIM_reg_bank__abc_33898_n9350) );
  OR2X2 OR2X2_4882 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9352), .B(REGFILE_SIM_reg_bank__abc_33898_n9353), .Y(REGFILE_SIM_reg_bank__abc_33898_n9354) );
  OR2X2 OR2X2_4883 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9354), .B(REGFILE_SIM_reg_bank__abc_33898_n9351), .Y(REGFILE_SIM_reg_bank__abc_33898_n9355) );
  OR2X2 OR2X2_4884 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9350), .B(REGFILE_SIM_reg_bank__abc_33898_n9355), .Y(REGFILE_SIM_reg_bank__abc_33898_n9356) );
  OR2X2 OR2X2_4885 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9357), .B(REGFILE_SIM_reg_bank__abc_33898_n9358), .Y(REGFILE_SIM_reg_bank__abc_33898_n9359) );
  OR2X2 OR2X2_4886 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9360), .B(REGFILE_SIM_reg_bank__abc_33898_n9361), .Y(REGFILE_SIM_reg_bank__abc_33898_n9362) );
  OR2X2 OR2X2_4887 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9362), .B(REGFILE_SIM_reg_bank__abc_33898_n9359), .Y(REGFILE_SIM_reg_bank__abc_33898_n9363) );
  OR2X2 OR2X2_4888 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9364), .B(REGFILE_SIM_reg_bank__abc_33898_n9365), .Y(REGFILE_SIM_reg_bank__abc_33898_n9366) );
  OR2X2 OR2X2_4889 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9367), .B(REGFILE_SIM_reg_bank__abc_33898_n9368), .Y(REGFILE_SIM_reg_bank__abc_33898_n9369) );
  OR2X2 OR2X2_489 ( .A(_abc_43815_n2054), .B(_abc_43815_n2053), .Y(_abc_43815_n2055_1) );
  OR2X2 OR2X2_4890 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9366), .B(REGFILE_SIM_reg_bank__abc_33898_n9369), .Y(REGFILE_SIM_reg_bank__abc_33898_n9370) );
  OR2X2 OR2X2_4891 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9363), .B(REGFILE_SIM_reg_bank__abc_33898_n9370), .Y(REGFILE_SIM_reg_bank__abc_33898_n9371) );
  OR2X2 OR2X2_4892 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9371), .B(REGFILE_SIM_reg_bank__abc_33898_n9356), .Y(REGFILE_SIM_reg_bank__abc_33898_n9372) );
  OR2X2 OR2X2_4893 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9343), .B(REGFILE_SIM_reg_bank__abc_33898_n9372), .Y(REGFILE_SIM_reg_bank_reg_ra_o_28_) );
  OR2X2 OR2X2_4894 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9374), .B(REGFILE_SIM_reg_bank__abc_33898_n9375), .Y(REGFILE_SIM_reg_bank__abc_33898_n9376) );
  OR2X2 OR2X2_4895 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9377), .B(REGFILE_SIM_reg_bank__abc_33898_n9378), .Y(REGFILE_SIM_reg_bank__abc_33898_n9379) );
  OR2X2 OR2X2_4896 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9379), .B(REGFILE_SIM_reg_bank__abc_33898_n9376), .Y(REGFILE_SIM_reg_bank__abc_33898_n9380) );
  OR2X2 OR2X2_4897 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9381), .B(REGFILE_SIM_reg_bank__abc_33898_n9382), .Y(REGFILE_SIM_reg_bank__abc_33898_n9383) );
  OR2X2 OR2X2_4898 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9384), .B(REGFILE_SIM_reg_bank__abc_33898_n9385), .Y(REGFILE_SIM_reg_bank__abc_33898_n9386) );
  OR2X2 OR2X2_4899 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9383), .B(REGFILE_SIM_reg_bank__abc_33898_n9386), .Y(REGFILE_SIM_reg_bank__abc_33898_n9387) );
  OR2X2 OR2X2_49 ( .A(_abc_43815_n796), .B(_abc_43815_n685), .Y(_abc_43815_n797) );
  OR2X2 OR2X2_490 ( .A(_abc_43815_n1431_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_43815_n2057) );
  OR2X2 OR2X2_4900 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9380), .B(REGFILE_SIM_reg_bank__abc_33898_n9387), .Y(REGFILE_SIM_reg_bank__abc_33898_n9388) );
  OR2X2 OR2X2_4901 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9389), .B(REGFILE_SIM_reg_bank__abc_33898_n9390), .Y(REGFILE_SIM_reg_bank__abc_33898_n9391) );
  OR2X2 OR2X2_4902 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9392), .B(REGFILE_SIM_reg_bank__abc_33898_n9393), .Y(REGFILE_SIM_reg_bank__abc_33898_n9394) );
  OR2X2 OR2X2_4903 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9391), .B(REGFILE_SIM_reg_bank__abc_33898_n9394), .Y(REGFILE_SIM_reg_bank__abc_33898_n9395) );
  OR2X2 OR2X2_4904 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9396), .B(REGFILE_SIM_reg_bank__abc_33898_n9397), .Y(REGFILE_SIM_reg_bank__abc_33898_n9398) );
  OR2X2 OR2X2_4905 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9399), .B(REGFILE_SIM_reg_bank__abc_33898_n9400), .Y(REGFILE_SIM_reg_bank__abc_33898_n9401) );
  OR2X2 OR2X2_4906 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9401), .B(REGFILE_SIM_reg_bank__abc_33898_n9398), .Y(REGFILE_SIM_reg_bank__abc_33898_n9402) );
  OR2X2 OR2X2_4907 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9395), .B(REGFILE_SIM_reg_bank__abc_33898_n9402), .Y(REGFILE_SIM_reg_bank__abc_33898_n9403) );
  OR2X2 OR2X2_4908 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9388), .B(REGFILE_SIM_reg_bank__abc_33898_n9403), .Y(REGFILE_SIM_reg_bank__abc_33898_n9404) );
  OR2X2 OR2X2_4909 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9405), .B(REGFILE_SIM_reg_bank__abc_33898_n9406), .Y(REGFILE_SIM_reg_bank__abc_33898_n9407) );
  OR2X2 OR2X2_491 ( .A(pc_q_17_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3), .Y(_abc_43815_n2058) );
  OR2X2 OR2X2_4910 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9408), .B(REGFILE_SIM_reg_bank__abc_33898_n9409), .Y(REGFILE_SIM_reg_bank__abc_33898_n9410) );
  OR2X2 OR2X2_4911 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9407), .B(REGFILE_SIM_reg_bank__abc_33898_n9410), .Y(REGFILE_SIM_reg_bank__abc_33898_n9411) );
  OR2X2 OR2X2_4912 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9413), .B(REGFILE_SIM_reg_bank__abc_33898_n9414), .Y(REGFILE_SIM_reg_bank__abc_33898_n9415) );
  OR2X2 OR2X2_4913 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9415), .B(REGFILE_SIM_reg_bank__abc_33898_n9412), .Y(REGFILE_SIM_reg_bank__abc_33898_n9416) );
  OR2X2 OR2X2_4914 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9411), .B(REGFILE_SIM_reg_bank__abc_33898_n9416), .Y(REGFILE_SIM_reg_bank__abc_33898_n9417) );
  OR2X2 OR2X2_4915 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9418), .B(REGFILE_SIM_reg_bank__abc_33898_n9419), .Y(REGFILE_SIM_reg_bank__abc_33898_n9420) );
  OR2X2 OR2X2_4916 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9421), .B(REGFILE_SIM_reg_bank__abc_33898_n9422), .Y(REGFILE_SIM_reg_bank__abc_33898_n9423) );
  OR2X2 OR2X2_4917 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9423), .B(REGFILE_SIM_reg_bank__abc_33898_n9420), .Y(REGFILE_SIM_reg_bank__abc_33898_n9424) );
  OR2X2 OR2X2_4918 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9425), .B(REGFILE_SIM_reg_bank__abc_33898_n9426), .Y(REGFILE_SIM_reg_bank__abc_33898_n9427) );
  OR2X2 OR2X2_4919 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9428), .B(REGFILE_SIM_reg_bank__abc_33898_n9429), .Y(REGFILE_SIM_reg_bank__abc_33898_n9430) );
  OR2X2 OR2X2_492 ( .A(_abc_43815_n2061), .B(_abc_43815_n2024), .Y(_abc_43815_n2062) );
  OR2X2 OR2X2_4920 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9427), .B(REGFILE_SIM_reg_bank__abc_33898_n9430), .Y(REGFILE_SIM_reg_bank__abc_33898_n9431) );
  OR2X2 OR2X2_4921 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9424), .B(REGFILE_SIM_reg_bank__abc_33898_n9431), .Y(REGFILE_SIM_reg_bank__abc_33898_n9432) );
  OR2X2 OR2X2_4922 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9432), .B(REGFILE_SIM_reg_bank__abc_33898_n9417), .Y(REGFILE_SIM_reg_bank__abc_33898_n9433) );
  OR2X2 OR2X2_4923 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9404), .B(REGFILE_SIM_reg_bank__abc_33898_n9433), .Y(REGFILE_SIM_reg_bank_reg_ra_o_29_) );
  OR2X2 OR2X2_4924 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9435), .B(REGFILE_SIM_reg_bank__abc_33898_n9436), .Y(REGFILE_SIM_reg_bank__abc_33898_n9437) );
  OR2X2 OR2X2_4925 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9438), .B(REGFILE_SIM_reg_bank__abc_33898_n9439), .Y(REGFILE_SIM_reg_bank__abc_33898_n9440) );
  OR2X2 OR2X2_4926 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9440), .B(REGFILE_SIM_reg_bank__abc_33898_n9437), .Y(REGFILE_SIM_reg_bank__abc_33898_n9441) );
  OR2X2 OR2X2_4927 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9442), .B(REGFILE_SIM_reg_bank__abc_33898_n9443), .Y(REGFILE_SIM_reg_bank__abc_33898_n9444) );
  OR2X2 OR2X2_4928 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9445), .B(REGFILE_SIM_reg_bank__abc_33898_n9446), .Y(REGFILE_SIM_reg_bank__abc_33898_n9447) );
  OR2X2 OR2X2_4929 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9444), .B(REGFILE_SIM_reg_bank__abc_33898_n9447), .Y(REGFILE_SIM_reg_bank__abc_33898_n9448) );
  OR2X2 OR2X2_493 ( .A(_abc_43815_n2028), .B(_abc_43815_n2062), .Y(_abc_43815_n2063) );
  OR2X2 OR2X2_4930 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9441), .B(REGFILE_SIM_reg_bank__abc_33898_n9448), .Y(REGFILE_SIM_reg_bank__abc_33898_n9449) );
  OR2X2 OR2X2_4931 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9450), .B(REGFILE_SIM_reg_bank__abc_33898_n9451), .Y(REGFILE_SIM_reg_bank__abc_33898_n9452) );
  OR2X2 OR2X2_4932 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9453), .B(REGFILE_SIM_reg_bank__abc_33898_n9454), .Y(REGFILE_SIM_reg_bank__abc_33898_n9455) );
  OR2X2 OR2X2_4933 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9452), .B(REGFILE_SIM_reg_bank__abc_33898_n9455), .Y(REGFILE_SIM_reg_bank__abc_33898_n9456) );
  OR2X2 OR2X2_4934 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9457), .B(REGFILE_SIM_reg_bank__abc_33898_n9458), .Y(REGFILE_SIM_reg_bank__abc_33898_n9459) );
  OR2X2 OR2X2_4935 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9460), .B(REGFILE_SIM_reg_bank__abc_33898_n9461), .Y(REGFILE_SIM_reg_bank__abc_33898_n9462) );
  OR2X2 OR2X2_4936 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9462), .B(REGFILE_SIM_reg_bank__abc_33898_n9459), .Y(REGFILE_SIM_reg_bank__abc_33898_n9463) );
  OR2X2 OR2X2_4937 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9456), .B(REGFILE_SIM_reg_bank__abc_33898_n9463), .Y(REGFILE_SIM_reg_bank__abc_33898_n9464) );
  OR2X2 OR2X2_4938 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9449), .B(REGFILE_SIM_reg_bank__abc_33898_n9464), .Y(REGFILE_SIM_reg_bank__abc_33898_n9465) );
  OR2X2 OR2X2_4939 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9466), .B(REGFILE_SIM_reg_bank__abc_33898_n9467), .Y(REGFILE_SIM_reg_bank__abc_33898_n9468) );
  OR2X2 OR2X2_494 ( .A(_abc_43815_n1428_bF_buf1), .B(_abc_43815_n2072), .Y(_abc_43815_n2073_1) );
  OR2X2 OR2X2_4940 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9469), .B(REGFILE_SIM_reg_bank__abc_33898_n9470), .Y(REGFILE_SIM_reg_bank__abc_33898_n9471) );
  OR2X2 OR2X2_4941 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9468), .B(REGFILE_SIM_reg_bank__abc_33898_n9471), .Y(REGFILE_SIM_reg_bank__abc_33898_n9472) );
  OR2X2 OR2X2_4942 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9474), .B(REGFILE_SIM_reg_bank__abc_33898_n9475), .Y(REGFILE_SIM_reg_bank__abc_33898_n9476) );
  OR2X2 OR2X2_4943 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9476), .B(REGFILE_SIM_reg_bank__abc_33898_n9473), .Y(REGFILE_SIM_reg_bank__abc_33898_n9477) );
  OR2X2 OR2X2_4944 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9472), .B(REGFILE_SIM_reg_bank__abc_33898_n9477), .Y(REGFILE_SIM_reg_bank__abc_33898_n9478) );
  OR2X2 OR2X2_4945 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9479), .B(REGFILE_SIM_reg_bank__abc_33898_n9480), .Y(REGFILE_SIM_reg_bank__abc_33898_n9481) );
  OR2X2 OR2X2_4946 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9482), .B(REGFILE_SIM_reg_bank__abc_33898_n9483), .Y(REGFILE_SIM_reg_bank__abc_33898_n9484) );
  OR2X2 OR2X2_4947 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9484), .B(REGFILE_SIM_reg_bank__abc_33898_n9481), .Y(REGFILE_SIM_reg_bank__abc_33898_n9485) );
  OR2X2 OR2X2_4948 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9486), .B(REGFILE_SIM_reg_bank__abc_33898_n9487), .Y(REGFILE_SIM_reg_bank__abc_33898_n9488) );
  OR2X2 OR2X2_4949 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9489), .B(REGFILE_SIM_reg_bank__abc_33898_n9490), .Y(REGFILE_SIM_reg_bank__abc_33898_n9491) );
  OR2X2 OR2X2_495 ( .A(_abc_43815_n2071), .B(_abc_43815_n2073_1), .Y(_abc_43815_n2074) );
  OR2X2 OR2X2_4950 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9488), .B(REGFILE_SIM_reg_bank__abc_33898_n9491), .Y(REGFILE_SIM_reg_bank__abc_33898_n9492) );
  OR2X2 OR2X2_4951 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9485), .B(REGFILE_SIM_reg_bank__abc_33898_n9492), .Y(REGFILE_SIM_reg_bank__abc_33898_n9493) );
  OR2X2 OR2X2_4952 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9493), .B(REGFILE_SIM_reg_bank__abc_33898_n9478), .Y(REGFILE_SIM_reg_bank__abc_33898_n9494) );
  OR2X2 OR2X2_4953 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9465), .B(REGFILE_SIM_reg_bank__abc_33898_n9494), .Y(REGFILE_SIM_reg_bank_reg_ra_o_30_) );
  OR2X2 OR2X2_4954 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9496), .B(REGFILE_SIM_reg_bank__abc_33898_n9497), .Y(REGFILE_SIM_reg_bank__abc_33898_n9498) );
  OR2X2 OR2X2_4955 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9499), .B(REGFILE_SIM_reg_bank__abc_33898_n9500), .Y(REGFILE_SIM_reg_bank__abc_33898_n9501) );
  OR2X2 OR2X2_4956 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9501), .B(REGFILE_SIM_reg_bank__abc_33898_n9498), .Y(REGFILE_SIM_reg_bank__abc_33898_n9502) );
  OR2X2 OR2X2_4957 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9503), .B(REGFILE_SIM_reg_bank__abc_33898_n9504), .Y(REGFILE_SIM_reg_bank__abc_33898_n9505) );
  OR2X2 OR2X2_4958 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9506), .B(REGFILE_SIM_reg_bank__abc_33898_n9507), .Y(REGFILE_SIM_reg_bank__abc_33898_n9508) );
  OR2X2 OR2X2_4959 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9505), .B(REGFILE_SIM_reg_bank__abc_33898_n9508), .Y(REGFILE_SIM_reg_bank__abc_33898_n9509) );
  OR2X2 OR2X2_496 ( .A(_abc_43815_n2075), .B(_abc_43815_n1473_bF_buf4), .Y(_abc_43815_n2076) );
  OR2X2 OR2X2_4960 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9502), .B(REGFILE_SIM_reg_bank__abc_33898_n9509), .Y(REGFILE_SIM_reg_bank__abc_33898_n9510) );
  OR2X2 OR2X2_4961 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9511), .B(REGFILE_SIM_reg_bank__abc_33898_n9512), .Y(REGFILE_SIM_reg_bank__abc_33898_n9513) );
  OR2X2 OR2X2_4962 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9514), .B(REGFILE_SIM_reg_bank__abc_33898_n9515), .Y(REGFILE_SIM_reg_bank__abc_33898_n9516) );
  OR2X2 OR2X2_4963 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9513), .B(REGFILE_SIM_reg_bank__abc_33898_n9516), .Y(REGFILE_SIM_reg_bank__abc_33898_n9517) );
  OR2X2 OR2X2_4964 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9518), .B(REGFILE_SIM_reg_bank__abc_33898_n9519), .Y(REGFILE_SIM_reg_bank__abc_33898_n9520) );
  OR2X2 OR2X2_4965 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9521), .B(REGFILE_SIM_reg_bank__abc_33898_n9522), .Y(REGFILE_SIM_reg_bank__abc_33898_n9523) );
  OR2X2 OR2X2_4966 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9523), .B(REGFILE_SIM_reg_bank__abc_33898_n9520), .Y(REGFILE_SIM_reg_bank__abc_33898_n9524) );
  OR2X2 OR2X2_4967 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9517), .B(REGFILE_SIM_reg_bank__abc_33898_n9524), .Y(REGFILE_SIM_reg_bank__abc_33898_n9525) );
  OR2X2 OR2X2_4968 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9510), .B(REGFILE_SIM_reg_bank__abc_33898_n9525), .Y(REGFILE_SIM_reg_bank__abc_33898_n9526) );
  OR2X2 OR2X2_4969 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9527), .B(REGFILE_SIM_reg_bank__abc_33898_n9528), .Y(REGFILE_SIM_reg_bank__abc_33898_n9529) );
  OR2X2 OR2X2_497 ( .A(_abc_43815_n2050), .B(_abc_43815_n1472_1_bF_buf3), .Y(_abc_43815_n2077) );
  OR2X2 OR2X2_4970 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9530), .B(REGFILE_SIM_reg_bank__abc_33898_n9531), .Y(REGFILE_SIM_reg_bank__abc_33898_n9532) );
  OR2X2 OR2X2_4971 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9529), .B(REGFILE_SIM_reg_bank__abc_33898_n9532), .Y(REGFILE_SIM_reg_bank__abc_33898_n9533) );
  OR2X2 OR2X2_4972 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9535), .B(REGFILE_SIM_reg_bank__abc_33898_n9536), .Y(REGFILE_SIM_reg_bank__abc_33898_n9537) );
  OR2X2 OR2X2_4973 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9537), .B(REGFILE_SIM_reg_bank__abc_33898_n9534), .Y(REGFILE_SIM_reg_bank__abc_33898_n9538) );
  OR2X2 OR2X2_4974 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9533), .B(REGFILE_SIM_reg_bank__abc_33898_n9538), .Y(REGFILE_SIM_reg_bank__abc_33898_n9539) );
  OR2X2 OR2X2_4975 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9540), .B(REGFILE_SIM_reg_bank__abc_33898_n9541), .Y(REGFILE_SIM_reg_bank__abc_33898_n9542) );
  OR2X2 OR2X2_4976 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9543), .B(REGFILE_SIM_reg_bank__abc_33898_n9544), .Y(REGFILE_SIM_reg_bank__abc_33898_n9545) );
  OR2X2 OR2X2_4977 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9545), .B(REGFILE_SIM_reg_bank__abc_33898_n9542), .Y(REGFILE_SIM_reg_bank__abc_33898_n9546) );
  OR2X2 OR2X2_4978 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9547), .B(REGFILE_SIM_reg_bank__abc_33898_n9548), .Y(REGFILE_SIM_reg_bank__abc_33898_n9549) );
  OR2X2 OR2X2_4979 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9550), .B(REGFILE_SIM_reg_bank__abc_33898_n9551), .Y(REGFILE_SIM_reg_bank__abc_33898_n9552) );
  OR2X2 OR2X2_498 ( .A(_abc_43815_n2079), .B(_abc_43815_n2056), .Y(_abc_43815_n2080) );
  OR2X2 OR2X2_4980 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9549), .B(REGFILE_SIM_reg_bank__abc_33898_n9552), .Y(REGFILE_SIM_reg_bank__abc_33898_n9553) );
  OR2X2 OR2X2_4981 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9546), .B(REGFILE_SIM_reg_bank__abc_33898_n9553), .Y(REGFILE_SIM_reg_bank__abc_33898_n9554) );
  OR2X2 OR2X2_4982 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9554), .B(REGFILE_SIM_reg_bank__abc_33898_n9539), .Y(REGFILE_SIM_reg_bank__abc_33898_n9555) );
  OR2X2 OR2X2_4983 ( .A(REGFILE_SIM_reg_bank__abc_33898_n9526), .B(REGFILE_SIM_reg_bank__abc_33898_n9555), .Y(REGFILE_SIM_reg_bank_reg_ra_o_31_) );
  OR2X2 OR2X2_4984 ( .A(alu__abc_41358_n173), .B(alu__abc_41358_n170), .Y(alu__abc_41358_n174) );
  OR2X2 OR2X2_4985 ( .A(alu__abc_41358_n253), .B(alu__abc_41358_n250), .Y(alu__abc_41358_n254) );
  OR2X2 OR2X2_4986 ( .A(alu__abc_41358_n274), .B(alu__abc_41358_n271), .Y(alu__abc_41358_n275) );
  OR2X2 OR2X2_4987 ( .A(alu__abc_41358_n288), .B(alu__abc_41358_n285), .Y(alu__abc_41358_n289) );
  OR2X2 OR2X2_4988 ( .A(alu__abc_41358_n295), .B(alu__abc_41358_n292), .Y(alu__abc_41358_n296) );
  OR2X2 OR2X2_4989 ( .A(alu__abc_41358_n300), .B(alu__abc_41358_n297), .Y(alu__abc_41358_n301) );
  OR2X2 OR2X2_499 ( .A(_abc_43815_n2081), .B(_abc_43815_n2052), .Y(_abc_43815_n2082) );
  OR2X2 OR2X2_4990 ( .A(alu__abc_41358_n390), .B(alu__abc_41358_n388), .Y(alu__abc_41358_n391) );
  OR2X2 OR2X2_4991 ( .A(alu__abc_41358_n399), .B(alu__abc_41358_n394), .Y(alu__abc_41358_n400) );
  OR2X2 OR2X2_4992 ( .A(alu__abc_41358_n393), .B(alu__abc_41358_n400), .Y(alu__abc_41358_n401) );
  OR2X2 OR2X2_4993 ( .A(alu__abc_41358_n258), .B(alu__abc_41358_n416), .Y(alu__abc_41358_n417) );
  OR2X2 OR2X2_4994 ( .A(alu__abc_41358_n418), .B(alu__abc_41358_n415), .Y(alu__abc_41358_n419) );
  OR2X2 OR2X2_4995 ( .A(alu__abc_41358_n420), .B(alu__abc_41358_n412), .Y(alu__abc_41358_n421) );
  OR2X2 OR2X2_4996 ( .A(alu__abc_41358_n422), .B(alu__abc_41358_n411), .Y(alu__abc_41358_n423) );
  OR2X2 OR2X2_4997 ( .A(alu__abc_41358_n424), .B(alu__abc_41358_n408), .Y(alu__abc_41358_n425) );
  OR2X2 OR2X2_4998 ( .A(alu__abc_41358_n426), .B(alu__abc_41358_n407), .Y(alu__abc_41358_n427) );
  OR2X2 OR2X2_4999 ( .A(alu__abc_41358_n428), .B(alu__abc_41358_n404), .Y(alu__abc_41358_n429) );
  OR2X2 OR2X2_5 ( .A(_abc_43815_n668), .B(_abc_43815_n664_1), .Y(_abc_43815_n669) );
  OR2X2 OR2X2_50 ( .A(_abc_43815_n797), .B(_abc_43815_n795_1), .Y(_abc_43815_n798) );
  OR2X2 OR2X2_500 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_17_), .Y(_abc_43815_n2083) );
  OR2X2 OR2X2_5000 ( .A(alu__abc_41358_n434), .B(alu__abc_41358_n435), .Y(alu__abc_41358_n436) );
  OR2X2 OR2X2_5001 ( .A(alu__abc_41358_n442), .B(alu__abc_41358_n440), .Y(alu__abc_41358_n443) );
  OR2X2 OR2X2_5002 ( .A(alu__abc_41358_n443), .B(alu__abc_41358_n439), .Y(alu__abc_41358_n444) );
  OR2X2 OR2X2_5003 ( .A(alu__abc_41358_n449), .B(alu__abc_41358_n450), .Y(alu__abc_41358_n451) );
  OR2X2 OR2X2_5004 ( .A(alu__abc_41358_n457), .B(alu__abc_41358_n455), .Y(alu__abc_41358_n458) );
  OR2X2 OR2X2_5005 ( .A(alu__abc_41358_n458), .B(alu__abc_41358_n454), .Y(alu__abc_41358_n459) );
  OR2X2 OR2X2_5006 ( .A(alu__abc_41358_n445), .B(alu__abc_41358_n459), .Y(alu__abc_41358_n460) );
  OR2X2 OR2X2_5007 ( .A(alu__abc_41358_n430), .B(alu__abc_41358_n460), .Y(alu__abc_41358_n461) );
  OR2X2 OR2X2_5008 ( .A(alu__abc_41358_n466), .B(alu__abc_41358_n467), .Y(alu__abc_41358_n468) );
  OR2X2 OR2X2_5009 ( .A(alu__abc_41358_n474), .B(alu__abc_41358_n472), .Y(alu__abc_41358_n475) );
  OR2X2 OR2X2_501 ( .A(_abc_43815_n2048), .B(pc_q_18_), .Y(_abc_43815_n2086) );
  OR2X2 OR2X2_5010 ( .A(alu__abc_41358_n475), .B(alu__abc_41358_n471), .Y(alu__abc_41358_n476) );
  OR2X2 OR2X2_5011 ( .A(alu__abc_41358_n481), .B(alu__abc_41358_n482), .Y(alu__abc_41358_n483) );
  OR2X2 OR2X2_5012 ( .A(alu__abc_41358_n489), .B(alu__abc_41358_n487), .Y(alu__abc_41358_n490) );
  OR2X2 OR2X2_5013 ( .A(alu__abc_41358_n490), .B(alu__abc_41358_n486), .Y(alu__abc_41358_n491) );
  OR2X2 OR2X2_5014 ( .A(alu__abc_41358_n477), .B(alu__abc_41358_n491), .Y(alu__abc_41358_n492) );
  OR2X2 OR2X2_5015 ( .A(alu__abc_41358_n462), .B(alu__abc_41358_n492), .Y(alu__abc_41358_n493) );
  OR2X2 OR2X2_5016 ( .A(alu__abc_41358_n494), .B(alu__abc_41358_n403), .Y(alu__abc_41358_n495) );
  OR2X2 OR2X2_5017 ( .A(alu__abc_41358_n502), .B(alu__abc_41358_n497), .Y(alu__abc_41358_n503) );
  OR2X2 OR2X2_5018 ( .A(alu__abc_41358_n496), .B(alu__abc_41358_n504), .Y(alu__abc_41358_n505) );
  OR2X2 OR2X2_5019 ( .A(alu__abc_41358_n511), .B(alu__abc_41358_n387), .Y(alu_less_than_signed_o) );
  OR2X2 OR2X2_502 ( .A(_abc_43815_n2090), .B(_abc_43815_n1278_bF_buf7), .Y(_abc_43815_n2091) );
  OR2X2 OR2X2_5020 ( .A(alu__abc_41358_n514), .B(alu__abc_41358_n114), .Y(alu__abc_41358_n515) );
  OR2X2 OR2X2_5021 ( .A(alu__abc_41358_n518), .B(alu__abc_41358_n135_1), .Y(alu__abc_41358_n519) );
  OR2X2 OR2X2_5022 ( .A(alu__abc_41358_n517), .B(alu__abc_41358_n519), .Y(alu__abc_41358_n520) );
  OR2X2 OR2X2_5023 ( .A(alu__abc_41358_n526), .B(alu__abc_41358_n157), .Y(alu__abc_41358_n527) );
  OR2X2 OR2X2_5024 ( .A(alu__abc_41358_n531), .B(alu__abc_41358_n170), .Y(alu__abc_41358_n532) );
  OR2X2 OR2X2_5025 ( .A(alu__abc_41358_n529), .B(alu__abc_41358_n532), .Y(alu__abc_41358_n533) );
  OR2X2 OR2X2_5026 ( .A(alu__abc_41358_n525), .B(alu__abc_41358_n533), .Y(alu__abc_41358_n534) );
  OR2X2 OR2X2_5027 ( .A(alu__abc_41358_n539), .B(alu__abc_41358_n242), .Y(alu__abc_41358_n540) );
  OR2X2 OR2X2_5028 ( .A(alu__abc_41358_n543), .B(alu__abc_41358_n225), .Y(alu__abc_41358_n544) );
  OR2X2 OR2X2_5029 ( .A(alu__abc_41358_n542), .B(alu__abc_41358_n545), .Y(alu__abc_41358_n546) );
  OR2X2 OR2X2_503 ( .A(_abc_43815_n1431_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_43815_n2092) );
  OR2X2 OR2X2_5030 ( .A(alu__abc_41358_n548), .B(alu__abc_41358_n207), .Y(alu__abc_41358_n549) );
  OR2X2 OR2X2_5031 ( .A(alu__abc_41358_n552), .B(alu__abc_41358_n186), .Y(alu__abc_41358_n553) );
  OR2X2 OR2X2_5032 ( .A(alu__abc_41358_n551), .B(alu__abc_41358_n553), .Y(alu__abc_41358_n554) );
  OR2X2 OR2X2_5033 ( .A(alu__abc_41358_n547), .B(alu__abc_41358_n554), .Y(alu__abc_41358_n555) );
  OR2X2 OR2X2_5034 ( .A(alu__abc_41358_n556), .B(alu__abc_41358_n330), .Y(alu__abc_41358_n557) );
  OR2X2 OR2X2_5035 ( .A(alu__abc_41358_n558), .B(alu__abc_41358_n313), .Y(alu__abc_41358_n559) );
  OR2X2 OR2X2_5036 ( .A(alu__abc_41358_n561), .B(alu__abc_41358_n557), .Y(alu__abc_41358_n562) );
  OR2X2 OR2X2_5037 ( .A(alu__abc_41358_n564), .B(alu__abc_41358_n369), .Y(alu__abc_41358_n565_1) );
  OR2X2 OR2X2_5038 ( .A(alu__abc_41358_n568), .B(alu__abc_41358_n348), .Y(alu__abc_41358_n569) );
  OR2X2 OR2X2_5039 ( .A(alu__abc_41358_n567), .B(alu__abc_41358_n569), .Y(alu__abc_41358_n570) );
  OR2X2 OR2X2_504 ( .A(pc_q_18_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(_abc_43815_n2096) );
  OR2X2 OR2X2_5040 ( .A(alu__abc_41358_n573), .B(alu__abc_41358_n562), .Y(alu__abc_41358_n574) );
  OR2X2 OR2X2_5041 ( .A(alu_a_i_1_), .B(alu_b_i_1_bF_buf5), .Y(alu__abc_41358_n576) );
  OR2X2 OR2X2_5042 ( .A(alu__abc_41358_n579), .B(alu__abc_41358_n250), .Y(alu__abc_41358_n580) );
  OR2X2 OR2X2_5043 ( .A(alu__abc_41358_n296), .B(alu__abc_41358_n301), .Y(alu__abc_41358_n581) );
  OR2X2 OR2X2_5044 ( .A(alu__abc_41358_n585), .B(alu__abc_41358_n292), .Y(alu__abc_41358_n586) );
  OR2X2 OR2X2_5045 ( .A(alu__abc_41358_n583), .B(alu__abc_41358_n586), .Y(alu__abc_41358_n587) );
  OR2X2 OR2X2_5046 ( .A(alu__abc_41358_n277), .B(alu__abc_41358_n285), .Y(alu__abc_41358_n595) );
  OR2X2 OR2X2_5047 ( .A(alu__abc_41358_n599), .B(alu__abc_41358_n271), .Y(alu__abc_41358_n600) );
  OR2X2 OR2X2_5048 ( .A(alu__abc_41358_n597), .B(alu__abc_41358_n600), .Y(alu__abc_41358_n601) );
  OR2X2 OR2X2_5049 ( .A(alu__abc_41358_n593), .B(alu__abc_41358_n601), .Y(alu__abc_41358_n602) );
  OR2X2 OR2X2_505 ( .A(_abc_43815_n2095), .B(_abc_43815_n2099), .Y(_abc_43815_n2102) );
  OR2X2 OR2X2_5050 ( .A(alu__abc_41358_n606), .B(alu__abc_41358_n574), .Y(alu__abc_41358_n607) );
  OR2X2 OR2X2_5051 ( .A(alu__abc_41358_n611), .B(alu__abc_41358_n555), .Y(alu__abc_41358_n612) );
  OR2X2 OR2X2_5052 ( .A(alu__abc_41358_n616), .B(alu__abc_41358_n534), .Y(alu__abc_41358_n617) );
  OR2X2 OR2X2_5053 ( .A(alu__abc_41358_n615), .B(alu__abc_41358_n520), .Y(alu__abc_41358_n618) );
  OR2X2 OR2X2_5054 ( .A(alu__abc_41358_n619), .B(alu__abc_41358_n528), .Y(alu__abc_41358_n620_1) );
  OR2X2 OR2X2_5055 ( .A(alu__abc_41358_n624), .B(alu__abc_41358_n522), .Y(alu__abc_41358_n625) );
  OR2X2 OR2X2_5056 ( .A(alu__abc_41358_n623), .B(alu__abc_41358_n174), .Y(alu__abc_41358_n626) );
  OR2X2 OR2X2_5057 ( .A(alu__abc_41358_n620_1), .B(alu__abc_41358_n168), .Y(alu__abc_41358_n628) );
  OR2X2 OR2X2_5058 ( .A(alu__abc_41358_n633), .B(alu__abc_41358_n159_1), .Y(alu__abc_41358_n634) );
  OR2X2 OR2X2_5059 ( .A(alu__abc_41358_n632), .B(alu__abc_41358_n160_1), .Y(alu__abc_41358_n635) );
  OR2X2 OR2X2_506 ( .A(_abc_43815_n1428_bF_buf0), .B(_abc_43815_n2105), .Y(_abc_43815_n2106) );
  OR2X2 OR2X2_5060 ( .A(alu__abc_41358_n609), .B(alu__abc_41358_n541), .Y(alu__abc_41358_n638) );
  OR2X2 OR2X2_5061 ( .A(alu__abc_41358_n639), .B(alu__abc_41358_n545), .Y(alu__abc_41358_n640) );
  OR2X2 OR2X2_5062 ( .A(alu__abc_41358_n641), .B(alu__abc_41358_n550), .Y(alu__abc_41358_n642) );
  OR2X2 OR2X2_5063 ( .A(alu__abc_41358_n647), .B(alu__abc_41358_n648), .Y(alu__abc_41358_n649) );
  OR2X2 OR2X2_5064 ( .A(alu__abc_41358_n614), .B(alu__abc_41358_n516), .Y(alu__abc_41358_n650) );
  OR2X2 OR2X2_5065 ( .A(alu__abc_41358_n654), .B(alu__abc_41358_n141), .Y(alu__abc_41358_n655) );
  OR2X2 OR2X2_5066 ( .A(alu__abc_41358_n653), .B(alu__abc_41358_n142), .Y(alu__abc_41358_n656) );
  OR2X2 OR2X2_5067 ( .A(alu__abc_41358_n650), .B(alu__abc_41358_n133), .Y(alu__abc_41358_n658) );
  OR2X2 OR2X2_5068 ( .A(alu__abc_41358_n663), .B(alu__abc_41358_n664), .Y(alu__abc_41358_n665) );
  OR2X2 OR2X2_5069 ( .A(alu__abc_41358_n612), .B(alu__abc_41358_n124_1), .Y(alu__abc_41358_n666) );
  OR2X2 OR2X2_507 ( .A(_abc_43815_n2104), .B(_abc_43815_n2106), .Y(_abc_43815_n2107) );
  OR2X2 OR2X2_5070 ( .A(alu__abc_41358_n642), .B(alu__abc_41358_n184), .Y(alu__abc_41358_n671) );
  OR2X2 OR2X2_5071 ( .A(alu__abc_41358_n640), .B(alu__abc_41358_n201), .Y(alu__abc_41358_n675) );
  OR2X2 OR2X2_5072 ( .A(alu__abc_41358_n681), .B(alu__abc_41358_n682), .Y(alu__abc_41358_n683) );
  OR2X2 OR2X2_5073 ( .A(alu__abc_41358_n638), .B(alu__abc_41358_n219), .Y(alu__abc_41358_n684) );
  OR2X2 OR2X2_5074 ( .A(alu__abc_41358_n691), .B(alu__abc_41358_n689), .Y(alu__abc_41358_n692) );
  OR2X2 OR2X2_5075 ( .A(alu__abc_41358_n607), .B(alu__abc_41358_n236), .Y(alu__abc_41358_n693) );
  OR2X2 OR2X2_5076 ( .A(alu__abc_41358_n695), .B(alu__abc_41358_n570), .Y(alu__abc_41358_n696) );
  OR2X2 OR2X2_5077 ( .A(alu__abc_41358_n697), .B(alu__abc_41358_n559), .Y(alu__abc_41358_n698) );
  OR2X2 OR2X2_5078 ( .A(alu__abc_41358_n699), .B(alu__abc_41358_n322), .Y(alu__abc_41358_n700) );
  OR2X2 OR2X2_5079 ( .A(alu__abc_41358_n702), .B(alu__abc_41358_n703), .Y(alu__abc_41358_n704_1) );
  OR2X2 OR2X2_508 ( .A(_abc_43815_n2108), .B(_abc_43815_n1473_bF_buf3), .Y(_abc_43815_n2109) );
  OR2X2 OR2X2_5080 ( .A(alu__abc_41358_n254), .B(alu__abc_41358_n706), .Y(alu__abc_41358_n707) );
  OR2X2 OR2X2_5081 ( .A(alu__abc_41358_n708), .B(alu__abc_41358_n581), .Y(alu__abc_41358_n709) );
  OR2X2 OR2X2_5082 ( .A(alu__abc_41358_n711), .B(alu__abc_41358_n712), .Y(alu__abc_41358_n713) );
  OR2X2 OR2X2_5083 ( .A(alu__abc_41358_n716), .B(alu__abc_41358_n705), .Y(alu__abc_41358_n717) );
  OR2X2 OR2X2_5084 ( .A(alu__abc_41358_n719), .B(alu__abc_41358_n596), .Y(alu__abc_41358_n720) );
  OR2X2 OR2X2_5085 ( .A(alu__abc_41358_n721), .B(alu__abc_41358_n263), .Y(alu__abc_41358_n722) );
  OR2X2 OR2X2_5086 ( .A(alu__abc_41358_n711), .B(alu__abc_41358_n725), .Y(alu__abc_41358_n726) );
  OR2X2 OR2X2_5087 ( .A(alu__abc_41358_n727), .B(alu__abc_41358_n270), .Y(alu__abc_41358_n728) );
  OR2X2 OR2X2_5088 ( .A(alu__abc_41358_n730), .B(alu__abc_41358_n723), .Y(alu__abc_41358_n731) );
  OR2X2 OR2X2_5089 ( .A(alu__abc_41358_n720), .B(alu__abc_41358_n269), .Y(alu__abc_41358_n732) );
  OR2X2 OR2X2_509 ( .A(_abc_43815_n2089), .B(_abc_43815_n1472_1_bF_buf2), .Y(_abc_43815_n2110) );
  OR2X2 OR2X2_5090 ( .A(alu__abc_41358_n734), .B(alu__abc_41358_n277), .Y(alu__abc_41358_n735) );
  OR2X2 OR2X2_5091 ( .A(alu__abc_41358_n711), .B(alu__abc_41358_n284), .Y(alu__abc_41358_n737) );
  OR2X2 OR2X2_5092 ( .A(alu__abc_41358_n739), .B(alu__abc_41358_n736), .Y(alu__abc_41358_n740) );
  OR2X2 OR2X2_5093 ( .A(alu__abc_41358_n708), .B(alu__abc_41358_n301), .Y(alu__abc_41358_n746) );
  OR2X2 OR2X2_5094 ( .A(alu__abc_41358_n580), .B(alu__abc_41358_n747), .Y(alu__abc_41358_n748) );
  OR2X2 OR2X2_5095 ( .A(alu__abc_41358_n755_1), .B(alu__abc_41358_n297), .Y(alu__abc_41358_n756) );
  OR2X2 OR2X2_5096 ( .A(alu__abc_41358_n754), .B(alu__abc_41358_n757), .Y(alu__abc_41358_n758) );
  OR2X2 OR2X2_5097 ( .A(alu__abc_41358_n587), .B(alu__abc_41358_n283), .Y(alu__abc_41358_n760) );
  OR2X2 OR2X2_5098 ( .A(alu__abc_41358_n715), .B(alu__abc_41358_n768), .Y(alu__abc_41358_n769) );
  OR2X2 OR2X2_5099 ( .A(alu__abc_41358_n770), .B(alu__abc_41358_n312), .Y(alu__abc_41358_n771) );
  OR2X2 OR2X2_51 ( .A(_abc_43815_n800_1), .B(_abc_43815_n799), .Y(_abc_43815_n801) );
  OR2X2 OR2X2_510 ( .A(_abc_43815_n2111), .B(_abc_43815_n1350_bF_buf3), .Y(_abc_43815_n2112) );
  OR2X2 OR2X2_5100 ( .A(alu__abc_41358_n696), .B(alu__abc_41358_n311), .Y(alu__abc_41358_n772) );
  OR2X2 OR2X2_5101 ( .A(alu__abc_41358_n715), .B(alu__abc_41358_n774), .Y(alu__abc_41358_n775) );
  OR2X2 OR2X2_5102 ( .A(alu__abc_41358_n776), .B(alu__abc_41358_n347), .Y(alu__abc_41358_n777) );
  OR2X2 OR2X2_5103 ( .A(alu__abc_41358_n778), .B(alu__abc_41358_n566), .Y(alu__abc_41358_n779) );
  OR2X2 OR2X2_5104 ( .A(alu__abc_41358_n779), .B(alu__abc_41358_n346), .Y(alu__abc_41358_n780) );
  OR2X2 OR2X2_5105 ( .A(alu__abc_41358_n705), .B(alu__abc_41358_n357), .Y(alu__abc_41358_n782) );
  OR2X2 OR2X2_5106 ( .A(alu__abc_41358_n715), .B(alu__abc_41358_n364), .Y(alu__abc_41358_n784) );
  OR2X2 OR2X2_5107 ( .A(alu__abc_41358_n786), .B(alu__abc_41358_n783), .Y(alu__abc_41358_n787_1) );
  OR2X2 OR2X2_5108 ( .A(alu__abc_41358_n791), .B(alu__abc_41358_n305), .Y(alu__abc_41358_n792) );
  OR2X2 OR2X2_5109 ( .A(alu__abc_41358_n795), .B(alu__abc_41358_n793), .Y(alu__abc_41358_n796) );
  OR2X2 OR2X2_511 ( .A(_abc_43815_n2114), .B(_abc_43815_n2113), .Y(_abc_43815_n2115_1) );
  OR2X2 OR2X2_5110 ( .A(alu__abc_41358_n698), .B(alu__abc_41358_n328), .Y(alu__abc_41358_n798) );
  OR2X2 OR2X2_5111 ( .A(alu__abc_41358_n802), .B(alu__abc_41358_n340), .Y(alu__abc_41358_n803) );
  OR2X2 OR2X2_5112 ( .A(alu__abc_41358_n801), .B(alu__abc_41358_n804), .Y(alu__abc_41358_n805) );
  OR2X2 OR2X2_5113 ( .A(alu__abc_41358_n819), .B(alu__abc_41358_n817), .Y(alu__abc_41358_n820) );
  OR2X2 OR2X2_5114 ( .A(alu__abc_41358_n618), .B(alu__abc_41358_n151), .Y(alu__abc_41358_n821) );
  OR2X2 OR2X2_5115 ( .A(alu__abc_41358_n829), .B(alu__abc_41358_n617), .Y(alu__abc_41358_n830) );
  OR2X2 OR2X2_5116 ( .A(alu__abc_41358_n259_bF_buf2), .B(alu_a_i_1_), .Y(alu__abc_41358_n834) );
  OR2X2 OR2X2_5117 ( .A(alu_a_i_2_), .B(alu_b_i_0_bF_buf1), .Y(alu__abc_41358_n837) );
  OR2X2 OR2X2_5118 ( .A(alu__abc_41358_n259_bF_buf1), .B(alu_a_i_3_), .Y(alu__abc_41358_n838) );
  OR2X2 OR2X2_5119 ( .A(alu__abc_41358_n840), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n841) );
  OR2X2 OR2X2_512 ( .A(_abc_43815_n1413_bF_buf1), .B(_abc_43815_n2115_1), .Y(_abc_43815_n2116) );
  OR2X2 OR2X2_5120 ( .A(alu__abc_41358_n841), .B(alu__abc_41358_n836), .Y(alu__abc_41358_n842) );
  OR2X2 OR2X2_5121 ( .A(alu_a_i_4_), .B(alu_b_i_0_bF_buf0), .Y(alu__abc_41358_n843) );
  OR2X2 OR2X2_5122 ( .A(alu__abc_41358_n259_bF_buf0), .B(alu_a_i_5_), .Y(alu__abc_41358_n844) );
  OR2X2 OR2X2_5123 ( .A(alu__abc_41358_n845), .B(alu_b_i_1_bF_buf3), .Y(alu__abc_41358_n846) );
  OR2X2 OR2X2_5124 ( .A(alu_a_i_6_), .B(alu_b_i_0_bF_buf4), .Y(alu__abc_41358_n847_1) );
  OR2X2 OR2X2_5125 ( .A(alu__abc_41358_n259_bF_buf4), .B(alu_a_i_7_), .Y(alu__abc_41358_n848) );
  OR2X2 OR2X2_5126 ( .A(alu__abc_41358_n849), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n850) );
  OR2X2 OR2X2_5127 ( .A(alu__abc_41358_n851), .B(alu__abc_41358_n299_bF_buf5), .Y(alu__abc_41358_n852) );
  OR2X2 OR2X2_5128 ( .A(alu__abc_41358_n853), .B(alu_b_i_3_bF_buf3), .Y(alu__abc_41358_n854) );
  OR2X2 OR2X2_5129 ( .A(alu_a_i_8_), .B(alu_b_i_0_bF_buf3), .Y(alu__abc_41358_n855) );
  OR2X2 OR2X2_513 ( .A(_abc_43815_n2118), .B(_abc_43815_n2091), .Y(_abc_43815_n2119) );
  OR2X2 OR2X2_5130 ( .A(alu__abc_41358_n259_bF_buf3), .B(alu_a_i_9_), .Y(alu__abc_41358_n856) );
  OR2X2 OR2X2_5131 ( .A(alu__abc_41358_n857), .B(alu_b_i_1_bF_buf2), .Y(alu__abc_41358_n858) );
  OR2X2 OR2X2_5132 ( .A(alu_a_i_10_), .B(alu_b_i_0_bF_buf2), .Y(alu__abc_41358_n859) );
  OR2X2 OR2X2_5133 ( .A(alu__abc_41358_n259_bF_buf2), .B(alu_a_i_11_), .Y(alu__abc_41358_n860) );
  OR2X2 OR2X2_5134 ( .A(alu__abc_41358_n861), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n862) );
  OR2X2 OR2X2_5135 ( .A(alu__abc_41358_n863), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n864) );
  OR2X2 OR2X2_5136 ( .A(alu_a_i_12_), .B(alu_b_i_0_bF_buf1), .Y(alu__abc_41358_n865) );
  OR2X2 OR2X2_5137 ( .A(alu__abc_41358_n259_bF_buf1), .B(alu_a_i_13_), .Y(alu__abc_41358_n866) );
  OR2X2 OR2X2_5138 ( .A(alu__abc_41358_n867), .B(alu_b_i_1_bF_buf1), .Y(alu__abc_41358_n868) );
  OR2X2 OR2X2_5139 ( .A(alu_a_i_14_), .B(alu_b_i_0_bF_buf0), .Y(alu__abc_41358_n869) );
  OR2X2 OR2X2_514 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_18_), .Y(_abc_43815_n2120) );
  OR2X2 OR2X2_5140 ( .A(alu__abc_41358_n259_bF_buf0), .B(alu_a_i_15_), .Y(alu__abc_41358_n870) );
  OR2X2 OR2X2_5141 ( .A(alu__abc_41358_n871), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n872_1) );
  OR2X2 OR2X2_5142 ( .A(alu__abc_41358_n873), .B(alu__abc_41358_n299_bF_buf4), .Y(alu__abc_41358_n874) );
  OR2X2 OR2X2_5143 ( .A(alu__abc_41358_n875), .B(alu__abc_41358_n294_bF_buf5), .Y(alu__abc_41358_n876) );
  OR2X2 OR2X2_5144 ( .A(alu__abc_41358_n877), .B(alu_b_i_4_bF_buf2), .Y(alu__abc_41358_n878) );
  OR2X2 OR2X2_5145 ( .A(alu_a_i_16_), .B(alu_b_i_0_bF_buf4), .Y(alu__abc_41358_n879) );
  OR2X2 OR2X2_5146 ( .A(alu__abc_41358_n259_bF_buf4), .B(alu_a_i_17_), .Y(alu__abc_41358_n880) );
  OR2X2 OR2X2_5147 ( .A(alu__abc_41358_n881), .B(alu_b_i_1_bF_buf0), .Y(alu__abc_41358_n882) );
  OR2X2 OR2X2_5148 ( .A(alu_a_i_18_), .B(alu_b_i_0_bF_buf3), .Y(alu__abc_41358_n883) );
  OR2X2 OR2X2_5149 ( .A(alu__abc_41358_n259_bF_buf3), .B(alu_a_i_19_), .Y(alu__abc_41358_n884) );
  OR2X2 OR2X2_515 ( .A(_abc_43815_n2087_1), .B(pc_q_19_), .Y(_abc_43815_n2123) );
  OR2X2 OR2X2_5150 ( .A(alu__abc_41358_n885), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n886) );
  OR2X2 OR2X2_5151 ( .A(alu__abc_41358_n887), .B(alu_b_i_2_bF_buf2), .Y(alu__abc_41358_n888) );
  OR2X2 OR2X2_5152 ( .A(alu_a_i_20_), .B(alu_b_i_0_bF_buf2), .Y(alu__abc_41358_n889) );
  OR2X2 OR2X2_5153 ( .A(alu__abc_41358_n259_bF_buf2), .B(alu_a_i_21_), .Y(alu__abc_41358_n890) );
  OR2X2 OR2X2_5154 ( .A(alu__abc_41358_n891), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n892) );
  OR2X2 OR2X2_5155 ( .A(alu_a_i_22_), .B(alu_b_i_0_bF_buf1), .Y(alu__abc_41358_n893) );
  OR2X2 OR2X2_5156 ( .A(alu__abc_41358_n259_bF_buf1), .B(alu_a_i_23_), .Y(alu__abc_41358_n894) );
  OR2X2 OR2X2_5157 ( .A(alu__abc_41358_n895), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n896) );
  OR2X2 OR2X2_5158 ( .A(alu__abc_41358_n897), .B(alu__abc_41358_n299_bF_buf3), .Y(alu__abc_41358_n898) );
  OR2X2 OR2X2_5159 ( .A(alu__abc_41358_n899), .B(alu_b_i_3_bF_buf2), .Y(alu__abc_41358_n900) );
  OR2X2 OR2X2_516 ( .A(_abc_43815_n2127), .B(_abc_43815_n1278_bF_buf6), .Y(_abc_43815_n2128) );
  OR2X2 OR2X2_5160 ( .A(alu_a_i_24_), .B(alu_b_i_0_bF_buf0), .Y(alu__abc_41358_n901) );
  OR2X2 OR2X2_5161 ( .A(alu__abc_41358_n259_bF_buf0), .B(alu_a_i_25_), .Y(alu__abc_41358_n902) );
  OR2X2 OR2X2_5162 ( .A(alu__abc_41358_n903_1), .B(alu_b_i_1_bF_buf6), .Y(alu__abc_41358_n904) );
  OR2X2 OR2X2_5163 ( .A(alu_a_i_26_), .B(alu_b_i_0_bF_buf4), .Y(alu__abc_41358_n905) );
  OR2X2 OR2X2_5164 ( .A(alu__abc_41358_n259_bF_buf4), .B(alu_a_i_27_), .Y(alu__abc_41358_n906) );
  OR2X2 OR2X2_5165 ( .A(alu__abc_41358_n907), .B(alu__abc_41358_n252_bF_buf5), .Y(alu__abc_41358_n908) );
  OR2X2 OR2X2_5166 ( .A(alu__abc_41358_n909), .B(alu_b_i_2_bF_buf1), .Y(alu__abc_41358_n910) );
  OR2X2 OR2X2_5167 ( .A(alu_a_i_28_), .B(alu_b_i_0_bF_buf3), .Y(alu__abc_41358_n911) );
  OR2X2 OR2X2_5168 ( .A(alu__abc_41358_n259_bF_buf3), .B(alu_a_i_29_), .Y(alu__abc_41358_n912) );
  OR2X2 OR2X2_5169 ( .A(alu__abc_41358_n913), .B(alu_b_i_1_bF_buf5), .Y(alu__abc_41358_n914) );
  OR2X2 OR2X2_517 ( .A(pc_q_19_), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(_abc_43815_n2131) );
  OR2X2 OR2X2_5170 ( .A(alu_a_i_30_), .B(alu_b_i_0_bF_buf2), .Y(alu__abc_41358_n915) );
  OR2X2 OR2X2_5171 ( .A(alu__abc_41358_n259_bF_buf2), .B(alu_a_i_31_), .Y(alu__abc_41358_n916) );
  OR2X2 OR2X2_5172 ( .A(alu__abc_41358_n917), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n918) );
  OR2X2 OR2X2_5173 ( .A(alu__abc_41358_n919), .B(alu__abc_41358_n299_bF_buf2), .Y(alu__abc_41358_n920) );
  OR2X2 OR2X2_5174 ( .A(alu__abc_41358_n921), .B(alu__abc_41358_n294_bF_buf4), .Y(alu__abc_41358_n922) );
  OR2X2 OR2X2_5175 ( .A(alu__abc_41358_n923), .B(alu__abc_41358_n279_bF_buf3), .Y(alu__abc_41358_n924) );
  OR2X2 OR2X2_5176 ( .A(alu__abc_41358_n930), .B(alu_op_i_3_), .Y(alu__abc_41358_n931) );
  OR2X2 OR2X2_5177 ( .A(alu__abc_41358_n938), .B(alu__abc_41358_n936), .Y(alu__abc_41358_n939) );
  OR2X2 OR2X2_5178 ( .A(alu__abc_41358_n933_1), .B(alu__abc_41358_n939), .Y(alu__abc_41358_n940) );
  OR2X2 OR2X2_5179 ( .A(alu__abc_41358_n743), .B(alu_c_i), .Y(alu__abc_41358_n944) );
  OR2X2 OR2X2_518 ( .A(_abc_43815_n2130), .B(_abc_43815_n2134), .Y(_abc_43815_n2135) );
  OR2X2 OR2X2_5180 ( .A(alu__abc_41358_n946), .B(alu__abc_41358_n952), .Y(alu__abc_41358_n953_1) );
  OR2X2 OR2X2_5181 ( .A(alu__abc_41358_n955), .B(alu__abc_41358_n954), .Y(alu__abc_41358_n956) );
  OR2X2 OR2X2_5182 ( .A(alu__abc_41358_n953_1), .B(alu__abc_41358_n957), .Y(alu__abc_41358_n958) );
  OR2X2 OR2X2_5183 ( .A(alu__abc_41358_n958), .B(alu__abc_41358_n940), .Y(alu__abc_41358_n959) );
  OR2X2 OR2X2_5184 ( .A(alu__abc_41358_n926), .B(alu__abc_41358_n959), .Y(alu_p_o_0_) );
  OR2X2 OR2X2_5185 ( .A(alu__abc_41358_n962), .B(alu__abc_41358_n963), .Y(alu__abc_41358_n964) );
  OR2X2 OR2X2_5186 ( .A(alu__abc_41358_n967), .B(alu__abc_41358_n966), .Y(alu__abc_41358_n968) );
  OR2X2 OR2X2_5187 ( .A(alu__abc_41358_n965), .B(alu__abc_41358_n969), .Y(alu__abc_41358_n970) );
  OR2X2 OR2X2_5188 ( .A(alu_a_i_25_), .B(alu_b_i_0_bF_buf0), .Y(alu__abc_41358_n972) );
  OR2X2 OR2X2_5189 ( .A(alu__abc_41358_n259_bF_buf4), .B(alu_a_i_26_), .Y(alu__abc_41358_n973) );
  OR2X2 OR2X2_519 ( .A(_abc_43815_n2129_1), .B(_abc_43815_n2136), .Y(_abc_43815_n2137) );
  OR2X2 OR2X2_5190 ( .A(alu__abc_41358_n974), .B(alu_b_i_1_bF_buf3), .Y(alu__abc_41358_n975_1) );
  OR2X2 OR2X2_5191 ( .A(alu_a_i_27_), .B(alu_b_i_0_bF_buf4), .Y(alu__abc_41358_n976) );
  OR2X2 OR2X2_5192 ( .A(alu__abc_41358_n259_bF_buf3), .B(alu_a_i_28_), .Y(alu__abc_41358_n977) );
  OR2X2 OR2X2_5193 ( .A(alu__abc_41358_n978), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n979) );
  OR2X2 OR2X2_5194 ( .A(alu__abc_41358_n971), .B(alu__abc_41358_n981), .Y(alu__abc_41358_n982) );
  OR2X2 OR2X2_5195 ( .A(alu_a_i_17_), .B(alu_b_i_0_bF_buf3), .Y(alu__abc_41358_n984) );
  OR2X2 OR2X2_5196 ( .A(alu__abc_41358_n259_bF_buf2), .B(alu_a_i_18_), .Y(alu__abc_41358_n985) );
  OR2X2 OR2X2_5197 ( .A(alu__abc_41358_n986), .B(alu_b_i_1_bF_buf2), .Y(alu__abc_41358_n987) );
  OR2X2 OR2X2_5198 ( .A(alu_a_i_19_), .B(alu_b_i_0_bF_buf2), .Y(alu__abc_41358_n988) );
  OR2X2 OR2X2_5199 ( .A(alu__abc_41358_n259_bF_buf1), .B(alu_a_i_20_), .Y(alu__abc_41358_n989) );
  OR2X2 OR2X2_52 ( .A(_abc_43815_n802), .B(_abc_43815_n803), .Y(_abc_43815_n804) );
  OR2X2 OR2X2_520 ( .A(_abc_43815_n1428_bF_buf4), .B(_abc_43815_n2140), .Y(_abc_43815_n2141) );
  OR2X2 OR2X2_5200 ( .A(alu__abc_41358_n990), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n991) );
  OR2X2 OR2X2_5201 ( .A(alu__abc_41358_n992), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n993) );
  OR2X2 OR2X2_5202 ( .A(alu_a_i_21_), .B(alu_b_i_0_bF_buf1), .Y(alu__abc_41358_n994) );
  OR2X2 OR2X2_5203 ( .A(alu__abc_41358_n259_bF_buf0), .B(alu_a_i_22_), .Y(alu__abc_41358_n995) );
  OR2X2 OR2X2_5204 ( .A(alu__abc_41358_n996), .B(alu_b_i_1_bF_buf1), .Y(alu__abc_41358_n997) );
  OR2X2 OR2X2_5205 ( .A(alu_a_i_23_), .B(alu_b_i_0_bF_buf0), .Y(alu__abc_41358_n998) );
  OR2X2 OR2X2_5206 ( .A(alu__abc_41358_n259_bF_buf4), .B(alu_a_i_24_), .Y(alu__abc_41358_n999) );
  OR2X2 OR2X2_5207 ( .A(alu__abc_41358_n1000), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n1001_1) );
  OR2X2 OR2X2_5208 ( .A(alu__abc_41358_n1002), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n1003) );
  OR2X2 OR2X2_5209 ( .A(alu__abc_41358_n983), .B(alu__abc_41358_n1005), .Y(alu__abc_41358_n1006) );
  OR2X2 OR2X2_521 ( .A(_abc_43815_n2139), .B(_abc_43815_n2141), .Y(_abc_43815_n2142) );
  OR2X2 OR2X2_5210 ( .A(alu__abc_41358_n1006), .B(alu__abc_41358_n279_bF_buf1), .Y(alu__abc_41358_n1007) );
  OR2X2 OR2X2_5211 ( .A(alu__abc_41358_n259_bF_buf3), .B(alu_a_i_2_), .Y(alu__abc_41358_n1008) );
  OR2X2 OR2X2_5212 ( .A(alu_a_i_1_), .B(alu_b_i_0_bF_buf4), .Y(alu__abc_41358_n1009) );
  OR2X2 OR2X2_5213 ( .A(alu_a_i_3_), .B(alu_b_i_0_bF_buf3), .Y(alu__abc_41358_n1012) );
  OR2X2 OR2X2_5214 ( .A(alu__abc_41358_n259_bF_buf2), .B(alu_a_i_4_), .Y(alu__abc_41358_n1013) );
  OR2X2 OR2X2_5215 ( .A(alu__abc_41358_n1015), .B(alu__abc_41358_n1011), .Y(alu__abc_41358_n1016) );
  OR2X2 OR2X2_5216 ( .A(alu__abc_41358_n1016), .B(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n1017) );
  OR2X2 OR2X2_5217 ( .A(alu_a_i_5_), .B(alu_b_i_0_bF_buf2), .Y(alu__abc_41358_n1018) );
  OR2X2 OR2X2_5218 ( .A(alu__abc_41358_n259_bF_buf1), .B(alu_a_i_6_), .Y(alu__abc_41358_n1019) );
  OR2X2 OR2X2_5219 ( .A(alu__abc_41358_n1020), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n1021) );
  OR2X2 OR2X2_522 ( .A(_abc_43815_n1431_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_43815_n2143_1) );
  OR2X2 OR2X2_5220 ( .A(alu_a_i_7_), .B(alu_b_i_0_bF_buf1), .Y(alu__abc_41358_n1022) );
  OR2X2 OR2X2_5221 ( .A(alu__abc_41358_n259_bF_buf0), .B(alu_a_i_8_), .Y(alu__abc_41358_n1023) );
  OR2X2 OR2X2_5222 ( .A(alu__abc_41358_n1024_1), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n1025) );
  OR2X2 OR2X2_5223 ( .A(alu__abc_41358_n1026), .B(alu__abc_41358_n299_bF_buf6), .Y(alu__abc_41358_n1027) );
  OR2X2 OR2X2_5224 ( .A(alu__abc_41358_n1028), .B(alu_b_i_3_bF_buf0), .Y(alu__abc_41358_n1029) );
  OR2X2 OR2X2_5225 ( .A(alu_a_i_9_), .B(alu_b_i_0_bF_buf0), .Y(alu__abc_41358_n1030) );
  OR2X2 OR2X2_5226 ( .A(alu__abc_41358_n259_bF_buf4), .B(alu_a_i_10_), .Y(alu__abc_41358_n1031) );
  OR2X2 OR2X2_5227 ( .A(alu__abc_41358_n1032), .B(alu_b_i_1_bF_buf6), .Y(alu__abc_41358_n1033) );
  OR2X2 OR2X2_5228 ( .A(alu_a_i_11_), .B(alu_b_i_0_bF_buf4), .Y(alu__abc_41358_n1034) );
  OR2X2 OR2X2_5229 ( .A(alu__abc_41358_n259_bF_buf3), .B(alu_a_i_12_), .Y(alu__abc_41358_n1035) );
  OR2X2 OR2X2_523 ( .A(_abc_43815_n2145), .B(_abc_43815_n2146), .Y(_abc_43815_n2147) );
  OR2X2 OR2X2_5230 ( .A(alu__abc_41358_n1036), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n1037) );
  OR2X2 OR2X2_5231 ( .A(alu__abc_41358_n1038), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n1039) );
  OR2X2 OR2X2_5232 ( .A(alu_a_i_13_), .B(alu_b_i_0_bF_buf3), .Y(alu__abc_41358_n1040) );
  OR2X2 OR2X2_5233 ( .A(alu__abc_41358_n259_bF_buf2), .B(alu_a_i_14_), .Y(alu__abc_41358_n1041) );
  OR2X2 OR2X2_5234 ( .A(alu__abc_41358_n1042), .B(alu_b_i_1_bF_buf5), .Y(alu__abc_41358_n1043) );
  OR2X2 OR2X2_5235 ( .A(alu_a_i_15_), .B(alu_b_i_0_bF_buf2), .Y(alu__abc_41358_n1044) );
  OR2X2 OR2X2_5236 ( .A(alu__abc_41358_n259_bF_buf1), .B(alu_a_i_16_), .Y(alu__abc_41358_n1045) );
  OR2X2 OR2X2_5237 ( .A(alu__abc_41358_n1046), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n1047) );
  OR2X2 OR2X2_5238 ( .A(alu__abc_41358_n1048), .B(alu__abc_41358_n299_bF_buf5), .Y(alu__abc_41358_n1049) );
  OR2X2 OR2X2_5239 ( .A(alu__abc_41358_n1050_1), .B(alu__abc_41358_n294_bF_buf1), .Y(alu__abc_41358_n1051) );
  OR2X2 OR2X2_524 ( .A(_abc_43815_n2147), .B(_abc_43815_n1350_bF_buf2), .Y(_abc_43815_n2148) );
  OR2X2 OR2X2_5240 ( .A(alu__abc_41358_n1052), .B(alu_b_i_4_bF_buf1), .Y(alu__abc_41358_n1053) );
  OR2X2 OR2X2_5241 ( .A(alu__abc_41358_n254), .B(alu__abc_41358_n257), .Y(alu__abc_41358_n1058) );
  OR2X2 OR2X2_5242 ( .A(alu__abc_41358_n577), .B(alu__abc_41358_n578), .Y(alu__abc_41358_n1062) );
  OR2X2 OR2X2_5243 ( .A(alu__abc_41358_n1064), .B(alu__abc_41358_n1068), .Y(alu__abc_41358_n1069) );
  OR2X2 OR2X2_5244 ( .A(alu__abc_41358_n1069), .B(alu__abc_41358_n1060), .Y(alu__abc_41358_n1070) );
  OR2X2 OR2X2_5245 ( .A(alu__abc_41358_n1063), .B(alu__abc_41358_n744), .Y(alu__abc_41358_n1071) );
  OR2X2 OR2X2_5246 ( .A(alu__abc_41358_n1079), .B(alu__abc_41358_n1080), .Y(alu__abc_41358_n1081) );
  OR2X2 OR2X2_5247 ( .A(alu__abc_41358_n1081), .B(alu__abc_41358_n1078), .Y(alu__abc_41358_n1082) );
  OR2X2 OR2X2_5248 ( .A(alu__abc_41358_n1082), .B(alu__abc_41358_n1074_1), .Y(alu__abc_41358_n1083) );
  OR2X2 OR2X2_5249 ( .A(alu__abc_41358_n1083), .B(alu__abc_41358_n1070), .Y(alu__abc_41358_n1084) );
  OR2X2 OR2X2_525 ( .A(_abc_43815_n2150), .B(_abc_43815_n2149), .Y(_abc_43815_n2151) );
  OR2X2 OR2X2_5250 ( .A(alu__abc_41358_n1055), .B(alu__abc_41358_n1084), .Y(alu_p_o_1_) );
  OR2X2 OR2X2_5251 ( .A(alu__abc_41358_n917), .B(alu_b_i_1_bF_buf4), .Y(alu__abc_41358_n1086) );
  OR2X2 OR2X2_5252 ( .A(alu__abc_41358_n962), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n1087) );
  OR2X2 OR2X2_5253 ( .A(alu__abc_41358_n907), .B(alu_b_i_1_bF_buf3), .Y(alu__abc_41358_n1090) );
  OR2X2 OR2X2_5254 ( .A(alu__abc_41358_n913), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n1091) );
  OR2X2 OR2X2_5255 ( .A(alu__abc_41358_n1089), .B(alu__abc_41358_n1093), .Y(alu__abc_41358_n1094) );
  OR2X2 OR2X2_5256 ( .A(alu__abc_41358_n885), .B(alu_b_i_1_bF_buf2), .Y(alu__abc_41358_n1096) );
  OR2X2 OR2X2_5257 ( .A(alu__abc_41358_n891), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n1097_1) );
  OR2X2 OR2X2_5258 ( .A(alu__abc_41358_n1098), .B(alu_b_i_2_bF_buf2), .Y(alu__abc_41358_n1099) );
  OR2X2 OR2X2_5259 ( .A(alu__abc_41358_n895), .B(alu_b_i_1_bF_buf1), .Y(alu__abc_41358_n1100) );
  OR2X2 OR2X2_526 ( .A(_abc_43815_n1413_bF_buf0), .B(_abc_43815_n2151), .Y(_abc_43815_n2152) );
  OR2X2 OR2X2_5260 ( .A(alu__abc_41358_n903_1), .B(alu__abc_41358_n252_bF_buf5), .Y(alu__abc_41358_n1101) );
  OR2X2 OR2X2_5261 ( .A(alu__abc_41358_n1102), .B(alu__abc_41358_n299_bF_buf2), .Y(alu__abc_41358_n1103) );
  OR2X2 OR2X2_5262 ( .A(alu__abc_41358_n1095), .B(alu__abc_41358_n1105), .Y(alu__abc_41358_n1106) );
  OR2X2 OR2X2_5263 ( .A(alu__abc_41358_n1106), .B(alu__abc_41358_n279_bF_buf0), .Y(alu__abc_41358_n1107) );
  OR2X2 OR2X2_5264 ( .A(alu__abc_41358_n1109), .B(alu_b_i_2_bF_buf1), .Y(alu__abc_41358_n1110) );
  OR2X2 OR2X2_5265 ( .A(alu__abc_41358_n1110), .B(alu__abc_41358_n1108), .Y(alu__abc_41358_n1111) );
  OR2X2 OR2X2_5266 ( .A(alu__abc_41358_n849), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n1112) );
  OR2X2 OR2X2_5267 ( .A(alu__abc_41358_n857), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n1113) );
  OR2X2 OR2X2_5268 ( .A(alu__abc_41358_n1114), .B(alu__abc_41358_n299_bF_buf1), .Y(alu__abc_41358_n1115) );
  OR2X2 OR2X2_5269 ( .A(alu__abc_41358_n861), .B(alu_b_i_1_bF_buf6), .Y(alu__abc_41358_n1118) );
  OR2X2 OR2X2_527 ( .A(_abc_43815_n2154), .B(_abc_43815_n2128), .Y(_abc_43815_n2155) );
  OR2X2 OR2X2_5270 ( .A(alu__abc_41358_n867), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n1119) );
  OR2X2 OR2X2_5271 ( .A(alu__abc_41358_n1120), .B(alu_b_i_2_bF_buf0), .Y(alu__abc_41358_n1121) );
  OR2X2 OR2X2_5272 ( .A(alu__abc_41358_n871), .B(alu_b_i_1_bF_buf5), .Y(alu__abc_41358_n1122) );
  OR2X2 OR2X2_5273 ( .A(alu__abc_41358_n881), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n1123) );
  OR2X2 OR2X2_5274 ( .A(alu__abc_41358_n1124), .B(alu__abc_41358_n299_bF_buf0), .Y(alu__abc_41358_n1125) );
  OR2X2 OR2X2_5275 ( .A(alu__abc_41358_n1127), .B(alu_b_i_4_bF_buf0), .Y(alu__abc_41358_n1128) );
  OR2X2 OR2X2_5276 ( .A(alu__abc_41358_n1128), .B(alu__abc_41358_n1117_1), .Y(alu__abc_41358_n1129) );
  OR2X2 OR2X2_5277 ( .A(alu__abc_41358_n417), .B(alu__abc_41358_n301), .Y(alu__abc_41358_n1138) );
  OR2X2 OR2X2_5278 ( .A(alu__abc_41358_n1141), .B(alu_b_i_1_bF_buf4), .Y(alu__abc_41358_n1142) );
  OR2X2 OR2X2_5279 ( .A(alu__abc_41358_n1140), .B(alu__abc_41358_n1148), .Y(alu__abc_41358_n1149) );
  OR2X2 OR2X2_528 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_19_), .Y(_abc_43815_n2156) );
  OR2X2 OR2X2_5280 ( .A(alu__abc_41358_n1149), .B(alu__abc_41358_n1136), .Y(alu__abc_41358_n1150) );
  OR2X2 OR2X2_5281 ( .A(alu__abc_41358_n749), .B(alu__abc_41358_n745), .Y(alu__abc_41358_n1152) );
  OR2X2 OR2X2_5282 ( .A(alu__abc_41358_n1156), .B(alu__abc_41358_n1157), .Y(alu__abc_41358_n1158_1) );
  OR2X2 OR2X2_5283 ( .A(alu__abc_41358_n1155), .B(alu__abc_41358_n1158_1), .Y(alu__abc_41358_n1159) );
  OR2X2 OR2X2_5284 ( .A(alu__abc_41358_n1154), .B(alu__abc_41358_n1159), .Y(alu__abc_41358_n1160) );
  OR2X2 OR2X2_5285 ( .A(alu__abc_41358_n1160), .B(alu__abc_41358_n1150), .Y(alu__abc_41358_n1161) );
  OR2X2 OR2X2_5286 ( .A(alu__abc_41358_n1161), .B(alu__abc_41358_n1131), .Y(alu_p_o_2_) );
  OR2X2 OR2X2_5287 ( .A(alu__abc_41358_n978), .B(alu_b_i_1_bF_buf2), .Y(alu__abc_41358_n1165) );
  OR2X2 OR2X2_5288 ( .A(alu__abc_41358_n968), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n1166) );
  OR2X2 OR2X2_5289 ( .A(alu__abc_41358_n1164), .B(alu__abc_41358_n1168), .Y(alu__abc_41358_n1169) );
  OR2X2 OR2X2_529 ( .A(_abc_43815_n2124), .B(pc_q_20_), .Y(_abc_43815_n2159) );
  OR2X2 OR2X2_5290 ( .A(alu__abc_41358_n990), .B(alu_b_i_1_bF_buf1), .Y(alu__abc_41358_n1171) );
  OR2X2 OR2X2_5291 ( .A(alu__abc_41358_n996), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n1172) );
  OR2X2 OR2X2_5292 ( .A(alu__abc_41358_n1173), .B(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n1174) );
  OR2X2 OR2X2_5293 ( .A(alu__abc_41358_n1000), .B(alu_b_i_1_bF_buf0), .Y(alu__abc_41358_n1175) );
  OR2X2 OR2X2_5294 ( .A(alu__abc_41358_n974), .B(alu__abc_41358_n252_bF_buf5), .Y(alu__abc_41358_n1176) );
  OR2X2 OR2X2_5295 ( .A(alu__abc_41358_n1177), .B(alu__abc_41358_n299_bF_buf5), .Y(alu__abc_41358_n1178) );
  OR2X2 OR2X2_5296 ( .A(alu__abc_41358_n1170), .B(alu__abc_41358_n1180), .Y(alu__abc_41358_n1181_1) );
  OR2X2 OR2X2_5297 ( .A(alu__abc_41358_n1181_1), .B(alu__abc_41358_n279_bF_buf5), .Y(alu__abc_41358_n1182) );
  OR2X2 OR2X2_5298 ( .A(alu__abc_41358_n1184), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n1185) );
  OR2X2 OR2X2_5299 ( .A(alu__abc_41358_n1185), .B(alu__abc_41358_n1183), .Y(alu__abc_41358_n1186) );
  OR2X2 OR2X2_53 ( .A(_abc_43815_n804), .B(_abc_43815_n801), .Y(_abc_43815_n805) );
  OR2X2 OR2X2_530 ( .A(_abc_43815_n2163), .B(_abc_43815_n1278_bF_buf5), .Y(_abc_43815_n2164) );
  OR2X2 OR2X2_5300 ( .A(alu__abc_41358_n1024_1), .B(alu_b_i_1_bF_buf6), .Y(alu__abc_41358_n1187) );
  OR2X2 OR2X2_5301 ( .A(alu__abc_41358_n1032), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n1188) );
  OR2X2 OR2X2_5302 ( .A(alu__abc_41358_n1189), .B(alu__abc_41358_n299_bF_buf4), .Y(alu__abc_41358_n1190) );
  OR2X2 OR2X2_5303 ( .A(alu__abc_41358_n1036), .B(alu_b_i_1_bF_buf5), .Y(alu__abc_41358_n1193) );
  OR2X2 OR2X2_5304 ( .A(alu__abc_41358_n1042), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n1194) );
  OR2X2 OR2X2_5305 ( .A(alu__abc_41358_n1195), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n1196) );
  OR2X2 OR2X2_5306 ( .A(alu__abc_41358_n1046), .B(alu_b_i_1_bF_buf4), .Y(alu__abc_41358_n1197) );
  OR2X2 OR2X2_5307 ( .A(alu__abc_41358_n986), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n1198) );
  OR2X2 OR2X2_5308 ( .A(alu__abc_41358_n1199), .B(alu__abc_41358_n299_bF_buf3), .Y(alu__abc_41358_n1200) );
  OR2X2 OR2X2_5309 ( .A(alu__abc_41358_n1202_1), .B(alu_b_i_4_bF_buf4), .Y(alu__abc_41358_n1203) );
  OR2X2 OR2X2_531 ( .A(_abc_43815_n2170), .B(_abc_43815_n2132), .Y(_abc_43815_n2171) );
  OR2X2 OR2X2_5310 ( .A(alu__abc_41358_n1203), .B(alu__abc_41358_n1192), .Y(alu__abc_41358_n1204) );
  OR2X2 OR2X2_5311 ( .A(alu__abc_41358_n758), .B(alu__abc_41358_n750), .Y(alu__abc_41358_n1207) );
  OR2X2 OR2X2_5312 ( .A(alu__abc_41358_n1212), .B(alu__abc_41358_n751), .Y(alu__abc_41358_n1213) );
  OR2X2 OR2X2_5313 ( .A(alu__abc_41358_n419), .B(alu__abc_41358_n296), .Y(alu__abc_41358_n1214) );
  OR2X2 OR2X2_5314 ( .A(alu__abc_41358_n1218), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n1219) );
  OR2X2 OR2X2_5315 ( .A(alu__abc_41358_n1220), .B(alu_b_i_1_bF_buf3), .Y(alu__abc_41358_n1221) );
  OR2X2 OR2X2_5316 ( .A(alu__abc_41358_n1230), .B(alu__abc_41358_n1231), .Y(alu__abc_41358_n1232) );
  OR2X2 OR2X2_5317 ( .A(alu__abc_41358_n1232), .B(alu__abc_41358_n1229), .Y(alu__abc_41358_n1233) );
  OR2X2 OR2X2_5318 ( .A(alu__abc_41358_n1225), .B(alu__abc_41358_n1233), .Y(alu__abc_41358_n1234) );
  OR2X2 OR2X2_5319 ( .A(alu__abc_41358_n1217), .B(alu__abc_41358_n1234), .Y(alu__abc_41358_n1235) );
  OR2X2 OR2X2_532 ( .A(_abc_43815_n2169), .B(_abc_43815_n2171), .Y(_abc_43815_n2172) );
  OR2X2 OR2X2_5320 ( .A(alu__abc_41358_n1235), .B(alu__abc_41358_n1216), .Y(alu__abc_41358_n1236) );
  OR2X2 OR2X2_5321 ( .A(alu__abc_41358_n1210), .B(alu__abc_41358_n1236), .Y(alu__abc_41358_n1237) );
  OR2X2 OR2X2_5322 ( .A(alu__abc_41358_n1237), .B(alu__abc_41358_n1206), .Y(alu_p_o_3_) );
  OR2X2 OR2X2_5323 ( .A(alu__abc_41358_n759), .B(alu__abc_41358_n761), .Y(alu__abc_41358_n1240) );
  OR2X2 OR2X2_5324 ( .A(alu__abc_41358_n851), .B(alu_b_i_2_bF_buf2), .Y(alu__abc_41358_n1243_1) );
  OR2X2 OR2X2_5325 ( .A(alu__abc_41358_n863), .B(alu__abc_41358_n299_bF_buf1), .Y(alu__abc_41358_n1244) );
  OR2X2 OR2X2_5326 ( .A(alu__abc_41358_n887), .B(alu__abc_41358_n299_bF_buf0), .Y(alu__abc_41358_n1247) );
  OR2X2 OR2X2_5327 ( .A(alu__abc_41358_n873), .B(alu_b_i_2_bF_buf1), .Y(alu__abc_41358_n1248) );
  OR2X2 OR2X2_5328 ( .A(alu__abc_41358_n1250), .B(alu__abc_41358_n1246), .Y(alu__abc_41358_n1251) );
  OR2X2 OR2X2_5329 ( .A(alu__abc_41358_n1251), .B(alu_b_i_4_bF_buf3), .Y(alu__abc_41358_n1252) );
  OR2X2 OR2X2_533 ( .A(_abc_43815_n2167), .B(_abc_43815_n2172), .Y(_abc_43815_n2173_1) );
  OR2X2 OR2X2_5330 ( .A(alu__abc_41358_n897), .B(alu_b_i_2_bF_buf0), .Y(alu__abc_41358_n1253) );
  OR2X2 OR2X2_5331 ( .A(alu__abc_41358_n909), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n1254) );
  OR2X2 OR2X2_5332 ( .A(alu__abc_41358_n1255), .B(alu_b_i_3_bF_buf1), .Y(alu__abc_41358_n1256) );
  OR2X2 OR2X2_5333 ( .A(alu__abc_41358_n1258), .B(alu__abc_41358_n1257), .Y(alu__abc_41358_n1259) );
  OR2X2 OR2X2_5334 ( .A(alu__abc_41358_n1259), .B(alu__abc_41358_n294_bF_buf0), .Y(alu__abc_41358_n1260) );
  OR2X2 OR2X2_5335 ( .A(alu__abc_41358_n1261), .B(alu__abc_41358_n279_bF_buf4), .Y(alu__abc_41358_n1262) );
  OR2X2 OR2X2_5336 ( .A(alu__abc_41358_n421), .B(alu__abc_41358_n284), .Y(alu__abc_41358_n1266) );
  OR2X2 OR2X2_5337 ( .A(alu__abc_41358_n949), .B(alu__abc_41358_n299_bF_buf5), .Y(alu__abc_41358_n1270) );
  OR2X2 OR2X2_5338 ( .A(alu__abc_41358_n1271), .B(alu_b_i_1_bF_buf2), .Y(alu__abc_41358_n1272) );
  OR2X2 OR2X2_5339 ( .A(alu__abc_41358_n1141), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n1273) );
  OR2X2 OR2X2_534 ( .A(pc_q_20_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(_abc_43815_n2174) );
  OR2X2 OR2X2_5340 ( .A(alu__abc_41358_n1274), .B(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n1275) );
  OR2X2 OR2X2_5341 ( .A(alu__abc_41358_n1284_1), .B(alu__abc_41358_n1280), .Y(alu__abc_41358_n1285) );
  OR2X2 OR2X2_5342 ( .A(alu__abc_41358_n1279), .B(alu__abc_41358_n1285), .Y(alu__abc_41358_n1286) );
  OR2X2 OR2X2_5343 ( .A(alu__abc_41358_n1278), .B(alu__abc_41358_n1286), .Y(alu__abc_41358_n1287) );
  OR2X2 OR2X2_5344 ( .A(alu__abc_41358_n1269), .B(alu__abc_41358_n1287), .Y(alu__abc_41358_n1288) );
  OR2X2 OR2X2_5345 ( .A(alu__abc_41358_n1268), .B(alu__abc_41358_n1288), .Y(alu__abc_41358_n1289) );
  OR2X2 OR2X2_5346 ( .A(alu__abc_41358_n1289), .B(alu__abc_41358_n1264_1), .Y(alu__abc_41358_n1290) );
  OR2X2 OR2X2_5347 ( .A(alu__abc_41358_n1290), .B(alu__abc_41358_n1242), .Y(alu_p_o_4_) );
  OR2X2 OR2X2_5348 ( .A(alu__abc_41358_n740), .B(alu__abc_41358_n762), .Y(alu__abc_41358_n1293) );
  OR2X2 OR2X2_5349 ( .A(alu__abc_41358_n1302), .B(alu_b_i_1_bF_buf1), .Y(alu__abc_41358_n1303) );
  OR2X2 OR2X2_535 ( .A(_abc_43815_n2173_1), .B(_abc_43815_n2177), .Y(_abc_43815_n2178) );
  OR2X2 OR2X2_5350 ( .A(alu__abc_41358_n1220), .B(alu__abc_41358_n252_bF_buf5), .Y(alu__abc_41358_n1304_1) );
  OR2X2 OR2X2_5351 ( .A(alu__abc_41358_n1306), .B(alu__abc_41358_n1301), .Y(alu__abc_41358_n1307) );
  OR2X2 OR2X2_5352 ( .A(alu__abc_41358_n1310), .B(alu__abc_41358_n1311), .Y(alu__abc_41358_n1312) );
  OR2X2 OR2X2_5353 ( .A(alu__abc_41358_n1309), .B(alu__abc_41358_n1312), .Y(alu__abc_41358_n1313) );
  OR2X2 OR2X2_5354 ( .A(alu__abc_41358_n1300), .B(alu__abc_41358_n1313), .Y(alu__abc_41358_n1314) );
  OR2X2 OR2X2_5355 ( .A(alu__abc_41358_n1314), .B(alu__abc_41358_n1299), .Y(alu__abc_41358_n1315) );
  OR2X2 OR2X2_5356 ( .A(alu__abc_41358_n1315), .B(alu__abc_41358_n1295), .Y(alu__abc_41358_n1316) );
  OR2X2 OR2X2_5357 ( .A(alu__abc_41358_n423), .B(alu__abc_41358_n289), .Y(alu__abc_41358_n1317) );
  OR2X2 OR2X2_5358 ( .A(alu__abc_41358_n1319), .B(alu__abc_41358_n590), .Y(alu__abc_41358_n1320) );
  OR2X2 OR2X2_5359 ( .A(alu__abc_41358_n1323_1), .B(alu__abc_41358_n1257), .Y(alu__abc_41358_n1324) );
  OR2X2 OR2X2_536 ( .A(_abc_43815_n1428_bF_buf3), .B(_abc_43815_n2183), .Y(_abc_43815_n2184) );
  OR2X2 OR2X2_5360 ( .A(alu__abc_41358_n1002), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n1326) );
  OR2X2 OR2X2_5361 ( .A(alu__abc_41358_n980), .B(alu__abc_41358_n299_bF_buf2), .Y(alu__abc_41358_n1327) );
  OR2X2 OR2X2_5362 ( .A(alu__abc_41358_n1325), .B(alu__abc_41358_n1329), .Y(alu__abc_41358_n1330) );
  OR2X2 OR2X2_5363 ( .A(alu__abc_41358_n1330), .B(alu__abc_41358_n279_bF_buf3), .Y(alu__abc_41358_n1331) );
  OR2X2 OR2X2_5364 ( .A(alu__abc_41358_n1333), .B(alu_b_i_3_bF_buf6), .Y(alu__abc_41358_n1334) );
  OR2X2 OR2X2_5365 ( .A(alu__abc_41358_n1334), .B(alu__abc_41358_n1332), .Y(alu__abc_41358_n1335) );
  OR2X2 OR2X2_5366 ( .A(alu__abc_41358_n1048), .B(alu_b_i_2_bF_buf1), .Y(alu__abc_41358_n1336) );
  OR2X2 OR2X2_5367 ( .A(alu__abc_41358_n992), .B(alu__abc_41358_n299_bF_buf0), .Y(alu__abc_41358_n1337) );
  OR2X2 OR2X2_5368 ( .A(alu__abc_41358_n1338), .B(alu__abc_41358_n294_bF_buf4), .Y(alu__abc_41358_n1339) );
  OR2X2 OR2X2_5369 ( .A(alu__abc_41358_n1340), .B(alu_b_i_4_bF_buf2), .Y(alu__abc_41358_n1341) );
  OR2X2 OR2X2_537 ( .A(_abc_43815_n2182), .B(_abc_43815_n2184), .Y(_abc_43815_n2185) );
  OR2X2 OR2X2_5370 ( .A(alu__abc_41358_n1322), .B(alu__abc_41358_n1343), .Y(alu__abc_41358_n1344_1) );
  OR2X2 OR2X2_5371 ( .A(alu__abc_41358_n1344_1), .B(alu__abc_41358_n1316), .Y(alu_p_o_5_) );
  OR2X2 OR2X2_5372 ( .A(alu__abc_41358_n425), .B(alu__abc_41358_n270), .Y(alu__abc_41358_n1346) );
  OR2X2 OR2X2_5373 ( .A(alu__abc_41358_n763), .B(alu__abc_41358_n733), .Y(alu__abc_41358_n1351) );
  OR2X2 OR2X2_5374 ( .A(alu__abc_41358_n1354), .B(alu__abc_41358_n1257), .Y(alu__abc_41358_n1355) );
  OR2X2 OR2X2_5375 ( .A(alu__abc_41358_n1355), .B(alu__abc_41358_n294_bF_buf3), .Y(alu__abc_41358_n1356) );
  OR2X2 OR2X2_5376 ( .A(alu__abc_41358_n1092), .B(alu__abc_41358_n299_bF_buf6), .Y(alu__abc_41358_n1357) );
  OR2X2 OR2X2_5377 ( .A(alu__abc_41358_n1102), .B(alu_b_i_2_bF_buf0), .Y(alu__abc_41358_n1358) );
  OR2X2 OR2X2_5378 ( .A(alu__abc_41358_n1359), .B(alu_b_i_3_bF_buf5), .Y(alu__abc_41358_n1360) );
  OR2X2 OR2X2_5379 ( .A(alu__abc_41358_n1361), .B(alu__abc_41358_n279_bF_buf2), .Y(alu__abc_41358_n1362_1) );
  OR2X2 OR2X2_538 ( .A(_abc_43815_n1431_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_43815_n2186) );
  OR2X2 OR2X2_5380 ( .A(alu__abc_41358_n1098), .B(alu__abc_41358_n299_bF_buf5), .Y(alu__abc_41358_n1363) );
  OR2X2 OR2X2_5381 ( .A(alu__abc_41358_n1124), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n1364) );
  OR2X2 OR2X2_5382 ( .A(alu__abc_41358_n1365), .B(alu__abc_41358_n294_bF_buf2), .Y(alu__abc_41358_n1366) );
  OR2X2 OR2X2_5383 ( .A(alu__abc_41358_n1114), .B(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n1367) );
  OR2X2 OR2X2_5384 ( .A(alu__abc_41358_n1120), .B(alu__abc_41358_n299_bF_buf4), .Y(alu__abc_41358_n1368) );
  OR2X2 OR2X2_5385 ( .A(alu__abc_41358_n1369), .B(alu_b_i_3_bF_buf4), .Y(alu__abc_41358_n1370) );
  OR2X2 OR2X2_5386 ( .A(alu__abc_41358_n1371), .B(alu_b_i_4_bF_buf1), .Y(alu__abc_41358_n1372) );
  OR2X2 OR2X2_5387 ( .A(alu__abc_41358_n1376), .B(alu_b_i_1_bF_buf0), .Y(alu__abc_41358_n1377) );
  OR2X2 OR2X2_5388 ( .A(alu__abc_41358_n1271), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n1378) );
  OR2X2 OR2X2_5389 ( .A(alu__abc_41358_n1379), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n1380) );
  OR2X2 OR2X2_539 ( .A(_abc_43815_n2188_1), .B(_abc_43815_n2189), .Y(_abc_43815_n2190) );
  OR2X2 OR2X2_5390 ( .A(alu__abc_41358_n1145), .B(alu__abc_41358_n299_bF_buf3), .Y(alu__abc_41358_n1381) );
  OR2X2 OR2X2_5391 ( .A(alu__abc_41358_n1390), .B(alu__abc_41358_n1386), .Y(alu__abc_41358_n1391) );
  OR2X2 OR2X2_5392 ( .A(alu__abc_41358_n1385), .B(alu__abc_41358_n1391), .Y(alu__abc_41358_n1392) );
  OR2X2 OR2X2_5393 ( .A(alu__abc_41358_n1384), .B(alu__abc_41358_n1392), .Y(alu__abc_41358_n1393) );
  OR2X2 OR2X2_5394 ( .A(alu__abc_41358_n1375), .B(alu__abc_41358_n1393), .Y(alu__abc_41358_n1394) );
  OR2X2 OR2X2_5395 ( .A(alu__abc_41358_n1394), .B(alu__abc_41358_n1374), .Y(alu__abc_41358_n1395) );
  OR2X2 OR2X2_5396 ( .A(alu__abc_41358_n1353), .B(alu__abc_41358_n1395), .Y(alu__abc_41358_n1396) );
  OR2X2 OR2X2_5397 ( .A(alu__abc_41358_n1396), .B(alu__abc_41358_n1349), .Y(alu_p_o_6_) );
  OR2X2 OR2X2_5398 ( .A(alu__abc_41358_n427), .B(alu__abc_41358_n275), .Y(alu__abc_41358_n1398) );
  OR2X2 OR2X2_5399 ( .A(alu__abc_41358_n1400), .B(alu__abc_41358_n588), .Y(alu__abc_41358_n1401_1) );
  OR2X2 OR2X2_54 ( .A(_abc_43815_n686_1_bF_buf3), .B(_abc_43815_n805), .Y(_abc_43815_n806) );
  OR2X2 OR2X2_540 ( .A(_abc_43815_n2190), .B(_abc_43815_n1350_bF_buf1), .Y(_abc_43815_n2191) );
  OR2X2 OR2X2_5400 ( .A(alu__abc_41358_n731), .B(alu__abc_41358_n764), .Y(alu__abc_41358_n1405) );
  OR2X2 OR2X2_5401 ( .A(alu__abc_41358_n1409), .B(alu__abc_41358_n1257), .Y(alu__abc_41358_n1410) );
  OR2X2 OR2X2_5402 ( .A(alu__abc_41358_n1410), .B(alu__abc_41358_n294_bF_buf0), .Y(alu__abc_41358_n1411) );
  OR2X2 OR2X2_5403 ( .A(alu__abc_41358_n1167), .B(alu__abc_41358_n299_bF_buf1), .Y(alu__abc_41358_n1412) );
  OR2X2 OR2X2_5404 ( .A(alu__abc_41358_n1177), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n1413) );
  OR2X2 OR2X2_5405 ( .A(alu__abc_41358_n1414), .B(alu_b_i_3_bF_buf3), .Y(alu__abc_41358_n1415) );
  OR2X2 OR2X2_5406 ( .A(alu__abc_41358_n1416), .B(alu__abc_41358_n279_bF_buf1), .Y(alu__abc_41358_n1417) );
  OR2X2 OR2X2_5407 ( .A(alu__abc_41358_n1173), .B(alu__abc_41358_n299_bF_buf0), .Y(alu__abc_41358_n1418) );
  OR2X2 OR2X2_5408 ( .A(alu__abc_41358_n1199), .B(alu_b_i_2_bF_buf2), .Y(alu__abc_41358_n1419_1) );
  OR2X2 OR2X2_5409 ( .A(alu__abc_41358_n1189), .B(alu_b_i_2_bF_buf1), .Y(alu__abc_41358_n1422) );
  OR2X2 OR2X2_541 ( .A(_abc_43815_n2193), .B(_abc_43815_n2192), .Y(_abc_43815_n2194) );
  OR2X2 OR2X2_5410 ( .A(alu__abc_41358_n1195), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n1423) );
  OR2X2 OR2X2_5411 ( .A(alu__abc_41358_n1425), .B(alu_b_i_4_bF_buf0), .Y(alu__abc_41358_n1426) );
  OR2X2 OR2X2_5412 ( .A(alu__abc_41358_n1426), .B(alu__abc_41358_n1421), .Y(alu__abc_41358_n1427) );
  OR2X2 OR2X2_5413 ( .A(alu__abc_41358_n1431), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n1432) );
  OR2X2 OR2X2_5414 ( .A(alu__abc_41358_n1302), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n1433) );
  OR2X2 OR2X2_5415 ( .A(alu__abc_41358_n1430), .B(alu__abc_41358_n1435_1), .Y(alu__abc_41358_n1436) );
  OR2X2 OR2X2_5416 ( .A(alu__abc_41358_n1444), .B(alu__abc_41358_n1440), .Y(alu__abc_41358_n1445) );
  OR2X2 OR2X2_5417 ( .A(alu__abc_41358_n1439), .B(alu__abc_41358_n1445), .Y(alu__abc_41358_n1446) );
  OR2X2 OR2X2_5418 ( .A(alu__abc_41358_n1438), .B(alu__abc_41358_n1446), .Y(alu__abc_41358_n1447) );
  OR2X2 OR2X2_5419 ( .A(alu__abc_41358_n1429), .B(alu__abc_41358_n1447), .Y(alu__abc_41358_n1448) );
  OR2X2 OR2X2_542 ( .A(_abc_43815_n1413_bF_buf4), .B(_abc_43815_n2194), .Y(_abc_43815_n2195) );
  OR2X2 OR2X2_5420 ( .A(alu__abc_41358_n1408), .B(alu__abc_41358_n1448), .Y(alu__abc_41358_n1449) );
  OR2X2 OR2X2_5421 ( .A(alu__abc_41358_n1407), .B(alu__abc_41358_n1449), .Y(alu__abc_41358_n1450) );
  OR2X2 OR2X2_5422 ( .A(alu__abc_41358_n1403), .B(alu__abc_41358_n1450), .Y(alu_p_o_7_) );
  OR2X2 OR2X2_5423 ( .A(alu__abc_41358_n429), .B(alu__abc_41358_n364), .Y(alu__abc_41358_n1454) );
  OR2X2 OR2X2_5424 ( .A(alu__abc_41358_n765), .B(alu__abc_41358_n718), .Y(alu__abc_41358_n1458) );
  OR2X2 OR2X2_5425 ( .A(alu__abc_41358_n875), .B(alu_b_i_3_bF_buf1), .Y(alu__abc_41358_n1462) );
  OR2X2 OR2X2_5426 ( .A(alu__abc_41358_n899), .B(alu__abc_41358_n294_bF_buf5), .Y(alu__abc_41358_n1463) );
  OR2X2 OR2X2_5427 ( .A(alu__abc_41358_n1464), .B(alu_b_i_4_bF_buf4), .Y(alu__abc_41358_n1465) );
  OR2X2 OR2X2_5428 ( .A(alu__abc_41358_n962), .B(alu__abc_41358_n294_bF_buf4), .Y(alu__abc_41358_n1466) );
  OR2X2 OR2X2_5429 ( .A(alu__abc_41358_n921), .B(alu_b_i_3_bF_buf0), .Y(alu__abc_41358_n1467) );
  OR2X2 OR2X2_543 ( .A(_abc_43815_n2197), .B(_abc_43815_n2164), .Y(_abc_43815_n2198) );
  OR2X2 OR2X2_5430 ( .A(alu__abc_41358_n1468), .B(alu__abc_41358_n279_bF_buf0), .Y(alu__abc_41358_n1469) );
  OR2X2 OR2X2_5431 ( .A(alu__abc_41358_n950), .B(alu__abc_41358_n294_bF_buf3), .Y(alu__abc_41358_n1472) );
  OR2X2 OR2X2_5432 ( .A(alu__abc_41358_n1473), .B(alu_b_i_1_bF_buf6), .Y(alu__abc_41358_n1474) );
  OR2X2 OR2X2_5433 ( .A(alu__abc_41358_n1376), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n1475) );
  OR2X2 OR2X2_5434 ( .A(alu__abc_41358_n1476), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n1477) );
  OR2X2 OR2X2_5435 ( .A(alu__abc_41358_n1274), .B(alu__abc_41358_n299_bF_buf5), .Y(alu__abc_41358_n1478) );
  OR2X2 OR2X2_5436 ( .A(alu__abc_41358_n1479), .B(alu_b_i_3_bF_buf6), .Y(alu__abc_41358_n1480) );
  OR2X2 OR2X2_5437 ( .A(alu__abc_41358_n1488), .B(alu__abc_41358_n1484), .Y(alu__abc_41358_n1489_1) );
  OR2X2 OR2X2_5438 ( .A(alu__abc_41358_n1483), .B(alu__abc_41358_n1489_1), .Y(alu__abc_41358_n1490_1) );
  OR2X2 OR2X2_5439 ( .A(alu__abc_41358_n1482), .B(alu__abc_41358_n1490_1), .Y(alu__abc_41358_n1491_1) );
  OR2X2 OR2X2_544 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_20_), .Y(_abc_43815_n2199) );
  OR2X2 OR2X2_5440 ( .A(alu__abc_41358_n1471), .B(alu__abc_41358_n1491_1), .Y(alu__abc_41358_n1492) );
  OR2X2 OR2X2_5441 ( .A(alu__abc_41358_n1492), .B(alu__abc_41358_n1461), .Y(alu__abc_41358_n1493) );
  OR2X2 OR2X2_5442 ( .A(alu__abc_41358_n1460), .B(alu__abc_41358_n1493), .Y(alu__abc_41358_n1494) );
  OR2X2 OR2X2_5443 ( .A(alu__abc_41358_n1456), .B(alu__abc_41358_n1494), .Y(alu_p_o_8_) );
  OR2X2 OR2X2_5444 ( .A(alu__abc_41358_n1497), .B(alu__abc_41358_n372), .Y(alu__abc_41358_n1498) );
  OR2X2 OR2X2_5445 ( .A(alu__abc_41358_n1496), .B(alu__abc_41358_n371), .Y(alu__abc_41358_n1499) );
  OR2X2 OR2X2_5446 ( .A(alu__abc_41358_n766), .B(alu__abc_41358_n787_1), .Y(alu__abc_41358_n1504) );
  OR2X2 OR2X2_5447 ( .A(alu__abc_41358_n1509), .B(alu__abc_41358_n1508), .Y(alu__abc_41358_n1510) );
  OR2X2 OR2X2_5448 ( .A(alu__abc_41358_n1510), .B(alu__abc_41358_n279_bF_buf5), .Y(alu__abc_41358_n1511) );
  OR2X2 OR2X2_5449 ( .A(alu__abc_41358_n1513), .B(alu_b_i_4_bF_buf3), .Y(alu__abc_41358_n1514) );
  OR2X2 OR2X2_545 ( .A(_abc_43815_n2160), .B(pc_q_21_), .Y(_abc_43815_n2202) );
  OR2X2 OR2X2_5450 ( .A(alu__abc_41358_n1514), .B(alu__abc_41358_n1512), .Y(alu__abc_41358_n1515) );
  OR2X2 OR2X2_5451 ( .A(alu__abc_41358_n1519), .B(alu_b_i_1_bF_buf5), .Y(alu__abc_41358_n1520) );
  OR2X2 OR2X2_5452 ( .A(alu__abc_41358_n1431), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n1521) );
  OR2X2 OR2X2_5453 ( .A(alu__abc_41358_n1522), .B(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n1523) );
  OR2X2 OR2X2_5454 ( .A(alu__abc_41358_n1305), .B(alu__abc_41358_n299_bF_buf4), .Y(alu__abc_41358_n1524) );
  OR2X2 OR2X2_5455 ( .A(alu__abc_41358_n1526), .B(alu__abc_41358_n1518), .Y(alu__abc_41358_n1527) );
  OR2X2 OR2X2_5456 ( .A(alu__abc_41358_n1533), .B(alu__abc_41358_n1534), .Y(alu__abc_41358_n1535) );
  OR2X2 OR2X2_5457 ( .A(alu__abc_41358_n1529), .B(alu__abc_41358_n1535), .Y(alu__abc_41358_n1536) );
  OR2X2 OR2X2_5458 ( .A(alu__abc_41358_n1528), .B(alu__abc_41358_n1536), .Y(alu__abc_41358_n1537) );
  OR2X2 OR2X2_5459 ( .A(alu__abc_41358_n1517), .B(alu__abc_41358_n1537), .Y(alu__abc_41358_n1538) );
  OR2X2 OR2X2_546 ( .A(_abc_43815_n2206), .B(_abc_43815_n1278_bF_buf4), .Y(_abc_43815_n2207) );
  OR2X2 OR2X2_5460 ( .A(alu__abc_41358_n1507), .B(alu__abc_41358_n1538), .Y(alu__abc_41358_n1539) );
  OR2X2 OR2X2_5461 ( .A(alu__abc_41358_n1506), .B(alu__abc_41358_n1539), .Y(alu__abc_41358_n1540) );
  OR2X2 OR2X2_5462 ( .A(alu__abc_41358_n1501), .B(alu__abc_41358_n1540), .Y(alu_p_o_9_) );
  OR2X2 OR2X2_5463 ( .A(alu__abc_41358_n1542), .B(alu__abc_41358_n438), .Y(alu__abc_41358_n1543) );
  OR2X2 OR2X2_5464 ( .A(alu__abc_41358_n1543), .B(alu__abc_41358_n347), .Y(alu__abc_41358_n1544) );
  OR2X2 OR2X2_5465 ( .A(alu__abc_41358_n1502), .B(alu__abc_41358_n781), .Y(alu__abc_41358_n1551) );
  OR2X2 OR2X2_5466 ( .A(alu__abc_41358_n1555), .B(alu__abc_41358_n1508), .Y(alu__abc_41358_n1556) );
  OR2X2 OR2X2_5467 ( .A(alu__abc_41358_n1556), .B(alu__abc_41358_n279_bF_buf4), .Y(alu__abc_41358_n1557) );
  OR2X2 OR2X2_5468 ( .A(alu__abc_41358_n1126), .B(alu_b_i_3_bF_buf2), .Y(alu__abc_41358_n1558) );
  OR2X2 OR2X2_5469 ( .A(alu__abc_41358_n1104), .B(alu__abc_41358_n294_bF_buf6), .Y(alu__abc_41358_n1559) );
  OR2X2 OR2X2_547 ( .A(_abc_43815_n1431_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_43815_n2208) );
  OR2X2 OR2X2_5470 ( .A(alu__abc_41358_n1560), .B(alu_b_i_4_bF_buf2), .Y(alu__abc_41358_n1561) );
  OR2X2 OR2X2_5471 ( .A(alu__abc_41358_n1565), .B(alu_b_i_1_bF_buf4), .Y(alu__abc_41358_n1566) );
  OR2X2 OR2X2_5472 ( .A(alu__abc_41358_n1473), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n1567) );
  OR2X2 OR2X2_5473 ( .A(alu__abc_41358_n1568), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n1569) );
  OR2X2 OR2X2_5474 ( .A(alu__abc_41358_n1379), .B(alu__abc_41358_n299_bF_buf3), .Y(alu__abc_41358_n1570) );
  OR2X2 OR2X2_5475 ( .A(alu__abc_41358_n1572), .B(alu__abc_41358_n1564), .Y(alu__abc_41358_n1573) );
  OR2X2 OR2X2_5476 ( .A(alu__abc_41358_n1579), .B(alu__abc_41358_n1580), .Y(alu__abc_41358_n1581) );
  OR2X2 OR2X2_5477 ( .A(alu__abc_41358_n1575), .B(alu__abc_41358_n1581), .Y(alu__abc_41358_n1582) );
  OR2X2 OR2X2_5478 ( .A(alu__abc_41358_n1574), .B(alu__abc_41358_n1582), .Y(alu__abc_41358_n1583) );
  OR2X2 OR2X2_5479 ( .A(alu__abc_41358_n1563), .B(alu__abc_41358_n1583), .Y(alu__abc_41358_n1584) );
  OR2X2 OR2X2_548 ( .A(pc_q_21_), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(_abc_43815_n2209) );
  OR2X2 OR2X2_5480 ( .A(alu__abc_41358_n1554), .B(alu__abc_41358_n1584), .Y(alu__abc_41358_n1585) );
  OR2X2 OR2X2_5481 ( .A(alu__abc_41358_n1553), .B(alu__abc_41358_n1585), .Y(alu__abc_41358_n1586) );
  OR2X2 OR2X2_5482 ( .A(alu__abc_41358_n1548), .B(alu__abc_41358_n1586), .Y(alu_p_o_10_) );
  OR2X2 OR2X2_5483 ( .A(alu__abc_41358_n1545), .B(alu__abc_41358_n441), .Y(alu__abc_41358_n1588) );
  OR2X2 OR2X2_5484 ( .A(alu__abc_41358_n1589), .B(alu__abc_41358_n354), .Y(alu__abc_41358_n1590) );
  OR2X2 OR2X2_5485 ( .A(alu__abc_41358_n1588), .B(alu__abc_41358_n355), .Y(alu__abc_41358_n1591) );
  OR2X2 OR2X2_5486 ( .A(alu__abc_41358_n1549), .B(alu__abc_41358_n805), .Y(alu__abc_41358_n1594) );
  OR2X2 OR2X2_5487 ( .A(alu__abc_41358_n1604), .B(alu__abc_41358_n1508), .Y(alu__abc_41358_n1605) );
  OR2X2 OR2X2_5488 ( .A(alu__abc_41358_n1605), .B(alu__abc_41358_n279_bF_buf3), .Y(alu__abc_41358_n1606) );
  OR2X2 OR2X2_5489 ( .A(alu__abc_41358_n1201), .B(alu_b_i_3_bF_buf0), .Y(alu__abc_41358_n1607) );
  OR2X2 OR2X2_549 ( .A(_abc_43815_n2212), .B(_abc_43815_n2175), .Y(_abc_43815_n2213) );
  OR2X2 OR2X2_5490 ( .A(alu__abc_41358_n1179), .B(alu__abc_41358_n294_bF_buf3), .Y(alu__abc_41358_n1608) );
  OR2X2 OR2X2_5491 ( .A(alu__abc_41358_n1609), .B(alu_b_i_4_bF_buf1), .Y(alu__abc_41358_n1610) );
  OR2X2 OR2X2_5492 ( .A(alu__abc_41358_n1614), .B(alu_b_i_1_bF_buf3), .Y(alu__abc_41358_n1615) );
  OR2X2 OR2X2_5493 ( .A(alu__abc_41358_n1519), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n1616) );
  OR2X2 OR2X2_5494 ( .A(alu__abc_41358_n1617), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n1618) );
  OR2X2 OR2X2_5495 ( .A(alu__abc_41358_n1434), .B(alu__abc_41358_n299_bF_buf2), .Y(alu__abc_41358_n1619) );
  OR2X2 OR2X2_5496 ( .A(alu__abc_41358_n1621), .B(alu__abc_41358_n1613), .Y(alu__abc_41358_n1622) );
  OR2X2 OR2X2_5497 ( .A(alu__abc_41358_n1624), .B(alu__abc_41358_n1625), .Y(alu__abc_41358_n1626) );
  OR2X2 OR2X2_5498 ( .A(alu__abc_41358_n1623), .B(alu__abc_41358_n1626), .Y(alu__abc_41358_n1627) );
  OR2X2 OR2X2_5499 ( .A(alu__abc_41358_n1612), .B(alu__abc_41358_n1627), .Y(alu__abc_41358_n1628) );
  OR2X2 OR2X2_55 ( .A(_abc_43815_n808), .B(_abc_43815_n794), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_) );
  OR2X2 OR2X2_550 ( .A(_abc_43815_n2179), .B(_abc_43815_n2213), .Y(_abc_43815_n2214) );
  OR2X2 OR2X2_5500 ( .A(alu__abc_41358_n1603), .B(alu__abc_41358_n1628), .Y(alu__abc_41358_n1629) );
  OR2X2 OR2X2_5501 ( .A(alu__abc_41358_n1629), .B(alu__abc_41358_n1602), .Y(alu__abc_41358_n1630) );
  OR2X2 OR2X2_5502 ( .A(alu__abc_41358_n1598), .B(alu__abc_41358_n1630), .Y(alu__abc_41358_n1631) );
  OR2X2 OR2X2_5503 ( .A(alu__abc_41358_n1593), .B(alu__abc_41358_n1631), .Y(alu_p_o_11_) );
  OR2X2 OR2X2_5504 ( .A(alu__abc_41358_n1633), .B(alu__abc_41358_n444), .Y(alu__abc_41358_n1634) );
  OR2X2 OR2X2_5505 ( .A(alu__abc_41358_n1634), .B(alu__abc_41358_n312), .Y(alu__abc_41358_n1635) );
  OR2X2 OR2X2_5506 ( .A(alu__abc_41358_n1595), .B(alu__abc_41358_n773), .Y(alu__abc_41358_n1642) );
  OR2X2 OR2X2_5507 ( .A(alu__abc_41358_n1249), .B(alu_b_i_3_bF_buf5), .Y(alu__abc_41358_n1646) );
  OR2X2 OR2X2_5508 ( .A(alu__abc_41358_n1255), .B(alu__abc_41358_n294_bF_buf1), .Y(alu__abc_41358_n1647) );
  OR2X2 OR2X2_5509 ( .A(alu__abc_41358_n1259), .B(alu_b_i_3_bF_buf4), .Y(alu__abc_41358_n1650) );
  OR2X2 OR2X2_551 ( .A(_abc_43815_n2216), .B(_abc_43815_n2217), .Y(_abc_43815_n2218) );
  OR2X2 OR2X2_5510 ( .A(alu__abc_41358_n1649), .B(alu__abc_41358_n1652), .Y(alu__abc_41358_n1653) );
  OR2X2 OR2X2_5511 ( .A(alu__abc_41358_n1276), .B(alu__abc_41358_n294_bF_buf0), .Y(alu__abc_41358_n1655) );
  OR2X2 OR2X2_5512 ( .A(alu__abc_41358_n1656), .B(alu_b_i_1_bF_buf2), .Y(alu__abc_41358_n1657) );
  OR2X2 OR2X2_5513 ( .A(alu__abc_41358_n1565), .B(alu__abc_41358_n252_bF_buf5), .Y(alu__abc_41358_n1658) );
  OR2X2 OR2X2_5514 ( .A(alu__abc_41358_n1659), .B(alu_b_i_2_bF_buf2), .Y(alu__abc_41358_n1660) );
  OR2X2 OR2X2_5515 ( .A(alu__abc_41358_n1476), .B(alu__abc_41358_n299_bF_buf1), .Y(alu__abc_41358_n1661) );
  OR2X2 OR2X2_5516 ( .A(alu__abc_41358_n1662), .B(alu_b_i_3_bF_buf3), .Y(alu__abc_41358_n1663) );
  OR2X2 OR2X2_5517 ( .A(alu__abc_41358_n1671), .B(alu__abc_41358_n1667), .Y(alu__abc_41358_n1672) );
  OR2X2 OR2X2_5518 ( .A(alu__abc_41358_n1666), .B(alu__abc_41358_n1672), .Y(alu__abc_41358_n1673) );
  OR2X2 OR2X2_5519 ( .A(alu__abc_41358_n1665), .B(alu__abc_41358_n1673), .Y(alu__abc_41358_n1674) );
  OR2X2 OR2X2_552 ( .A(_abc_43815_n1428_bF_buf2), .B(_abc_43815_n2222_1), .Y(_abc_43815_n2223) );
  OR2X2 OR2X2_5520 ( .A(alu__abc_41358_n1654), .B(alu__abc_41358_n1674), .Y(alu__abc_41358_n1675) );
  OR2X2 OR2X2_5521 ( .A(alu__abc_41358_n1645), .B(alu__abc_41358_n1675), .Y(alu__abc_41358_n1676) );
  OR2X2 OR2X2_5522 ( .A(alu__abc_41358_n1644), .B(alu__abc_41358_n1676), .Y(alu__abc_41358_n1677) );
  OR2X2 OR2X2_5523 ( .A(alu__abc_41358_n1639), .B(alu__abc_41358_n1677), .Y(alu_p_o_12_) );
  OR2X2 OR2X2_5524 ( .A(alu__abc_41358_n1679), .B(alu__abc_41358_n319), .Y(alu__abc_41358_n1680) );
  OR2X2 OR2X2_5525 ( .A(alu__abc_41358_n1681), .B(alu__abc_41358_n320), .Y(alu__abc_41358_n1682) );
  OR2X2 OR2X2_5526 ( .A(alu__abc_41358_n1640), .B(alu__abc_41358_n796), .Y(alu__abc_41358_n1687) );
  OR2X2 OR2X2_5527 ( .A(alu__abc_41358_n1338), .B(alu_b_i_3_bF_buf2), .Y(alu__abc_41358_n1691) );
  OR2X2 OR2X2_5528 ( .A(alu__abc_41358_n1328), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n1692) );
  OR2X2 OR2X2_5529 ( .A(alu__abc_41358_n1695), .B(alu__abc_41358_n1508), .Y(alu__abc_41358_n1696) );
  OR2X2 OR2X2_553 ( .A(_abc_43815_n2221), .B(_abc_43815_n2223), .Y(_abc_43815_n2224) );
  OR2X2 OR2X2_5530 ( .A(alu__abc_41358_n1697), .B(alu__abc_41358_n1694), .Y(alu__abc_41358_n1698) );
  OR2X2 OR2X2_5531 ( .A(alu__abc_41358_n1700), .B(alu_b_i_1_bF_buf1), .Y(alu__abc_41358_n1701) );
  OR2X2 OR2X2_5532 ( .A(alu__abc_41358_n1614), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n1702) );
  OR2X2 OR2X2_5533 ( .A(alu__abc_41358_n1703), .B(alu_b_i_2_bF_buf1), .Y(alu__abc_41358_n1704) );
  OR2X2 OR2X2_5534 ( .A(alu__abc_41358_n1522), .B(alu__abc_41358_n299_bF_buf0), .Y(alu__abc_41358_n1705) );
  OR2X2 OR2X2_5535 ( .A(alu__abc_41358_n1706), .B(alu_b_i_3_bF_buf1), .Y(alu__abc_41358_n1707) );
  OR2X2 OR2X2_5536 ( .A(alu__abc_41358_n1307), .B(alu__abc_41358_n294_bF_buf5), .Y(alu__abc_41358_n1708) );
  OR2X2 OR2X2_5537 ( .A(alu__abc_41358_n1716), .B(alu__abc_41358_n1712), .Y(alu__abc_41358_n1717) );
  OR2X2 OR2X2_5538 ( .A(alu__abc_41358_n1711), .B(alu__abc_41358_n1717), .Y(alu__abc_41358_n1718) );
  OR2X2 OR2X2_5539 ( .A(alu__abc_41358_n1710), .B(alu__abc_41358_n1718), .Y(alu__abc_41358_n1719) );
  OR2X2 OR2X2_554 ( .A(_abc_43815_n2225), .B(_abc_43815_n1473_bF_buf0), .Y(_abc_43815_n2226) );
  OR2X2 OR2X2_5540 ( .A(alu__abc_41358_n1699), .B(alu__abc_41358_n1719), .Y(alu__abc_41358_n1720) );
  OR2X2 OR2X2_5541 ( .A(alu__abc_41358_n1690), .B(alu__abc_41358_n1720), .Y(alu__abc_41358_n1721) );
  OR2X2 OR2X2_5542 ( .A(alu__abc_41358_n1689), .B(alu__abc_41358_n1721), .Y(alu__abc_41358_n1722) );
  OR2X2 OR2X2_5543 ( .A(alu__abc_41358_n1684), .B(alu__abc_41358_n1722), .Y(alu_p_o_13_) );
  OR2X2 OR2X2_5544 ( .A(alu__abc_41358_n1724), .B(alu__abc_41358_n453), .Y(alu__abc_41358_n1725) );
  OR2X2 OR2X2_5545 ( .A(alu__abc_41358_n1725), .B(alu__abc_41358_n329_1), .Y(alu__abc_41358_n1726) );
  OR2X2 OR2X2_5546 ( .A(alu__abc_41358_n1685), .B(alu__abc_41358_n799), .Y(alu__abc_41358_n1731) );
  OR2X2 OR2X2_5547 ( .A(alu__abc_41358_n1736), .B(alu__abc_41358_n1737), .Y(alu__abc_41358_n1738) );
  OR2X2 OR2X2_5548 ( .A(alu__abc_41358_n1365), .B(alu_b_i_3_bF_buf0), .Y(alu__abc_41358_n1740) );
  OR2X2 OR2X2_5549 ( .A(alu__abc_41358_n1359), .B(alu__abc_41358_n294_bF_buf4), .Y(alu__abc_41358_n1741) );
  OR2X2 OR2X2_555 ( .A(_abc_43815_n2205), .B(_abc_43815_n1472_1_bF_buf4), .Y(_abc_43815_n2227) );
  OR2X2 OR2X2_5550 ( .A(alu__abc_41358_n1744), .B(alu__abc_41358_n1508), .Y(alu__abc_41358_n1745) );
  OR2X2 OR2X2_5551 ( .A(alu__abc_41358_n1746), .B(alu__abc_41358_n1743), .Y(alu__abc_41358_n1747) );
  OR2X2 OR2X2_5552 ( .A(alu__abc_41358_n1749), .B(alu_b_i_1_bF_buf0), .Y(alu__abc_41358_n1750) );
  OR2X2 OR2X2_5553 ( .A(alu__abc_41358_n1656), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n1751) );
  OR2X2 OR2X2_5554 ( .A(alu__abc_41358_n1752), .B(alu_b_i_2_bF_buf0), .Y(alu__abc_41358_n1753) );
  OR2X2 OR2X2_5555 ( .A(alu__abc_41358_n1568), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n1754) );
  OR2X2 OR2X2_5556 ( .A(alu__abc_41358_n1755), .B(alu_b_i_3_bF_buf6), .Y(alu__abc_41358_n1756) );
  OR2X2 OR2X2_5557 ( .A(alu__abc_41358_n1382_1), .B(alu__abc_41358_n294_bF_buf2), .Y(alu__abc_41358_n1757) );
  OR2X2 OR2X2_5558 ( .A(alu__abc_41358_n1765), .B(alu__abc_41358_n1761), .Y(alu__abc_41358_n1766) );
  OR2X2 OR2X2_5559 ( .A(alu__abc_41358_n1760), .B(alu__abc_41358_n1766), .Y(alu__abc_41358_n1767) );
  OR2X2 OR2X2_556 ( .A(_abc_43815_n2228), .B(_abc_43815_n1350_bF_buf0), .Y(_abc_43815_n2229) );
  OR2X2 OR2X2_5560 ( .A(alu__abc_41358_n1759), .B(alu__abc_41358_n1767), .Y(alu__abc_41358_n1768) );
  OR2X2 OR2X2_5561 ( .A(alu__abc_41358_n1748), .B(alu__abc_41358_n1768), .Y(alu__abc_41358_n1769) );
  OR2X2 OR2X2_5562 ( .A(alu__abc_41358_n1739), .B(alu__abc_41358_n1769), .Y(alu__abc_41358_n1770) );
  OR2X2 OR2X2_5563 ( .A(alu__abc_41358_n1730), .B(alu__abc_41358_n1770), .Y(alu_p_o_14_) );
  OR2X2 OR2X2_5564 ( .A(alu__abc_41358_n1727), .B(alu__abc_41358_n456), .Y(alu__abc_41358_n1772) );
  OR2X2 OR2X2_5565 ( .A(alu__abc_41358_n1773), .B(alu__abc_41358_n336), .Y(alu__abc_41358_n1774) );
  OR2X2 OR2X2_5566 ( .A(alu__abc_41358_n1772), .B(alu__abc_41358_n337), .Y(alu__abc_41358_n1775) );
  OR2X2 OR2X2_5567 ( .A(alu__abc_41358_n1734), .B(alu__abc_41358_n704_1), .Y(alu__abc_41358_n1780) );
  OR2X2 OR2X2_5568 ( .A(alu__abc_41358_n1420), .B(alu_b_i_3_bF_buf5), .Y(alu__abc_41358_n1788) );
  OR2X2 OR2X2_5569 ( .A(alu__abc_41358_n1414), .B(alu__abc_41358_n294_bF_buf1), .Y(alu__abc_41358_n1789) );
  OR2X2 OR2X2_557 ( .A(_abc_43815_n2231), .B(_abc_43815_n2230), .Y(_abc_43815_n2232_1) );
  OR2X2 OR2X2_5570 ( .A(alu__abc_41358_n1792), .B(alu__abc_41358_n1508), .Y(alu__abc_41358_n1793) );
  OR2X2 OR2X2_5571 ( .A(alu__abc_41358_n1794), .B(alu__abc_41358_n1791), .Y(alu__abc_41358_n1795) );
  OR2X2 OR2X2_5572 ( .A(alu__abc_41358_n1798), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n1799) );
  OR2X2 OR2X2_5573 ( .A(alu__abc_41358_n1700), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n1800) );
  OR2X2 OR2X2_5574 ( .A(alu__abc_41358_n1801), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n1802) );
  OR2X2 OR2X2_5575 ( .A(alu__abc_41358_n1617), .B(alu__abc_41358_n299_bF_buf6), .Y(alu__abc_41358_n1803) );
  OR2X2 OR2X2_5576 ( .A(alu__abc_41358_n1797), .B(alu__abc_41358_n1805), .Y(alu__abc_41358_n1806) );
  OR2X2 OR2X2_5577 ( .A(alu__abc_41358_n1808), .B(alu__abc_41358_n1809), .Y(alu__abc_41358_n1810) );
  OR2X2 OR2X2_5578 ( .A(alu__abc_41358_n1807), .B(alu__abc_41358_n1810), .Y(alu__abc_41358_n1811) );
  OR2X2 OR2X2_5579 ( .A(alu__abc_41358_n1796), .B(alu__abc_41358_n1811), .Y(alu__abc_41358_n1812) );
  OR2X2 OR2X2_558 ( .A(_abc_43815_n1413_bF_buf3), .B(_abc_43815_n2232_1), .Y(_abc_43815_n2233) );
  OR2X2 OR2X2_5580 ( .A(alu__abc_41358_n1787), .B(alu__abc_41358_n1812), .Y(alu__abc_41358_n1813) );
  OR2X2 OR2X2_5581 ( .A(alu__abc_41358_n1813), .B(alu__abc_41358_n1786), .Y(alu__abc_41358_n1814) );
  OR2X2 OR2X2_5582 ( .A(alu__abc_41358_n1782), .B(alu__abc_41358_n1814), .Y(alu__abc_41358_n1815) );
  OR2X2 OR2X2_5583 ( .A(alu__abc_41358_n1777), .B(alu__abc_41358_n1815), .Y(alu_p_o_15_) );
  OR2X2 OR2X2_5584 ( .A(alu__abc_41358_n1778), .B(alu__abc_41358_n694), .Y(alu__abc_41358_n1817) );
  OR2X2 OR2X2_5585 ( .A(alu__abc_41358_n461), .B(alu__abc_41358_n237), .Y(alu__abc_41358_n1822) );
  OR2X2 OR2X2_5586 ( .A(alu__abc_41358_n923), .B(alu_b_i_4_bF_buf1), .Y(alu__abc_41358_n1828) );
  OR2X2 OR2X2_5587 ( .A(alu__abc_41358_n961), .B(alu__abc_41358_n279_bF_buf4), .Y(alu__abc_41358_n1829) );
  OR2X2 OR2X2_5588 ( .A(alu__abc_41358_n1659), .B(alu__abc_41358_n299_bF_buf5), .Y(alu__abc_41358_n1833) );
  OR2X2 OR2X2_5589 ( .A(alu__abc_41358_n1749), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n1834) );
  OR2X2 OR2X2_559 ( .A(_abc_43815_n2235), .B(_abc_43815_n2207), .Y(_abc_43815_n2236) );
  OR2X2 OR2X2_5590 ( .A(alu__abc_41358_n1835), .B(alu_b_i_1_bF_buf6), .Y(alu__abc_41358_n1836) );
  OR2X2 OR2X2_5591 ( .A(alu__abc_41358_n1837), .B(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n1838) );
  OR2X2 OR2X2_5592 ( .A(alu__abc_41358_n1832), .B(alu__abc_41358_n1840), .Y(alu__abc_41358_n1841) );
  OR2X2 OR2X2_5593 ( .A(alu__abc_41358_n1848), .B(alu__abc_41358_n1844), .Y(alu__abc_41358_n1849) );
  OR2X2 OR2X2_5594 ( .A(alu__abc_41358_n1849), .B(alu__abc_41358_n1851), .Y(alu__abc_41358_n1852) );
  OR2X2 OR2X2_5595 ( .A(alu__abc_41358_n1852), .B(alu__abc_41358_n1843), .Y(alu__abc_41358_n1853) );
  OR2X2 OR2X2_5596 ( .A(alu__abc_41358_n1842), .B(alu__abc_41358_n1853), .Y(alu__abc_41358_n1854) );
  OR2X2 OR2X2_5597 ( .A(alu__abc_41358_n1854), .B(alu__abc_41358_n1831), .Y(alu__abc_41358_n1855) );
  OR2X2 OR2X2_5598 ( .A(alu__abc_41358_n1827), .B(alu__abc_41358_n1855), .Y(alu__abc_41358_n1856) );
  OR2X2 OR2X2_5599 ( .A(alu__abc_41358_n1826), .B(alu__abc_41358_n1856), .Y(alu__abc_41358_n1857) );
  OR2X2 OR2X2_56 ( .A(_abc_43815_n810), .B(_abc_43815_n811), .Y(_abc_43815_n812) );
  OR2X2 OR2X2_560 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_21_), .Y(_abc_43815_n2237) );
  OR2X2 OR2X2_5600 ( .A(alu__abc_41358_n1857), .B(alu__abc_41358_n1821), .Y(alu_p_o_16_) );
  OR2X2 OR2X2_5601 ( .A(alu__abc_41358_n1860), .B(alu__abc_41358_n245), .Y(alu__abc_41358_n1861) );
  OR2X2 OR2X2_5602 ( .A(alu__abc_41358_n1859), .B(alu__abc_41358_n244), .Y(alu__abc_41358_n1862) );
  OR2X2 OR2X2_5603 ( .A(alu__abc_41358_n1818), .B(alu__abc_41358_n692), .Y(alu__abc_41358_n1865) );
  OR2X2 OR2X2_5604 ( .A(alu__abc_41358_n1870), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n1872) );
  OR2X2 OR2X2_5605 ( .A(alu__abc_41358_n1874), .B(alu_b_i_1_bF_buf5), .Y(alu__abc_41358_n1875) );
  OR2X2 OR2X2_5606 ( .A(alu__abc_41358_n1798), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n1876) );
  OR2X2 OR2X2_5607 ( .A(alu__abc_41358_n1877), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n1878) );
  OR2X2 OR2X2_5608 ( .A(alu__abc_41358_n1703), .B(alu__abc_41358_n299_bF_buf4), .Y(alu__abc_41358_n1879) );
  OR2X2 OR2X2_5609 ( .A(alu__abc_41358_n1882), .B(alu_b_i_4_bF_buf3), .Y(alu__abc_41358_n1883) );
  OR2X2 OR2X2_561 ( .A(_abc_43815_n2203_1), .B(pc_q_22_), .Y(_abc_43815_n2240) );
  OR2X2 OR2X2_5610 ( .A(alu__abc_41358_n1883), .B(alu__abc_41358_n1881), .Y(alu__abc_41358_n1884) );
  OR2X2 OR2X2_5611 ( .A(alu__abc_41358_n1077), .B(alu__abc_41358_n279_bF_buf2), .Y(alu__abc_41358_n1885) );
  OR2X2 OR2X2_5612 ( .A(alu__abc_41358_n1893), .B(alu__abc_41358_n1889), .Y(alu__abc_41358_n1894) );
  OR2X2 OR2X2_5613 ( .A(alu__abc_41358_n1888), .B(alu__abc_41358_n1894), .Y(alu__abc_41358_n1895) );
  OR2X2 OR2X2_5614 ( .A(alu__abc_41358_n1887), .B(alu__abc_41358_n1895), .Y(alu__abc_41358_n1896) );
  OR2X2 OR2X2_5615 ( .A(alu__abc_41358_n1873), .B(alu__abc_41358_n1896), .Y(alu__abc_41358_n1897) );
  OR2X2 OR2X2_5616 ( .A(alu__abc_41358_n1869), .B(alu__abc_41358_n1897), .Y(alu__abc_41358_n1898) );
  OR2X2 OR2X2_5617 ( .A(alu__abc_41358_n1868), .B(alu__abc_41358_n1898), .Y(alu__abc_41358_n1899) );
  OR2X2 OR2X2_5618 ( .A(alu__abc_41358_n1899), .B(alu__abc_41358_n1864), .Y(alu_p_o_17_) );
  OR2X2 OR2X2_5619 ( .A(alu__abc_41358_n811), .B(alu__abc_41358_n685), .Y(alu__abc_41358_n1904) );
  OR2X2 OR2X2_562 ( .A(_abc_43815_n2244), .B(_abc_43815_n1278_bF_buf3), .Y(_abc_43815_n2245) );
  OR2X2 OR2X2_5620 ( .A(alu__abc_41358_n1907), .B(alu__abc_41358_n470), .Y(alu__abc_41358_n1908) );
  OR2X2 OR2X2_5621 ( .A(alu__abc_41358_n1908), .B(alu__abc_41358_n220), .Y(alu__abc_41358_n1909) );
  OR2X2 OR2X2_5622 ( .A(alu__abc_41358_n1915), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n1916) );
  OR2X2 OR2X2_5623 ( .A(alu__abc_41358_n1918), .B(alu_b_i_1_bF_buf4), .Y(alu__abc_41358_n1919) );
  OR2X2 OR2X2_5624 ( .A(alu__abc_41358_n1835), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n1920) );
  OR2X2 OR2X2_5625 ( .A(alu__abc_41358_n1921), .B(alu_b_i_2_bF_buf3), .Y(alu__abc_41358_n1922) );
  OR2X2 OR2X2_5626 ( .A(alu__abc_41358_n1752), .B(alu__abc_41358_n299_bF_buf3), .Y(alu__abc_41358_n1923) );
  OR2X2 OR2X2_5627 ( .A(alu__abc_41358_n1926), .B(alu_b_i_4_bF_buf2), .Y(alu__abc_41358_n1927) );
  OR2X2 OR2X2_5628 ( .A(alu__abc_41358_n1927), .B(alu__abc_41358_n1925), .Y(alu__abc_41358_n1928) );
  OR2X2 OR2X2_5629 ( .A(alu__abc_41358_n1147), .B(alu__abc_41358_n279_bF_buf0), .Y(alu__abc_41358_n1929) );
  OR2X2 OR2X2_563 ( .A(_abc_43815_n2243), .B(_abc_43815_n1472_1_bF_buf3), .Y(_abc_43815_n2246) );
  OR2X2 OR2X2_5630 ( .A(alu__abc_41358_n1937), .B(alu__abc_41358_n1933), .Y(alu__abc_41358_n1938) );
  OR2X2 OR2X2_5631 ( .A(alu__abc_41358_n1932), .B(alu__abc_41358_n1938), .Y(alu__abc_41358_n1939) );
  OR2X2 OR2X2_5632 ( .A(alu__abc_41358_n1931), .B(alu__abc_41358_n1939), .Y(alu__abc_41358_n1940) );
  OR2X2 OR2X2_5633 ( .A(alu__abc_41358_n1917), .B(alu__abc_41358_n1940), .Y(alu__abc_41358_n1941) );
  OR2X2 OR2X2_5634 ( .A(alu__abc_41358_n1914), .B(alu__abc_41358_n1941), .Y(alu__abc_41358_n1942) );
  OR2X2 OR2X2_5635 ( .A(alu__abc_41358_n1913), .B(alu__abc_41358_n1942), .Y(alu__abc_41358_n1943) );
  OR2X2 OR2X2_5636 ( .A(alu__abc_41358_n1943), .B(alu__abc_41358_n1906), .Y(alu_p_o_18_) );
  OR2X2 OR2X2_5637 ( .A(alu__abc_41358_n1910), .B(alu__abc_41358_n473), .Y(alu__abc_41358_n1945) );
  OR2X2 OR2X2_5638 ( .A(alu__abc_41358_n1945), .B(alu__abc_41358_n228), .Y(alu__abc_41358_n1946) );
  OR2X2 OR2X2_5639 ( .A(alu__abc_41358_n1947), .B(alu__abc_41358_n227), .Y(alu__abc_41358_n1948) );
  OR2X2 OR2X2_564 ( .A(pc_q_22_), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(_abc_43815_n2249) );
  OR2X2 OR2X2_5640 ( .A(alu__abc_41358_n1902), .B(alu__abc_41358_n683), .Y(alu__abc_41358_n1951) );
  OR2X2 OR2X2_5641 ( .A(alu__abc_41358_n1957), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n1958) );
  OR2X2 OR2X2_5642 ( .A(alu__abc_41358_n1960), .B(alu_b_i_1_bF_buf3), .Y(alu__abc_41358_n1961) );
  OR2X2 OR2X2_5643 ( .A(alu__abc_41358_n1874), .B(alu__abc_41358_n252_bF_buf5), .Y(alu__abc_41358_n1962) );
  OR2X2 OR2X2_5644 ( .A(alu__abc_41358_n1963), .B(alu_b_i_2_bF_buf2), .Y(alu__abc_41358_n1964) );
  OR2X2 OR2X2_5645 ( .A(alu__abc_41358_n1801), .B(alu__abc_41358_n299_bF_buf2), .Y(alu__abc_41358_n1965) );
  OR2X2 OR2X2_5646 ( .A(alu__abc_41358_n1968), .B(alu_b_i_4_bF_buf1), .Y(alu__abc_41358_n1969) );
  OR2X2 OR2X2_5647 ( .A(alu__abc_41358_n1969), .B(alu__abc_41358_n1967), .Y(alu__abc_41358_n1970) );
  OR2X2 OR2X2_5648 ( .A(alu__abc_41358_n1224), .B(alu__abc_41358_n279_bF_buf4), .Y(alu__abc_41358_n1971) );
  OR2X2 OR2X2_5649 ( .A(alu__abc_41358_n1979), .B(alu__abc_41358_n1975), .Y(alu__abc_41358_n1980) );
  OR2X2 OR2X2_565 ( .A(_abc_43815_n2248), .B(_abc_43815_n2252_1), .Y(_abc_43815_n2255) );
  OR2X2 OR2X2_5650 ( .A(alu__abc_41358_n1974), .B(alu__abc_41358_n1980), .Y(alu__abc_41358_n1981) );
  OR2X2 OR2X2_5651 ( .A(alu__abc_41358_n1973), .B(alu__abc_41358_n1981), .Y(alu__abc_41358_n1982) );
  OR2X2 OR2X2_5652 ( .A(alu__abc_41358_n1959), .B(alu__abc_41358_n1982), .Y(alu__abc_41358_n1983) );
  OR2X2 OR2X2_5653 ( .A(alu__abc_41358_n1956), .B(alu__abc_41358_n1983), .Y(alu__abc_41358_n1984) );
  OR2X2 OR2X2_5654 ( .A(alu__abc_41358_n1955), .B(alu__abc_41358_n1984), .Y(alu__abc_41358_n1985) );
  OR2X2 OR2X2_5655 ( .A(alu__abc_41358_n1950), .B(alu__abc_41358_n1985), .Y(alu_p_o_19_) );
  OR2X2 OR2X2_5656 ( .A(alu__abc_41358_n1952), .B(alu__abc_41358_n676), .Y(alu__abc_41358_n1987) );
  OR2X2 OR2X2_5657 ( .A(alu__abc_41358_n1992), .B(alu__abc_41358_n476), .Y(alu__abc_41358_n1993) );
  OR2X2 OR2X2_5658 ( .A(alu__abc_41358_n1993), .B(alu__abc_41358_n202), .Y(alu__abc_41358_n1996) );
  OR2X2 OR2X2_5659 ( .A(alu__abc_41358_n1261), .B(alu_b_i_4_bF_buf0), .Y(alu__abc_41358_n2000) );
  OR2X2 OR2X2_566 ( .A(_abc_43815_n1428_bF_buf1), .B(_abc_43815_n2258), .Y(_abc_43815_n2259) );
  OR2X2 OR2X2_5660 ( .A(alu__abc_41358_n1837), .B(alu__abc_41358_n299_bF_buf1), .Y(alu__abc_41358_n2003) );
  OR2X2 OR2X2_5661 ( .A(alu__abc_41358_n1918), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n2004) );
  OR2X2 OR2X2_5662 ( .A(alu__abc_41358_n2005), .B(alu_b_i_1_bF_buf2), .Y(alu__abc_41358_n2006) );
  OR2X2 OR2X2_5663 ( .A(alu__abc_41358_n2007), .B(alu_b_i_2_bF_buf1), .Y(alu__abc_41358_n2008) );
  OR2X2 OR2X2_5664 ( .A(alu__abc_41358_n2002), .B(alu__abc_41358_n2010), .Y(alu__abc_41358_n2011) );
  OR2X2 OR2X2_5665 ( .A(alu__abc_41358_n2018), .B(alu__abc_41358_n2019), .Y(alu__abc_41358_n2020) );
  OR2X2 OR2X2_5666 ( .A(alu__abc_41358_n2014), .B(alu__abc_41358_n2020), .Y(alu__abc_41358_n2021) );
  OR2X2 OR2X2_5667 ( .A(alu__abc_41358_n2013), .B(alu__abc_41358_n2021), .Y(alu__abc_41358_n2022) );
  OR2X2 OR2X2_5668 ( .A(alu__abc_41358_n2012), .B(alu__abc_41358_n2022), .Y(alu__abc_41358_n2023) );
  OR2X2 OR2X2_5669 ( .A(alu__abc_41358_n2023), .B(alu__abc_41358_n2001), .Y(alu__abc_41358_n2024) );
  OR2X2 OR2X2_567 ( .A(_abc_43815_n2257), .B(_abc_43815_n2259), .Y(_abc_43815_n2260) );
  OR2X2 OR2X2_5670 ( .A(alu__abc_41358_n1999), .B(alu__abc_41358_n2024), .Y(alu__abc_41358_n2025) );
  OR2X2 OR2X2_5671 ( .A(alu__abc_41358_n1998), .B(alu__abc_41358_n2025), .Y(alu__abc_41358_n2026) );
  OR2X2 OR2X2_5672 ( .A(alu__abc_41358_n2026), .B(alu__abc_41358_n1991), .Y(alu_p_o_20_) );
  OR2X2 OR2X2_5673 ( .A(alu__abc_41358_n1988), .B(alu__abc_41358_n820), .Y(alu__abc_41358_n2028) );
  OR2X2 OR2X2_5674 ( .A(alu__abc_41358_n2034), .B(alu__abc_41358_n210), .Y(alu__abc_41358_n2035) );
  OR2X2 OR2X2_5675 ( .A(alu__abc_41358_n2033), .B(alu__abc_41358_n209), .Y(alu__abc_41358_n2036) );
  OR2X2 OR2X2_5676 ( .A(alu__abc_41358_n2040), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2041) );
  OR2X2 OR2X2_5677 ( .A(alu__abc_41358_n1308), .B(alu__abc_41358_n279_bF_buf2), .Y(alu__abc_41358_n2043) );
  OR2X2 OR2X2_5678 ( .A(alu__abc_41358_n1706), .B(alu__abc_41358_n294_bF_buf1), .Y(alu__abc_41358_n2044) );
  OR2X2 OR2X2_5679 ( .A(alu__abc_41358_n2045), .B(alu_b_i_1_bF_buf1), .Y(alu__abc_41358_n2046) );
  OR2X2 OR2X2_568 ( .A(_abc_43815_n1431_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_43815_n2261) );
  OR2X2 OR2X2_5680 ( .A(alu__abc_41358_n1960), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n2047) );
  OR2X2 OR2X2_5681 ( .A(alu__abc_41358_n2048), .B(alu_b_i_2_bF_buf0), .Y(alu__abc_41358_n2049) );
  OR2X2 OR2X2_5682 ( .A(alu__abc_41358_n1877), .B(alu__abc_41358_n299_bF_buf0), .Y(alu__abc_41358_n2050) );
  OR2X2 OR2X2_5683 ( .A(alu_b_i_4_bF_buf4), .B(alu_b_i_3_bF_buf5), .Y(alu__abc_41358_n2052) );
  OR2X2 OR2X2_5684 ( .A(alu__abc_41358_n2051), .B(alu__abc_41358_n2052), .Y(alu__abc_41358_n2053) );
  OR2X2 OR2X2_5685 ( .A(alu__abc_41358_n2061), .B(alu__abc_41358_n2062), .Y(alu__abc_41358_n2063) );
  OR2X2 OR2X2_5686 ( .A(alu__abc_41358_n2057), .B(alu__abc_41358_n2063), .Y(alu__abc_41358_n2064) );
  OR2X2 OR2X2_5687 ( .A(alu__abc_41358_n2056), .B(alu__abc_41358_n2064), .Y(alu__abc_41358_n2065) );
  OR2X2 OR2X2_5688 ( .A(alu__abc_41358_n2042), .B(alu__abc_41358_n2065), .Y(alu__abc_41358_n2066) );
  OR2X2 OR2X2_5689 ( .A(alu__abc_41358_n2039), .B(alu__abc_41358_n2066), .Y(alu__abc_41358_n2067) );
  OR2X2 OR2X2_569 ( .A(_abc_43815_n2262_1), .B(_abc_43815_n1473_bF_buf4), .Y(_abc_43815_n2263) );
  OR2X2 OR2X2_5690 ( .A(alu__abc_41358_n2038), .B(alu__abc_41358_n2067), .Y(alu__abc_41358_n2068) );
  OR2X2 OR2X2_5691 ( .A(alu__abc_41358_n2068), .B(alu__abc_41358_n2032), .Y(alu_p_o_21_) );
  OR2X2 OR2X2_5692 ( .A(alu__abc_41358_n2029), .B(alu__abc_41358_n672), .Y(alu__abc_41358_n2070) );
  OR2X2 OR2X2_5693 ( .A(alu__abc_41358_n2075), .B(alu__abc_41358_n485), .Y(alu__abc_41358_n2076) );
  OR2X2 OR2X2_5694 ( .A(alu__abc_41358_n2076), .B(alu__abc_41358_n185), .Y(alu__abc_41358_n2077) );
  OR2X2 OR2X2_5695 ( .A(alu__abc_41358_n2082), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2083) );
  OR2X2 OR2X2_5696 ( .A(alu__abc_41358_n2085), .B(alu_b_i_1_bF_buf0), .Y(alu__abc_41358_n2086) );
  OR2X2 OR2X2_5697 ( .A(alu__abc_41358_n2005), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n2087) );
  OR2X2 OR2X2_5698 ( .A(alu__abc_41358_n2088), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n2089) );
  OR2X2 OR2X2_5699 ( .A(alu__abc_41358_n1921), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n2090) );
  OR2X2 OR2X2_57 ( .A(_abc_43815_n813), .B(_abc_43815_n814), .Y(_abc_43815_n815) );
  OR2X2 OR2X2_570 ( .A(_abc_43815_n2264), .B(_abc_43815_n1350_bF_buf4), .Y(_abc_43815_n2265) );
  OR2X2 OR2X2_5700 ( .A(alu__abc_41358_n2093), .B(alu_b_i_4_bF_buf3), .Y(alu__abc_41358_n2094) );
  OR2X2 OR2X2_5701 ( .A(alu__abc_41358_n2094), .B(alu__abc_41358_n2092), .Y(alu__abc_41358_n2095) );
  OR2X2 OR2X2_5702 ( .A(alu__abc_41358_n1383), .B(alu__abc_41358_n279_bF_buf0), .Y(alu__abc_41358_n2096) );
  OR2X2 OR2X2_5703 ( .A(alu__abc_41358_n2104), .B(alu__abc_41358_n2100), .Y(alu__abc_41358_n2105) );
  OR2X2 OR2X2_5704 ( .A(alu__abc_41358_n2099), .B(alu__abc_41358_n2105), .Y(alu__abc_41358_n2106) );
  OR2X2 OR2X2_5705 ( .A(alu__abc_41358_n2098), .B(alu__abc_41358_n2106), .Y(alu__abc_41358_n2107) );
  OR2X2 OR2X2_5706 ( .A(alu__abc_41358_n2084), .B(alu__abc_41358_n2107), .Y(alu__abc_41358_n2108) );
  OR2X2 OR2X2_5707 ( .A(alu__abc_41358_n2109), .B(alu__abc_41358_n2108), .Y(alu__abc_41358_n2110) );
  OR2X2 OR2X2_5708 ( .A(alu__abc_41358_n2081), .B(alu__abc_41358_n2110), .Y(alu__abc_41358_n2111) );
  OR2X2 OR2X2_5709 ( .A(alu__abc_41358_n2111), .B(alu__abc_41358_n2074), .Y(alu_p_o_22_) );
  OR2X2 OR2X2_571 ( .A(_abc_43815_n2267), .B(_abc_43815_n2266), .Y(_abc_43815_n2268) );
  OR2X2 OR2X2_5710 ( .A(alu__abc_41358_n2071), .B(alu__abc_41358_n649), .Y(alu__abc_41358_n2113) );
  OR2X2 OR2X2_5711 ( .A(alu__abc_41358_n2078), .B(alu__abc_41358_n488), .Y(alu__abc_41358_n2118) );
  OR2X2 OR2X2_5712 ( .A(alu__abc_41358_n2119), .B(alu__abc_41358_n192_1), .Y(alu__abc_41358_n2120) );
  OR2X2 OR2X2_5713 ( .A(alu__abc_41358_n2118), .B(alu__abc_41358_n193), .Y(alu__abc_41358_n2121) );
  OR2X2 OR2X2_5714 ( .A(alu__abc_41358_n2124), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2125) );
  OR2X2 OR2X2_5715 ( .A(alu__abc_41358_n2127), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n2128) );
  OR2X2 OR2X2_5716 ( .A(alu__abc_41358_n2045), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n2129) );
  OR2X2 OR2X2_5717 ( .A(alu__abc_41358_n2130), .B(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n2131) );
  OR2X2 OR2X2_5718 ( .A(alu__abc_41358_n1963), .B(alu__abc_41358_n299_bF_buf6), .Y(alu__abc_41358_n2132) );
  OR2X2 OR2X2_5719 ( .A(alu__abc_41358_n2135), .B(alu_b_i_4_bF_buf2), .Y(alu__abc_41358_n2136) );
  OR2X2 OR2X2_572 ( .A(_abc_43815_n1413_bF_buf2), .B(_abc_43815_n2268), .Y(_abc_43815_n2269) );
  OR2X2 OR2X2_5720 ( .A(alu__abc_41358_n2136), .B(alu__abc_41358_n2134), .Y(alu__abc_41358_n2137) );
  OR2X2 OR2X2_5721 ( .A(alu__abc_41358_n1437), .B(alu__abc_41358_n279_bF_buf4), .Y(alu__abc_41358_n2138) );
  OR2X2 OR2X2_5722 ( .A(alu__abc_41358_n2145), .B(alu__abc_41358_n2146), .Y(alu__abc_41358_n2147) );
  OR2X2 OR2X2_5723 ( .A(alu__abc_41358_n2141), .B(alu__abc_41358_n2147), .Y(alu__abc_41358_n2148) );
  OR2X2 OR2X2_5724 ( .A(alu__abc_41358_n2140), .B(alu__abc_41358_n2148), .Y(alu__abc_41358_n2149) );
  OR2X2 OR2X2_5725 ( .A(alu__abc_41358_n2149), .B(alu__abc_41358_n2126), .Y(alu__abc_41358_n2150) );
  OR2X2 OR2X2_5726 ( .A(alu__abc_41358_n2151), .B(alu__abc_41358_n2150), .Y(alu__abc_41358_n2152) );
  OR2X2 OR2X2_5727 ( .A(alu__abc_41358_n2123), .B(alu__abc_41358_n2152), .Y(alu__abc_41358_n2153) );
  OR2X2 OR2X2_5728 ( .A(alu__abc_41358_n2153), .B(alu__abc_41358_n2117), .Y(alu_p_o_23_) );
  OR2X2 OR2X2_5729 ( .A(alu__abc_41358_n2114), .B(alu__abc_41358_n667), .Y(alu__abc_41358_n2157) );
  OR2X2 OR2X2_573 ( .A(_abc_43815_n2271), .B(_abc_43815_n2245), .Y(_abc_43815_n2272_1) );
  OR2X2 OR2X2_5730 ( .A(alu__abc_41358_n493), .B(alu__abc_41358_n125_1), .Y(alu__abc_41358_n2160) );
  OR2X2 OR2X2_5731 ( .A(alu__abc_41358_n1468), .B(alu_b_i_4_bF_buf1), .Y(alu__abc_41358_n2166) );
  OR2X2 OR2X2_5732 ( .A(alu__abc_41358_n1839), .B(alu__abc_41358_n294_bF_buf6), .Y(alu__abc_41358_n2169) );
  OR2X2 OR2X2_5733 ( .A(alu__abc_41358_n2085), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n2170) );
  OR2X2 OR2X2_5734 ( .A(alu__abc_41358_n2171), .B(alu_b_i_1_bF_buf6), .Y(alu__abc_41358_n2172) );
  OR2X2 OR2X2_5735 ( .A(alu__abc_41358_n2173), .B(alu_b_i_2_bF_buf4), .Y(alu__abc_41358_n2174) );
  OR2X2 OR2X2_5736 ( .A(alu__abc_41358_n2007), .B(alu__abc_41358_n299_bF_buf5), .Y(alu__abc_41358_n2175) );
  OR2X2 OR2X2_5737 ( .A(alu__abc_41358_n2176), .B(alu_b_i_3_bF_buf2), .Y(alu__abc_41358_n2177) );
  OR2X2 OR2X2_5738 ( .A(alu__abc_41358_n2184), .B(alu__abc_41358_n2185), .Y(alu__abc_41358_n2186) );
  OR2X2 OR2X2_5739 ( .A(alu__abc_41358_n2186), .B(alu__abc_41358_n2183), .Y(alu__abc_41358_n2187) );
  OR2X2 OR2X2_574 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_22_), .Y(_abc_43815_n2273) );
  OR2X2 OR2X2_5740 ( .A(alu__abc_41358_n2179), .B(alu__abc_41358_n2187), .Y(alu__abc_41358_n2188) );
  OR2X2 OR2X2_5741 ( .A(alu__abc_41358_n2188), .B(alu__abc_41358_n2168), .Y(alu__abc_41358_n2189) );
  OR2X2 OR2X2_5742 ( .A(alu__abc_41358_n2189), .B(alu__abc_41358_n2167), .Y(alu__abc_41358_n2190) );
  OR2X2 OR2X2_5743 ( .A(alu__abc_41358_n2165), .B(alu__abc_41358_n2190), .Y(alu__abc_41358_n2191) );
  OR2X2 OR2X2_5744 ( .A(alu__abc_41358_n2164), .B(alu__abc_41358_n2191), .Y(alu__abc_41358_n2192) );
  OR2X2 OR2X2_5745 ( .A(alu__abc_41358_n2159), .B(alu__abc_41358_n2192), .Y(alu_p_o_24_) );
  OR2X2 OR2X2_5746 ( .A(alu__abc_41358_n2155), .B(alu__abc_41358_n665), .Y(alu__abc_41358_n2194) );
  OR2X2 OR2X2_5747 ( .A(alu__abc_41358_n2200), .B(alu__abc_41358_n117), .Y(alu__abc_41358_n2201) );
  OR2X2 OR2X2_5748 ( .A(alu__abc_41358_n2199), .B(alu__abc_41358_n116), .Y(alu__abc_41358_n2202) );
  OR2X2 OR2X2_5749 ( .A(alu__abc_41358_n2206), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2207) );
  OR2X2 OR2X2_575 ( .A(_abc_43815_n2241), .B(pc_q_23_), .Y(_abc_43815_n2276) );
  OR2X2 OR2X2_5750 ( .A(alu__abc_41358_n2210), .B(alu_b_i_1_bF_buf5), .Y(alu__abc_41358_n2211) );
  OR2X2 OR2X2_5751 ( .A(alu__abc_41358_n2127), .B(alu__abc_41358_n252_bF_buf6), .Y(alu__abc_41358_n2212) );
  OR2X2 OR2X2_5752 ( .A(alu__abc_41358_n2215), .B(alu_b_i_3_bF_buf1), .Y(alu__abc_41358_n2216) );
  OR2X2 OR2X2_5753 ( .A(alu__abc_41358_n2216), .B(alu__abc_41358_n2214), .Y(alu__abc_41358_n2217) );
  OR2X2 OR2X2_5754 ( .A(alu__abc_41358_n1880), .B(alu__abc_41358_n294_bF_buf5), .Y(alu__abc_41358_n2218) );
  OR2X2 OR2X2_5755 ( .A(alu__abc_41358_n2225), .B(alu__abc_41358_n2226), .Y(alu__abc_41358_n2227) );
  OR2X2 OR2X2_5756 ( .A(alu__abc_41358_n2221), .B(alu__abc_41358_n2227), .Y(alu__abc_41358_n2228) );
  OR2X2 OR2X2_5757 ( .A(alu__abc_41358_n2220), .B(alu__abc_41358_n2228), .Y(alu__abc_41358_n2229) );
  OR2X2 OR2X2_5758 ( .A(alu__abc_41358_n2229), .B(alu__abc_41358_n2209), .Y(alu__abc_41358_n2230) );
  OR2X2 OR2X2_5759 ( .A(alu__abc_41358_n2208), .B(alu__abc_41358_n2230), .Y(alu__abc_41358_n2231) );
  OR2X2 OR2X2_576 ( .A(_abc_43815_n2280), .B(_abc_43815_n1278_bF_buf2), .Y(_abc_43815_n2281) );
  OR2X2 OR2X2_5760 ( .A(alu__abc_41358_n2205), .B(alu__abc_41358_n2231), .Y(alu__abc_41358_n2232) );
  OR2X2 OR2X2_5761 ( .A(alu__abc_41358_n2204), .B(alu__abc_41358_n2232), .Y(alu__abc_41358_n2233) );
  OR2X2 OR2X2_5762 ( .A(alu__abc_41358_n2198), .B(alu__abc_41358_n2233), .Y(alu_p_o_25_) );
  OR2X2 OR2X2_5763 ( .A(alu__abc_41358_n2195), .B(alu__abc_41358_n659), .Y(alu__abc_41358_n2235) );
  OR2X2 OR2X2_5764 ( .A(alu__abc_41358_n2240), .B(alu__abc_41358_n394), .Y(alu__abc_41358_n2241) );
  OR2X2 OR2X2_5765 ( .A(alu__abc_41358_n2242), .B(alu__abc_41358_n134), .Y(alu__abc_41358_n2243) );
  OR2X2 OR2X2_5766 ( .A(alu__abc_41358_n2249), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2250) );
  OR2X2 OR2X2_5767 ( .A(alu__abc_41358_n2088), .B(alu__abc_41358_n299_bF_buf3), .Y(alu__abc_41358_n2253) );
  OR2X2 OR2X2_5768 ( .A(alu__abc_41358_n2254), .B(alu_b_i_1_bF_buf4), .Y(alu__abc_41358_n2255) );
  OR2X2 OR2X2_5769 ( .A(alu__abc_41358_n2171), .B(alu__abc_41358_n252_bF_buf5), .Y(alu__abc_41358_n2256) );
  OR2X2 OR2X2_577 ( .A(_abc_43815_n2253), .B(_abc_43815_n2250), .Y(_abc_43815_n2282_1) );
  OR2X2 OR2X2_5770 ( .A(alu__abc_41358_n2257), .B(alu_b_i_2_bF_buf2), .Y(alu__abc_41358_n2258) );
  OR2X2 OR2X2_5771 ( .A(alu__abc_41358_n2259), .B(alu_b_i_3_bF_buf0), .Y(alu__abc_41358_n2260) );
  OR2X2 OR2X2_5772 ( .A(alu__abc_41358_n1924), .B(alu__abc_41358_n294_bF_buf4), .Y(alu__abc_41358_n2261) );
  OR2X2 OR2X2_5773 ( .A(alu__abc_41358_n2269), .B(alu__abc_41358_n2265), .Y(alu__abc_41358_n2270) );
  OR2X2 OR2X2_5774 ( .A(alu__abc_41358_n2264), .B(alu__abc_41358_n2270), .Y(alu__abc_41358_n2271) );
  OR2X2 OR2X2_5775 ( .A(alu__abc_41358_n2263), .B(alu__abc_41358_n2271), .Y(alu__abc_41358_n2272) );
  OR2X2 OR2X2_5776 ( .A(alu__abc_41358_n2272), .B(alu__abc_41358_n2252), .Y(alu__abc_41358_n2273) );
  OR2X2 OR2X2_5777 ( .A(alu__abc_41358_n2251), .B(alu__abc_41358_n2273), .Y(alu__abc_41358_n2274) );
  OR2X2 OR2X2_5778 ( .A(alu__abc_41358_n2248), .B(alu__abc_41358_n2274), .Y(alu__abc_41358_n2275) );
  OR2X2 OR2X2_5779 ( .A(alu__abc_41358_n2247), .B(alu__abc_41358_n2275), .Y(alu__abc_41358_n2276) );
  OR2X2 OR2X2_578 ( .A(opcode_q_21_), .B(pc_q_23_), .Y(_abc_43815_n2284) );
  OR2X2 OR2X2_5780 ( .A(alu__abc_41358_n2239), .B(alu__abc_41358_n2276), .Y(alu_p_o_26_) );
  OR2X2 OR2X2_5781 ( .A(alu__abc_41358_n2236), .B(alu__abc_41358_n657), .Y(alu__abc_41358_n2278) );
  OR2X2 OR2X2_5782 ( .A(alu__abc_41358_n2244), .B(alu__abc_41358_n389), .Y(alu__abc_41358_n2283) );
  OR2X2 OR2X2_5783 ( .A(alu__abc_41358_n2284), .B(alu__abc_41358_n141), .Y(alu__abc_41358_n2285) );
  OR2X2 OR2X2_5784 ( .A(alu__abc_41358_n2283), .B(alu__abc_41358_n142), .Y(alu__abc_41358_n2286) );
  OR2X2 OR2X2_5785 ( .A(alu__abc_41358_n2290), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2291) );
  OR2X2 OR2X2_5786 ( .A(alu__abc_41358_n2293), .B(alu_b_i_1_bF_buf3), .Y(alu__abc_41358_n2294) );
  OR2X2 OR2X2_5787 ( .A(alu__abc_41358_n2210), .B(alu__abc_41358_n252_bF_buf4), .Y(alu__abc_41358_n2295) );
  OR2X2 OR2X2_5788 ( .A(alu__abc_41358_n2296), .B(alu_b_i_2_bF_buf1), .Y(alu__abc_41358_n2297) );
  OR2X2 OR2X2_5789 ( .A(alu__abc_41358_n2130), .B(alu__abc_41358_n299_bF_buf2), .Y(alu__abc_41358_n2298) );
  OR2X2 OR2X2_579 ( .A(_abc_43815_n2283), .B(_abc_43815_n2288), .Y(_abc_43815_n2289) );
  OR2X2 OR2X2_5790 ( .A(alu__abc_41358_n2299), .B(alu_b_i_3_bF_buf6), .Y(alu__abc_41358_n2300) );
  OR2X2 OR2X2_5791 ( .A(alu__abc_41358_n1966), .B(alu__abc_41358_n294_bF_buf3), .Y(alu__abc_41358_n2301) );
  OR2X2 OR2X2_5792 ( .A(alu__abc_41358_n2310), .B(alu__abc_41358_n2306), .Y(alu__abc_41358_n2311) );
  OR2X2 OR2X2_5793 ( .A(alu__abc_41358_n2305), .B(alu__abc_41358_n2311), .Y(alu__abc_41358_n2312) );
  OR2X2 OR2X2_5794 ( .A(alu__abc_41358_n2304), .B(alu__abc_41358_n2312), .Y(alu__abc_41358_n2313) );
  OR2X2 OR2X2_5795 ( .A(alu__abc_41358_n2313), .B(alu__abc_41358_n2303), .Y(alu__abc_41358_n2314) );
  OR2X2 OR2X2_5796 ( .A(alu__abc_41358_n2292), .B(alu__abc_41358_n2314), .Y(alu__abc_41358_n2315) );
  OR2X2 OR2X2_5797 ( .A(alu__abc_41358_n2289), .B(alu__abc_41358_n2315), .Y(alu__abc_41358_n2316) );
  OR2X2 OR2X2_5798 ( .A(alu__abc_41358_n2288), .B(alu__abc_41358_n2316), .Y(alu__abc_41358_n2317) );
  OR2X2 OR2X2_5799 ( .A(alu__abc_41358_n2282), .B(alu__abc_41358_n2317), .Y(alu_p_o_27_) );
  OR2X2 OR2X2_58 ( .A(_abc_43815_n812), .B(_abc_43815_n815), .Y(_abc_43815_n816_1) );
  OR2X2 OR2X2_580 ( .A(_abc_43815_n2282_1), .B(_abc_43815_n2287), .Y(_abc_43815_n2290) );
  OR2X2 OR2X2_5800 ( .A(alu__abc_41358_n2279), .B(alu__abc_41358_n822), .Y(alu__abc_41358_n2319) );
  OR2X2 OR2X2_5801 ( .A(alu__abc_41358_n495), .B(alu__abc_41358_n152), .Y(alu__abc_41358_n2324) );
  OR2X2 OR2X2_5802 ( .A(alu__abc_41358_n1651), .B(alu_b_i_4_bF_buf0), .Y(alu__abc_41358_n2330) );
  OR2X2 OR2X2_5803 ( .A(alu__abc_41358_n2009), .B(alu__abc_41358_n294_bF_buf2), .Y(alu__abc_41358_n2332) );
  OR2X2 OR2X2_5804 ( .A(alu__abc_41358_n2254), .B(alu__abc_41358_n252_bF_buf3), .Y(alu__abc_41358_n2333) );
  OR2X2 OR2X2_5805 ( .A(alu__abc_41358_n2334), .B(alu_b_i_1_bF_buf2), .Y(alu__abc_41358_n2335) );
  OR2X2 OR2X2_5806 ( .A(alu__abc_41358_n2336), .B(alu_b_i_2_bF_buf0), .Y(alu__abc_41358_n2337) );
  OR2X2 OR2X2_5807 ( .A(alu__abc_41358_n2173), .B(alu__abc_41358_n299_bF_buf1), .Y(alu__abc_41358_n2338) );
  OR2X2 OR2X2_5808 ( .A(alu__abc_41358_n2339), .B(alu_b_i_3_bF_buf5), .Y(alu__abc_41358_n2340) );
  OR2X2 OR2X2_5809 ( .A(alu__abc_41358_n2348), .B(alu__abc_41358_n2349), .Y(alu__abc_41358_n2350) );
  OR2X2 OR2X2_581 ( .A(_abc_43815_n1428_bF_buf0), .B(_abc_43815_n2293), .Y(_abc_43815_n2294) );
  OR2X2 OR2X2_5810 ( .A(alu__abc_41358_n2350), .B(alu__abc_41358_n2347), .Y(alu__abc_41358_n2351) );
  OR2X2 OR2X2_5811 ( .A(alu__abc_41358_n2343), .B(alu__abc_41358_n2351), .Y(alu__abc_41358_n2352) );
  OR2X2 OR2X2_5812 ( .A(alu__abc_41358_n2352), .B(alu__abc_41358_n2342), .Y(alu__abc_41358_n2353) );
  OR2X2 OR2X2_5813 ( .A(alu__abc_41358_n2353), .B(alu__abc_41358_n2331), .Y(alu__abc_41358_n2354) );
  OR2X2 OR2X2_5814 ( .A(alu__abc_41358_n2329), .B(alu__abc_41358_n2354), .Y(alu__abc_41358_n2355) );
  OR2X2 OR2X2_5815 ( .A(alu__abc_41358_n2328), .B(alu__abc_41358_n2355), .Y(alu__abc_41358_n2356) );
  OR2X2 OR2X2_5816 ( .A(alu__abc_41358_n2323), .B(alu__abc_41358_n2356), .Y(alu_p_o_28_) );
  OR2X2 OR2X2_5817 ( .A(alu__abc_41358_n2321), .B(alu__abc_41358_n636), .Y(alu__abc_41358_n2358) );
  OR2X2 OR2X2_5818 ( .A(alu__abc_41358_n2363), .B(alu__abc_41358_n159_1), .Y(alu__abc_41358_n2364) );
  OR2X2 OR2X2_5819 ( .A(alu__abc_41358_n2365), .B(alu__abc_41358_n160_1), .Y(alu__abc_41358_n2366) );
  OR2X2 OR2X2_582 ( .A(_abc_43815_n2292_1), .B(_abc_43815_n2294), .Y(_abc_43815_n2295) );
  OR2X2 OR2X2_5820 ( .A(alu__abc_41358_n2370), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2371) );
  OR2X2 OR2X2_5821 ( .A(alu__abc_41358_n1709), .B(alu__abc_41358_n279_bF_buf5), .Y(alu__abc_41358_n2373) );
  OR2X2 OR2X2_5822 ( .A(alu_a_i_29_), .B(alu_b_i_0_bF_buf1), .Y(alu__abc_41358_n2374) );
  OR2X2 OR2X2_5823 ( .A(alu__abc_41358_n2375), .B(alu_b_i_1_bF_buf1), .Y(alu__abc_41358_n2376) );
  OR2X2 OR2X2_5824 ( .A(alu__abc_41358_n2293), .B(alu__abc_41358_n252_bF_buf2), .Y(alu__abc_41358_n2377) );
  OR2X2 OR2X2_5825 ( .A(alu__abc_41358_n2378), .B(alu_b_i_2_bF_buf6), .Y(alu__abc_41358_n2379) );
  OR2X2 OR2X2_5826 ( .A(alu__abc_41358_n2213), .B(alu__abc_41358_n299_bF_buf0), .Y(alu__abc_41358_n2380) );
  OR2X2 OR2X2_5827 ( .A(alu__abc_41358_n2383), .B(alu_b_i_4_bF_buf4), .Y(alu__abc_41358_n2384) );
  OR2X2 OR2X2_5828 ( .A(alu__abc_41358_n2384), .B(alu__abc_41358_n2382), .Y(alu__abc_41358_n2385) );
  OR2X2 OR2X2_5829 ( .A(alu__abc_41358_n2392), .B(alu__abc_41358_n2393), .Y(alu__abc_41358_n2394) );
  OR2X2 OR2X2_583 ( .A(_abc_43815_n1431_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_43815_n2296) );
  OR2X2 OR2X2_5830 ( .A(alu__abc_41358_n2394), .B(alu__abc_41358_n2391), .Y(alu__abc_41358_n2395) );
  OR2X2 OR2X2_5831 ( .A(alu__abc_41358_n2387), .B(alu__abc_41358_n2395), .Y(alu__abc_41358_n2396) );
  OR2X2 OR2X2_5832 ( .A(alu__abc_41358_n2372), .B(alu__abc_41358_n2396), .Y(alu__abc_41358_n2397) );
  OR2X2 OR2X2_5833 ( .A(alu__abc_41358_n2369), .B(alu__abc_41358_n2397), .Y(alu__abc_41358_n2398) );
  OR2X2 OR2X2_5834 ( .A(alu__abc_41358_n2368), .B(alu__abc_41358_n2398), .Y(alu__abc_41358_n2399) );
  OR2X2 OR2X2_5835 ( .A(alu__abc_41358_n2362), .B(alu__abc_41358_n2399), .Y(alu_p_o_29_) );
  OR2X2 OR2X2_5836 ( .A(alu__abc_41358_n2359), .B(alu__abc_41358_n629), .Y(alu__abc_41358_n2403) );
  OR2X2 OR2X2_5837 ( .A(alu__abc_41358_n505), .B(alu__abc_41358_n169), .Y(alu__abc_41358_n2406) );
  OR2X2 OR2X2_5838 ( .A(alu__abc_41358_n2410), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2411) );
  OR2X2 OR2X2_5839 ( .A(alu__abc_41358_n2413), .B(alu_b_i_1_bF_buf0), .Y(alu__abc_41358_n2414) );
  OR2X2 OR2X2_584 ( .A(_abc_43815_n2297), .B(_abc_43815_n1473_bF_buf3), .Y(_abc_43815_n2298) );
  OR2X2 OR2X2_5840 ( .A(alu__abc_41358_n2334), .B(alu__abc_41358_n252_bF_buf1), .Y(alu__abc_41358_n2415) );
  OR2X2 OR2X2_5841 ( .A(alu__abc_41358_n2416), .B(alu_b_i_2_bF_buf5), .Y(alu__abc_41358_n2417) );
  OR2X2 OR2X2_5842 ( .A(alu__abc_41358_n2257), .B(alu__abc_41358_n299_bF_buf7), .Y(alu__abc_41358_n2418) );
  OR2X2 OR2X2_5843 ( .A(alu__abc_41358_n2419), .B(alu_b_i_3_bF_buf3), .Y(alu__abc_41358_n2420) );
  OR2X2 OR2X2_5844 ( .A(alu__abc_41358_n2091), .B(alu__abc_41358_n294_bF_buf0), .Y(alu__abc_41358_n2421) );
  OR2X2 OR2X2_5845 ( .A(alu__abc_41358_n2429), .B(alu__abc_41358_n2430), .Y(alu__abc_41358_n2431) );
  OR2X2 OR2X2_5846 ( .A(alu__abc_41358_n2425), .B(alu__abc_41358_n2431), .Y(alu__abc_41358_n2432) );
  OR2X2 OR2X2_5847 ( .A(alu__abc_41358_n2424), .B(alu__abc_41358_n2432), .Y(alu__abc_41358_n2433) );
  OR2X2 OR2X2_5848 ( .A(alu__abc_41358_n2433), .B(alu__abc_41358_n2423), .Y(alu__abc_41358_n2434) );
  OR2X2 OR2X2_5849 ( .A(alu__abc_41358_n2412), .B(alu__abc_41358_n2434), .Y(alu__abc_41358_n2435) );
  OR2X2 OR2X2_585 ( .A(_abc_43815_n2279), .B(_abc_43815_n1472_1_bF_buf2), .Y(_abc_43815_n2299) );
  OR2X2 OR2X2_5850 ( .A(alu__abc_41358_n2409), .B(alu__abc_41358_n2435), .Y(alu__abc_41358_n2436) );
  OR2X2 OR2X2_5851 ( .A(alu__abc_41358_n2408), .B(alu__abc_41358_n2436), .Y(alu__abc_41358_n2437) );
  OR2X2 OR2X2_5852 ( .A(alu__abc_41358_n2405), .B(alu__abc_41358_n2437), .Y(alu_p_o_30_) );
  OR2X2 OR2X2_5853 ( .A(alu__abc_41358_n2401), .B(alu__abc_41358_n627), .Y(alu__abc_41358_n2439) );
  OR2X2 OR2X2_5854 ( .A(alu__abc_41358_n963), .B(alu__abc_41358_n966), .Y(alu__abc_41358_n2443) );
  OR2X2 OR2X2_5855 ( .A(alu__abc_41358_n2443), .B(alu_b_i_1_bF_buf7), .Y(alu__abc_41358_n2444) );
  OR2X2 OR2X2_5856 ( .A(alu__abc_41358_n2375), .B(alu__abc_41358_n252_bF_buf0), .Y(alu__abc_41358_n2445) );
  OR2X2 OR2X2_5857 ( .A(alu__abc_41358_n2448), .B(alu_b_i_3_bF_buf2), .Y(alu__abc_41358_n2449) );
  OR2X2 OR2X2_5858 ( .A(alu__abc_41358_n2449), .B(alu__abc_41358_n2447), .Y(alu__abc_41358_n2450) );
  OR2X2 OR2X2_5859 ( .A(alu__abc_41358_n2133), .B(alu__abc_41358_n294_bF_buf7), .Y(alu__abc_41358_n2451) );
  OR2X2 OR2X2_586 ( .A(_abc_43815_n2300), .B(_abc_43815_n1350_bF_buf3), .Y(_abc_43815_n2301) );
  OR2X2 OR2X2_5860 ( .A(alu__abc_41358_n506), .B(alu__abc_41358_n508), .Y(alu__abc_41358_n2455) );
  OR2X2 OR2X2_5861 ( .A(alu__abc_41358_n511), .B(alu__abc_41358_n2456), .Y(alu__abc_41358_n2457) );
  OR2X2 OR2X2_5862 ( .A(alu__abc_41358_n2459), .B(alu__abc_41358_n1871), .Y(alu__abc_41358_n2460) );
  OR2X2 OR2X2_5863 ( .A(alu__abc_41358_n2467), .B(alu__abc_41358_n2468), .Y(alu__abc_41358_n2469) );
  OR2X2 OR2X2_5864 ( .A(alu__abc_41358_n2463), .B(alu__abc_41358_n2469), .Y(alu__abc_41358_n2470) );
  OR2X2 OR2X2_5865 ( .A(alu__abc_41358_n2462), .B(alu__abc_41358_n2470), .Y(alu__abc_41358_n2471) );
  OR2X2 OR2X2_5866 ( .A(alu__abc_41358_n2461), .B(alu__abc_41358_n2471), .Y(alu__abc_41358_n2472) );
  OR2X2 OR2X2_5867 ( .A(alu__abc_41358_n2458), .B(alu__abc_41358_n2472), .Y(alu__abc_41358_n2473) );
  OR2X2 OR2X2_5868 ( .A(alu__abc_41358_n2473), .B(alu__abc_41358_n2454), .Y(alu__abc_41358_n2474) );
  OR2X2 OR2X2_5869 ( .A(alu__abc_41358_n2474), .B(alu__abc_41358_n2453), .Y(alu__abc_41358_n2475) );
  OR2X2 OR2X2_587 ( .A(_abc_43815_n2303), .B(_abc_43815_n2302_1), .Y(_abc_43815_n2304) );
  OR2X2 OR2X2_5870 ( .A(alu__abc_41358_n2442), .B(alu__abc_41358_n2475), .Y(alu_p_o_31_) );
  OR2X2 OR2X2_5871 ( .A(alu__abc_41358_n949), .B(alu_a_i_1_), .Y(alu__abc_41358_n2477) );
  OR2X2 OR2X2_5872 ( .A(alu__abc_41358_n2482), .B(alu__abc_41358_n405), .Y(alu__abc_41358_n2483) );
  OR2X2 OR2X2_5873 ( .A(alu__abc_41358_n2485), .B(alu__abc_41358_n409), .Y(alu__abc_41358_n2486) );
  OR2X2 OR2X2_5874 ( .A(alu__abc_41358_n2487), .B(alu__abc_41358_n2483), .Y(alu__abc_41358_n2488) );
  OR2X2 OR2X2_5875 ( .A(alu__abc_41358_n2490), .B(alu__abc_41358_n413), .Y(alu__abc_41358_n2491) );
  OR2X2 OR2X2_5876 ( .A(alu__abc_41358_n2488), .B(alu__abc_41358_n2492), .Y(alu__abc_41358_n2493) );
  OR2X2 OR2X2_5877 ( .A(alu__abc_41358_n2493), .B(alu__abc_41358_n2480), .Y(alu__abc_41358_n2494) );
  OR2X2 OR2X2_5878 ( .A(alu__abc_41358_n2498), .B(alu__abc_41358_n2496), .Y(alu__abc_41358_n2499) );
  OR2X2 OR2X2_5879 ( .A(alu__abc_41358_n435), .B(alu__abc_41358_n2500), .Y(alu__abc_41358_n2501) );
  OR2X2 OR2X2_588 ( .A(_abc_43815_n1413_bF_buf1), .B(_abc_43815_n2304), .Y(_abc_43815_n2305) );
  OR2X2 OR2X2_5880 ( .A(alu__abc_41358_n2499), .B(alu__abc_41358_n2503), .Y(alu__abc_41358_n2504) );
  OR2X2 OR2X2_5881 ( .A(alu__abc_41358_n2508), .B(alu__abc_41358_n2506), .Y(alu__abc_41358_n2509) );
  OR2X2 OR2X2_5882 ( .A(alu__abc_41358_n450), .B(alu__abc_41358_n2510), .Y(alu__abc_41358_n2511) );
  OR2X2 OR2X2_5883 ( .A(alu__abc_41358_n2509), .B(alu__abc_41358_n2513), .Y(alu__abc_41358_n2514) );
  OR2X2 OR2X2_5884 ( .A(alu__abc_41358_n2505), .B(alu__abc_41358_n2514), .Y(alu__abc_41358_n2515) );
  OR2X2 OR2X2_5885 ( .A(alu__abc_41358_n2495), .B(alu__abc_41358_n2515), .Y(alu__abc_41358_n2516) );
  OR2X2 OR2X2_5886 ( .A(alu__abc_41358_n2520), .B(alu__abc_41358_n2518), .Y(alu__abc_41358_n2521) );
  OR2X2 OR2X2_5887 ( .A(alu__abc_41358_n394), .B(alu__abc_41358_n2522), .Y(alu__abc_41358_n2523) );
  OR2X2 OR2X2_5888 ( .A(alu__abc_41358_n2521), .B(alu__abc_41358_n2525), .Y(alu__abc_41358_n2526) );
  OR2X2 OR2X2_5889 ( .A(alu__abc_41358_n2529), .B(alu__abc_41358_n2530), .Y(alu__abc_41358_n2531) );
  OR2X2 OR2X2_589 ( .A(_abc_43815_n2307), .B(_abc_43815_n2281), .Y(_abc_43815_n2308) );
  OR2X2 OR2X2_5890 ( .A(alu__abc_41358_n497), .B(alu__abc_41358_n2532), .Y(alu__abc_41358_n2533) );
  OR2X2 OR2X2_5891 ( .A(alu__abc_41358_n2535), .B(alu__abc_41358_n2531), .Y(alu__abc_41358_n2536) );
  OR2X2 OR2X2_5892 ( .A(alu__abc_41358_n2527), .B(alu__abc_41358_n2536), .Y(alu__abc_41358_n2537) );
  OR2X2 OR2X2_5893 ( .A(alu__abc_41358_n2540), .B(alu__abc_41358_n2538), .Y(alu__abc_41358_n2541) );
  OR2X2 OR2X2_5894 ( .A(alu__abc_41358_n467), .B(alu__abc_41358_n2542), .Y(alu__abc_41358_n2543) );
  OR2X2 OR2X2_5895 ( .A(alu__abc_41358_n2541), .B(alu__abc_41358_n2545), .Y(alu__abc_41358_n2546) );
  OR2X2 OR2X2_5896 ( .A(alu__abc_41358_n2550), .B(alu__abc_41358_n2548), .Y(alu__abc_41358_n2551) );
  OR2X2 OR2X2_5897 ( .A(alu__abc_41358_n482), .B(alu__abc_41358_n2552), .Y(alu__abc_41358_n2553) );
  OR2X2 OR2X2_5898 ( .A(alu__abc_41358_n2551), .B(alu__abc_41358_n2555), .Y(alu__abc_41358_n2556) );
  OR2X2 OR2X2_5899 ( .A(alu__abc_41358_n2547), .B(alu__abc_41358_n2556), .Y(alu__abc_41358_n2557) );
  OR2X2 OR2X2_59 ( .A(_abc_43815_n686_1_bF_buf2), .B(_abc_43815_n816_1), .Y(_abc_43815_n817_1) );
  OR2X2 OR2X2_590 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_23_), .Y(_abc_43815_n2309) );
  OR2X2 OR2X2_5900 ( .A(alu__abc_41358_n2558), .B(alu__abc_41358_n2537), .Y(alu__abc_41358_n2559) );
  OR2X2 OR2X2_5901 ( .A(alu__abc_41358_n2517), .B(alu__abc_41358_n2559), .Y(alu__abc_41358_n2560) );
  OR2X2 OR2X2_591 ( .A(_abc_43815_n2277), .B(pc_q_24_), .Y(_abc_43815_n2312_1) );
  OR2X2 OR2X2_592 ( .A(_abc_43815_n2316), .B(_abc_43815_n1278_bF_buf1), .Y(_abc_43815_n2317) );
  OR2X2 OR2X2_593 ( .A(_abc_43815_n2217), .B(_abc_43815_n2210), .Y(_abc_43815_n2318) );
  OR2X2 OR2X2_594 ( .A(_abc_43815_n2321), .B(_abc_43815_n2285), .Y(_abc_43815_n2322_1) );
  OR2X2 OR2X2_595 ( .A(_abc_43815_n2320), .B(_abc_43815_n2322_1), .Y(_abc_43815_n2323) );
  OR2X2 OR2X2_596 ( .A(_abc_43815_n2325), .B(_abc_43815_n2323), .Y(_abc_43815_n2326) );
  OR2X2 OR2X2_597 ( .A(opcode_q_22_), .B(pc_q_24_), .Y(_abc_43815_n2327) );
  OR2X2 OR2X2_598 ( .A(_abc_43815_n2326), .B(_abc_43815_n2330), .Y(_abc_43815_n2333) );
  OR2X2 OR2X2_599 ( .A(_abc_43815_n1428_bF_buf4), .B(_abc_43815_n2336), .Y(_abc_43815_n2337) );
  OR2X2 OR2X2_6 ( .A(_abc_43815_n672), .B(_abc_43815_n635), .Y(_abc_27555_n288) );
  OR2X2 OR2X2_60 ( .A(_abc_43815_n819), .B(_abc_43815_n818), .Y(_abc_43815_n820) );
  OR2X2 OR2X2_600 ( .A(_abc_43815_n2335), .B(_abc_43815_n2337), .Y(_abc_43815_n2338) );
  OR2X2 OR2X2_601 ( .A(_abc_43815_n1431_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_43815_n2339) );
  OR2X2 OR2X2_602 ( .A(_abc_43815_n2340), .B(_abc_43815_n1473_bF_buf2), .Y(_abc_43815_n2341) );
  OR2X2 OR2X2_603 ( .A(_abc_43815_n2315), .B(_abc_43815_n1472_1_bF_buf1), .Y(_abc_43815_n2342_1) );
  OR2X2 OR2X2_604 ( .A(_abc_43815_n2343), .B(_abc_43815_n1350_bF_buf2), .Y(_abc_43815_n2344) );
  OR2X2 OR2X2_605 ( .A(_abc_43815_n2346), .B(_abc_43815_n2345), .Y(_abc_43815_n2347) );
  OR2X2 OR2X2_606 ( .A(_abc_43815_n1413_bF_buf0), .B(_abc_43815_n2347), .Y(_abc_43815_n2348) );
  OR2X2 OR2X2_607 ( .A(_abc_43815_n2350), .B(_abc_43815_n2317), .Y(_abc_43815_n2351) );
  OR2X2 OR2X2_608 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_24_), .Y(_abc_43815_n2352_1) );
  OR2X2 OR2X2_609 ( .A(_abc_43815_n2313), .B(pc_q_25_), .Y(_abc_43815_n2355) );
  OR2X2 OR2X2_61 ( .A(_abc_43815_n820), .B(_abc_43815_n685), .Y(_abc_43815_n821) );
  OR2X2 OR2X2_610 ( .A(_abc_43815_n2359), .B(_abc_43815_n1278_bF_buf0), .Y(_abc_43815_n2360) );
  OR2X2 OR2X2_611 ( .A(opcode_q_23_), .B(pc_q_25_), .Y(_abc_43815_n2361) );
  OR2X2 OR2X2_612 ( .A(_abc_43815_n2364), .B(_abc_43815_n2328), .Y(_abc_43815_n2365) );
  OR2X2 OR2X2_613 ( .A(_abc_43815_n2331), .B(_abc_43815_n2365), .Y(_abc_43815_n2366) );
  OR2X2 OR2X2_614 ( .A(_abc_43815_n1428_bF_buf3), .B(_abc_43815_n2375), .Y(_abc_43815_n2376) );
  OR2X2 OR2X2_615 ( .A(_abc_43815_n2374), .B(_abc_43815_n2376), .Y(_abc_43815_n2377) );
  OR2X2 OR2X2_616 ( .A(_abc_43815_n1431_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_43815_n2378) );
  OR2X2 OR2X2_617 ( .A(_abc_43815_n2379), .B(_abc_43815_n1473_bF_buf1), .Y(_abc_43815_n2380) );
  OR2X2 OR2X2_618 ( .A(_abc_43815_n2358), .B(_abc_43815_n1472_1_bF_buf0), .Y(_abc_43815_n2381) );
  OR2X2 OR2X2_619 ( .A(_abc_43815_n2382), .B(_abc_43815_n1350_bF_buf1), .Y(_abc_43815_n2383) );
  OR2X2 OR2X2_62 ( .A(_abc_43815_n822), .B(_abc_43815_n682), .Y(_abc_43815_n823) );
  OR2X2 OR2X2_620 ( .A(_abc_43815_n2385), .B(_abc_43815_n2384), .Y(_abc_43815_n2386) );
  OR2X2 OR2X2_621 ( .A(_abc_43815_n1413_bF_buf4), .B(_abc_43815_n2386), .Y(_abc_43815_n2387) );
  OR2X2 OR2X2_622 ( .A(_abc_43815_n2389), .B(_abc_43815_n2360), .Y(_abc_43815_n2390) );
  OR2X2 OR2X2_623 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_25_), .Y(_abc_43815_n2391) );
  OR2X2 OR2X2_624 ( .A(_abc_43815_n2356), .B(pc_q_26_), .Y(_abc_43815_n2394) );
  OR2X2 OR2X2_625 ( .A(_abc_43815_n2398), .B(_abc_43815_n1278_bF_buf7), .Y(_abc_43815_n2399) );
  OR2X2 OR2X2_626 ( .A(opcode_q_24_), .B(pc_q_26_), .Y(_abc_43815_n2403) );
  OR2X2 OR2X2_627 ( .A(_abc_43815_n2402), .B(_abc_43815_n2406), .Y(_abc_43815_n2409) );
  OR2X2 OR2X2_628 ( .A(_abc_43815_n1428_bF_buf2), .B(_abc_43815_n2412), .Y(_abc_43815_n2413) );
  OR2X2 OR2X2_629 ( .A(_abc_43815_n2411), .B(_abc_43815_n2413), .Y(_abc_43815_n2414) );
  OR2X2 OR2X2_63 ( .A(state_q_1_bF_buf4), .B(alu_p_o_7_), .Y(_abc_43815_n824) );
  OR2X2 OR2X2_630 ( .A(_abc_43815_n1431_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_43815_n2415) );
  OR2X2 OR2X2_631 ( .A(_abc_43815_n2416), .B(_abc_43815_n1473_bF_buf0), .Y(_abc_43815_n2417) );
  OR2X2 OR2X2_632 ( .A(_abc_43815_n2397), .B(_abc_43815_n1472_1_bF_buf4), .Y(_abc_43815_n2418) );
  OR2X2 OR2X2_633 ( .A(_abc_43815_n2419), .B(_abc_43815_n1350_bF_buf0), .Y(_abc_43815_n2420_1) );
  OR2X2 OR2X2_634 ( .A(_abc_43815_n2422), .B(_abc_43815_n2421), .Y(_abc_43815_n2423) );
  OR2X2 OR2X2_635 ( .A(_abc_43815_n1413_bF_buf3), .B(_abc_43815_n2423), .Y(_abc_43815_n2424) );
  OR2X2 OR2X2_636 ( .A(_abc_43815_n2426), .B(_abc_43815_n2399), .Y(_abc_43815_n2427) );
  OR2X2 OR2X2_637 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_26_), .Y(_abc_43815_n2428) );
  OR2X2 OR2X2_638 ( .A(_abc_43815_n2395), .B(pc_q_27_), .Y(_abc_43815_n2431) );
  OR2X2 OR2X2_639 ( .A(_abc_43815_n2435), .B(_abc_43815_n1278_bF_buf6), .Y(_abc_43815_n2436) );
  OR2X2 OR2X2_64 ( .A(state_q_1_bF_buf3), .B(alu_p_o_8_), .Y(_abc_43815_n826) );
  OR2X2 OR2X2_640 ( .A(opcode_q_25_), .B(pc_q_27_), .Y(_abc_43815_n2437) );
  OR2X2 OR2X2_641 ( .A(_abc_43815_n2440), .B(_abc_43815_n2404), .Y(_abc_43815_n2441) );
  OR2X2 OR2X2_642 ( .A(_abc_43815_n2407), .B(_abc_43815_n2441), .Y(_abc_43815_n2442) );
  OR2X2 OR2X2_643 ( .A(_abc_43815_n2401), .B(_abc_43815_n2444), .Y(_abc_43815_n2445_1) );
  OR2X2 OR2X2_644 ( .A(_abc_43815_n1428_bF_buf1), .B(_abc_43815_n2451), .Y(_abc_43815_n2452) );
  OR2X2 OR2X2_645 ( .A(_abc_43815_n2450), .B(_abc_43815_n2452), .Y(_abc_43815_n2453) );
  OR2X2 OR2X2_646 ( .A(_abc_43815_n1431_1_bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_43815_n2454) );
  OR2X2 OR2X2_647 ( .A(_abc_43815_n2455), .B(_abc_43815_n1473_bF_buf4), .Y(_abc_43815_n2456) );
  OR2X2 OR2X2_648 ( .A(_abc_43815_n2434), .B(_abc_43815_n1472_1_bF_buf3), .Y(_abc_43815_n2457) );
  OR2X2 OR2X2_649 ( .A(_abc_43815_n2458), .B(_abc_43815_n1350_bF_buf4), .Y(_abc_43815_n2459) );
  OR2X2 OR2X2_65 ( .A(_abc_43815_n693), .B(\mem_dat_i[8] ), .Y(_abc_43815_n827) );
  OR2X2 OR2X2_650 ( .A(_abc_43815_n2461), .B(_abc_43815_n2460), .Y(_abc_43815_n2462) );
  OR2X2 OR2X2_651 ( .A(_abc_43815_n1413_bF_buf2), .B(_abc_43815_n2462), .Y(_abc_43815_n2463) );
  OR2X2 OR2X2_652 ( .A(_abc_43815_n2465), .B(_abc_43815_n2436), .Y(_abc_43815_n2466) );
  OR2X2 OR2X2_653 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_27_), .Y(_abc_43815_n2467) );
  OR2X2 OR2X2_654 ( .A(_abc_43815_n2432), .B(pc_q_28_), .Y(_abc_43815_n2470) );
  OR2X2 OR2X2_655 ( .A(_abc_43815_n2474), .B(_abc_43815_n1278_bF_buf5), .Y(_abc_43815_n2475) );
  OR2X2 OR2X2_656 ( .A(_abc_43815_n2400), .B(_abc_43815_n2444), .Y(_abc_43815_n2477) );
  OR2X2 OR2X2_657 ( .A(_abc_43815_n2481), .B(_abc_43815_n2479), .Y(_abc_43815_n2482) );
  OR2X2 OR2X2_658 ( .A(opcode_q_25_), .B(pc_q_28_), .Y(_abc_43815_n2483) );
  OR2X2 OR2X2_659 ( .A(_abc_43815_n2482), .B(_abc_43815_n2486), .Y(_abc_43815_n2489) );
  OR2X2 OR2X2_66 ( .A(_abc_43815_n692_bF_buf1), .B(_abc_43815_n703), .Y(_abc_43815_n828) );
  OR2X2 OR2X2_660 ( .A(_abc_43815_n1428_bF_buf0), .B(_abc_43815_n2492), .Y(_abc_43815_n2493_1) );
  OR2X2 OR2X2_661 ( .A(_abc_43815_n2491), .B(_abc_43815_n2493_1), .Y(_abc_43815_n2494) );
  OR2X2 OR2X2_662 ( .A(_abc_43815_n1431_1_bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_43815_n2495) );
  OR2X2 OR2X2_663 ( .A(_abc_43815_n2496), .B(_abc_43815_n1473_bF_buf3), .Y(_abc_43815_n2497) );
  OR2X2 OR2X2_664 ( .A(_abc_43815_n2473), .B(_abc_43815_n1472_1_bF_buf2), .Y(_abc_43815_n2498) );
  OR2X2 OR2X2_665 ( .A(_abc_43815_n2499), .B(_abc_43815_n1350_bF_buf3), .Y(_abc_43815_n2500) );
  OR2X2 OR2X2_666 ( .A(_abc_43815_n2502), .B(_abc_43815_n2501), .Y(_abc_43815_n2503) );
  OR2X2 OR2X2_667 ( .A(_abc_43815_n1413_bF_buf1), .B(_abc_43815_n2503), .Y(_abc_43815_n2504) );
  OR2X2 OR2X2_668 ( .A(_abc_43815_n2506), .B(_abc_43815_n2475), .Y(_abc_43815_n2507) );
  OR2X2 OR2X2_669 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_28_), .Y(_abc_43815_n2508) );
  OR2X2 OR2X2_67 ( .A(_abc_43815_n831), .B(_abc_43815_n682), .Y(_abc_43815_n832_1) );
  OR2X2 OR2X2_670 ( .A(_abc_43815_n2471), .B(pc_q_29_), .Y(_abc_43815_n2511) );
  OR2X2 OR2X2_671 ( .A(_abc_43815_n2515), .B(_abc_43815_n1278_bF_buf4), .Y(_abc_43815_n2516) );
  OR2X2 OR2X2_672 ( .A(_abc_43815_n2487), .B(_abc_43815_n2484), .Y(_abc_43815_n2517_1) );
  OR2X2 OR2X2_673 ( .A(opcode_q_25_), .B(pc_q_29_), .Y(_abc_43815_n2519) );
  OR2X2 OR2X2_674 ( .A(_abc_43815_n2518), .B(_abc_43815_n2523), .Y(_abc_43815_n2524) );
  OR2X2 OR2X2_675 ( .A(_abc_43815_n2517_1), .B(_abc_43815_n2522), .Y(_abc_43815_n2525) );
  OR2X2 OR2X2_676 ( .A(_abc_43815_n1428_bF_buf4), .B(_abc_43815_n2528), .Y(_abc_43815_n2529) );
  OR2X2 OR2X2_677 ( .A(_abc_43815_n2527), .B(_abc_43815_n2529), .Y(_abc_43815_n2530) );
  OR2X2 OR2X2_678 ( .A(_abc_43815_n1431_1_bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_43815_n2531) );
  OR2X2 OR2X2_679 ( .A(_abc_43815_n2532), .B(_abc_43815_n1473_bF_buf2), .Y(_abc_43815_n2533) );
  OR2X2 OR2X2_68 ( .A(_abc_43815_n830), .B(_abc_43815_n832_1_bF_buf3), .Y(_abc_43815_n833) );
  OR2X2 OR2X2_680 ( .A(_abc_43815_n2514), .B(_abc_43815_n1472_1_bF_buf1), .Y(_abc_43815_n2534) );
  OR2X2 OR2X2_681 ( .A(_abc_43815_n2535), .B(_abc_43815_n1350_bF_buf2), .Y(_abc_43815_n2536) );
  OR2X2 OR2X2_682 ( .A(_abc_43815_n2538), .B(_abc_43815_n2537), .Y(_abc_43815_n2539) );
  OR2X2 OR2X2_683 ( .A(_abc_43815_n1413_bF_buf0), .B(_abc_43815_n2539), .Y(_abc_43815_n2540) );
  OR2X2 OR2X2_684 ( .A(_abc_43815_n2542), .B(_abc_43815_n2516), .Y(_abc_43815_n2543) );
  OR2X2 OR2X2_685 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_29_), .Y(_abc_43815_n2544) );
  OR2X2 OR2X2_686 ( .A(_abc_43815_n2512), .B(pc_q_30_), .Y(_abc_43815_n2547) );
  OR2X2 OR2X2_687 ( .A(_abc_43815_n2551), .B(_abc_43815_n1278_bF_buf3), .Y(_abc_43815_n2552) );
  OR2X2 OR2X2_688 ( .A(_abc_43815_n2554), .B(_abc_43815_n2556), .Y(_abc_43815_n2557) );
  OR2X2 OR2X2_689 ( .A(opcode_q_25_), .B(pc_q_30_), .Y(_abc_43815_n2558) );
  OR2X2 OR2X2_69 ( .A(_abc_43815_n835), .B(_abc_43815_n836), .Y(_abc_43815_n837) );
  OR2X2 OR2X2_690 ( .A(_abc_43815_n2557), .B(_abc_43815_n2561), .Y(_abc_43815_n2564) );
  OR2X2 OR2X2_691 ( .A(_abc_43815_n1428_bF_buf3), .B(_abc_43815_n2567), .Y(_abc_43815_n2568) );
  OR2X2 OR2X2_692 ( .A(_abc_43815_n2566), .B(_abc_43815_n2568), .Y(_abc_43815_n2569) );
  OR2X2 OR2X2_693 ( .A(_abc_43815_n1431_1_bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_43815_n2570) );
  OR2X2 OR2X2_694 ( .A(_abc_43815_n2571), .B(_abc_43815_n1473_bF_buf1), .Y(_abc_43815_n2572) );
  OR2X2 OR2X2_695 ( .A(_abc_43815_n2550), .B(_abc_43815_n1472_1_bF_buf0), .Y(_abc_43815_n2573) );
  OR2X2 OR2X2_696 ( .A(_abc_43815_n2574), .B(_abc_43815_n1350_bF_buf1), .Y(_abc_43815_n2575) );
  OR2X2 OR2X2_697 ( .A(_abc_43815_n2577), .B(_abc_43815_n2576), .Y(_abc_43815_n2578) );
  OR2X2 OR2X2_698 ( .A(_abc_43815_n1413_bF_buf4), .B(_abc_43815_n2578), .Y(_abc_43815_n2579) );
  OR2X2 OR2X2_699 ( .A(_abc_43815_n2581), .B(_abc_43815_n2552), .Y(_abc_43815_n2582) );
  OR2X2 OR2X2_7 ( .A(_abc_43815_n675), .B(state_q_3_bF_buf5), .Y(_abc_27555_n343) );
  OR2X2 OR2X2_70 ( .A(_abc_43815_n838), .B(_abc_43815_n832_1_bF_buf2), .Y(_abc_43815_n839) );
  OR2X2 OR2X2_700 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_30_), .Y(_abc_43815_n2583) );
  OR2X2 OR2X2_701 ( .A(_abc_43815_n2548), .B(pc_q_31_), .Y(_abc_43815_n2586) );
  OR2X2 OR2X2_702 ( .A(_abc_43815_n2590), .B(_abc_43815_n1278_bF_buf2), .Y(_abc_43815_n2591) );
  OR2X2 OR2X2_703 ( .A(_abc_43815_n2562), .B(_abc_43815_n2559), .Y(_abc_43815_n2592) );
  OR2X2 OR2X2_704 ( .A(_abc_43815_n621), .B(pc_q_31_), .Y(_abc_43815_n2594) );
  OR2X2 OR2X2_705 ( .A(_abc_43815_n2595), .B(opcode_q_25_), .Y(_abc_43815_n2596) );
  OR2X2 OR2X2_706 ( .A(_abc_43815_n2593), .B(_abc_43815_n2597), .Y(_abc_43815_n2598) );
  OR2X2 OR2X2_707 ( .A(_abc_43815_n2592), .B(_abc_43815_n2599), .Y(_abc_43815_n2600) );
  OR2X2 OR2X2_708 ( .A(_abc_43815_n1428_bF_buf2), .B(_abc_43815_n2603), .Y(_abc_43815_n2604) );
  OR2X2 OR2X2_709 ( .A(_abc_43815_n2602), .B(_abc_43815_n2604), .Y(_abc_43815_n2605) );
  OR2X2 OR2X2_71 ( .A(state_q_1_bF_buf2), .B(alu_p_o_9_), .Y(_abc_43815_n840) );
  OR2X2 OR2X2_710 ( .A(_abc_43815_n1431_1_bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_43815_n2606) );
  OR2X2 OR2X2_711 ( .A(_abc_43815_n2607), .B(_abc_43815_n1473_bF_buf0), .Y(_abc_43815_n2608) );
  OR2X2 OR2X2_712 ( .A(_abc_43815_n2589_1), .B(_abc_43815_n1472_1_bF_buf4), .Y(_abc_43815_n2609) );
  OR2X2 OR2X2_713 ( .A(_abc_43815_n2610), .B(_abc_43815_n1350_bF_buf0), .Y(_abc_43815_n2611) );
  OR2X2 OR2X2_714 ( .A(_abc_43815_n2613), .B(_abc_43815_n2612), .Y(_abc_43815_n2614_1) );
  OR2X2 OR2X2_715 ( .A(_abc_43815_n1413_bF_buf3), .B(_abc_43815_n2614_1), .Y(_abc_43815_n2615) );
  OR2X2 OR2X2_716 ( .A(_abc_43815_n2617), .B(_abc_43815_n2591), .Y(_abc_43815_n2618) );
  OR2X2 OR2X2_717 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_31_), .Y(_abc_43815_n2619) );
  OR2X2 OR2X2_718 ( .A(_abc_43815_n2623), .B(_abc_43815_n2622), .Y(_abc_43815_n2624) );
  OR2X2 OR2X2_719 ( .A(_abc_43815_n2627), .B(_abc_43815_n2626), .Y(_abc_43815_n2628) );
  OR2X2 OR2X2_72 ( .A(state_q_1_bF_buf1), .B(alu_p_o_10_), .Y(_abc_43815_n842) );
  OR2X2 OR2X2_720 ( .A(_abc_43815_n2630), .B(_abc_43815_n2631), .Y(_abc_43815_n2632) );
  OR2X2 OR2X2_721 ( .A(_abc_43815_n2634), .B(_abc_43815_n2635), .Y(_abc_43815_n2636) );
  OR2X2 OR2X2_722 ( .A(_abc_43815_n2638_1), .B(_abc_43815_n2639), .Y(_abc_43815_n2640) );
  OR2X2 OR2X2_723 ( .A(_abc_43815_n2642), .B(_abc_43815_n2643), .Y(_abc_43815_n2644) );
  OR2X2 OR2X2_724 ( .A(_abc_43815_n2646), .B(_abc_43815_n2647), .Y(_abc_43815_n2648) );
  OR2X2 OR2X2_725 ( .A(_abc_43815_n2651), .B(_abc_43815_n2650), .Y(_abc_43815_n2652) );
  OR2X2 OR2X2_726 ( .A(_abc_43815_n1348), .B(_abc_43815_n1273), .Y(_abc_43815_n2654) );
  OR2X2 OR2X2_727 ( .A(_abc_43815_n1718), .B(_abc_43815_n2654), .Y(_abc_43815_n2655) );
  OR2X2 OR2X2_728 ( .A(_abc_43815_n2657), .B(_abc_43815_n634), .Y(_abc_43815_n2658) );
  OR2X2 OR2X2_729 ( .A(_abc_43815_n2656), .B(_abc_43815_n2658), .Y(pc_q_8__FF_INPUT) );
  OR2X2 OR2X2_73 ( .A(_abc_43815_n693), .B(\mem_dat_i[10] ), .Y(_abc_43815_n843) );
  OR2X2 OR2X2_730 ( .A(_abc_43815_n1761), .B(_abc_43815_n1413_bF_buf2), .Y(_abc_43815_n2660) );
  OR2X2 OR2X2_731 ( .A(_abc_43815_n2662_1), .B(_abc_43815_n1190), .Y(_abc_43815_n2663) );
  OR2X2 OR2X2_732 ( .A(_abc_43815_n2663), .B(_abc_43815_n1278_bF_buf0), .Y(_abc_43815_n2664) );
  OR2X2 OR2X2_733 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(pc_q_9_), .Y(_abc_43815_n2665) );
  OR2X2 OR2X2_734 ( .A(_abc_43815_n2668), .B(_abc_43815_n1273), .Y(_abc_43815_n2669) );
  OR2X2 OR2X2_735 ( .A(_abc_43815_n2670), .B(_abc_43815_n2671), .Y(_abc_43815_n2672) );
  OR2X2 OR2X2_736 ( .A(_abc_43815_n2676), .B(_abc_43815_n1278_bF_buf6), .Y(_abc_43815_n2677) );
  OR2X2 OR2X2_737 ( .A(_abc_43815_n2674), .B(_abc_43815_n2677), .Y(_abc_43815_n2678) );
  OR2X2 OR2X2_738 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(pc_q_11_), .Y(_abc_43815_n2679) );
  OR2X2 OR2X2_739 ( .A(_abc_43815_n2682), .B(_abc_43815_n2683), .Y(_abc_43815_n2684) );
  OR2X2 OR2X2_74 ( .A(_abc_43815_n692_bF_buf0), .B(_abc_43815_n737), .Y(_abc_43815_n844) );
  OR2X2 OR2X2_740 ( .A(_abc_43815_n2686_1), .B(_abc_43815_n2687), .Y(_abc_43815_n2688) );
  OR2X2 OR2X2_741 ( .A(_abc_43815_n2690), .B(_abc_43815_n2691), .Y(_abc_43815_n2692) );
  OR2X2 OR2X2_742 ( .A(_abc_43815_n2694), .B(_abc_43815_n2695), .Y(_abc_43815_n2696) );
  OR2X2 OR2X2_743 ( .A(_abc_43815_n2698), .B(_abc_43815_n2699), .Y(_abc_43815_n2700) );
  OR2X2 OR2X2_744 ( .A(_abc_43815_n2702), .B(_abc_43815_n2703), .Y(_abc_43815_n2704) );
  OR2X2 OR2X2_745 ( .A(_abc_43815_n2706), .B(_abc_43815_n2707), .Y(_abc_43815_n2708) );
  OR2X2 OR2X2_746 ( .A(_abc_43815_n2710_1), .B(_abc_43815_n2711), .Y(_abc_43815_n2712) );
  OR2X2 OR2X2_747 ( .A(_abc_43815_n2714), .B(_abc_43815_n2715), .Y(_abc_43815_n2716) );
  OR2X2 OR2X2_748 ( .A(_abc_43815_n2718), .B(_abc_43815_n2719), .Y(_abc_43815_n2720) );
  OR2X2 OR2X2_749 ( .A(_abc_43815_n2722), .B(_abc_43815_n2723), .Y(_abc_43815_n2724) );
  OR2X2 OR2X2_75 ( .A(_abc_43815_n846), .B(_abc_43815_n832_1_bF_buf1), .Y(_abc_43815_n847) );
  OR2X2 OR2X2_750 ( .A(_abc_43815_n2726), .B(_abc_43815_n2727), .Y(_abc_43815_n2728) );
  OR2X2 OR2X2_751 ( .A(_abc_43815_n2730), .B(_abc_43815_n2731), .Y(_abc_43815_n2732) );
  OR2X2 OR2X2_752 ( .A(_abc_43815_n2734_1), .B(_abc_43815_n2735), .Y(_abc_43815_n2736) );
  OR2X2 OR2X2_753 ( .A(_abc_43815_n2738), .B(_abc_43815_n2739), .Y(_abc_43815_n2740) );
  OR2X2 OR2X2_754 ( .A(_abc_43815_n2742), .B(_abc_43815_n2743), .Y(_abc_43815_n2744) );
  OR2X2 OR2X2_755 ( .A(_abc_43815_n2746), .B(_abc_43815_n2747), .Y(_abc_43815_n2748) );
  OR2X2 OR2X2_756 ( .A(_abc_43815_n2750), .B(_abc_43815_n2751), .Y(_abc_43815_n2752) );
  OR2X2 OR2X2_757 ( .A(_abc_43815_n2755), .B(_abc_43815_n2754), .Y(_abc_43815_n2756) );
  OR2X2 OR2X2_758 ( .A(_abc_43815_n2758_1), .B(_abc_43815_n2759_1), .Y(_abc_43815_n2760) );
  OR2X2 OR2X2_759 ( .A(_abc_43815_n1177), .B(_abc_43815_n1183), .Y(_abc_43815_n2763) );
  OR2X2 OR2X2_76 ( .A(state_q_1_bF_buf0), .B(alu_p_o_11_), .Y(_abc_43815_n849_1) );
  OR2X2 OR2X2_760 ( .A(_abc_43815_n2763), .B(_abc_43815_n1171_bF_buf4), .Y(_abc_43815_n2764) );
  OR2X2 OR2X2_761 ( .A(_abc_43815_n2762), .B(_abc_43815_n2764), .Y(_abc_43815_n2765) );
  OR2X2 OR2X2_762 ( .A(_abc_43815_n2766), .B(_abc_43815_n2767), .Y(_abc_43815_n2768) );
  OR2X2 OR2X2_763 ( .A(_abc_43815_n2772), .B(_abc_43815_n1050), .Y(_abc_43815_n2773) );
  OR2X2 OR2X2_764 ( .A(_abc_43815_n1056), .B(_abc_43815_n1134), .Y(_abc_43815_n2774) );
  OR2X2 OR2X2_765 ( .A(_abc_43815_n1044), .B(_abc_43815_n1060_bF_buf2), .Y(_abc_43815_n2776) );
  OR2X2 OR2X2_766 ( .A(_abc_43815_n2776), .B(_abc_43815_n2775), .Y(_abc_43815_n2777) );
  OR2X2 OR2X2_767 ( .A(_abc_43815_n2777), .B(_abc_43815_n2774), .Y(_abc_43815_n2778) );
  OR2X2 OR2X2_768 ( .A(_abc_43815_n2778), .B(_abc_43815_n2773), .Y(_abc_43815_n2779) );
  OR2X2 OR2X2_769 ( .A(_abc_43815_n2765), .B(_abc_43815_n2779), .Y(_abc_43815_n2780) );
  OR2X2 OR2X2_77 ( .A(_abc_43815_n693), .B(\mem_dat_i[11] ), .Y(_abc_43815_n850) );
  OR2X2 OR2X2_770 ( .A(_abc_43815_n2785_1), .B(_abc_43815_n2783), .Y(_abc_43815_n2786) );
  OR2X2 OR2X2_771 ( .A(_abc_43815_n1124), .B(_abc_43815_n1138), .Y(_abc_43815_n2789) );
  OR2X2 OR2X2_772 ( .A(_abc_43815_n2790), .B(_abc_43815_n1159), .Y(_abc_43815_n2791) );
  OR2X2 OR2X2_773 ( .A(_abc_43815_n2791), .B(_abc_43815_n2788), .Y(_abc_43815_n2792) );
  OR2X2 OR2X2_774 ( .A(_abc_43815_n2792), .B(_abc_43815_n2786), .Y(_abc_43815_n2793) );
  OR2X2 OR2X2_775 ( .A(_abc_43815_n1264), .B(_abc_43815_n1239), .Y(_abc_43815_n2794) );
  OR2X2 OR2X2_776 ( .A(_abc_43815_n2794), .B(_abc_43815_n1417), .Y(_abc_43815_n2795) );
  OR2X2 OR2X2_777 ( .A(_abc_43815_n2796), .B(_abc_43815_n2793), .Y(_abc_43815_n2797) );
  OR2X2 OR2X2_778 ( .A(_abc_43815_n2780), .B(_abc_43815_n2797), .Y(_abc_43815_n2798) );
  OR2X2 OR2X2_779 ( .A(_abc_43815_n2799), .B(_abc_43815_n1171_bF_buf3), .Y(ex_rd_q_0__FF_INPUT) );
  OR2X2 OR2X2_78 ( .A(_abc_43815_n692_bF_buf3), .B(_abc_43815_n753_1), .Y(_abc_43815_n851) );
  OR2X2 OR2X2_780 ( .A(_abc_43815_n2805), .B(_abc_43815_n1171_bF_buf2), .Y(ex_rd_q_3__FF_INPUT) );
  OR2X2 OR2X2_781 ( .A(_abc_43815_n1183), .B(_abc_43815_n2775), .Y(_abc_43815_n2809) );
  OR2X2 OR2X2_782 ( .A(_abc_43815_n1056), .B(_abc_43815_n1044), .Y(_abc_43815_n2810_1) );
  OR2X2 OR2X2_783 ( .A(_abc_43815_n984), .B(_abc_43815_n1050), .Y(_abc_43815_n2811_1) );
  OR2X2 OR2X2_784 ( .A(_abc_43815_n2810_1), .B(_abc_43815_n2811_1), .Y(_abc_43815_n2812) );
  OR2X2 OR2X2_785 ( .A(_abc_43815_n2812), .B(_abc_43815_n2809), .Y(_abc_43815_n2813) );
  OR2X2 OR2X2_786 ( .A(_abc_43815_n2815), .B(_abc_43815_n1177), .Y(_abc_43815_n2816) );
  OR2X2 OR2X2_787 ( .A(_abc_43815_n2816), .B(_abc_43815_n986_bF_buf3), .Y(_abc_43815_n2817) );
  OR2X2 OR2X2_788 ( .A(_abc_43815_n2793), .B(_abc_43815_n2817), .Y(_abc_43815_n2818) );
  OR2X2 OR2X2_789 ( .A(_abc_43815_n2819), .B(_abc_43815_n2814), .Y(alu_input_b_r_0_) );
  OR2X2 OR2X2_79 ( .A(_abc_43815_n853), .B(_abc_43815_n832_1_bF_buf0), .Y(_abc_43815_n854) );
  OR2X2 OR2X2_790 ( .A(_abc_43815_n2822), .B(_abc_43815_n2821), .Y(alu_input_b_r_1_) );
  OR2X2 OR2X2_791 ( .A(_abc_43815_n2825), .B(_abc_43815_n2824), .Y(alu_input_b_r_2_) );
  OR2X2 OR2X2_792 ( .A(_abc_43815_n2828), .B(_abc_43815_n2827), .Y(alu_input_b_r_3_) );
  OR2X2 OR2X2_793 ( .A(_abc_43815_n2831), .B(_abc_43815_n2830), .Y(alu_input_b_r_4_) );
  OR2X2 OR2X2_794 ( .A(_abc_43815_n2834), .B(_abc_43815_n2833), .Y(alu_input_b_r_5_) );
  OR2X2 OR2X2_795 ( .A(_abc_43815_n2837_1), .B(_abc_43815_n2836_1), .Y(_abc_43815_n2838) );
  OR2X2 OR2X2_796 ( .A(_abc_43815_n2786), .B(_abc_43815_n1159), .Y(_abc_43815_n2839) );
  OR2X2 OR2X2_797 ( .A(_abc_43815_n2839), .B(_abc_43815_n2816), .Y(_abc_43815_n2840) );
  OR2X2 OR2X2_798 ( .A(_abc_43815_n2841), .B(_abc_43815_n2838), .Y(alu_input_b_r_6_) );
  OR2X2 OR2X2_799 ( .A(_abc_43815_n2844), .B(_abc_43815_n2843), .Y(_abc_43815_n2845) );
  OR2X2 OR2X2_8 ( .A(_abc_43815_n680_1_bF_buf4), .B(_abc_43815_n677), .Y(_abc_27555_n353) );
  OR2X2 OR2X2_80 ( .A(state_q_1_bF_buf4), .B(alu_p_o_12_), .Y(_abc_43815_n856) );
  OR2X2 OR2X2_800 ( .A(_abc_43815_n2846), .B(_abc_43815_n2845), .Y(alu_input_b_r_7_) );
  OR2X2 OR2X2_801 ( .A(_abc_43815_n2849), .B(_abc_43815_n2848), .Y(_abc_43815_n2850) );
  OR2X2 OR2X2_802 ( .A(_abc_43815_n2851), .B(_abc_43815_n2850), .Y(alu_input_b_r_8_) );
  OR2X2 OR2X2_803 ( .A(_abc_43815_n2854), .B(_abc_43815_n2853), .Y(_abc_43815_n2855) );
  OR2X2 OR2X2_804 ( .A(_abc_43815_n2856), .B(_abc_43815_n2855), .Y(alu_input_b_r_9_) );
  OR2X2 OR2X2_805 ( .A(_abc_43815_n2859), .B(_abc_43815_n2858), .Y(_abc_43815_n2860) );
  OR2X2 OR2X2_806 ( .A(_abc_43815_n2861), .B(_abc_43815_n2860), .Y(alu_input_b_r_10_) );
  OR2X2 OR2X2_807 ( .A(_abc_43815_n2864), .B(_abc_43815_n2863_1), .Y(_abc_43815_n2865) );
  OR2X2 OR2X2_808 ( .A(_abc_43815_n2866), .B(_abc_43815_n2865), .Y(alu_input_b_r_11_) );
  OR2X2 OR2X2_809 ( .A(_abc_43815_n2869), .B(_abc_43815_n2868), .Y(_abc_43815_n2870) );
  OR2X2 OR2X2_81 ( .A(_abc_43815_n693), .B(\mem_dat_i[12] ), .Y(_abc_43815_n857) );
  OR2X2 OR2X2_810 ( .A(_abc_43815_n2871), .B(_abc_43815_n2870), .Y(alu_input_b_r_12_) );
  OR2X2 OR2X2_811 ( .A(_abc_43815_n2874), .B(_abc_43815_n2873), .Y(_abc_43815_n2875) );
  OR2X2 OR2X2_812 ( .A(_abc_43815_n2876), .B(_abc_43815_n2875), .Y(alu_input_b_r_13_) );
  OR2X2 OR2X2_813 ( .A(_abc_43815_n2879), .B(_abc_43815_n2878), .Y(_abc_43815_n2880) );
  OR2X2 OR2X2_814 ( .A(_abc_43815_n2881), .B(_abc_43815_n2880), .Y(alu_input_b_r_14_) );
  OR2X2 OR2X2_815 ( .A(_abc_43815_n2884), .B(_abc_43815_n2883), .Y(_abc_43815_n2885) );
  OR2X2 OR2X2_816 ( .A(_abc_43815_n2886), .B(_abc_43815_n2885), .Y(alu_input_b_r_15_) );
  OR2X2 OR2X2_817 ( .A(_abc_43815_n2890), .B(_abc_43815_n984), .Y(_abc_43815_n2891) );
  OR2X2 OR2X2_818 ( .A(_abc_43815_n2891), .B(_abc_43815_n2889_1), .Y(_abc_43815_n2892) );
  OR2X2 OR2X2_819 ( .A(_abc_43815_n2893), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2), .Y(_abc_43815_n2894) );
  OR2X2 OR2X2_82 ( .A(_abc_43815_n692_bF_buf2), .B(_abc_43815_n769), .Y(_abc_43815_n858) );
  OR2X2 OR2X2_820 ( .A(_abc_43815_n2895), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2896) );
  OR2X2 OR2X2_821 ( .A(_abc_43815_n2897), .B(_abc_43815_n2896), .Y(alu_input_b_r_16_) );
  OR2X2 OR2X2_822 ( .A(_abc_43815_n2891), .B(_abc_43815_n2899), .Y(_abc_43815_n2900) );
  OR2X2 OR2X2_823 ( .A(_abc_43815_n2901), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2902) );
  OR2X2 OR2X2_824 ( .A(_abc_43815_n2903), .B(_abc_43815_n2902), .Y(alu_input_b_r_17_) );
  OR2X2 OR2X2_825 ( .A(_abc_43815_n2891), .B(_abc_43815_n2905), .Y(_abc_43815_n2906) );
  OR2X2 OR2X2_826 ( .A(_abc_43815_n2907), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2908) );
  OR2X2 OR2X2_827 ( .A(_abc_43815_n2909), .B(_abc_43815_n2908), .Y(alu_input_b_r_18_) );
  OR2X2 OR2X2_828 ( .A(_abc_43815_n2891), .B(_abc_43815_n2911), .Y(_abc_43815_n2912) );
  OR2X2 OR2X2_829 ( .A(_abc_43815_n2913), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2914_1) );
  OR2X2 OR2X2_83 ( .A(_abc_43815_n860), .B(_abc_43815_n832_1_bF_buf3), .Y(_abc_43815_n861) );
  OR2X2 OR2X2_830 ( .A(_abc_43815_n2915_1), .B(_abc_43815_n2914_1), .Y(alu_input_b_r_19_) );
  OR2X2 OR2X2_831 ( .A(_abc_43815_n2891), .B(_abc_43815_n2917), .Y(_abc_43815_n2918) );
  OR2X2 OR2X2_832 ( .A(_abc_43815_n2919), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2920) );
  OR2X2 OR2X2_833 ( .A(_abc_43815_n2921), .B(_abc_43815_n2920), .Y(alu_input_b_r_20_) );
  OR2X2 OR2X2_834 ( .A(_abc_43815_n2891), .B(_abc_43815_n2923), .Y(_abc_43815_n2924) );
  OR2X2 OR2X2_835 ( .A(_abc_43815_n2925), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2926) );
  OR2X2 OR2X2_836 ( .A(_abc_43815_n2927), .B(_abc_43815_n2926), .Y(alu_input_b_r_21_) );
  OR2X2 OR2X2_837 ( .A(_abc_43815_n2891), .B(_abc_43815_n2929), .Y(_abc_43815_n2930) );
  OR2X2 OR2X2_838 ( .A(_abc_43815_n2931), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2932) );
  OR2X2 OR2X2_839 ( .A(_abc_43815_n2933), .B(_abc_43815_n2932), .Y(alu_input_b_r_22_) );
  OR2X2 OR2X2_84 ( .A(state_q_1_bF_buf3), .B(alu_p_o_13_), .Y(_abc_43815_n863) );
  OR2X2 OR2X2_840 ( .A(_abc_43815_n2891), .B(_abc_43815_n2935), .Y(_abc_43815_n2936) );
  OR2X2 OR2X2_841 ( .A(_abc_43815_n2937), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2938) );
  OR2X2 OR2X2_842 ( .A(_abc_43815_n2939), .B(_abc_43815_n2938), .Y(alu_input_b_r_23_) );
  OR2X2 OR2X2_843 ( .A(_abc_43815_n2891), .B(_abc_43815_n2941_1), .Y(_abc_43815_n2942) );
  OR2X2 OR2X2_844 ( .A(_abc_43815_n2943), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2944) );
  OR2X2 OR2X2_845 ( .A(_abc_43815_n2945), .B(_abc_43815_n2944), .Y(alu_input_b_r_24_) );
  OR2X2 OR2X2_846 ( .A(_abc_43815_n2891), .B(_abc_43815_n2947), .Y(_abc_43815_n2948) );
  OR2X2 OR2X2_847 ( .A(_abc_43815_n2949), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2950) );
  OR2X2 OR2X2_848 ( .A(_abc_43815_n2951), .B(_abc_43815_n2950), .Y(alu_input_b_r_25_) );
  OR2X2 OR2X2_849 ( .A(_abc_43815_n2891), .B(_abc_43815_n2953), .Y(_abc_43815_n2954) );
  OR2X2 OR2X2_85 ( .A(_abc_43815_n693), .B(\mem_dat_i[13] ), .Y(_abc_43815_n864) );
  OR2X2 OR2X2_850 ( .A(_abc_43815_n2955), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2956) );
  OR2X2 OR2X2_851 ( .A(_abc_43815_n2957), .B(_abc_43815_n2956), .Y(alu_input_b_r_26_) );
  OR2X2 OR2X2_852 ( .A(_abc_43815_n2891), .B(_abc_43815_n2959), .Y(_abc_43815_n2960) );
  OR2X2 OR2X2_853 ( .A(_abc_43815_n2961), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2962) );
  OR2X2 OR2X2_854 ( .A(_abc_43815_n2963), .B(_abc_43815_n2962), .Y(alu_input_b_r_27_) );
  OR2X2 OR2X2_855 ( .A(_abc_43815_n2891), .B(_abc_43815_n2965), .Y(_abc_43815_n2966_1) );
  OR2X2 OR2X2_856 ( .A(_abc_43815_n2967_1), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2968) );
  OR2X2 OR2X2_857 ( .A(_abc_43815_n2969), .B(_abc_43815_n2968), .Y(alu_input_b_r_28_) );
  OR2X2 OR2X2_858 ( .A(_abc_43815_n2891), .B(_abc_43815_n2971), .Y(_abc_43815_n2972) );
  OR2X2 OR2X2_859 ( .A(_abc_43815_n2973), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2974) );
  OR2X2 OR2X2_86 ( .A(_abc_43815_n692_bF_buf1), .B(_abc_43815_n785), .Y(_abc_43815_n865_1) );
  OR2X2 OR2X2_860 ( .A(_abc_43815_n2975), .B(_abc_43815_n2974), .Y(alu_input_b_r_29_) );
  OR2X2 OR2X2_861 ( .A(_abc_43815_n2891), .B(_abc_43815_n2977), .Y(_abc_43815_n2978) );
  OR2X2 OR2X2_862 ( .A(_abc_43815_n2979), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2980) );
  OR2X2 OR2X2_863 ( .A(_abc_43815_n2981), .B(_abc_43815_n2980), .Y(alu_input_b_r_30_) );
  OR2X2 OR2X2_864 ( .A(_abc_43815_n2891), .B(_abc_43815_n2983), .Y(_abc_43815_n2984) );
  OR2X2 OR2X2_865 ( .A(_abc_43815_n2985), .B(_abc_43815_n2888_1), .Y(_abc_43815_n2986) );
  OR2X2 OR2X2_866 ( .A(_abc_43815_n2987), .B(_abc_43815_n2986), .Y(alu_input_b_r_31_) );
  OR2X2 OR2X2_867 ( .A(_abc_43815_n1044), .B(_abc_43815_n1050), .Y(_abc_43815_n2989) );
  OR2X2 OR2X2_868 ( .A(_abc_43815_n987), .B(_abc_43815_n2989), .Y(_abc_43815_n2990) );
  OR2X2 OR2X2_869 ( .A(_abc_43815_n2990), .B(_abc_43815_n2809), .Y(_abc_43815_n2991) );
  OR2X2 OR2X2_87 ( .A(_abc_43815_n867), .B(_abc_43815_n832_1_bF_buf2), .Y(_abc_43815_n868_1) );
  OR2X2 OR2X2_870 ( .A(_abc_43815_n2994), .B(_abc_43815_n1171_bF_buf1), .Y(_abc_43815_n2995) );
  OR2X2 OR2X2_871 ( .A(_abc_43815_n2995), .B(_abc_43815_n2992_1), .Y(_abc_43815_n2996) );
  OR2X2 OR2X2_872 ( .A(_abc_43815_n1172_1_bF_buf4), .B(next_pc_r_0_), .Y(_abc_43815_n2997) );
  OR2X2 OR2X2_873 ( .A(_abc_43815_n2786), .B(_abc_43815_n2774), .Y(alu_func_r_2_) );
  OR2X2 OR2X2_874 ( .A(_abc_43815_n2792), .B(_abc_43815_n1177), .Y(_abc_43815_n3001) );
  OR2X2 OR2X2_875 ( .A(_abc_43815_n3001), .B(alu_func_r_2_), .Y(_abc_43815_n3002) );
  OR2X2 OR2X2_876 ( .A(_abc_43815_n2999), .B(_abc_43815_n3003), .Y(alu_input_a_r_0_) );
  OR2X2 OR2X2_877 ( .A(_abc_43815_n3006), .B(_abc_43815_n1171_bF_buf0), .Y(_abc_43815_n3007) );
  OR2X2 OR2X2_878 ( .A(_abc_43815_n3007), .B(_abc_43815_n3005), .Y(_abc_43815_n3008) );
  OR2X2 OR2X2_879 ( .A(_abc_43815_n1172_1_bF_buf3), .B(next_pc_r_1_), .Y(_abc_43815_n3009) );
  OR2X2 OR2X2_88 ( .A(_abc_43815_n870), .B(_abc_43815_n871), .Y(_abc_43815_n872) );
  OR2X2 OR2X2_880 ( .A(_abc_43815_n3011), .B(_abc_43815_n3012), .Y(alu_input_a_r_1_) );
  OR2X2 OR2X2_881 ( .A(_abc_43815_n3014), .B(_abc_43815_n1171_bF_buf5), .Y(_abc_43815_n3015) );
  OR2X2 OR2X2_882 ( .A(_abc_43815_n3017), .B(_abc_43815_n3018_1), .Y(_abc_43815_n3019_1) );
  OR2X2 OR2X2_883 ( .A(_abc_43815_n3016), .B(_abc_43815_n3019_1), .Y(_abc_43815_n3020) );
  OR2X2 OR2X2_884 ( .A(_abc_43815_n3021), .B(_abc_43815_n3015), .Y(_abc_43815_n3022) );
  OR2X2 OR2X2_885 ( .A(_abc_43815_n1172_1_bF_buf2), .B(_abc_43815_n1485), .Y(_abc_43815_n3023) );
  OR2X2 OR2X2_886 ( .A(_abc_43815_n3024), .B(_abc_43815_n3025), .Y(alu_input_a_r_2_) );
  OR2X2 OR2X2_887 ( .A(_abc_43815_n3028), .B(_abc_43815_n1171_bF_buf4), .Y(_abc_43815_n3029) );
  OR2X2 OR2X2_888 ( .A(_abc_43815_n3029), .B(_abc_43815_n3027), .Y(_abc_43815_n3030) );
  OR2X2 OR2X2_889 ( .A(_abc_43815_n1172_1_bF_buf1), .B(_abc_43815_n1526), .Y(_abc_43815_n3031) );
  OR2X2 OR2X2_89 ( .A(_abc_43815_n873), .B(_abc_43815_n832_1_bF_buf1), .Y(_abc_43815_n874) );
  OR2X2 OR2X2_890 ( .A(_abc_43815_n3033), .B(_abc_43815_n3034), .Y(alu_input_a_r_3_) );
  OR2X2 OR2X2_891 ( .A(_abc_43815_n3037), .B(_abc_43815_n1171_bF_buf3), .Y(_abc_43815_n3038) );
  OR2X2 OR2X2_892 ( .A(_abc_43815_n3038), .B(_abc_43815_n3036), .Y(_abc_43815_n3039) );
  OR2X2 OR2X2_893 ( .A(_abc_43815_n1172_1_bF_buf0), .B(_abc_43815_n1563), .Y(_abc_43815_n3040) );
  OR2X2 OR2X2_894 ( .A(_abc_43815_n3042), .B(_abc_43815_n3043), .Y(alu_input_a_r_4_) );
  OR2X2 OR2X2_895 ( .A(_abc_43815_n3046), .B(_abc_43815_n1171_bF_buf2), .Y(_abc_43815_n3047) );
  OR2X2 OR2X2_896 ( .A(_abc_43815_n3047), .B(_abc_43815_n3045_1), .Y(_abc_43815_n3048) );
  OR2X2 OR2X2_897 ( .A(_abc_43815_n1172_1_bF_buf4), .B(_abc_43815_n1603_1), .Y(_abc_43815_n3049) );
  OR2X2 OR2X2_898 ( .A(_abc_43815_n3051), .B(_abc_43815_n3052), .Y(alu_input_a_r_5_) );
  OR2X2 OR2X2_899 ( .A(_abc_43815_n3055), .B(_abc_43815_n1171_bF_buf1), .Y(_abc_43815_n3056) );
  OR2X2 OR2X2_9 ( .A(_abc_43815_n684), .B(_abc_43815_n660), .Y(_abc_43815_n685) );
  OR2X2 OR2X2_90 ( .A(state_q_1_bF_buf2), .B(alu_p_o_14_), .Y(_abc_43815_n875) );
  OR2X2 OR2X2_900 ( .A(_abc_43815_n3056), .B(_abc_43815_n3054), .Y(_abc_43815_n3057) );
  OR2X2 OR2X2_901 ( .A(_abc_43815_n1635_1), .B(_abc_43815_n1172_1_bF_buf3), .Y(_abc_43815_n3058) );
  OR2X2 OR2X2_902 ( .A(_abc_43815_n3060), .B(_abc_43815_n3061), .Y(alu_input_a_r_6_) );
  OR2X2 OR2X2_903 ( .A(_abc_43815_n3064), .B(_abc_43815_n1171_bF_buf0), .Y(_abc_43815_n3065) );
  OR2X2 OR2X2_904 ( .A(_abc_43815_n3065), .B(_abc_43815_n3063), .Y(_abc_43815_n3066) );
  OR2X2 OR2X2_905 ( .A(_abc_43815_n1680), .B(_abc_43815_n1172_1_bF_buf2), .Y(_abc_43815_n3067) );
  OR2X2 OR2X2_906 ( .A(_abc_43815_n3069), .B(_abc_43815_n3070_1), .Y(alu_input_a_r_7_) );
  OR2X2 OR2X2_907 ( .A(_abc_43815_n3072), .B(_abc_43815_n3073), .Y(_abc_43815_n3074) );
  OR2X2 OR2X2_908 ( .A(_abc_43815_n3074), .B(_abc_43815_n3075), .Y(_abc_43815_n3076) );
  OR2X2 OR2X2_909 ( .A(_abc_43815_n3077), .B(_abc_43815_n3076), .Y(alu_input_a_r_8_) );
  OR2X2 OR2X2_91 ( .A(state_q_1_bF_buf1), .B(alu_p_o_15_), .Y(_abc_43815_n877) );
  OR2X2 OR2X2_910 ( .A(_abc_43815_n3079), .B(_abc_43815_n1171_bF_buf4), .Y(_abc_43815_n3080) );
  OR2X2 OR2X2_911 ( .A(_abc_43815_n3082), .B(_abc_43815_n3083), .Y(_abc_43815_n3084) );
  OR2X2 OR2X2_912 ( .A(_abc_43815_n3081), .B(_abc_43815_n3084), .Y(_abc_43815_n3085) );
  OR2X2 OR2X2_913 ( .A(_abc_43815_n3086), .B(_abc_43815_n3080), .Y(_abc_43815_n3087) );
  OR2X2 OR2X2_914 ( .A(_abc_43815_n1733), .B(_abc_43815_n1172_1_bF_buf1), .Y(_abc_43815_n3088) );
  OR2X2 OR2X2_915 ( .A(_abc_43815_n3089), .B(_abc_43815_n3090), .Y(alu_input_a_r_9_) );
  OR2X2 OR2X2_916 ( .A(_abc_43815_n3092), .B(_abc_43815_n1171_bF_buf3), .Y(_abc_43815_n3093) );
  OR2X2 OR2X2_917 ( .A(_abc_43815_n3095), .B(_abc_43815_n3096_1), .Y(_abc_43815_n3097_1) );
  OR2X2 OR2X2_918 ( .A(_abc_43815_n3094), .B(_abc_43815_n3097_1), .Y(_abc_43815_n3098) );
  OR2X2 OR2X2_919 ( .A(_abc_43815_n3099), .B(_abc_43815_n3093), .Y(_abc_43815_n3100) );
  OR2X2 OR2X2_92 ( .A(_abc_43815_n693), .B(\mem_dat_i[15] ), .Y(_abc_43815_n878) );
  OR2X2 OR2X2_920 ( .A(_abc_43815_n1772), .B(_abc_43815_n1172_1_bF_buf0), .Y(_abc_43815_n3101) );
  OR2X2 OR2X2_921 ( .A(_abc_43815_n3102), .B(_abc_43815_n3103), .Y(alu_input_a_r_10_) );
  OR2X2 OR2X2_922 ( .A(_abc_43815_n3105), .B(_abc_43815_n3106), .Y(_abc_43815_n3107) );
  OR2X2 OR2X2_923 ( .A(_abc_43815_n3108), .B(_abc_43815_n3107), .Y(_abc_43815_n3109) );
  OR2X2 OR2X2_924 ( .A(_abc_43815_n3109), .B(_abc_43815_n3110), .Y(alu_input_a_r_11_) );
  OR2X2 OR2X2_925 ( .A(_abc_43815_n3112), .B(_abc_43815_n3113), .Y(_abc_43815_n3114) );
  OR2X2 OR2X2_926 ( .A(_abc_43815_n3115), .B(_abc_43815_n3114), .Y(_abc_43815_n3116) );
  OR2X2 OR2X2_927 ( .A(_abc_43815_n3116), .B(_abc_43815_n3117), .Y(alu_input_a_r_12_) );
  OR2X2 OR2X2_928 ( .A(_abc_43815_n3119), .B(_abc_43815_n3120), .Y(_abc_43815_n3121) );
  OR2X2 OR2X2_929 ( .A(_abc_43815_n3122_1), .B(_abc_43815_n3121), .Y(_abc_43815_n3123_1) );
  OR2X2 OR2X2_93 ( .A(_abc_43815_n692_bF_buf0), .B(_abc_43815_n812), .Y(_abc_43815_n879) );
  OR2X2 OR2X2_930 ( .A(_abc_43815_n3123_1), .B(_abc_43815_n3124), .Y(alu_input_a_r_13_) );
  OR2X2 OR2X2_931 ( .A(_abc_43815_n3126), .B(_abc_43815_n3127), .Y(_abc_43815_n3128) );
  OR2X2 OR2X2_932 ( .A(_abc_43815_n3129), .B(_abc_43815_n3128), .Y(_abc_43815_n3130) );
  OR2X2 OR2X2_933 ( .A(_abc_43815_n3130), .B(_abc_43815_n3131), .Y(alu_input_a_r_14_) );
  OR2X2 OR2X2_934 ( .A(_abc_43815_n1969), .B(_abc_43815_n1172_1_bF_buf4), .Y(_abc_43815_n3133) );
  OR2X2 OR2X2_935 ( .A(_abc_43815_n3135), .B(_abc_43815_n1171_bF_buf4), .Y(_abc_43815_n3136) );
  OR2X2 OR2X2_936 ( .A(_abc_43815_n3136), .B(_abc_43815_n3134), .Y(_abc_43815_n3137) );
  OR2X2 OR2X2_937 ( .A(_abc_43815_n3138), .B(_abc_43815_n3139), .Y(alu_input_a_r_15_) );
  OR2X2 OR2X2_938 ( .A(_abc_43815_n2005), .B(_abc_43815_n1172_1_bF_buf3), .Y(_abc_43815_n3141) );
  OR2X2 OR2X2_939 ( .A(_abc_43815_n1171_bF_buf3), .B(_abc_43815_n3144), .Y(_abc_43815_n3145) );
  OR2X2 OR2X2_94 ( .A(_abc_43815_n881), .B(_abc_43815_n832_1_bF_buf0), .Y(_abc_43815_n882) );
  OR2X2 OR2X2_940 ( .A(_abc_43815_n3143), .B(_abc_43815_n3145), .Y(_abc_43815_n3146) );
  OR2X2 OR2X2_941 ( .A(_abc_43815_n3146), .B(_abc_43815_n3142), .Y(_abc_43815_n3147) );
  OR2X2 OR2X2_942 ( .A(_abc_43815_n3148_1), .B(_abc_43815_n3149_1), .Y(alu_input_a_r_16_) );
  OR2X2 OR2X2_943 ( .A(_abc_43815_n2050), .B(_abc_43815_n1172_1_bF_buf2), .Y(_abc_43815_n3151) );
  OR2X2 OR2X2_944 ( .A(_abc_43815_n1171_bF_buf2), .B(_abc_43815_n3154), .Y(_abc_43815_n3155) );
  OR2X2 OR2X2_945 ( .A(_abc_43815_n3153), .B(_abc_43815_n3155), .Y(_abc_43815_n3156) );
  OR2X2 OR2X2_946 ( .A(_abc_43815_n3156), .B(_abc_43815_n3152), .Y(_abc_43815_n3157) );
  OR2X2 OR2X2_947 ( .A(_abc_43815_n3158), .B(_abc_43815_n3159), .Y(alu_input_a_r_17_) );
  OR2X2 OR2X2_948 ( .A(_abc_43815_n3161), .B(_abc_43815_n3162), .Y(_abc_43815_n3163) );
  OR2X2 OR2X2_949 ( .A(_abc_43815_n3163), .B(_abc_43815_n3164), .Y(_abc_43815_n3165) );
  OR2X2 OR2X2_95 ( .A(_abc_43815_n886), .B(_abc_43815_n885_1), .Y(_abc_43815_n887) );
  OR2X2 OR2X2_950 ( .A(_abc_43815_n3166), .B(_abc_43815_n3165), .Y(_abc_43815_n3167) );
  OR2X2 OR2X2_951 ( .A(_abc_43815_n3167), .B(_abc_43815_n3168), .Y(alu_input_a_r_18_) );
  OR2X2 OR2X2_952 ( .A(_abc_43815_n3172), .B(_abc_43815_n3171), .Y(_abc_43815_n3173) );
  OR2X2 OR2X2_953 ( .A(_abc_43815_n3173), .B(_abc_43815_n3170), .Y(_abc_43815_n3174_1) );
  OR2X2 OR2X2_954 ( .A(_abc_43815_n3175), .B(_abc_43815_n3174_1), .Y(_abc_43815_n3176) );
  OR2X2 OR2X2_955 ( .A(_abc_43815_n3176), .B(_abc_43815_n3177), .Y(alu_input_a_r_19_) );
  OR2X2 OR2X2_956 ( .A(_abc_43815_n2162), .B(_abc_43815_n1172_1_bF_buf1), .Y(_abc_43815_n3179) );
  OR2X2 OR2X2_957 ( .A(_abc_43815_n1171_bF_buf5), .B(_abc_43815_n3182), .Y(_abc_43815_n3183) );
  OR2X2 OR2X2_958 ( .A(_abc_43815_n3181), .B(_abc_43815_n3183), .Y(_abc_43815_n3184) );
  OR2X2 OR2X2_959 ( .A(_abc_43815_n3184), .B(_abc_43815_n3180), .Y(_abc_43815_n3185) );
  OR2X2 OR2X2_96 ( .A(_abc_43815_n888), .B(_abc_43815_n832_1_bF_buf3), .Y(_abc_43815_n889) );
  OR2X2 OR2X2_960 ( .A(_abc_43815_n3186), .B(_abc_43815_n3187), .Y(alu_input_a_r_20_) );
  OR2X2 OR2X2_961 ( .A(_abc_43815_n2205), .B(_abc_43815_n1172_1_bF_buf0), .Y(_abc_43815_n3189) );
  OR2X2 OR2X2_962 ( .A(_abc_43815_n1171_bF_buf4), .B(_abc_43815_n3192), .Y(_abc_43815_n3193_1) );
  OR2X2 OR2X2_963 ( .A(_abc_43815_n3191), .B(_abc_43815_n3193_1), .Y(_abc_43815_n3194) );
  OR2X2 OR2X2_964 ( .A(_abc_43815_n3194), .B(_abc_43815_n3190), .Y(_abc_43815_n3195) );
  OR2X2 OR2X2_965 ( .A(_abc_43815_n3196), .B(_abc_43815_n3197), .Y(alu_input_a_r_21_) );
  OR2X2 OR2X2_966 ( .A(_abc_43815_n2243), .B(_abc_43815_n1172_1_bF_buf4), .Y(_abc_43815_n3199) );
  OR2X2 OR2X2_967 ( .A(_abc_43815_n1171_bF_buf3), .B(_abc_43815_n3202), .Y(_abc_43815_n3203) );
  OR2X2 OR2X2_968 ( .A(_abc_43815_n3201), .B(_abc_43815_n3203), .Y(_abc_43815_n3204) );
  OR2X2 OR2X2_969 ( .A(_abc_43815_n3204), .B(_abc_43815_n3200), .Y(_abc_43815_n3205) );
  OR2X2 OR2X2_97 ( .A(state_q_1_bF_buf0), .B(alu_p_o_16_), .Y(_abc_43815_n890) );
  OR2X2 OR2X2_970 ( .A(_abc_43815_n3206), .B(_abc_43815_n3207), .Y(alu_input_a_r_22_) );
  OR2X2 OR2X2_971 ( .A(_abc_43815_n2279), .B(_abc_43815_n1172_1_bF_buf3), .Y(_abc_43815_n3209_1) );
  OR2X2 OR2X2_972 ( .A(_abc_43815_n1171_bF_buf2), .B(_abc_43815_n3212), .Y(_abc_43815_n3213) );
  OR2X2 OR2X2_973 ( .A(_abc_43815_n3211), .B(_abc_43815_n3213), .Y(_abc_43815_n3214) );
  OR2X2 OR2X2_974 ( .A(_abc_43815_n3214), .B(_abc_43815_n3210), .Y(_abc_43815_n3215) );
  OR2X2 OR2X2_975 ( .A(_abc_43815_n3216), .B(_abc_43815_n3217_1), .Y(alu_input_a_r_23_) );
  OR2X2 OR2X2_976 ( .A(_abc_43815_n2315), .B(_abc_43815_n1172_1_bF_buf2), .Y(_abc_43815_n3219) );
  OR2X2 OR2X2_977 ( .A(_abc_43815_n1171_bF_buf1), .B(_abc_43815_n3222), .Y(_abc_43815_n3223) );
  OR2X2 OR2X2_978 ( .A(_abc_43815_n3221), .B(_abc_43815_n3223), .Y(_abc_43815_n3224) );
  OR2X2 OR2X2_979 ( .A(_abc_43815_n3224), .B(_abc_43815_n3220), .Y(_abc_43815_n3225) );
  OR2X2 OR2X2_98 ( .A(_abc_43815_n892), .B(_abc_43815_n885_1), .Y(_abc_43815_n893) );
  OR2X2 OR2X2_980 ( .A(_abc_43815_n3226), .B(_abc_43815_n3227), .Y(alu_input_a_r_24_) );
  OR2X2 OR2X2_981 ( .A(_abc_43815_n2358), .B(_abc_43815_n1172_1_bF_buf1), .Y(_abc_43815_n3229) );
  OR2X2 OR2X2_982 ( .A(_abc_43815_n1171_bF_buf0), .B(_abc_43815_n3232), .Y(_abc_43815_n3233) );
  OR2X2 OR2X2_983 ( .A(_abc_43815_n3231), .B(_abc_43815_n3233), .Y(_abc_43815_n3234) );
  OR2X2 OR2X2_984 ( .A(_abc_43815_n3234), .B(_abc_43815_n3230), .Y(_abc_43815_n3235_1) );
  OR2X2 OR2X2_985 ( .A(_abc_43815_n3236), .B(_abc_43815_n3237), .Y(alu_input_a_r_25_) );
  OR2X2 OR2X2_986 ( .A(_abc_43815_n2397), .B(_abc_43815_n1172_1_bF_buf0), .Y(_abc_43815_n3239) );
  OR2X2 OR2X2_987 ( .A(_abc_43815_n1171_bF_buf5), .B(_abc_43815_n3242), .Y(_abc_43815_n3243) );
  OR2X2 OR2X2_988 ( .A(_abc_43815_n3241), .B(_abc_43815_n3243), .Y(_abc_43815_n3244_1) );
  OR2X2 OR2X2_989 ( .A(_abc_43815_n3244_1), .B(_abc_43815_n3240), .Y(_abc_43815_n3245) );
  OR2X2 OR2X2_99 ( .A(_abc_43815_n894), .B(_abc_43815_n832_1_bF_buf2), .Y(_abc_43815_n895) );
  OR2X2 OR2X2_990 ( .A(_abc_43815_n3246_1), .B(_abc_43815_n3247), .Y(alu_input_a_r_26_) );
  OR2X2 OR2X2_991 ( .A(_abc_43815_n2434), .B(_abc_43815_n1172_1_bF_buf4), .Y(_abc_43815_n3249) );
  OR2X2 OR2X2_992 ( .A(_abc_43815_n1171_bF_buf4), .B(_abc_43815_n3252_1), .Y(_abc_43815_n3253) );
  OR2X2 OR2X2_993 ( .A(_abc_43815_n3251), .B(_abc_43815_n3253), .Y(_abc_43815_n3254_1) );
  OR2X2 OR2X2_994 ( .A(_abc_43815_n3254_1), .B(_abc_43815_n3250_1), .Y(_abc_43815_n3255) );
  OR2X2 OR2X2_995 ( .A(_abc_43815_n3256_1), .B(_abc_43815_n3257), .Y(alu_input_a_r_27_) );
  OR2X2 OR2X2_996 ( .A(_abc_43815_n2473), .B(_abc_43815_n1172_1_bF_buf3), .Y(_abc_43815_n3259) );
  OR2X2 OR2X2_997 ( .A(_abc_43815_n1171_bF_buf3), .B(_abc_43815_n3262_1), .Y(_abc_43815_n3263) );
  OR2X2 OR2X2_998 ( .A(_abc_43815_n3261), .B(_abc_43815_n3263), .Y(_abc_43815_n3264_1) );
  OR2X2 OR2X2_999 ( .A(_abc_43815_n3264_1), .B(_abc_43815_n3260_1), .Y(_abc_43815_n3265) );
endmodule
